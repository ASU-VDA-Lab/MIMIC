module fake_netlist_1_5120_n_35 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_35);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_35;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
BUFx2_ASAP7_75t_L g10 ( .A(n_1), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
INVx5_ASAP7_75t_L g12 ( .A(n_2), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_1), .Y(n_13) );
BUFx3_ASAP7_75t_L g14 ( .A(n_9), .Y(n_14) );
AOI22xp33_ASAP7_75t_L g15 ( .A1(n_11), .A2(n_0), .B1(n_2), .B2(n_3), .Y(n_15) );
NAND2xp5_ASAP7_75t_SL g16 ( .A(n_12), .B(n_0), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_14), .Y(n_17) );
BUFx2_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
AO21x2_ASAP7_75t_L g19 ( .A1(n_16), .A2(n_13), .B(n_11), .Y(n_19) );
INVx2_ASAP7_75t_SL g20 ( .A(n_18), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_19), .Y(n_21) );
AND2x2_ASAP7_75t_SL g22 ( .A(n_21), .B(n_10), .Y(n_22) );
INVx1_ASAP7_75t_SL g23 ( .A(n_20), .Y(n_23) );
OAI221xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_15), .B1(n_10), .B2(n_21), .C(n_13), .Y(n_24) );
O2A1O1Ixp33_ASAP7_75t_L g25 ( .A1(n_22), .A2(n_17), .B(n_19), .C(n_14), .Y(n_25) );
AOI22xp5_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_22), .B1(n_19), .B2(n_14), .Y(n_26) );
AOI22xp5_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_22), .B1(n_12), .B2(n_5), .Y(n_27) );
AOI21xp33_ASAP7_75t_L g28 ( .A1(n_25), .A2(n_12), .B(n_4), .Y(n_28) );
OAI211xp5_ASAP7_75t_SL g29 ( .A1(n_27), .A2(n_12), .B(n_4), .C(n_5), .Y(n_29) );
AND4x1_ASAP7_75t_L g30 ( .A(n_26), .B(n_3), .C(n_6), .D(n_7), .Y(n_30) );
NAND3xp33_ASAP7_75t_L g31 ( .A(n_28), .B(n_12), .C(n_7), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_29), .Y(n_33) );
NAND2xp5_ASAP7_75t_L g34 ( .A(n_32), .B(n_12), .Y(n_34) );
OAI22xp33_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_33), .B1(n_31), .B2(n_8), .Y(n_35) );
endmodule