module fake_jpeg_28393_n_297 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_175;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx6_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_7),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_19),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_17),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_21),
.B1(n_22),
.B2(n_30),
.Y(n_64)
);

AO22x1_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_16),
.B1(n_21),
.B2(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_49),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_16),
.B1(n_23),
.B2(n_27),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_48),
.A2(n_53),
.B1(n_62),
.B2(n_31),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_22),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_22),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_51),
.B(n_55),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_16),
.B1(n_23),
.B2(n_27),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_36),
.B(n_30),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_22),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_58),
.Y(n_66)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_39),
.A2(n_16),
.B1(n_23),
.B2(n_27),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_48),
.Y(n_89)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_54),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_68),
.Y(n_92)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_69),
.B(n_72),
.Y(n_111)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_45),
.A2(n_21),
.B1(n_20),
.B2(n_26),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_76),
.B1(n_31),
.B2(n_45),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_43),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_53),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_86),
.B(n_58),
.Y(n_94)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_88),
.B1(n_61),
.B2(n_60),
.Y(n_112)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_89),
.A2(n_28),
.B1(n_18),
.B2(n_17),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_80),
.B1(n_84),
.B2(n_75),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_91),
.A2(n_114),
.B1(n_63),
.B2(n_59),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_94),
.B(n_97),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_91),
.B1(n_114),
.B2(n_106),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_43),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_32),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_79),
.B(n_58),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_73),
.B(n_43),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_101),
.A2(n_109),
.B(n_0),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_104),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_20),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_47),
.C(n_50),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_82),
.C(n_78),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_80),
.A2(n_64),
.B(n_44),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_74),
.A2(n_30),
.B(n_24),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_110),
.A2(n_32),
.B(n_25),
.Y(n_140)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_44),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_85),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_65),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_70),
.B1(n_87),
.B2(n_88),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_115),
.A2(n_130),
.B1(n_137),
.B2(n_98),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_138),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_100),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_90),
.B(n_85),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_118),
.A2(n_120),
.B(n_105),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_93),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_119),
.Y(n_144)
);

OA21x2_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_68),
.B(n_40),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_121),
.A2(n_126),
.B1(n_98),
.B2(n_107),
.Y(n_161)
);

OAI32xp33_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_26),
.A3(n_24),
.B1(n_22),
.B2(n_32),
.Y(n_122)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_124),
.B(n_133),
.Y(n_163)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_131),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_111),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_129),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_94),
.A2(n_24),
.B1(n_17),
.B2(n_29),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_25),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_140),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_90),
.A2(n_81),
.B1(n_29),
.B2(n_28),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_81),
.C(n_32),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_110),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_139),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_32),
.C(n_25),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_142),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_146),
.Y(n_177)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_151),
.Y(n_178)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_153),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_120),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_154),
.B(n_155),
.Y(n_197)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_157),
.A2(n_127),
.B1(n_123),
.B2(n_134),
.Y(n_176)
);

XNOR2x1_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_89),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_160),
.A2(n_172),
.B(n_100),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_162),
.B1(n_29),
.B2(n_28),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_123),
.A2(n_106),
.B1(n_97),
.B2(n_109),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_104),
.C(n_25),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_156),
.Y(n_184)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_105),
.Y(n_169)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_170),
.A2(n_99),
.B(n_107),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_128),
.Y(n_171)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_116),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_124),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_186),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_176),
.A2(n_183),
.B1(n_198),
.B2(n_5),
.Y(n_220)
);

OA22x2_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_131),
.B1(n_142),
.B2(n_140),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_179),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_136),
.C(n_141),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_148),
.C(n_156),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_168),
.A2(n_129),
.B1(n_132),
.B2(n_125),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_184),
.B(n_165),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_143),
.A2(n_146),
.B1(n_153),
.B2(n_168),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_185),
.A2(n_191),
.B1(n_155),
.B2(n_159),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_128),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_144),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_159),
.Y(n_208)
);

INVxp33_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_188),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_193),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_190),
.A2(n_192),
.B(n_169),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_143),
.A2(n_99),
.B1(n_102),
.B2(n_29),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_102),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_148),
.B(n_25),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_194),
.A2(n_158),
.B1(n_165),
.B2(n_18),
.Y(n_211)
);

OAI32xp33_ASAP7_75t_L g196 ( 
.A1(n_158),
.A2(n_28),
.A3(n_18),
.B1(n_17),
.B2(n_8),
.Y(n_196)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_196),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_147),
.A2(n_18),
.B1(n_7),
.B2(n_8),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_192),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_209),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_202),
.A2(n_217),
.B(n_183),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_151),
.Y(n_203)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_204),
.A2(n_214),
.B1(n_220),
.B2(n_181),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_219),
.C(n_12),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_178),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_160),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_213),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_191),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_212),
.B(n_193),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_166),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_176),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_6),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_218),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_6),
.B(n_14),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_177),
.B(n_6),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_15),
.C(n_5),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_14),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_205),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_199),
.Y(n_223)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_223),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_200),
.A2(n_190),
.B(n_188),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_225),
.A2(n_231),
.B(n_211),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_226),
.A2(n_230),
.B1(n_234),
.B2(n_239),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_235),
.Y(n_245)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_228),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_204),
.A2(n_173),
.B1(n_197),
.B2(n_175),
.Y(n_230)
);

AO21x1_ASAP7_75t_L g231 ( 
.A1(n_215),
.A2(n_179),
.B(n_185),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_205),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_233),
.B(n_10),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_207),
.A2(n_179),
.B1(n_196),
.B2(n_2),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_179),
.Y(n_235)
);

INVxp33_ASAP7_75t_SL g236 ( 
.A(n_199),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_214),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_219),
.C(n_221),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_240),
.B(n_232),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_247),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_206),
.C(n_201),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_251),
.C(n_237),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_224),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_231),
.A2(n_213),
.B(n_210),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_253),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_223),
.A2(n_201),
.B1(n_1),
.B2(n_2),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_249),
.A2(n_230),
.B1(n_3),
.B2(n_4),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_250),
.A2(n_238),
.B1(n_226),
.B2(n_229),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_10),
.C(n_11),
.Y(n_251)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_251),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_235),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_257),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_258),
.B(n_263),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_252),
.A2(n_234),
.B(n_225),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_260),
.A2(n_248),
.B(n_227),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_262),
.A2(n_249),
.B1(n_246),
.B2(n_242),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_245),
.C(n_240),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_244),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_267),
.A2(n_272),
.B(n_256),
.Y(n_280)
);

INVxp33_ASAP7_75t_L g276 ( 
.A(n_268),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_261),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_258),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_275),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_259),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_274),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_264),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_273),
.A2(n_265),
.B(n_260),
.Y(n_277)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_277),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_280),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_263),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_282),
.B(n_279),
.Y(n_286)
);

NOR2xp67_ASAP7_75t_R g283 ( 
.A(n_267),
.B(n_257),
.Y(n_283)
);

NOR2x1_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_266),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_287),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_271),
.Y(n_288)
);

AOI21x1_ASAP7_75t_SL g289 ( 
.A1(n_288),
.A2(n_276),
.B(n_281),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_289),
.Y(n_292)
);

NAND2x1_ASAP7_75t_SL g291 ( 
.A(n_284),
.B(n_266),
.Y(n_291)
);

NAND4xp25_ASAP7_75t_SL g293 ( 
.A(n_292),
.B(n_288),
.C(n_291),
.D(n_290),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_293),
.A2(n_285),
.B(n_281),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_0),
.B(n_3),
.Y(n_295)
);

NAND3xp33_ASAP7_75t_SL g296 ( 
.A(n_295),
.B(n_3),
.C(n_4),
.Y(n_296)
);

BUFx24_ASAP7_75t_SL g297 ( 
.A(n_296),
.Y(n_297)
);


endmodule