module fake_netlist_1_5144_n_16 (n_1, n_2, n_0, n_16);
input n_1;
input n_2;
input n_0;
output n_16;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_10;
wire n_15;
wire n_7;
wire n_8;
INVx1_ASAP7_75t_L g3 ( .A(n_0), .Y(n_3) );
INVx1_ASAP7_75t_SL g4 ( .A(n_2), .Y(n_4) );
INVx2_ASAP7_75t_L g5 ( .A(n_2), .Y(n_5) );
INVx1_ASAP7_75t_L g6 ( .A(n_3), .Y(n_6) );
A2O1A1Ixp33_ASAP7_75t_L g7 ( .A1(n_3), .A2(n_0), .B(n_1), .C(n_2), .Y(n_7) );
OA21x2_ASAP7_75t_L g8 ( .A1(n_5), .A2(n_0), .B(n_1), .Y(n_8) );
NAND2xp5_ASAP7_75t_L g9 ( .A(n_6), .B(n_4), .Y(n_9) );
HB1xp67_ASAP7_75t_L g10 ( .A(n_6), .Y(n_10) );
NAND2xp5_ASAP7_75t_SL g11 ( .A(n_10), .B(n_6), .Y(n_11) );
OAI22xp5_ASAP7_75t_L g12 ( .A1(n_9), .A2(n_7), .B1(n_5), .B2(n_8), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_11), .Y(n_13) );
NAND4xp25_ASAP7_75t_L g14 ( .A(n_12), .B(n_7), .C(n_0), .D(n_2), .Y(n_14) );
OAI22xp5_ASAP7_75t_L g15 ( .A1(n_14), .A2(n_1), .B1(n_8), .B2(n_9), .Y(n_15) );
AOI22xp33_ASAP7_75t_L g16 ( .A1(n_15), .A2(n_8), .B1(n_13), .B2(n_11), .Y(n_16) );
endmodule