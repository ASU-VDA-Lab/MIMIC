module fake_jpeg_24926_n_326 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_10),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_20),
.B(n_8),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

NAND2x1_ASAP7_75t_SL g65 ( 
.A(n_47),
.B(n_23),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_22),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_35),
.B1(n_27),
.B2(n_28),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_50),
.A2(n_30),
.B1(n_34),
.B2(n_33),
.Y(n_87)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

BUFx2_ASAP7_75t_SL g88 ( 
.A(n_51),
.Y(n_88)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_61),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_53),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_35),
.B1(n_29),
.B2(n_28),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_55),
.A2(n_74),
.B1(n_75),
.B2(n_82),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_58),
.B(n_66),
.Y(n_94)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_60),
.B(n_21),
.Y(n_119)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NAND2xp33_ASAP7_75t_SL g108 ( 
.A(n_65),
.B(n_76),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_49),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_72),
.B(n_78),
.Y(n_106)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_41),
.A2(n_29),
.B1(n_32),
.B2(n_24),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_41),
.A2(n_29),
.B1(n_32),
.B2(n_24),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_40),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_27),
.Y(n_77)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_49),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_49),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_33),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_41),
.A2(n_32),
.B1(n_24),
.B2(n_22),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_41),
.A2(n_22),
.B1(n_30),
.B2(n_26),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_34),
.B1(n_36),
.B2(n_31),
.Y(n_93)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_85),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_41),
.A2(n_30),
.B1(n_20),
.B2(n_26),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_86),
.A2(n_25),
.B1(n_21),
.B2(n_20),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_87),
.A2(n_98),
.B1(n_101),
.B2(n_57),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_17),
.B1(n_19),
.B2(n_27),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_90),
.A2(n_95),
.B1(n_117),
.B2(n_68),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_93),
.A2(n_102),
.B1(n_104),
.B2(n_115),
.Y(n_143)
);

AO22x1_ASAP7_75t_SL g95 ( 
.A1(n_65),
.A2(n_78),
.B1(n_81),
.B2(n_66),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_97),
.B(n_9),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_60),
.A2(n_84),
.B1(n_80),
.B2(n_61),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_65),
.A2(n_18),
.B1(n_23),
.B2(n_33),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_54),
.A2(n_31),
.B1(n_26),
.B2(n_25),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_36),
.B1(n_31),
.B2(n_25),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_18),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_109),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_62),
.B(n_18),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_18),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_64),
.Y(n_127)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_114),
.Y(n_149)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_L g117 ( 
.A1(n_69),
.A2(n_19),
.B1(n_23),
.B2(n_18),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_119),
.B(n_23),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_63),
.A2(n_21),
.B1(n_19),
.B2(n_13),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_120),
.A2(n_63),
.B1(n_84),
.B2(n_57),
.Y(n_130)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_16),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_126),
.Y(n_164)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_125),
.B(n_133),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_97),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_150),
.Y(n_159)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_128),
.B(n_129),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_106),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_130),
.A2(n_152),
.B1(n_153),
.B2(n_156),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_95),
.B(n_23),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_131),
.B(n_144),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_SL g132 ( 
.A1(n_91),
.A2(n_18),
.B(n_23),
.C(n_19),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_SL g168 ( 
.A1(n_132),
.A2(n_110),
.B(n_116),
.C(n_105),
.Y(n_168)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_134),
.A2(n_16),
.B1(n_7),
.B2(n_9),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_95),
.A2(n_73),
.B1(n_79),
.B2(n_85),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_135),
.A2(n_141),
.B1(n_110),
.B2(n_100),
.Y(n_160)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_136),
.B(n_142),
.Y(n_188)
);

O2A1O1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_87),
.A2(n_70),
.B(n_67),
.C(n_51),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_137),
.A2(n_154),
.B(n_1),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_138),
.A2(n_140),
.B1(n_100),
.B2(n_111),
.Y(n_171)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_139),
.B(n_145),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_108),
.A2(n_68),
.B1(n_52),
.B2(n_18),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_107),
.A2(n_23),
.B1(n_56),
.B2(n_53),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_119),
.B(n_9),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_147),
.Y(n_173)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_0),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_117),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_151),
.B(n_155),
.Y(n_161)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_92),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_101),
.A2(n_0),
.B(n_1),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_90),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_167),
.Y(n_194)
);

AO21x2_ASAP7_75t_SL g158 ( 
.A1(n_135),
.A2(n_101),
.B(n_122),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_158),
.A2(n_184),
.B(n_137),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_160),
.A2(n_168),
.B1(n_176),
.B2(n_143),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_101),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_165),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_103),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_118),
.C(n_121),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_186),
.C(n_141),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_171),
.A2(n_189),
.B1(n_190),
.B2(n_183),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_111),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_174),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_123),
.B(n_126),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_125),
.A2(n_118),
.B1(n_113),
.B2(n_89),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_116),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_185),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_124),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_180),
.Y(n_196)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_128),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_136),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_148),
.A2(n_89),
.B1(n_12),
.B2(n_3),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_129),
.B(n_1),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_1),
.C(n_2),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_138),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_158),
.A2(n_168),
.B1(n_151),
.B2(n_156),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_192),
.A2(n_210),
.B1(n_217),
.B2(n_218),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_187),
.B(n_134),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_202),
.Y(n_227)
);

INVx11_ASAP7_75t_L g195 ( 
.A(n_157),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_197),
.Y(n_221)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

INVx13_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_206),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_154),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_199),
.A2(n_200),
.B(n_204),
.Y(n_241)
);

AND2x6_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_146),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_158),
.B(n_132),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_205),
.B(n_211),
.Y(n_243)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_164),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_208),
.A2(n_160),
.B1(n_176),
.B2(n_168),
.Y(n_222)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_209),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_132),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_172),
.Y(n_212)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_165),
.B(n_142),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_213),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_174),
.B(n_142),
.Y(n_214)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_180),
.Y(n_215)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_159),
.B(n_145),
.Y(n_216)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_169),
.A2(n_132),
.B(n_7),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_184),
.Y(n_225)
);

BUFx12_ASAP7_75t_L g220 ( 
.A(n_167),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_219),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_210),
.A2(n_171),
.B1(n_166),
.B2(n_189),
.Y(n_223)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_193),
.B(n_170),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_224),
.B(n_211),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_191),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_159),
.C(n_175),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_235),
.C(n_239),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_204),
.A2(n_168),
.B1(n_188),
.B2(n_186),
.Y(n_229)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_229),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_196),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_232),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_194),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_233),
.B(n_237),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_201),
.B(n_173),
.C(n_162),
.Y(n_235)
);

FAx1_ASAP7_75t_SL g237 ( 
.A(n_191),
.B(n_185),
.CI(n_132),
.CON(n_237),
.SN(n_237)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_161),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_255),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_247),
.A2(n_248),
.B1(n_263),
.B2(n_207),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_243),
.A2(n_212),
.B(n_217),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_211),
.C(n_216),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_228),
.C(n_234),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_203),
.Y(n_251)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_251),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_220),
.Y(n_252)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_221),
.B(n_220),
.Y(n_254)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_203),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_260),
.Y(n_271)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_242),
.Y(n_257)
);

INVxp33_ASAP7_75t_SL g270 ( 
.A(n_257),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_227),
.B(n_199),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_223),
.Y(n_278)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_241),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_262),
.B(n_264),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_243),
.A2(n_207),
.B(n_200),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_233),
.B(n_197),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_262),
.A2(n_241),
.B1(n_222),
.B2(n_231),
.Y(n_265)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_265),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_257),
.Y(n_266)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_266),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_248),
.Y(n_267)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_267),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_269),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_278),
.C(n_255),
.Y(n_286)
);

AOI211xp5_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_225),
.B(n_208),
.C(n_229),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_274),
.A2(n_260),
.B1(n_249),
.B2(n_258),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_227),
.C(n_239),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_277),
.C(n_250),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_235),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_261),
.B(n_218),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_279),
.B(n_261),
.Y(n_282)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_282),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_286),
.C(n_288),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_245),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_284),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_245),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_253),
.C(n_251),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_290),
.C(n_294),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_253),
.C(n_249),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_271),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_278),
.C(n_277),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_292),
.A2(n_285),
.B1(n_291),
.B2(n_275),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_296),
.A2(n_298),
.B1(n_226),
.B2(n_240),
.Y(n_306)
);

NOR2xp67_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_274),
.Y(n_297)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_297),
.Y(n_311)
);

OAI322xp33_ASAP7_75t_L g300 ( 
.A1(n_283),
.A2(n_246),
.A3(n_271),
.B1(n_281),
.B2(n_265),
.C1(n_294),
.C2(n_214),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_213),
.C(n_237),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_290),
.A2(n_281),
.B(n_280),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_301),
.A2(n_298),
.B(n_302),
.Y(n_307)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_287),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_246),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_304),
.A2(n_270),
.B1(n_195),
.B2(n_206),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_305),
.A2(n_307),
.B(n_309),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_306),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_312),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_296),
.A2(n_237),
.B1(n_205),
.B2(n_199),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_310),
.A2(n_205),
.B1(n_301),
.B2(n_303),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_198),
.C(n_220),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_313),
.A2(n_308),
.B1(n_309),
.B2(n_311),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_198),
.Y(n_316)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_316),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_320),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_315),
.A2(n_299),
.B1(n_312),
.B2(n_295),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_319),
.B(n_295),
.C(n_317),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_314),
.C(n_313),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);

OAI21xp33_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_322),
.B(n_7),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_6),
.Y(n_326)
);


endmodule