module real_jpeg_18802_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_0),
.Y(n_116)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_1),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_2),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_2),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_2),
.B(n_126),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_3),
.Y(n_124)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_5),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_5),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_5),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_5),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_6),
.B(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_6),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_6),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_6),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_6),
.B(n_109),
.Y(n_108)
);

AND2x4_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_17),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_7),
.B(n_41),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_7),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_7),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_7),
.B(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_8),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_9),
.B(n_124),
.Y(n_123)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_10),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_10),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_95),
.Y(n_11)
);

AOI21x1_ASAP7_75t_SL g12 ( 
.A1(n_13),
.A2(n_60),
.B(n_94),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_50),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_14),
.B(n_50),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_31),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_15),
.B(n_32),
.C(n_43),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_21),
.Y(n_15)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_16),
.Y(n_101)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_20),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_22),
.B(n_27),
.C(n_101),
.Y(n_100)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_42),
.B2(n_43),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_38),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_SL g52 ( 
.A(n_34),
.B(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AO22x1_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_43)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_47),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_47),
.B(n_48),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_53),
.C(n_55),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_51),
.A2(n_52),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_53),
.A2(n_55),
.B1(n_56),
.B2(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_75),
.B(n_93),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_71),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_71),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_68),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_64),
.B1(n_68),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_64),
.B(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_85),
.B(n_92),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_83),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_128),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_98),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_119),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_102),
.Y(n_99)
);

XOR2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_107),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_113),
.B1(n_117),
.B2(n_118),
.Y(n_107)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_113),
.Y(n_117)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_125),
.Y(n_121)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);


endmodule