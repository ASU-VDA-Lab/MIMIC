module fake_jpeg_18584_n_325 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_325);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

BUFx24_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_30),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_28),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_20),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_32),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_20),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_20),
.Y(n_33)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_26),
.A2(n_22),
.B1(n_16),
.B2(n_23),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_42),
.B1(n_28),
.B2(n_33),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_26),
.A2(n_22),
.B1(n_16),
.B2(n_13),
.Y(n_42)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_31),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_56),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_25),
.Y(n_48)
);

NOR2x1_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_57),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_14),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_52),
.Y(n_77)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_45),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_31),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_14),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_31),
.Y(n_57)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_59),
.A2(n_37),
.B1(n_36),
.B2(n_44),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_30),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_43),
.B1(n_33),
.B2(n_30),
.Y(n_63)
);

INVxp67_ASAP7_75t_R g62 ( 
.A(n_52),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_62),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_66),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_61),
.B1(n_56),
.B2(n_47),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_56),
.B1(n_48),
.B2(n_54),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_74),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_46),
.A2(n_37),
.B1(n_36),
.B2(n_25),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_26),
.B1(n_33),
.B2(n_28),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_27),
.B(n_28),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_76),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_50),
.A2(n_26),
.B1(n_33),
.B2(n_28),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_53),
.A2(n_41),
.B1(n_36),
.B2(n_42),
.Y(n_78)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_79),
.B(n_27),
.Y(n_87)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_89),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_80),
.B(n_30),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_82),
.B(n_83),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_30),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_92),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_32),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_27),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_68),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_98),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_32),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_27),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_76),
.Y(n_110)
);

BUFx24_ASAP7_75t_SL g101 ( 
.A(n_92),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_101),
.B(n_126),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_95),
.A2(n_62),
.B(n_67),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_103),
.A2(n_99),
.B(n_85),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

AO21x2_ASAP7_75t_L g106 ( 
.A1(n_100),
.A2(n_62),
.B(n_63),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g149 ( 
.A1(n_106),
.A2(n_51),
.B1(n_38),
.B2(n_34),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_94),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_107),
.B(n_116),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_84),
.A2(n_62),
.B1(n_79),
.B2(n_67),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_114),
.B1(n_99),
.B2(n_85),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_111),
.Y(n_130)
);

OAI32xp33_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_67),
.A3(n_77),
.B1(n_70),
.B2(n_74),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_75),
.B(n_70),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_112),
.A2(n_125),
.B(n_24),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_75),
.B1(n_78),
.B2(n_73),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_87),
.B(n_32),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_78),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_129),
.C(n_127),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_86),
.A2(n_39),
.B1(n_41),
.B2(n_32),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_120),
.A2(n_121),
.B1(n_127),
.B2(n_25),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_41),
.B1(n_59),
.B2(n_53),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_58),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_123),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_58),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_13),
.B(n_17),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_81),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_85),
.A2(n_59),
.B1(n_65),
.B2(n_71),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_72),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_128),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_99),
.B(n_13),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_138),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_133),
.A2(n_145),
.B(n_149),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_120),
.A2(n_93),
.B1(n_22),
.B2(n_16),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_135),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_123),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_137),
.B(n_143),
.Y(n_167)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_103),
.A2(n_15),
.B(n_21),
.C(n_19),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_90),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_147),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_148),
.B1(n_158),
.B2(n_165),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_125),
.Y(n_177)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_25),
.C(n_58),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_146),
.C(n_129),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_118),
.A2(n_15),
.B(n_19),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_25),
.C(n_58),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_23),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_114),
.A2(n_46),
.B1(n_51),
.B2(n_38),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_113),
.A2(n_19),
.B1(n_15),
.B2(n_21),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_72),
.Y(n_151)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_153),
.A2(n_49),
.B(n_8),
.Y(n_194)
);

INVxp33_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_155),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_156),
.A2(n_106),
.B(n_102),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_111),
.A2(n_21),
.B1(n_17),
.B2(n_34),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_110),
.Y(n_160)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_105),
.Y(n_161)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_161),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_107),
.B(n_72),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_162),
.B(n_164),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_106),
.B(n_12),
.Y(n_163)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_105),
.B(n_49),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_106),
.A2(n_17),
.B1(n_34),
.B2(n_24),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_171),
.B(n_177),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_161),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_173),
.B(n_179),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_141),
.A2(n_109),
.B1(n_106),
.B2(n_115),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_176),
.A2(n_159),
.B1(n_143),
.B2(n_138),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_178),
.A2(n_181),
.B(n_172),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_140),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_133),
.A2(n_106),
.B(n_121),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_151),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_187),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_134),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_139),
.Y(n_189)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_139),
.Y(n_190)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_152),
.Y(n_191)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

OA22x2_ASAP7_75t_L g192 ( 
.A1(n_136),
.A2(n_34),
.B1(n_24),
.B2(n_29),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_192),
.A2(n_194),
.B(n_149),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_149),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_149),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_196),
.A2(n_216),
.B(n_194),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_195),
.A2(n_130),
.B1(n_158),
.B2(n_163),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_197),
.A2(n_200),
.B1(n_213),
.B2(n_166),
.Y(n_233)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_167),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_199),
.B(n_206),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_188),
.A2(n_130),
.B1(n_131),
.B2(n_136),
.Y(n_200)
);

AND2x6_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_142),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_201),
.A2(n_215),
.B(n_49),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_144),
.C(n_146),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_211),
.C(n_212),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_147),
.Y(n_207)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_191),
.Y(n_209)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_169),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_210),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_156),
.C(n_160),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_148),
.C(n_132),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_188),
.A2(n_165),
.B1(n_153),
.B2(n_152),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_184),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_174),
.B1(n_170),
.B2(n_193),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_145),
.Y(n_219)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_220),
.A2(n_168),
.B1(n_190),
.B2(n_189),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_181),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_222),
.B(n_236),
.C(n_238),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_224),
.A2(n_227),
.B1(n_235),
.B2(n_243),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_217),
.A2(n_174),
.B1(n_183),
.B2(n_193),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_172),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_228),
.B(n_240),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_166),
.B1(n_176),
.B2(n_183),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_233),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_198),
.A2(n_200),
.B1(n_216),
.B2(n_197),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_234),
.A2(n_205),
.B1(n_220),
.B2(n_214),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_202),
.A2(n_175),
.B1(n_184),
.B2(n_180),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_175),
.C(n_180),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_237),
.A2(n_196),
.B(n_208),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_154),
.C(n_192),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_192),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_192),
.C(n_49),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_241),
.B(n_213),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_242),
.A2(n_34),
.B(n_24),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_202),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_244),
.B(n_253),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_246),
.A2(n_255),
.B1(n_259),
.B2(n_243),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_203),
.Y(n_247)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

BUFx24_ASAP7_75t_SL g251 ( 
.A(n_221),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_262),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_252),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_205),
.B(n_214),
.Y(n_253)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_233),
.A2(n_219),
.B1(n_1),
.B2(n_2),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_49),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_256),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_226),
.A2(n_18),
.B1(n_8),
.B2(n_10),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_257),
.A2(n_258),
.B1(n_7),
.B2(n_6),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_239),
.A2(n_18),
.B1(n_8),
.B2(n_10),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_234),
.A2(n_223),
.B1(n_228),
.B2(n_227),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_34),
.Y(n_273)
);

NOR3xp33_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_232),
.C(n_236),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_232),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_263),
.B(n_271),
.Y(n_278)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_264),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_244),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_268),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_L g268 ( 
.A1(n_249),
.A2(n_224),
.B1(n_235),
.B2(n_240),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_222),
.C(n_29),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_250),
.C(n_248),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_245),
.A2(n_18),
.B1(n_7),
.B2(n_9),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_246),
.Y(n_281)
);

A2O1A1O1Ixp25_ASAP7_75t_L g275 ( 
.A1(n_253),
.A2(n_7),
.B(n_6),
.C(n_12),
.D(n_3),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_275),
.A2(n_247),
.B(n_255),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_276),
.A2(n_267),
.B1(n_266),
.B2(n_265),
.Y(n_284)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_279),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_281),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_259),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_282),
.B(n_287),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_285),
.Y(n_297)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_284),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_277),
.A2(n_248),
.B1(n_6),
.B2(n_7),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_29),
.C(n_12),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_272),
.B(n_0),
.Y(n_288)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_288),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_274),
.B(n_0),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_289),
.B(n_0),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_269),
.A2(n_24),
.B(n_1),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_291),
.B(n_0),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_273),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_294),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_281),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_286),
.A2(n_275),
.B1(n_29),
.B2(n_12),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_299),
.Y(n_308)
);

FAx1_ASAP7_75t_SL g310 ( 
.A(n_296),
.B(n_3),
.CI(n_4),
.CON(n_310),
.SN(n_310)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_290),
.A2(n_29),
.B1(n_12),
.B2(n_2),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_1),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_278),
.B(n_283),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_304),
.A2(n_305),
.B(n_296),
.Y(n_316)
);

MAJx2_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_291),
.C(n_287),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_306),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_3),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_307),
.A2(n_302),
.B(n_308),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_311),
.C(n_312),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_300),
.C(n_301),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_29),
.C(n_4),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_315),
.B(n_316),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_308),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_318),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_314),
.Y(n_320)
);

NAND3xp33_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_309),
.C(n_317),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_310),
.B(n_4),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_322),
.B(n_5),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_3),
.C(n_5),
.Y(n_325)
);


endmodule