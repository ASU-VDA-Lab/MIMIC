module fake_jpeg_26304_n_225 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_225);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_213;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_3),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_39),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_42),
.B(n_50),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_22),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_44),
.B(n_49),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_19),
.B(n_0),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_51),
.B(n_2),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_34),
.B1(n_30),
.B2(n_35),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_52),
.A2(n_63),
.B1(n_8),
.B2(n_12),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_17),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_72),
.Y(n_90)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_35),
.B1(n_25),
.B2(n_27),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_74),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_47),
.A2(n_25),
.B1(n_23),
.B2(n_33),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_57),
.A2(n_73),
.B1(n_7),
.B2(n_8),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_33),
.B(n_23),
.C(n_22),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_32),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_68),
.Y(n_93)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_75),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_67),
.Y(n_92)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_17),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_32),
.B1(n_19),
.B2(n_20),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_48),
.B(n_18),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_27),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_32),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_2),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_38),
.A2(n_32),
.B1(n_29),
.B2(n_20),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_68),
.A2(n_50),
.B1(n_42),
.B2(n_18),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_78),
.A2(n_80),
.B1(n_65),
.B2(n_62),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_66),
.A2(n_20),
.B1(n_29),
.B2(n_4),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_79),
.A2(n_82),
.B1(n_74),
.B2(n_61),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_66),
.A2(n_41),
.B1(n_46),
.B2(n_45),
.Y(n_80)
);

AOI32xp33_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_46),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_81),
.A2(n_53),
.B(n_72),
.C(n_56),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_61),
.A2(n_62),
.B1(n_60),
.B2(n_69),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_71),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_98),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_64),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_96),
.B(n_97),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_11),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_99),
.B(n_104),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_105),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_59),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_101),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_6),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_103),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_6),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_10),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_56),
.Y(n_121)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_60),
.Y(n_122)
);

INVx3_ASAP7_75t_SL g108 ( 
.A(n_88),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_108),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_125),
.B(n_90),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_121),
.B1(n_126),
.B2(n_80),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_122),
.Y(n_146)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_128),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_56),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_53),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_89),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_12),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_72),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_100),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_55),
.Y(n_148)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_132),
.B(n_136),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_115),
.A2(n_98),
.B1(n_83),
.B2(n_87),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_133),
.A2(n_138),
.B1(n_124),
.B2(n_110),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_150),
.Y(n_170)
);

AOI211xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_83),
.B(n_102),
.C(n_87),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_135),
.A2(n_141),
.B(n_145),
.Y(n_164)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_112),
.B(n_96),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_137),
.B(n_152),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_115),
.A2(n_87),
.B1(n_90),
.B2(n_106),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_144),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_129),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_142),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_119),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_143),
.Y(n_169)
);

INVxp33_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_86),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_125),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_94),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_92),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_118),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_124),
.B(n_99),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_161),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_125),
.B(n_111),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_159),
.A2(n_111),
.B(n_121),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_163),
.Y(n_174)
);

NOR3xp33_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_117),
.C(n_81),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_152),
.B(n_110),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_166),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_134),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_123),
.Y(n_167)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_167),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_111),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_114),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_146),
.Y(n_172)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

OAI221xp5_ASAP7_75t_L g173 ( 
.A1(n_155),
.A2(n_149),
.B1(n_136),
.B2(n_137),
.C(n_135),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_78),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

INVxp33_ASAP7_75t_L g192 ( 
.A(n_176),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_133),
.B(n_145),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_177),
.A2(n_178),
.B(n_166),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_132),
.B1(n_121),
.B2(n_138),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_181),
.A2(n_164),
.B1(n_159),
.B2(n_171),
.Y(n_188)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_184),
.Y(n_194)
);

NOR2x1_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_146),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_185),
.B(n_186),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_114),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_168),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_188),
.A2(n_177),
.B1(n_181),
.B2(n_178),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_195),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_170),
.C(n_163),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_180),
.C(n_185),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_175),
.A2(n_168),
.B(n_154),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_191),
.B(n_198),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_193),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_170),
.Y(n_195)
);

NAND4xp25_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_169),
.C(n_165),
.D(n_120),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_186),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_201),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_180),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_206),
.C(n_188),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_197),
.A2(n_179),
.B1(n_182),
.B2(n_158),
.Y(n_205)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_205),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_192),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_210),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_203),
.A2(n_194),
.B(n_198),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_208),
.A2(n_212),
.B(n_140),
.Y(n_217)
);

NAND4xp25_ASAP7_75t_SL g210 ( 
.A(n_206),
.B(n_158),
.C(n_192),
.D(n_8),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_SL g213 ( 
.A1(n_211),
.A2(n_189),
.B(n_190),
.C(n_199),
.Y(n_213)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g220 ( 
.A1(n_213),
.A2(n_215),
.B(n_216),
.C(n_13),
.D(n_15),
.Y(n_220)
);

AOI21x1_ASAP7_75t_L g215 ( 
.A1(n_207),
.A2(n_199),
.B(n_204),
.Y(n_215)
);

AOI31xp67_ASAP7_75t_L g216 ( 
.A1(n_209),
.A2(n_13),
.A3(n_14),
.B(n_15),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_217),
.A2(n_153),
.B1(n_143),
.B2(n_119),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_218),
.Y(n_221)
);

NOR2x1_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_153),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_219),
.A2(n_220),
.B1(n_85),
.B2(n_95),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_219),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_223),
.A2(n_221),
.B(n_85),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_55),
.Y(n_225)
);


endmodule