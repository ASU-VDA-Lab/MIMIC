module fake_netlist_1_12354_n_733 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_733);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_733;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_638;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_711;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_SL g108 ( .A(n_18), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_8), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_90), .Y(n_110) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_59), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_63), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_62), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_15), .Y(n_114) );
CKINVDCx14_ASAP7_75t_R g115 ( .A(n_99), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_97), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_1), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_89), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_105), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_32), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_29), .Y(n_121) );
XOR2xp5_ASAP7_75t_L g122 ( .A(n_42), .B(n_58), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_40), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_88), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_24), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_9), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_102), .Y(n_127) );
BUFx3_ASAP7_75t_L g128 ( .A(n_19), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_37), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_48), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_5), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_41), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_98), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_31), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_47), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_96), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_56), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_27), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_10), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_69), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_103), .Y(n_141) );
BUFx3_ASAP7_75t_L g142 ( .A(n_104), .Y(n_142) );
BUFx3_ASAP7_75t_L g143 ( .A(n_87), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_6), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_91), .Y(n_145) );
OR2x2_ASAP7_75t_L g146 ( .A(n_15), .B(n_14), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_65), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_22), .Y(n_148) );
OR2x2_ASAP7_75t_L g149 ( .A(n_35), .B(n_20), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_60), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_1), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_81), .Y(n_152) );
BUFx3_ASAP7_75t_L g153 ( .A(n_55), .Y(n_153) );
INVx2_ASAP7_75t_SL g154 ( .A(n_142), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_128), .Y(n_155) );
NAND2xp33_ASAP7_75t_L g156 ( .A(n_110), .B(n_107), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_111), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_115), .B(n_128), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_138), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_111), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_111), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_111), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_117), .B(n_0), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_112), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_113), .Y(n_165) );
INVx2_ASAP7_75t_SL g166 ( .A(n_142), .Y(n_166) );
OAI22xp5_ASAP7_75t_L g167 ( .A1(n_140), .A2(n_0), .B1(n_2), .B2(n_3), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_114), .B(n_2), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_129), .Y(n_169) );
INVxp67_ASAP7_75t_L g170 ( .A(n_126), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_129), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_129), .Y(n_172) );
AND2x4_ASAP7_75t_L g173 ( .A(n_143), .B(n_3), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_159), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_158), .B(n_116), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_159), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_160), .Y(n_177) );
INVx1_ASAP7_75t_SL g178 ( .A(n_158), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_173), .Y(n_179) );
NOR2xp33_ASAP7_75t_SL g180 ( .A(n_173), .B(n_140), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_170), .B(n_114), .Y(n_181) );
INVx3_ASAP7_75t_L g182 ( .A(n_173), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_173), .Y(n_183) );
AO22x2_ASAP7_75t_L g184 ( .A1(n_167), .A2(n_122), .B1(n_146), .B2(n_108), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_164), .B(n_138), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_159), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_160), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_160), .Y(n_188) );
AOI22xp33_ASAP7_75t_SL g189 ( .A1(n_167), .A2(n_109), .B1(n_139), .B2(n_144), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_159), .Y(n_190) );
NAND3xp33_ASAP7_75t_L g191 ( .A(n_164), .B(n_134), .C(n_123), .Y(n_191) );
AND2x6_ASAP7_75t_L g192 ( .A(n_168), .B(n_143), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_160), .Y(n_193) );
INVx2_ASAP7_75t_SL g194 ( .A(n_154), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_160), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_157), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_155), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_165), .B(n_120), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_157), .Y(n_199) );
BUFx3_ASAP7_75t_L g200 ( .A(n_154), .Y(n_200) );
OR2x2_ASAP7_75t_L g201 ( .A(n_181), .B(n_168), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_192), .A2(n_165), .B1(n_154), .B2(n_166), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_178), .B(n_166), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_178), .B(n_166), .Y(n_204) );
INVx8_ASAP7_75t_L g205 ( .A(n_192), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_181), .B(n_163), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_197), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_197), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_175), .B(n_163), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_197), .Y(n_210) );
AND2x2_ASAP7_75t_L g211 ( .A(n_185), .B(n_155), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_197), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_179), .B(n_156), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g214 ( .A1(n_189), .A2(n_139), .B1(n_109), .B2(n_151), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_196), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_179), .A2(n_141), .B(n_121), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_179), .B(n_110), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_179), .B(n_127), .Y(n_218) );
BUFx3_ASAP7_75t_L g219 ( .A(n_192), .Y(n_219) );
AOI22xp5_ASAP7_75t_L g220 ( .A1(n_180), .A2(n_192), .B1(n_182), .B2(n_183), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_192), .A2(n_144), .B1(n_124), .B2(n_145), .Y(n_221) );
INVx3_ASAP7_75t_L g222 ( .A(n_182), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_192), .B(n_127), .Y(n_223) );
AOI221xp5_ASAP7_75t_L g224 ( .A1(n_184), .A2(n_131), .B1(n_147), .B2(n_150), .C(n_152), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_192), .A2(n_132), .B1(n_135), .B2(n_153), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_192), .B(n_147), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_180), .A2(n_150), .B1(n_152), .B2(n_125), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_196), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_199), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g230 ( .A1(n_192), .A2(n_148), .B1(n_119), .B2(n_130), .Y(n_230) );
AOI221xp5_ASAP7_75t_L g231 ( .A1(n_184), .A2(n_118), .B1(n_133), .B2(n_136), .C(n_137), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_185), .B(n_153), .Y(n_232) );
INVxp67_ASAP7_75t_L g233 ( .A(n_184), .Y(n_233) );
INVx2_ASAP7_75t_SL g234 ( .A(n_182), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_182), .B(n_141), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_222), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_213), .A2(n_183), .B(n_194), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_209), .A2(n_183), .B(n_198), .C(n_191), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_220), .B(n_183), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_206), .B(n_200), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_220), .B(n_200), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_235), .A2(n_194), .B(n_200), .Y(n_242) );
OA22x2_ASAP7_75t_L g243 ( .A1(n_233), .A2(n_184), .B1(n_189), .B2(n_174), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_206), .B(n_211), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_211), .B(n_174), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_201), .B(n_194), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_201), .B(n_176), .Y(n_247) );
NOR2xp67_ASAP7_75t_L g248 ( .A(n_214), .B(n_191), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_219), .B(n_176), .Y(n_249) );
BUFx4f_ASAP7_75t_L g250 ( .A(n_205), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_214), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_235), .A2(n_186), .B(n_190), .Y(n_252) );
O2A1O1Ixp5_ASAP7_75t_L g253 ( .A1(n_216), .A2(n_186), .B(n_190), .C(n_149), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_232), .B(n_184), .Y(n_254) );
OAI21xp5_ASAP7_75t_L g255 ( .A1(n_207), .A2(n_199), .B(n_195), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_207), .A2(n_195), .B(n_193), .Y(n_256) );
INVx4_ASAP7_75t_L g257 ( .A(n_205), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_208), .A2(n_195), .B(n_193), .Y(n_258) );
AOI21x1_ASAP7_75t_L g259 ( .A1(n_208), .A2(n_193), .B(n_188), .Y(n_259) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_210), .A2(n_188), .B(n_187), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_L g261 ( .A1(n_203), .A2(n_172), .B(n_171), .C(n_162), .Y(n_261) );
INVx4_ASAP7_75t_L g262 ( .A(n_205), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_232), .B(n_4), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_222), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_210), .A2(n_188), .B(n_187), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_234), .A2(n_187), .B(n_177), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_224), .B(n_4), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_244), .B(n_222), .Y(n_268) );
BUFx3_ASAP7_75t_L g269 ( .A(n_250), .Y(n_269) );
AOI21xp5_ASAP7_75t_SL g270 ( .A1(n_241), .A2(n_219), .B(n_205), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_245), .B(n_215), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_240), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_250), .Y(n_273) );
OAI22x1_ASAP7_75t_L g274 ( .A1(n_251), .A2(n_227), .B1(n_230), .B2(n_231), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_254), .B(n_227), .Y(n_275) );
OAI21x1_ASAP7_75t_L g276 ( .A1(n_259), .A2(n_202), .B(n_225), .Y(n_276) );
O2A1O1Ixp33_ASAP7_75t_L g277 ( .A1(n_238), .A2(n_204), .B(n_226), .C(n_223), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_243), .A2(n_267), .B1(n_248), .B2(n_246), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_246), .B(n_230), .Y(n_279) );
OA21x2_ASAP7_75t_L g280 ( .A1(n_253), .A2(n_221), .B(n_212), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_L g281 ( .A1(n_238), .A2(n_217), .B(n_218), .C(n_234), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_236), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_257), .B(n_205), .Y(n_283) );
AO31x2_ASAP7_75t_L g284 ( .A1(n_237), .A2(n_171), .A3(n_157), .B(n_162), .Y(n_284) );
BUFx3_ASAP7_75t_L g285 ( .A(n_257), .Y(n_285) );
AO31x2_ASAP7_75t_L g286 ( .A1(n_263), .A2(n_171), .A3(n_162), .B(n_172), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_247), .B(n_212), .Y(n_287) );
OAI21x1_ASAP7_75t_L g288 ( .A1(n_242), .A2(n_229), .B(n_228), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_243), .B(n_215), .Y(n_289) );
BUFx2_ASAP7_75t_L g290 ( .A(n_262), .Y(n_290) );
INVx3_ASAP7_75t_SL g291 ( .A(n_262), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_239), .A2(n_229), .B(n_228), .Y(n_292) );
BUFx2_ASAP7_75t_L g293 ( .A(n_271), .Y(n_293) );
OAI21x1_ASAP7_75t_L g294 ( .A1(n_288), .A2(n_241), .B(n_239), .Y(n_294) );
OA21x2_ASAP7_75t_L g295 ( .A1(n_288), .A2(n_255), .B(n_260), .Y(n_295) );
OAI21x1_ASAP7_75t_L g296 ( .A1(n_292), .A2(n_266), .B(n_265), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_271), .B(n_264), .Y(n_297) );
OA21x2_ASAP7_75t_L g298 ( .A1(n_281), .A2(n_252), .B(n_258), .Y(n_298) );
AOI21x1_ASAP7_75t_L g299 ( .A1(n_292), .A2(n_256), .B(n_172), .Y(n_299) );
NOR2x1_ASAP7_75t_SL g300 ( .A(n_285), .B(n_249), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_272), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_278), .B(n_249), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_272), .Y(n_303) );
OAI21xp5_ASAP7_75t_L g304 ( .A1(n_277), .A2(n_261), .B(n_177), .Y(n_304) );
OAI21x1_ASAP7_75t_L g305 ( .A1(n_277), .A2(n_177), .B(n_169), .Y(n_305) );
OA21x2_ASAP7_75t_L g306 ( .A1(n_276), .A2(n_169), .B(n_161), .Y(n_306) );
OR2x6_ASAP7_75t_L g307 ( .A(n_270), .B(n_129), .Y(n_307) );
NAND2x1p5_ASAP7_75t_L g308 ( .A(n_285), .B(n_160), .Y(n_308) );
OAI21x1_ASAP7_75t_SL g309 ( .A1(n_287), .A2(n_5), .B(n_6), .Y(n_309) );
BUFx2_ASAP7_75t_R g310 ( .A(n_291), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_282), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_268), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_290), .B(n_291), .Y(n_313) );
OAI21xp5_ASAP7_75t_L g314 ( .A1(n_276), .A2(n_169), .B(n_161), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_306), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_301), .B(n_275), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_301), .Y(n_317) );
AO21x2_ASAP7_75t_L g318 ( .A1(n_314), .A2(n_289), .B(n_279), .Y(n_318) );
OAI21x1_ASAP7_75t_L g319 ( .A1(n_305), .A2(n_270), .B(n_289), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_303), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_311), .Y(n_321) );
AOI21x1_ASAP7_75t_L g322 ( .A1(n_299), .A2(n_280), .B(n_287), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_303), .Y(n_323) );
OR2x6_ASAP7_75t_L g324 ( .A(n_307), .B(n_290), .Y(n_324) );
OAI21x1_ASAP7_75t_L g325 ( .A1(n_305), .A2(n_299), .B(n_314), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_311), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_311), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_312), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_312), .Y(n_329) );
INVx3_ASAP7_75t_L g330 ( .A(n_307), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_310), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_293), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_293), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_306), .Y(n_334) );
AOI21xp33_ASAP7_75t_SL g335 ( .A1(n_313), .A2(n_274), .B(n_291), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_309), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_309), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_305), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_297), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_310), .Y(n_340) );
INVx2_ASAP7_75t_SL g341 ( .A(n_308), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_315), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_339), .B(n_302), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_326), .B(n_294), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_326), .B(n_294), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_327), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_332), .B(n_302), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_317), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_324), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_327), .B(n_294), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_339), .B(n_297), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_317), .B(n_307), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_320), .B(n_307), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_320), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_315), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_315), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_332), .B(n_286), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_333), .B(n_286), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_323), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_323), .B(n_321), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_321), .B(n_307), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_333), .B(n_286), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_328), .B(n_286), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_328), .B(n_286), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_329), .B(n_284), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_329), .B(n_286), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_334), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_318), .B(n_284), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_318), .B(n_284), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_316), .A2(n_274), .B1(n_285), .B2(n_298), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_318), .B(n_284), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_334), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_341), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_340), .A2(n_298), .B1(n_280), .B2(n_268), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_334), .B(n_284), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_336), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_336), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_337), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_337), .B(n_284), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_338), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_338), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_330), .B(n_306), .Y(n_382) );
NOR2x1_ASAP7_75t_SL g383 ( .A(n_324), .B(n_269), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_322), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_324), .A2(n_295), .B1(n_308), .B2(n_298), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_346), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_351), .B(n_335), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_351), .B(n_335), .Y(n_388) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_373), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_342), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_348), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_348), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_354), .B(n_341), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_354), .Y(n_394) );
INVx1_ASAP7_75t_SL g395 ( .A(n_360), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_359), .B(n_331), .Y(n_396) );
INVx5_ASAP7_75t_L g397 ( .A(n_349), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_379), .B(n_330), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_342), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_347), .B(n_330), .Y(n_400) );
NOR2x1_ASAP7_75t_L g401 ( .A(n_364), .B(n_324), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_379), .B(n_330), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_342), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_343), .B(n_7), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_368), .B(n_319), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_368), .B(n_319), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_359), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_360), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_376), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_376), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_369), .B(n_325), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_377), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_377), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_343), .B(n_324), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_356), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_378), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_356), .Y(n_417) );
NAND2x1p5_ASAP7_75t_L g418 ( .A(n_349), .B(n_306), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_378), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_355), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_369), .B(n_325), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_355), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_371), .B(n_322), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_356), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_371), .B(n_295), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_372), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_372), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_367), .Y(n_428) );
INVxp67_ASAP7_75t_SL g429 ( .A(n_367), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_372), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_347), .B(n_7), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_365), .Y(n_432) );
OR2x6_ASAP7_75t_L g433 ( .A(n_385), .B(n_352), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_363), .B(n_295), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_363), .B(n_300), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_357), .B(n_298), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_384), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_384), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_366), .B(n_295), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_364), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_365), .Y(n_441) );
AND2x4_ASAP7_75t_L g442 ( .A(n_352), .B(n_300), .Y(n_442) );
AND2x4_ASAP7_75t_L g443 ( .A(n_382), .B(n_296), .Y(n_443) );
AND2x4_ASAP7_75t_L g444 ( .A(n_382), .B(n_296), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_366), .B(n_295), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_357), .B(n_8), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_353), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_380), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_380), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_344), .B(n_345), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_358), .B(n_9), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_344), .B(n_304), .Y(n_452) );
BUFx3_ASAP7_75t_L g453 ( .A(n_389), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_386), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_450), .B(n_345), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_395), .B(n_358), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_450), .B(n_350), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_391), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_396), .B(n_362), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_391), .Y(n_460) );
INVx3_ASAP7_75t_L g461 ( .A(n_418), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_390), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_392), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_392), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_411), .B(n_350), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_394), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_440), .B(n_362), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_394), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_407), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_407), .Y(n_470) );
AND2x2_ASAP7_75t_SL g471 ( .A(n_420), .B(n_353), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_390), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_408), .B(n_370), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_408), .B(n_375), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_432), .B(n_375), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_432), .B(n_374), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_441), .B(n_361), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_411), .B(n_385), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_409), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_399), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_399), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_422), .B(n_381), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_421), .B(n_381), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_409), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_410), .Y(n_485) );
NOR2x1_ASAP7_75t_L g486 ( .A(n_401), .B(n_361), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_403), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_410), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_421), .B(n_384), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_447), .B(n_10), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_412), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_423), .B(n_405), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_423), .B(n_383), .Y(n_493) );
A2O1A1O1Ixp25_ASAP7_75t_L g494 ( .A1(n_431), .A2(n_11), .B(n_12), .C(n_13), .D(n_14), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_441), .B(n_383), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_405), .B(n_161), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_436), .B(n_161), .Y(n_497) );
BUFx3_ASAP7_75t_L g498 ( .A(n_397), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_412), .Y(n_499) );
NOR2xp67_ASAP7_75t_L g500 ( .A(n_397), .B(n_11), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_387), .B(n_12), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_406), .B(n_161), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_406), .B(n_161), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_425), .B(n_169), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_388), .B(n_13), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_425), .B(n_169), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_446), .B(n_16), .Y(n_507) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_429), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_398), .B(n_169), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_403), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_400), .B(n_16), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_398), .B(n_304), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_402), .B(n_296), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_413), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_415), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_413), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_416), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_451), .B(n_17), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_402), .B(n_308), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_434), .B(n_17), .Y(n_520) );
NOR3xp33_ASAP7_75t_L g521 ( .A(n_404), .B(n_283), .C(n_282), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_416), .Y(n_522) );
INVxp67_ASAP7_75t_L g523 ( .A(n_401), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_419), .Y(n_524) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_428), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_434), .B(n_439), .Y(n_526) );
INVx3_ASAP7_75t_L g527 ( .A(n_418), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_439), .B(n_18), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_445), .B(n_19), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_445), .B(n_280), .Y(n_530) );
NAND2x1p5_ASAP7_75t_L g531 ( .A(n_397), .B(n_442), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_419), .B(n_280), .Y(n_532) );
AND2x4_ASAP7_75t_L g533 ( .A(n_433), .B(n_21), .Y(n_533) );
INVx1_ASAP7_75t_SL g534 ( .A(n_400), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_428), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_452), .B(n_282), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_525), .Y(n_537) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_533), .A2(n_397), .B(n_442), .C(n_435), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_454), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_526), .B(n_433), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_508), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_533), .B(n_397), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_526), .B(n_433), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_483), .B(n_448), .Y(n_544) );
INVx2_ASAP7_75t_SL g545 ( .A(n_453), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_458), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_460), .Y(n_547) );
NOR2x1p5_ASAP7_75t_L g548 ( .A(n_533), .B(n_414), .Y(n_548) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_453), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_492), .B(n_455), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_483), .B(n_448), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_504), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_492), .B(n_433), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_478), .A2(n_442), .B1(n_443), .B2(n_444), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_497), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_504), .B(n_449), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_456), .B(n_436), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_463), .Y(n_558) );
INVx5_ASAP7_75t_L g559 ( .A(n_461), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_497), .Y(n_560) );
INVx1_ASAP7_75t_SL g561 ( .A(n_493), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_455), .B(n_430), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_457), .B(n_443), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_506), .B(n_449), .Y(n_564) );
AND2x4_ASAP7_75t_SL g565 ( .A(n_493), .B(n_443), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_464), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_466), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_457), .B(n_443), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_468), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_506), .B(n_465), .Y(n_570) );
AOI21xp33_ASAP7_75t_L g571 ( .A1(n_501), .A2(n_393), .B(n_438), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_465), .B(n_444), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_467), .B(n_430), .Y(n_573) );
NAND2x2_ASAP7_75t_L g574 ( .A(n_498), .B(n_397), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_471), .B(n_444), .Y(n_575) );
INVxp33_ASAP7_75t_L g576 ( .A(n_520), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_471), .B(n_444), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_489), .B(n_452), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_469), .Y(n_579) );
INVxp67_ASAP7_75t_L g580 ( .A(n_496), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_470), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_479), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_534), .B(n_424), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_478), .B(n_424), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_484), .Y(n_585) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_489), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_500), .B(n_415), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_505), .B(n_427), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_485), .Y(n_589) );
INVx1_ASAP7_75t_SL g590 ( .A(n_520), .Y(n_590) );
NOR2x1p5_ASAP7_75t_L g591 ( .A(n_498), .B(n_427), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_488), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_459), .B(n_426), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_535), .B(n_426), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_477), .B(n_417), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_491), .Y(n_596) );
NOR2x1_ASAP7_75t_L g597 ( .A(n_490), .B(n_438), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_499), .B(n_417), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_514), .B(n_437), .Y(n_599) );
NOR4xp25_ASAP7_75t_L g600 ( .A(n_507), .B(n_437), .C(n_418), .D(n_26), .Y(n_600) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_496), .Y(n_601) );
OAI22xp33_ASAP7_75t_SL g602 ( .A1(n_523), .A2(n_273), .B1(n_269), .B2(n_28), .Y(n_602) );
AOI21x1_ASAP7_75t_L g603 ( .A1(n_528), .A2(n_23), .B(n_25), .Y(n_603) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_502), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_516), .Y(n_605) );
A2O1A1Ixp33_ASAP7_75t_L g606 ( .A1(n_459), .A2(n_269), .B(n_273), .C(n_34), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_513), .B(n_30), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_517), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_474), .B(n_33), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_522), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_528), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_524), .B(n_36), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_482), .Y(n_613) );
NAND2x1_ASAP7_75t_SL g614 ( .A(n_461), .B(n_38), .Y(n_614) );
OAI31xp33_ASAP7_75t_L g615 ( .A1(n_602), .A2(n_531), .A3(n_521), .B(n_511), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_541), .B(n_502), .Y(n_616) );
AOI32xp33_ASAP7_75t_L g617 ( .A1(n_576), .A2(n_486), .A3(n_503), .B1(n_461), .B2(n_527), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_591), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_578), .B(n_503), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_537), .Y(n_620) );
AND2x4_ASAP7_75t_L g621 ( .A(n_565), .B(n_509), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_604), .B(n_509), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_562), .B(n_482), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_544), .Y(n_624) );
AOI21xp33_ASAP7_75t_SL g625 ( .A1(n_549), .A2(n_531), .B(n_495), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_544), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_578), .B(n_476), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_551), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_571), .A2(n_518), .B1(n_529), .B2(n_473), .C(n_513), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_545), .B(n_475), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_604), .Y(n_631) );
AND2x4_ASAP7_75t_L g632 ( .A(n_549), .B(n_580), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_580), .A2(n_512), .B1(n_519), .B2(n_527), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_590), .A2(n_527), .B1(n_519), .B2(n_536), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_593), .B(n_512), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_540), .B(n_487), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_551), .Y(n_637) );
OAI21xp33_ASAP7_75t_L g638 ( .A1(n_554), .A2(n_530), .B(n_487), .Y(n_638) );
OR2x2_ASAP7_75t_L g639 ( .A(n_557), .B(n_515), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_543), .B(n_515), .Y(n_640) );
AOI22xp33_ASAP7_75t_SL g641 ( .A1(n_575), .A2(n_480), .B1(n_510), .B2(n_481), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_552), .Y(n_642) );
OR2x2_ASAP7_75t_L g643 ( .A(n_586), .B(n_510), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_570), .Y(n_644) );
OAI221xp5_ASAP7_75t_L g645 ( .A1(n_571), .A2(n_494), .B1(n_481), .B2(n_480), .C(n_472), .Y(n_645) );
AOI222xp33_ASAP7_75t_L g646 ( .A1(n_611), .A2(n_472), .B1(n_462), .B2(n_532), .C1(n_273), .C2(n_46), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_570), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_553), .B(n_462), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_613), .B(n_106), .Y(n_649) );
OAI31xp33_ASAP7_75t_L g650 ( .A1(n_548), .A2(n_39), .A3(n_43), .B(n_44), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_546), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_572), .B(n_45), .Y(n_652) );
NAND2x1_ASAP7_75t_L g653 ( .A(n_577), .B(n_49), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_539), .B(n_50), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_550), .B(n_51), .Y(n_655) );
NAND2xp33_ASAP7_75t_SL g656 ( .A(n_542), .B(n_52), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_601), .B(n_53), .Y(n_657) );
NAND3xp33_ASAP7_75t_SL g658 ( .A(n_600), .B(n_606), .C(n_538), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_547), .Y(n_659) );
O2A1O1Ixp33_ASAP7_75t_SL g660 ( .A1(n_561), .A2(n_54), .B(n_57), .C(n_61), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_558), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_555), .Y(n_662) );
BUFx2_ASAP7_75t_L g663 ( .A(n_597), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_560), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_566), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_619), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_658), .A2(n_588), .B1(n_574), .B2(n_607), .Y(n_667) );
AOI21xp5_ASAP7_75t_L g668 ( .A1(n_615), .A2(n_587), .B(n_556), .Y(n_668) );
NAND2x2_ASAP7_75t_L g669 ( .A(n_653), .B(n_603), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_619), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_624), .Y(n_671) );
OAI221xp5_ASAP7_75t_SL g672 ( .A1(n_615), .A2(n_556), .B1(n_564), .B2(n_573), .C(n_609), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_646), .A2(n_564), .B1(n_584), .B2(n_559), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_629), .A2(n_634), .B1(n_638), .B2(n_627), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_643), .Y(n_675) );
AOI221xp5_ASAP7_75t_L g676 ( .A1(n_634), .A2(n_589), .B1(n_567), .B2(n_610), .C(n_608), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_627), .A2(n_585), .B1(n_569), .B2(n_605), .C(n_579), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_633), .A2(n_568), .B1(n_563), .B2(n_581), .Y(n_678) );
BUFx2_ASAP7_75t_L g679 ( .A(n_632), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_645), .A2(n_596), .B1(n_592), .B2(n_582), .C(n_583), .Y(n_680) );
OAI321xp33_ASAP7_75t_L g681 ( .A1(n_617), .A2(n_612), .A3(n_599), .B1(n_598), .B2(n_594), .C(n_595), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_625), .A2(n_559), .B1(n_598), .B2(n_594), .Y(n_682) );
NAND3xp33_ASAP7_75t_L g683 ( .A(n_646), .B(n_612), .C(n_599), .Y(n_683) );
OAI221xp5_ASAP7_75t_L g684 ( .A1(n_641), .A2(n_614), .B1(n_559), .B2(n_67), .C(n_68), .Y(n_684) );
OAI221xp5_ASAP7_75t_L g685 ( .A1(n_663), .A2(n_559), .B1(n_66), .B2(n_70), .C(n_71), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_626), .B(n_64), .Y(n_686) );
OAI21xp5_ASAP7_75t_L g687 ( .A1(n_656), .A2(n_72), .B(n_73), .Y(n_687) );
A2O1A1Ixp33_ASAP7_75t_L g688 ( .A1(n_650), .A2(n_632), .B(n_621), .C(n_630), .Y(n_688) );
O2A1O1Ixp33_ASAP7_75t_L g689 ( .A1(n_620), .A2(n_74), .B(n_75), .C(n_76), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g690 ( .A1(n_660), .A2(n_77), .B(n_78), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_628), .Y(n_691) );
AOI321xp33_ASAP7_75t_L g692 ( .A1(n_644), .A2(n_79), .A3(n_80), .B1(n_82), .B2(n_83), .C(n_84), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_631), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_680), .B(n_647), .Y(n_694) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_688), .B(n_621), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_666), .B(n_637), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_679), .B(n_618), .Y(n_697) );
OAI211xp5_ASAP7_75t_L g698 ( .A1(n_667), .A2(n_650), .B(n_655), .C(n_657), .Y(n_698) );
O2A1O1Ixp5_ASAP7_75t_L g699 ( .A1(n_672), .A2(n_665), .B(n_651), .C(n_659), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_673), .A2(n_623), .B1(n_622), .B2(n_635), .Y(n_700) );
NOR3xp33_ASAP7_75t_L g701 ( .A(n_681), .B(n_649), .C(n_654), .Y(n_701) );
NOR3xp33_ASAP7_75t_L g702 ( .A(n_681), .B(n_652), .C(n_616), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_674), .B(n_661), .Y(n_703) );
NOR4xp25_ASAP7_75t_L g704 ( .A(n_683), .B(n_642), .C(n_662), .D(n_664), .Y(n_704) );
O2A1O1Ixp33_ASAP7_75t_L g705 ( .A1(n_668), .A2(n_639), .B(n_640), .C(n_648), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_670), .Y(n_706) );
OAI21xp5_ASAP7_75t_SL g707 ( .A1(n_684), .A2(n_636), .B(n_86), .Y(n_707) );
AOI21xp33_ASAP7_75t_SL g708 ( .A1(n_682), .A2(n_85), .B(n_92), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_695), .A2(n_676), .B1(n_669), .B2(n_677), .Y(n_709) );
XNOR2x1_ASAP7_75t_L g710 ( .A(n_700), .B(n_687), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_697), .A2(n_678), .B1(n_691), .B2(n_671), .Y(n_711) );
A2O1A1Ixp33_ASAP7_75t_L g712 ( .A1(n_699), .A2(n_687), .B(n_690), .C(n_689), .Y(n_712) );
NOR3xp33_ASAP7_75t_L g713 ( .A(n_707), .B(n_685), .C(n_686), .Y(n_713) );
NAND3xp33_ASAP7_75t_SL g714 ( .A(n_704), .B(n_692), .C(n_693), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_703), .B(n_675), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_715), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_709), .B(n_703), .Y(n_717) );
NAND3xp33_ASAP7_75t_L g718 ( .A(n_710), .B(n_705), .C(n_701), .Y(n_718) );
AND2x4_ASAP7_75t_L g719 ( .A(n_713), .B(n_706), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_716), .Y(n_720) );
NOR3xp33_ASAP7_75t_L g721 ( .A(n_718), .B(n_714), .C(n_712), .Y(n_721) );
NOR4xp75_ASAP7_75t_SL g722 ( .A(n_717), .B(n_694), .C(n_696), .D(n_711), .Y(n_722) );
INVx2_ASAP7_75t_L g723 ( .A(n_720), .Y(n_723) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_721), .Y(n_724) );
NOR3x1_ASAP7_75t_L g725 ( .A(n_724), .B(n_722), .C(n_698), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_723), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_726), .Y(n_727) );
AOI21xp33_ASAP7_75t_L g728 ( .A1(n_725), .A2(n_719), .B(n_708), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_727), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_729), .A2(n_728), .B(n_702), .Y(n_730) );
NAND2xp33_ASAP7_75t_L g731 ( .A(n_730), .B(n_93), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_731), .B(n_94), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_732), .A2(n_95), .B1(n_100), .B2(n_101), .Y(n_733) );
endmodule