module fake_jpeg_9237_n_122 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_122);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_122;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_31),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_30),
.B(n_37),
.Y(n_46)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_0),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_35),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_34),
.B(n_16),
.Y(n_51)
);

OR2x4_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_15),
.B(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_47),
.Y(n_58)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_50),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_56),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_35),
.C(n_21),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_57),
.C(n_14),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_55),
.B(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_50),
.B(n_33),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_27),
.B(n_26),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_68),
.B(n_69),
.Y(n_73)
);

XNOR2x1_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_21),
.Y(n_60)
);

XOR2x1_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_17),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_31),
.B1(n_29),
.B2(n_25),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_25),
.B1(n_22),
.B2(n_16),
.Y(n_76)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_66),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_27),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_21),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_74),
.C(n_79),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_17),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_78),
.B1(n_84),
.B2(n_61),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_83),
.B(n_57),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_54),
.A2(n_22),
.B1(n_28),
.B2(n_14),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_20),
.B(n_23),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_54),
.A2(n_23),
.B1(n_19),
.B2(n_32),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_85),
.B(n_86),
.Y(n_99)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_89),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_80),
.B(n_65),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_91),
.Y(n_100)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_57),
.C(n_69),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_73),
.C(n_83),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_93),
.B(n_95),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_55),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_58),
.B(n_19),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_90),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_90),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_103),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_73),
.C(n_84),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_100),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_104),
.B(n_108),
.Y(n_113)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_107),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_94),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_103),
.B(n_102),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_109),
.A2(n_92),
.B(n_101),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_109),
.C(n_108),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_81),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_110),
.Y(n_116)
);

AOI322xp5_ASAP7_75t_L g115 ( 
.A1(n_112),
.A2(n_82),
.A3(n_24),
.B1(n_6),
.B2(n_8),
.C1(n_9),
.C2(n_4),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_115),
.A2(n_111),
.B(n_6),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_117),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_5),
.Y(n_118)
);

OA21x2_ASAP7_75t_L g120 ( 
.A1(n_118),
.A2(n_5),
.B(n_10),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_67),
.B1(n_13),
.B2(n_12),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_121),
.B(n_119),
.Y(n_122)
);


endmodule