module fake_jpeg_12235_n_472 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_472);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_472;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx4f_ASAP7_75t_SL g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_26),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_51),
.B(n_82),
.Y(n_102)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_15),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_53),
.B(n_55),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_15),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

BUFx24_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g105 ( 
.A(n_58),
.Y(n_105)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_60),
.Y(n_97)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_61),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_32),
.B(n_8),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_62),
.B(n_70),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_32),
.B(n_8),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_63),
.B(n_64),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_14),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_67),
.Y(n_124)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_36),
.B(n_7),
.Y(n_70)
);

INVx6_ASAP7_75t_SL g71 ( 
.A(n_40),
.Y(n_71)
);

INVx6_ASAP7_75t_SL g143 ( 
.A(n_71),
.Y(n_143)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_40),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_72),
.Y(n_93)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_73),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

BUFx10_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_16),
.B(n_14),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_76),
.B(n_12),
.Y(n_142)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

AND2x4_ASAP7_75t_L g80 ( 
.A(n_42),
.B(n_14),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_80),
.A2(n_11),
.B(n_13),
.Y(n_135)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_20),
.B(n_7),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_16),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_16),
.Y(n_86)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_37),
.B(n_6),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_87),
.B(n_89),
.Y(n_144)
);

BUFx24_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_88),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_43),
.B(n_6),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_60),
.B(n_35),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_94),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_52),
.B1(n_92),
.B2(n_90),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_104),
.A2(n_86),
.B1(n_79),
.B2(n_54),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_85),
.A2(n_30),
.B1(n_29),
.B2(n_23),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_118),
.A2(n_34),
.B1(n_23),
.B2(n_29),
.Y(n_173)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_45),
.Y(n_127)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_88),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_41),
.Y(n_149)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_49),
.Y(n_131)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_131),
.Y(n_180)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_133),
.Y(n_185)
);

NAND3xp33_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_142),
.C(n_11),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_66),
.B(n_41),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_137),
.B(n_139),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_66),
.B(n_41),
.Y(n_139)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_50),
.Y(n_145)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_145),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_146),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_138),
.A2(n_77),
.B1(n_88),
.B2(n_91),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_147),
.A2(n_156),
.B1(n_160),
.B2(n_189),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_80),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_148),
.B(n_157),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_149),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_80),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_153),
.B(n_154),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_117),
.A2(n_83),
.B1(n_56),
.B2(n_20),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_102),
.B(n_38),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_143),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_168),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_117),
.A2(n_20),
.B1(n_39),
.B2(n_27),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_161),
.Y(n_217)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_98),
.Y(n_162)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_162),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_94),
.B(n_38),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_163),
.B(n_177),
.Y(n_210)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_123),
.Y(n_164)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_164),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_113),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_165),
.Y(n_212)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_166),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_176),
.B1(n_184),
.B2(n_99),
.Y(n_194)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_119),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_169),
.Y(n_215)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

INVxp33_ASAP7_75t_L g221 ( 
.A(n_170),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_119),
.Y(n_171)
);

BUFx24_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_178),
.Y(n_198)
);

AO21x2_ASAP7_75t_L g192 ( 
.A1(n_173),
.A2(n_58),
.B(n_177),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_174),
.Y(n_191)
);

O2A1O1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_58),
.B(n_75),
.C(n_61),
.Y(n_175)
);

O2A1O1Ixp33_ASAP7_75t_L g206 ( 
.A1(n_175),
.A2(n_105),
.B(n_72),
.C(n_22),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_144),
.A2(n_74),
.B1(n_29),
.B2(n_34),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_124),
.B(n_21),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_93),
.Y(n_178)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_96),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_182),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_103),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_181),
.Y(n_204)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_93),
.Y(n_182)
);

BUFx10_ASAP7_75t_L g183 ( 
.A(n_105),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_183),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_L g184 ( 
.A1(n_101),
.A2(n_48),
.B1(n_75),
.B2(n_29),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_95),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_187),
.Y(n_214)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_107),
.Y(n_187)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_106),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_115),
.A2(n_27),
.B1(n_39),
.B2(n_38),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_190),
.A2(n_21),
.B1(n_110),
.B2(n_39),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_192),
.A2(n_196),
.B1(n_197),
.B2(n_225),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_194),
.A2(n_30),
.B1(n_34),
.B2(n_125),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_159),
.A2(n_101),
.B1(n_111),
.B2(n_108),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_159),
.A2(n_111),
.B1(n_108),
.B2(n_99),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_163),
.A2(n_97),
.B(n_122),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_205),
.A2(n_219),
.B(n_128),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_134),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_184),
.A2(n_109),
.B1(n_132),
.B2(n_112),
.Y(n_209)
);

AO21x2_ASAP7_75t_L g238 ( 
.A1(n_209),
.A2(n_183),
.B(n_21),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_148),
.B(n_130),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_211),
.B(n_172),
.C(n_168),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_153),
.A2(n_188),
.B(n_157),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_175),
.A2(n_96),
.B1(n_132),
.B2(n_109),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_223),
.A2(n_171),
.B1(n_181),
.B2(n_169),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_162),
.A2(n_112),
.B1(n_121),
.B2(n_100),
.Y(n_225)
);

AOI32xp33_ASAP7_75t_L g227 ( 
.A1(n_210),
.A2(n_181),
.A3(n_183),
.B1(n_116),
.B2(n_152),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_227),
.B(n_255),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_164),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_250),
.Y(n_258)
);

INVxp33_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_229),
.B(n_235),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_230),
.A2(n_236),
.B1(n_238),
.B2(n_239),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_192),
.A2(n_179),
.B1(n_170),
.B2(n_150),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_231),
.A2(n_243),
.B1(n_245),
.B2(n_206),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_182),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_232),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_223),
.A2(n_183),
.B1(n_178),
.B2(n_165),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_233),
.A2(n_204),
.B1(n_215),
.B2(n_218),
.Y(n_257)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_234),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_214),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_192),
.A2(n_161),
.B1(n_189),
.B2(n_151),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_237),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_192),
.A2(n_151),
.B1(n_166),
.B2(n_187),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_206),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_192),
.A2(n_186),
.B1(n_155),
.B2(n_180),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_242),
.A2(n_209),
.B1(n_194),
.B2(n_197),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_192),
.A2(n_100),
.B1(n_134),
.B2(n_185),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_244),
.B(n_198),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_200),
.B(n_125),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_246),
.B(n_204),
.Y(n_270)
);

MAJx2_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_110),
.C(n_27),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_249),
.C(n_196),
.Y(n_267)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_214),
.Y(n_248)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_211),
.B(n_116),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_200),
.B(n_30),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_192),
.A2(n_34),
.B1(n_30),
.B2(n_146),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_251),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_205),
.B(n_12),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_208),
.Y(n_264)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_198),
.Y(n_254)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_203),
.Y(n_256)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_257),
.A2(n_268),
.B(n_218),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_260),
.A2(n_281),
.B1(n_282),
.B2(n_241),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_263),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_264),
.B(n_228),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_267),
.B(n_284),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_235),
.B(n_202),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_285),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_270),
.Y(n_287)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_234),
.Y(n_274)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_274),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_226),
.A2(n_213),
.B1(n_221),
.B2(n_215),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_275),
.A2(n_280),
.B1(n_240),
.B2(n_238),
.Y(n_296)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_237),
.Y(n_278)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_278),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_242),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_236),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_226),
.A2(n_213),
.B1(n_215),
.B2(n_208),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_255),
.A2(n_216),
.B1(n_193),
.B2(n_207),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_248),
.A2(n_193),
.B1(n_207),
.B2(n_225),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_254),
.Y(n_283)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_283),
.Y(n_315)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_239),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_249),
.Y(n_298)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_288),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_289),
.B(n_293),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_269),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_290),
.B(n_292),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_281),
.A2(n_241),
.B(n_240),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_284),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_276),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_294),
.B(n_299),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_295),
.A2(n_301),
.B1(n_309),
.B2(n_277),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_296),
.A2(n_305),
.B1(n_273),
.B2(n_266),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_250),
.Y(n_297)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_297),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_298),
.B(n_258),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_276),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_244),
.Y(n_300)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_300),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_279),
.A2(n_231),
.B1(n_243),
.B2(n_227),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_261),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_304),
.B(n_310),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_280),
.A2(n_253),
.B1(n_238),
.B2(n_230),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_283),
.B(n_195),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_306),
.B(n_282),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_247),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_312),
.C(n_317),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_261),
.A2(n_238),
.B1(n_252),
.B2(n_199),
.Y(n_309)
);

NAND2xp33_ASAP7_75t_L g310 ( 
.A(n_265),
.B(n_238),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_311),
.B(n_313),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_267),
.B(n_201),
.C(n_217),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_268),
.B(n_252),
.Y(n_313)
);

OAI32xp33_ASAP7_75t_L g314 ( 
.A1(n_265),
.A2(n_201),
.A3(n_217),
.B1(n_224),
.B2(n_222),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_263),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_270),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_316),
.B(n_264),
.Y(n_318)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_318),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_319),
.B(n_323),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_320),
.A2(n_324),
.B1(n_343),
.B2(n_301),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_317),
.B(n_258),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_322),
.B(n_331),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_307),
.B(n_271),
.Y(n_323)
);

AOI22x1_ASAP7_75t_SL g324 ( 
.A1(n_296),
.A2(n_285),
.B1(n_275),
.B2(n_260),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_325),
.B(n_314),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_308),
.A2(n_277),
.B1(n_257),
.B2(n_238),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_327),
.A2(n_329),
.B1(n_332),
.B2(n_345),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_312),
.B(n_278),
.C(n_274),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_330),
.B(n_346),
.C(n_303),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_298),
.B(n_262),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_308),
.A2(n_262),
.B1(n_259),
.B2(n_266),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_293),
.B(n_259),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_334),
.B(n_342),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_338),
.A2(n_336),
.B1(n_335),
.B2(n_333),
.Y(n_357)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_315),
.Y(n_341)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_341),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_293),
.B(n_273),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_308),
.A2(n_199),
.B1(n_256),
.B2(n_222),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_300),
.B(n_224),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_344),
.B(n_302),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_295),
.A2(n_199),
.B1(n_218),
.B2(n_212),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_291),
.B(n_191),
.C(n_203),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_330),
.B(n_299),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g377 ( 
.A(n_347),
.Y(n_377)
);

FAx1_ASAP7_75t_L g348 ( 
.A(n_334),
.B(n_292),
.CI(n_311),
.CON(n_348),
.SN(n_348)
);

FAx1_ASAP7_75t_L g393 ( 
.A(n_348),
.B(n_355),
.CI(n_35),
.CON(n_393),
.SN(n_393)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_349),
.B(n_350),
.C(n_352),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_321),
.B(n_291),
.C(n_313),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_340),
.A2(n_294),
.B(n_313),
.Y(n_351)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_351),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_321),
.B(n_316),
.C(n_304),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_353),
.A2(n_357),
.B1(n_24),
.B2(n_10),
.Y(n_389)
);

AO22x1_ASAP7_75t_L g355 ( 
.A1(n_328),
.A2(n_287),
.B1(n_315),
.B2(n_305),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_324),
.A2(n_309),
.B1(n_297),
.B2(n_303),
.Y(n_356)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_356),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_331),
.B(n_302),
.C(n_191),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_361),
.B(n_364),
.C(n_19),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_SL g373 ( 
.A(n_362),
.B(n_344),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_363),
.B(n_367),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_322),
.B(n_203),
.C(n_41),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_333),
.Y(n_365)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_365),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_326),
.A2(n_203),
.B(n_22),
.Y(n_366)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_366),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_319),
.B(n_203),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_335),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_368),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_325),
.A2(n_41),
.B1(n_19),
.B2(n_22),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_369),
.A2(n_370),
.B1(n_339),
.B2(n_346),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_337),
.A2(n_22),
.B1(n_19),
.B2(n_2),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_373),
.B(n_376),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_372),
.B(n_323),
.Y(n_376)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_380),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_358),
.A2(n_338),
.B1(n_326),
.B2(n_339),
.Y(n_381)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_381),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_358),
.A2(n_342),
.B1(n_345),
.B2(n_327),
.Y(n_383)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_383),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_372),
.B(n_332),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_384),
.B(n_389),
.Y(n_409)
);

NOR2xp67_ASAP7_75t_SL g413 ( 
.A(n_387),
.B(n_395),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_355),
.A2(n_10),
.B1(n_13),
.B2(n_12),
.Y(n_388)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_388),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_349),
.B(n_28),
.C(n_42),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_390),
.B(n_395),
.Y(n_407)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_354),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_391),
.B(n_394),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_357),
.B(n_9),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_392),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_393),
.Y(n_408)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_359),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_350),
.B(n_28),
.C(n_35),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_378),
.A2(n_352),
.B(n_348),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_398),
.A2(n_383),
.B(n_393),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_381),
.B(n_369),
.Y(n_401)
);

XNOR2x1_ASAP7_75t_L g424 ( 
.A(n_401),
.B(n_371),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_385),
.B(n_361),
.C(n_362),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_404),
.B(n_411),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_385),
.B(n_360),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_405),
.B(n_413),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_379),
.A2(n_360),
.B(n_348),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_410),
.A2(n_393),
.B(n_386),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_384),
.B(n_367),
.C(n_364),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_377),
.A2(n_371),
.B(n_370),
.Y(n_412)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_412),
.Y(n_421)
);

BUFx24_ASAP7_75t_SL g414 ( 
.A(n_382),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_414),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_417),
.B(n_424),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_418),
.A2(n_428),
.B(n_429),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_400),
.A2(n_389),
.B1(n_392),
.B2(n_374),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_419),
.B(n_420),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_404),
.B(n_376),
.C(n_375),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_403),
.A2(n_388),
.B1(n_387),
.B2(n_390),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_422),
.B(n_425),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_402),
.A2(n_380),
.B1(n_375),
.B2(n_373),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_423),
.A2(n_427),
.B1(n_408),
.B2(n_410),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_405),
.B(n_409),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_399),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_426),
.B(n_0),
.Y(n_443)
);

OAI321xp33_ASAP7_75t_L g427 ( 
.A1(n_406),
.A2(n_9),
.A3(n_13),
.B1(n_11),
.B2(n_10),
.C(n_6),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_411),
.B(n_28),
.C(n_35),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_396),
.B(n_9),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_415),
.B(n_398),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_431),
.B(n_443),
.Y(n_450)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_434),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_425),
.B(n_409),
.C(n_401),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_435),
.B(n_438),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_416),
.B(n_408),
.Y(n_436)
);

AOI21xp33_ASAP7_75t_L g451 ( 
.A1(n_436),
.A2(n_0),
.B(n_1),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_421),
.A2(n_407),
.B(n_401),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_437),
.A2(n_439),
.B(n_441),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_416),
.B(n_397),
.C(n_28),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_420),
.A2(n_418),
.B(n_417),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_423),
.B(n_424),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_440),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_428),
.A2(n_397),
.B(n_24),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_444),
.A2(n_419),
.B(n_429),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_448),
.A2(n_453),
.B(n_432),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_442),
.B(n_430),
.C(n_28),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_449),
.B(n_435),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_451),
.A2(n_454),
.B(n_432),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_436),
.A2(n_24),
.B(n_35),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g454 ( 
.A(n_434),
.B(n_0),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_433),
.A2(n_24),
.B1(n_2),
.B2(n_3),
.Y(n_455)
);

OA21x2_ASAP7_75t_L g462 ( 
.A1(n_455),
.A2(n_1),
.B(n_3),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_450),
.B(n_449),
.Y(n_456)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_456),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_446),
.A2(n_445),
.B(n_447),
.Y(n_457)
);

AOI21x1_ASAP7_75t_L g464 ( 
.A1(n_457),
.A2(n_458),
.B(n_460),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_459),
.A2(n_462),
.B1(n_454),
.B2(n_4),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_452),
.B(n_440),
.Y(n_461)
);

NOR3xp33_ASAP7_75t_L g463 ( 
.A(n_461),
.B(n_447),
.C(n_438),
.Y(n_463)
);

NAND3xp33_ASAP7_75t_L g467 ( 
.A(n_463),
.B(n_459),
.C(n_4),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_465),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_467),
.B(n_466),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_469),
.B(n_464),
.C(n_468),
.Y(n_470)
);

AO21x1_ASAP7_75t_L g471 ( 
.A1(n_470),
.A2(n_24),
.B(n_3),
.Y(n_471)
);

NAND2x1_ASAP7_75t_L g472 ( 
.A(n_471),
.B(n_4),
.Y(n_472)
);


endmodule