module real_aes_7310_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_502;
wire n_527;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_288;
wire n_147;
wire n_404;
wire n_598;
wire n_756;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g448 ( .A(n_0), .Y(n_448) );
INVx1_ASAP7_75t_L g492 ( .A(n_1), .Y(n_492) );
INVx1_ASAP7_75t_L g189 ( .A(n_2), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_3), .A2(n_37), .B1(n_150), .B2(n_522), .Y(n_537) );
AOI21xp33_ASAP7_75t_L g157 ( .A1(n_4), .A2(n_131), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_5), .B(n_124), .Y(n_505) );
AND2x6_ASAP7_75t_L g136 ( .A(n_6), .B(n_137), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_7), .A2(n_239), .B(n_240), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_8), .B(n_38), .Y(n_449) );
INVx1_ASAP7_75t_L g164 ( .A(n_9), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_10), .B(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g129 ( .A(n_11), .Y(n_129) );
INVx1_ASAP7_75t_L g486 ( .A(n_12), .Y(n_486) );
INVx1_ASAP7_75t_L g245 ( .A(n_13), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_14), .B(n_172), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_15), .B(n_125), .Y(n_563) );
AO32x2_ASAP7_75t_L g535 ( .A1(n_16), .A2(n_124), .A3(n_169), .B1(n_514), .B2(n_536), .Y(n_535) );
OAI22xp5_ASAP7_75t_SL g112 ( .A1(n_17), .A2(n_62), .B1(n_113), .B2(n_114), .Y(n_112) );
INVx1_ASAP7_75t_L g114 ( .A(n_17), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_18), .B(n_150), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_19), .B(n_145), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_20), .B(n_125), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_21), .A2(n_50), .B1(n_150), .B2(n_522), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_22), .B(n_131), .Y(n_201) );
AOI22xp33_ASAP7_75t_SL g523 ( .A1(n_23), .A2(n_79), .B1(n_150), .B2(n_172), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_24), .B(n_150), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_25), .B(n_153), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_26), .A2(n_243), .B(n_244), .C(n_246), .Y(n_242) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_27), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_28), .B(n_166), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_29), .B(n_162), .Y(n_191) );
INVx1_ASAP7_75t_L g178 ( .A(n_30), .Y(n_178) );
OAI22xp5_ASAP7_75t_SL g106 ( .A1(n_31), .A2(n_32), .B1(n_107), .B2(n_108), .Y(n_106) );
INVx1_ASAP7_75t_L g108 ( .A(n_31), .Y(n_108) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_32), .A2(n_104), .B1(n_451), .B2(n_459), .C1(n_769), .C2(n_774), .Y(n_103) );
INVxp67_ASAP7_75t_L g107 ( .A(n_32), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_32), .B(n_166), .Y(n_552) );
INVx2_ASAP7_75t_L g134 ( .A(n_33), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_34), .B(n_150), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_35), .B(n_166), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_36), .A2(n_136), .B(n_140), .C(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g176 ( .A(n_39), .Y(n_176) );
OAI22xp5_ASAP7_75t_SL g464 ( .A1(n_40), .A2(n_465), .B1(n_468), .B2(n_469), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_40), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_41), .B(n_162), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_42), .B(n_150), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_43), .A2(n_89), .B1(n_208), .B2(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_44), .B(n_150), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_45), .B(n_150), .Y(n_487) );
CKINVDCx16_ASAP7_75t_R g179 ( .A(n_46), .Y(n_179) );
OAI22xp5_ASAP7_75t_L g465 ( .A1(n_47), .A2(n_69), .B1(n_466), .B2(n_467), .Y(n_465) );
CKINVDCx16_ASAP7_75t_R g467 ( .A(n_47), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_48), .B(n_491), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_49), .B(n_131), .Y(n_233) );
AOI22xp33_ASAP7_75t_SL g561 ( .A1(n_51), .A2(n_60), .B1(n_150), .B2(n_172), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_52), .A2(n_140), .B1(n_172), .B2(n_174), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_53), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_54), .B(n_150), .Y(n_513) );
CKINVDCx16_ASAP7_75t_R g186 ( .A(n_55), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_56), .B(n_150), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g160 ( .A1(n_57), .A2(n_149), .B(n_161), .C(n_163), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_58), .Y(n_221) );
INVx1_ASAP7_75t_L g159 ( .A(n_59), .Y(n_159) );
INVx1_ASAP7_75t_L g137 ( .A(n_61), .Y(n_137) );
INVx1_ASAP7_75t_L g113 ( .A(n_62), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_63), .B(n_150), .Y(n_493) );
INVx1_ASAP7_75t_L g128 ( .A(n_64), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_65), .Y(n_455) );
AO32x2_ASAP7_75t_L g519 ( .A1(n_66), .A2(n_124), .A3(n_225), .B1(n_514), .B2(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g512 ( .A(n_67), .Y(n_512) );
INVx1_ASAP7_75t_L g547 ( .A(n_68), .Y(n_547) );
INVx1_ASAP7_75t_L g466 ( .A(n_69), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_SL g144 ( .A1(n_70), .A2(n_145), .B(n_146), .C(n_149), .Y(n_144) );
INVxp67_ASAP7_75t_L g147 ( .A(n_71), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_72), .B(n_172), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_73), .A2(n_463), .B1(n_464), .B2(n_470), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_73), .Y(n_463) );
INVx1_ASAP7_75t_L g458 ( .A(n_74), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_75), .B(n_444), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_76), .A2(n_446), .B1(n_461), .B2(n_766), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_77), .Y(n_182) );
INVx1_ASAP7_75t_L g214 ( .A(n_78), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_80), .A2(n_136), .B(n_140), .C(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_81), .B(n_522), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_82), .B(n_172), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_83), .B(n_190), .Y(n_204) );
INVx2_ASAP7_75t_L g126 ( .A(n_84), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_85), .B(n_145), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_86), .B(n_172), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_L g187 ( .A1(n_87), .A2(n_136), .B(n_140), .C(n_188), .Y(n_187) );
OR2x2_ASAP7_75t_L g445 ( .A(n_88), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g472 ( .A(n_88), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_90), .A2(n_102), .B1(n_172), .B2(n_173), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_91), .B(n_166), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_92), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_93), .A2(n_136), .B(n_140), .C(n_228), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_94), .Y(n_235) );
INVx1_ASAP7_75t_L g143 ( .A(n_95), .Y(n_143) );
CKINVDCx16_ASAP7_75t_R g241 ( .A(n_96), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_97), .B(n_190), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_98), .B(n_172), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_99), .B(n_124), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g130 ( .A1(n_100), .A2(n_131), .B(n_138), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_101), .B(n_458), .Y(n_457) );
OAI21xp5_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_442), .B(n_450), .Y(n_104) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_109), .B1(n_110), .B2(n_441), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_106), .Y(n_441) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OAI22xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_112), .B1(n_115), .B2(n_440), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g440 ( .A(n_115), .Y(n_440) );
AOI22xp5_ASAP7_75t_SL g471 ( .A1(n_115), .A2(n_472), .B1(n_473), .B2(n_765), .Y(n_471) );
INVx3_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND4x1_ASAP7_75t_L g116 ( .A(n_117), .B(n_358), .C(n_405), .D(n_425), .Y(n_116) );
NOR3xp33_ASAP7_75t_SL g117 ( .A(n_118), .B(n_288), .C(n_313), .Y(n_117) );
OAI211xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_196), .B(n_248), .C(n_278), .Y(n_118) );
INVxp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_121), .B(n_167), .Y(n_120) );
INVx3_ASAP7_75t_SL g330 ( .A(n_121), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_121), .B(n_261), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_121), .B(n_183), .Y(n_411) );
AND2x2_ASAP7_75t_L g434 ( .A(n_121), .B(n_300), .Y(n_434) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_155), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g252 ( .A(n_123), .B(n_156), .Y(n_252) );
INVx3_ASAP7_75t_L g265 ( .A(n_123), .Y(n_265) );
AND2x2_ASAP7_75t_L g270 ( .A(n_123), .B(n_155), .Y(n_270) );
OR2x2_ASAP7_75t_L g321 ( .A(n_123), .B(n_262), .Y(n_321) );
BUFx2_ASAP7_75t_L g341 ( .A(n_123), .Y(n_341) );
AND2x2_ASAP7_75t_L g351 ( .A(n_123), .B(n_262), .Y(n_351) );
AND2x2_ASAP7_75t_L g357 ( .A(n_123), .B(n_168), .Y(n_357) );
OA21x2_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_130), .B(n_152), .Y(n_123) );
INVx4_ASAP7_75t_L g154 ( .A(n_124), .Y(n_154) );
OA21x2_ASAP7_75t_L g497 ( .A1(n_124), .A2(n_498), .B(n_505), .Y(n_497) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g169 ( .A(n_125), .Y(n_169) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
AND2x2_ASAP7_75t_SL g166 ( .A(n_126), .B(n_127), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
BUFx2_ASAP7_75t_L g239 ( .A(n_131), .Y(n_239) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_136), .Y(n_131) );
NAND2x1p5_ASAP7_75t_L g180 ( .A(n_132), .B(n_136), .Y(n_180) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
INVx1_ASAP7_75t_L g491 ( .A(n_133), .Y(n_491) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g141 ( .A(n_134), .Y(n_141) );
INVx1_ASAP7_75t_L g173 ( .A(n_134), .Y(n_173) );
INVx1_ASAP7_75t_L g142 ( .A(n_135), .Y(n_142) );
INVx1_ASAP7_75t_L g145 ( .A(n_135), .Y(n_145) );
INVx3_ASAP7_75t_L g148 ( .A(n_135), .Y(n_148) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_135), .Y(n_162) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_135), .Y(n_175) );
INVx4_ASAP7_75t_SL g151 ( .A(n_136), .Y(n_151) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_136), .A2(n_485), .B(n_489), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_136), .A2(n_499), .B(n_502), .Y(n_498) );
BUFx3_ASAP7_75t_L g514 ( .A(n_136), .Y(n_514) );
OAI21xp5_ASAP7_75t_L g526 ( .A1(n_136), .A2(n_527), .B(n_531), .Y(n_526) );
OAI21xp5_ASAP7_75t_L g545 ( .A1(n_136), .A2(n_546), .B(n_549), .Y(n_545) );
O2A1O1Ixp33_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_143), .B(n_144), .C(n_151), .Y(n_138) );
O2A1O1Ixp33_ASAP7_75t_L g158 ( .A1(n_139), .A2(n_151), .B(n_159), .C(n_160), .Y(n_158) );
O2A1O1Ixp33_ASAP7_75t_L g240 ( .A1(n_139), .A2(n_151), .B(n_241), .C(n_242), .Y(n_240) );
INVx5_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_141), .Y(n_150) );
BUFx3_ASAP7_75t_L g208 ( .A(n_141), .Y(n_208) );
INVx1_ASAP7_75t_L g522 ( .A(n_141), .Y(n_522) );
INVx1_ASAP7_75t_L g530 ( .A(n_145), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_148), .B(n_164), .Y(n_163) );
INVx5_ASAP7_75t_L g190 ( .A(n_148), .Y(n_190) );
OAI22xp5_ASAP7_75t_SL g520 ( .A1(n_148), .A2(n_162), .B1(n_521), .B2(n_523), .Y(n_520) );
O2A1O1Ixp5_ASAP7_75t_SL g546 ( .A1(n_149), .A2(n_190), .B(n_547), .C(n_548), .Y(n_546) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_150), .Y(n_232) );
OAI22xp33_ASAP7_75t_L g170 ( .A1(n_151), .A2(n_171), .B1(n_179), .B2(n_180), .Y(n_170) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_153), .A2(n_157), .B(n_165), .Y(n_156) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NOR2xp33_ASAP7_75t_SL g210 ( .A(n_154), .B(n_211), .Y(n_210) );
AO21x1_ASAP7_75t_L g558 ( .A1(n_154), .A2(n_559), .B(n_562), .Y(n_558) );
NAND3xp33_ASAP7_75t_L g577 ( .A(n_154), .B(n_514), .C(n_559), .Y(n_577) );
INVx1_ASAP7_75t_SL g155 ( .A(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_156), .B(n_262), .Y(n_276) );
INVx2_ASAP7_75t_L g286 ( .A(n_156), .Y(n_286) );
AND2x2_ASAP7_75t_L g299 ( .A(n_156), .B(n_265), .Y(n_299) );
OR2x2_ASAP7_75t_L g310 ( .A(n_156), .B(n_262), .Y(n_310) );
AND2x2_ASAP7_75t_SL g356 ( .A(n_156), .B(n_357), .Y(n_356) );
BUFx2_ASAP7_75t_L g368 ( .A(n_156), .Y(n_368) );
AND2x2_ASAP7_75t_L g414 ( .A(n_156), .B(n_168), .Y(n_414) );
O2A1O1Ixp5_ASAP7_75t_L g511 ( .A1(n_161), .A2(n_490), .B(n_512), .C(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_161), .A2(n_532), .B(n_533), .Y(n_531) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx4_ASAP7_75t_L g231 ( .A(n_162), .Y(n_231) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_162), .A2(n_494), .B1(n_537), .B2(n_538), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_162), .A2(n_494), .B1(n_560), .B2(n_561), .Y(n_559) );
INVx1_ASAP7_75t_L g195 ( .A(n_166), .Y(n_195) );
INVx2_ASAP7_75t_L g225 ( .A(n_166), .Y(n_225) );
OA21x2_ASAP7_75t_L g237 ( .A1(n_166), .A2(n_238), .B(n_247), .Y(n_237) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_166), .A2(n_526), .B(n_534), .Y(n_525) );
OA21x2_ASAP7_75t_L g544 ( .A1(n_166), .A2(n_545), .B(n_552), .Y(n_544) );
INVx3_ASAP7_75t_SL g287 ( .A(n_167), .Y(n_287) );
OR2x2_ASAP7_75t_L g340 ( .A(n_167), .B(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_183), .Y(n_167) );
INVx3_ASAP7_75t_L g262 ( .A(n_168), .Y(n_262) );
AND2x2_ASAP7_75t_L g329 ( .A(n_168), .B(n_184), .Y(n_329) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_168), .Y(n_397) );
AOI33xp33_ASAP7_75t_L g401 ( .A1(n_168), .A2(n_330), .A3(n_337), .B1(n_346), .B2(n_402), .B3(n_403), .Y(n_401) );
AO21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_181), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_169), .B(n_182), .Y(n_181) );
AO21x2_ASAP7_75t_L g184 ( .A1(n_169), .A2(n_185), .B(n_193), .Y(n_184) );
INVx2_ASAP7_75t_L g209 ( .A(n_169), .Y(n_209) );
INVx2_ASAP7_75t_L g192 ( .A(n_172), .Y(n_192) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
OAI22xp5_ASAP7_75t_SL g174 ( .A1(n_175), .A2(n_176), .B1(n_177), .B2(n_178), .Y(n_174) );
INVx2_ASAP7_75t_L g177 ( .A(n_175), .Y(n_177) );
INVx4_ASAP7_75t_L g243 ( .A(n_175), .Y(n_243) );
OAI21xp5_ASAP7_75t_L g185 ( .A1(n_180), .A2(n_186), .B(n_187), .Y(n_185) );
OAI21xp5_ASAP7_75t_L g213 ( .A1(n_180), .A2(n_214), .B(n_215), .Y(n_213) );
INVx1_ASAP7_75t_L g250 ( .A(n_183), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_183), .B(n_265), .Y(n_264) );
NOR3xp33_ASAP7_75t_L g324 ( .A(n_183), .B(n_325), .C(n_327), .Y(n_324) );
AND2x2_ASAP7_75t_L g350 ( .A(n_183), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_183), .B(n_357), .Y(n_360) );
AND2x2_ASAP7_75t_L g413 ( .A(n_183), .B(n_414), .Y(n_413) );
INVx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx3_ASAP7_75t_L g269 ( .A(n_184), .Y(n_269) );
OR2x2_ASAP7_75t_L g363 ( .A(n_184), .B(n_262), .Y(n_363) );
O2A1O1Ixp33_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_191), .C(n_192), .Y(n_188) );
INVx2_ASAP7_75t_L g494 ( .A(n_190), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_190), .A2(n_500), .B(n_501), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_190), .A2(n_509), .B(n_510), .Y(n_508) );
O2A1O1Ixp33_ASAP7_75t_L g485 ( .A1(n_192), .A2(n_486), .B(n_487), .C(n_488), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_195), .B(n_221), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_195), .B(n_235), .Y(n_234) );
OR2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_222), .Y(n_196) );
AOI32xp33_ASAP7_75t_L g314 ( .A1(n_197), .A2(n_315), .A3(n_317), .B1(n_319), .B2(n_322), .Y(n_314) );
NOR2xp67_ASAP7_75t_L g387 ( .A(n_197), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g417 ( .A(n_197), .Y(n_417) );
INVx4_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g349 ( .A(n_198), .B(n_333), .Y(n_349) );
AND2x2_ASAP7_75t_L g369 ( .A(n_198), .B(n_295), .Y(n_369) );
AND2x2_ASAP7_75t_L g437 ( .A(n_198), .B(n_355), .Y(n_437) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_212), .Y(n_198) );
INVx3_ASAP7_75t_L g258 ( .A(n_199), .Y(n_258) );
AND2x2_ASAP7_75t_L g272 ( .A(n_199), .B(n_256), .Y(n_272) );
OR2x2_ASAP7_75t_L g277 ( .A(n_199), .B(n_255), .Y(n_277) );
INVx1_ASAP7_75t_L g284 ( .A(n_199), .Y(n_284) );
AND2x2_ASAP7_75t_L g292 ( .A(n_199), .B(n_266), .Y(n_292) );
AND2x2_ASAP7_75t_L g294 ( .A(n_199), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_199), .B(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g347 ( .A(n_199), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_199), .B(n_432), .Y(n_431) );
OR2x6_ASAP7_75t_L g199 ( .A(n_200), .B(n_210), .Y(n_199) );
AOI21xp5_ASAP7_75t_SL g200 ( .A1(n_201), .A2(n_202), .B(n_209), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_206), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_206), .A2(n_217), .B(n_218), .Y(n_216) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g246 ( .A(n_208), .Y(n_246) );
INVx1_ASAP7_75t_L g219 ( .A(n_209), .Y(n_219) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_209), .A2(n_484), .B(n_495), .Y(n_483) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_209), .A2(n_507), .B(n_515), .Y(n_506) );
INVx2_ASAP7_75t_L g256 ( .A(n_212), .Y(n_256) );
AND2x2_ASAP7_75t_L g302 ( .A(n_212), .B(n_223), .Y(n_302) );
AND2x2_ASAP7_75t_L g312 ( .A(n_212), .B(n_237), .Y(n_312) );
AO21x2_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_219), .B(n_220), .Y(n_212) );
INVx2_ASAP7_75t_L g432 ( .A(n_222), .Y(n_432) );
OR2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_236), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_223), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g273 ( .A(n_223), .Y(n_273) );
AND2x2_ASAP7_75t_L g317 ( .A(n_223), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g333 ( .A(n_223), .B(n_296), .Y(n_333) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g281 ( .A(n_224), .Y(n_281) );
AND2x2_ASAP7_75t_L g295 ( .A(n_224), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g346 ( .A(n_224), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_224), .B(n_256), .Y(n_378) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_234), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_227), .B(n_233), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_232), .Y(n_228) );
AND2x2_ASAP7_75t_L g257 ( .A(n_236), .B(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g318 ( .A(n_236), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_236), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g355 ( .A(n_236), .Y(n_355) );
INVx1_ASAP7_75t_L g388 ( .A(n_236), .Y(n_388) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g266 ( .A(n_237), .B(n_256), .Y(n_266) );
INVx1_ASAP7_75t_L g296 ( .A(n_237), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_243), .B(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g488 ( .A(n_243), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_243), .A2(n_550), .B(n_551), .Y(n_549) );
AOI221xp5_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_253), .B1(n_259), .B2(n_266), .C(n_267), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_250), .B(n_270), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_250), .B(n_333), .Y(n_410) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_252), .B(n_300), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_252), .B(n_261), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_252), .B(n_275), .Y(n_404) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_257), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g326 ( .A(n_256), .Y(n_326) );
AND2x2_ASAP7_75t_L g301 ( .A(n_257), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g379 ( .A(n_257), .Y(n_379) );
AND2x2_ASAP7_75t_L g311 ( .A(n_258), .B(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_258), .B(n_281), .Y(n_327) );
AND2x2_ASAP7_75t_L g391 ( .A(n_258), .B(n_317), .Y(n_391) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
BUFx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g300 ( .A(n_262), .B(n_269), .Y(n_300) );
AND2x2_ASAP7_75t_L g396 ( .A(n_263), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_265), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_266), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_266), .B(n_273), .Y(n_361) );
AND2x2_ASAP7_75t_L g381 ( .A(n_266), .B(n_281), .Y(n_381) );
AND2x2_ASAP7_75t_L g402 ( .A(n_266), .B(n_346), .Y(n_402) );
OAI32xp33_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_271), .A3(n_273), .B1(n_274), .B2(n_277), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx1_ASAP7_75t_SL g275 ( .A(n_269), .Y(n_275) );
NAND2x1_ASAP7_75t_L g316 ( .A(n_269), .B(n_299), .Y(n_316) );
OR2x2_ASAP7_75t_L g320 ( .A(n_269), .B(n_321), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_269), .B(n_368), .Y(n_421) );
INVx1_ASAP7_75t_L g289 ( .A(n_270), .Y(n_289) );
OAI221xp5_ASAP7_75t_SL g407 ( .A1(n_271), .A2(n_362), .B1(n_408), .B2(n_411), .C(n_412), .Y(n_407) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g279 ( .A(n_272), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g322 ( .A(n_272), .B(n_295), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_272), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g400 ( .A(n_272), .B(n_333), .Y(n_400) );
INVxp67_ASAP7_75t_L g336 ( .A(n_273), .Y(n_336) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
AND2x2_ASAP7_75t_L g406 ( .A(n_275), .B(n_393), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_275), .B(n_356), .Y(n_429) );
INVx1_ASAP7_75t_L g304 ( .A(n_277), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g385 ( .A(n_277), .B(n_386), .Y(n_385) );
OR2x2_ASAP7_75t_L g422 ( .A(n_277), .B(n_423), .Y(n_422) );
OAI21xp5_ASAP7_75t_SL g278 ( .A1(n_279), .A2(n_282), .B(n_285), .Y(n_278) );
AND2x2_ASAP7_75t_L g291 ( .A(n_280), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g375 ( .A(n_284), .B(n_295), .Y(n_375) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
AND2x2_ASAP7_75t_L g393 ( .A(n_286), .B(n_351), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_286), .B(n_350), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_287), .B(n_299), .Y(n_373) );
OAI211xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_290), .B(n_293), .C(n_303), .Y(n_288) );
AOI221xp5_ASAP7_75t_L g323 ( .A1(n_289), .A2(n_324), .B1(n_328), .B2(n_331), .C(n_334), .Y(n_323) );
AOI31xp33_ASAP7_75t_L g418 ( .A1(n_289), .A2(n_419), .A3(n_420), .B(n_422), .Y(n_418) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AOI22xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_297), .B1(n_299), .B2(n_301), .Y(n_293) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx1_ASAP7_75t_L g419 ( .A(n_299), .Y(n_419) );
INVx1_ASAP7_75t_L g382 ( .A(n_300), .Y(n_382) );
O2A1O1Ixp33_ASAP7_75t_L g425 ( .A1(n_302), .A2(n_426), .B(n_428), .C(n_430), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_305), .B1(n_307), .B2(n_311), .Y(n_303) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_308), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OAI221xp5_ASAP7_75t_SL g398 ( .A1(n_310), .A2(n_344), .B1(n_363), .B2(n_399), .C(n_401), .Y(n_398) );
INVx1_ASAP7_75t_L g394 ( .A(n_311), .Y(n_394) );
INVx1_ASAP7_75t_L g348 ( .A(n_312), .Y(n_348) );
NAND3xp33_ASAP7_75t_SL g313 ( .A(n_314), .B(n_323), .C(n_338), .Y(n_313) );
OAI21xp33_ASAP7_75t_L g364 ( .A1(n_315), .A2(n_365), .B(n_369), .Y(n_364) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_317), .B(n_417), .Y(n_416) );
INVxp67_ASAP7_75t_L g424 ( .A(n_318), .Y(n_424) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g362 ( .A(n_325), .B(n_345), .Y(n_362) );
INVx1_ASAP7_75t_L g337 ( .A(n_326), .Y(n_337) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g335 ( .A(n_329), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_329), .B(n_367), .Y(n_366) );
NOR4xp25_ASAP7_75t_L g334 ( .A(n_330), .B(n_335), .C(n_336), .D(n_337), .Y(n_334) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AOI222xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_343), .B1(n_349), .B2(n_350), .C1(n_352), .C2(n_356), .Y(n_338) );
NAND2xp5_ASAP7_75t_SL g339 ( .A(n_340), .B(n_342), .Y(n_339) );
INVx1_ASAP7_75t_L g436 ( .A(n_340), .Y(n_436) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_348), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_352), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OAI21xp5_ASAP7_75t_SL g412 ( .A1(n_357), .A2(n_413), .B(n_415), .Y(n_412) );
NOR4xp25_ASAP7_75t_L g358 ( .A(n_359), .B(n_370), .C(n_383), .D(n_398), .Y(n_358) );
OAI221xp5_ASAP7_75t_SL g359 ( .A1(n_360), .A2(n_361), .B1(n_362), .B2(n_363), .C(n_364), .Y(n_359) );
INVx1_ASAP7_75t_L g439 ( .A(n_360), .Y(n_439) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_367), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
OAI222xp33_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_374), .B1(n_376), .B2(n_377), .C1(n_380), .C2(n_382), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AOI211xp5_ASAP7_75t_L g405 ( .A1(n_375), .A2(n_406), .B(n_407), .C(n_418), .Y(n_405) );
OR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx1_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
OAI222xp33_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_389), .B1(n_390), .B2(n_392), .C1(n_394), .C2(n_395), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVxp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_400), .A2(n_403), .B1(n_436), .B2(n_437), .Y(n_435) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OAI211xp5_ASAP7_75t_SL g430 ( .A1(n_431), .A2(n_433), .B(n_435), .C(n_438), .Y(n_430) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_SL g773 ( .A(n_445), .Y(n_773) );
BUFx2_ASAP7_75t_L g776 ( .A(n_445), .Y(n_776) );
NOR2x2_ASAP7_75t_L g768 ( .A(n_446), .B(n_472), .Y(n_768) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_456), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NOR2xp33_ASAP7_75t_SL g771 ( .A(n_455), .B(n_457), .Y(n_771) );
OA21x2_ASAP7_75t_L g775 ( .A1(n_455), .A2(n_456), .B(n_776), .Y(n_775) );
INVx1_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
INVxp67_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
XNOR2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_471), .Y(n_461) );
INVx1_ASAP7_75t_L g470 ( .A(n_464), .Y(n_470) );
INVx1_ASAP7_75t_L g468 ( .A(n_465), .Y(n_468) );
INVx2_ASAP7_75t_L g765 ( .A(n_472), .Y(n_765) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_SL g474 ( .A(n_475), .B(n_731), .Y(n_474) );
NOR3xp33_ASAP7_75t_L g475 ( .A(n_476), .B(n_635), .C(n_719), .Y(n_475) );
NAND4xp25_ASAP7_75t_L g476 ( .A(n_477), .B(n_578), .C(n_600), .D(n_616), .Y(n_476) );
AOI221xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_516), .B1(n_539), .B2(n_557), .C(n_564), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_496), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_480), .B(n_557), .Y(n_590) );
NAND4xp25_ASAP7_75t_L g630 ( .A(n_480), .B(n_618), .C(n_631), .D(n_633), .Y(n_630) );
INVxp67_ASAP7_75t_L g747 ( .A(n_480), .Y(n_747) );
INVx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OR2x2_ASAP7_75t_L g629 ( .A(n_481), .B(n_567), .Y(n_629) );
AND2x2_ASAP7_75t_L g653 ( .A(n_481), .B(n_496), .Y(n_653) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g620 ( .A(n_482), .B(n_556), .Y(n_620) );
AND2x2_ASAP7_75t_L g660 ( .A(n_482), .B(n_641), .Y(n_660) );
AND2x2_ASAP7_75t_L g677 ( .A(n_482), .B(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_482), .B(n_497), .Y(n_701) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g555 ( .A(n_483), .B(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g572 ( .A(n_483), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g584 ( .A(n_483), .B(n_497), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_483), .B(n_506), .Y(n_606) );
O2A1O1Ixp33_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_492), .B(n_493), .C(n_494), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_494), .A2(n_503), .B(n_504), .Y(n_502) );
AND2x2_ASAP7_75t_L g587 ( .A(n_496), .B(n_588), .Y(n_587) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_496), .A2(n_637), .B1(n_640), .B2(n_642), .C(n_646), .Y(n_636) );
AND2x2_ASAP7_75t_L g695 ( .A(n_496), .B(n_660), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_496), .B(n_677), .Y(n_729) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_506), .Y(n_496) );
INVx3_ASAP7_75t_L g556 ( .A(n_497), .Y(n_556) );
AND2x2_ASAP7_75t_L g604 ( .A(n_497), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g658 ( .A(n_497), .B(n_573), .Y(n_658) );
AND2x2_ASAP7_75t_L g716 ( .A(n_497), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g557 ( .A(n_506), .B(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g573 ( .A(n_506), .Y(n_573) );
INVx1_ASAP7_75t_L g628 ( .A(n_506), .Y(n_628) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_506), .Y(n_634) );
AND2x2_ASAP7_75t_L g679 ( .A(n_506), .B(n_556), .Y(n_679) );
OR2x2_ASAP7_75t_L g718 ( .A(n_506), .B(n_558), .Y(n_718) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_511), .B(n_514), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_516), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_524), .Y(n_516) );
AND2x2_ASAP7_75t_L g714 ( .A(n_517), .B(n_711), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_517), .B(n_696), .Y(n_746) );
BUFx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g645 ( .A(n_518), .B(n_569), .Y(n_645) );
AND2x2_ASAP7_75t_L g694 ( .A(n_518), .B(n_542), .Y(n_694) );
INVx1_ASAP7_75t_L g740 ( .A(n_518), .Y(n_740) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_519), .Y(n_554) );
AND2x2_ASAP7_75t_L g595 ( .A(n_519), .B(n_569), .Y(n_595) );
INVx1_ASAP7_75t_L g612 ( .A(n_519), .Y(n_612) );
AND2x2_ASAP7_75t_L g618 ( .A(n_519), .B(n_535), .Y(n_618) );
AND2x2_ASAP7_75t_L g686 ( .A(n_524), .B(n_594), .Y(n_686) );
INVx2_ASAP7_75t_L g751 ( .A(n_524), .Y(n_751) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_535), .Y(n_524) );
AND2x2_ASAP7_75t_L g568 ( .A(n_525), .B(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g581 ( .A(n_525), .B(n_543), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_525), .B(n_542), .Y(n_609) );
INVx1_ASAP7_75t_L g615 ( .A(n_525), .Y(n_615) );
INVx1_ASAP7_75t_L g632 ( .A(n_525), .Y(n_632) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_525), .Y(n_644) );
INVx2_ASAP7_75t_L g712 ( .A(n_525), .Y(n_712) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_529), .B(n_530), .Y(n_527) );
INVx2_ASAP7_75t_L g569 ( .A(n_535), .Y(n_569) );
BUFx2_ASAP7_75t_L g666 ( .A(n_535), .Y(n_666) );
AND2x2_ASAP7_75t_L g711 ( .A(n_535), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_553), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_541), .B(n_648), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_541), .A2(n_710), .B(n_724), .Y(n_734) );
AND2x2_ASAP7_75t_L g759 ( .A(n_541), .B(n_645), .Y(n_759) );
BUFx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g681 ( .A(n_543), .Y(n_681) );
AND2x2_ASAP7_75t_L g710 ( .A(n_543), .B(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_544), .Y(n_594) );
INVx2_ASAP7_75t_L g613 ( .A(n_544), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_544), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
INVx2_ASAP7_75t_L g567 ( .A(n_554), .Y(n_567) );
OR2x2_ASAP7_75t_L g580 ( .A(n_554), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g648 ( .A(n_554), .B(n_644), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_554), .B(n_744), .Y(n_743) );
OR2x2_ASAP7_75t_L g749 ( .A(n_554), .B(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_554), .B(n_686), .Y(n_761) );
AND2x2_ASAP7_75t_L g640 ( .A(n_555), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g663 ( .A(n_555), .B(n_557), .Y(n_663) );
INVx2_ASAP7_75t_L g575 ( .A(n_556), .Y(n_575) );
AND2x2_ASAP7_75t_L g603 ( .A(n_556), .B(n_576), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_556), .B(n_628), .Y(n_684) );
AND2x2_ASAP7_75t_L g598 ( .A(n_557), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g745 ( .A(n_557), .Y(n_745) );
AND2x2_ASAP7_75t_L g757 ( .A(n_557), .B(n_620), .Y(n_757) );
AND2x2_ASAP7_75t_L g583 ( .A(n_558), .B(n_573), .Y(n_583) );
INVx1_ASAP7_75t_L g678 ( .A(n_558), .Y(n_678) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x4_ASAP7_75t_L g576 ( .A(n_563), .B(n_577), .Y(n_576) );
INVxp67_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_570), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_567), .B(n_614), .Y(n_623) );
OR2x2_ASAP7_75t_L g755 ( .A(n_567), .B(n_756), .Y(n_755) );
AND2x2_ASAP7_75t_L g672 ( .A(n_568), .B(n_613), .Y(n_672) );
AND2x2_ASAP7_75t_L g680 ( .A(n_568), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g739 ( .A(n_568), .B(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g763 ( .A(n_568), .B(n_610), .Y(n_763) );
NOR2xp67_ASAP7_75t_L g721 ( .A(n_569), .B(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g750 ( .A(n_569), .B(n_613), .Y(n_750) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2x1p5_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
AND2x2_ASAP7_75t_L g602 ( .A(n_572), .B(n_603), .Y(n_602) );
INVxp67_ASAP7_75t_L g764 ( .A(n_572), .Y(n_764) );
NOR2x1_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
INVx1_ASAP7_75t_L g599 ( .A(n_575), .Y(n_599) );
AND2x2_ASAP7_75t_L g650 ( .A(n_575), .B(n_583), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_575), .B(n_718), .Y(n_744) );
INVx2_ASAP7_75t_L g589 ( .A(n_576), .Y(n_589) );
INVx3_ASAP7_75t_L g641 ( .A(n_576), .Y(n_641) );
OR2x2_ASAP7_75t_L g669 ( .A(n_576), .B(n_670), .Y(n_669) );
AOI311xp33_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_582), .A3(n_584), .B(n_585), .C(n_596), .Y(n_578) );
O2A1O1Ixp33_ASAP7_75t_L g616 ( .A1(n_579), .A2(n_617), .B(n_619), .C(n_621), .Y(n_616) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx2_ASAP7_75t_SL g601 ( .A(n_581), .Y(n_601) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g619 ( .A(n_583), .B(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_583), .B(n_599), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_583), .B(n_584), .Y(n_752) );
AND2x2_ASAP7_75t_L g674 ( .A(n_584), .B(n_588), .Y(n_674) );
AOI21xp33_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_590), .B(n_591), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g732 ( .A(n_588), .B(n_620), .Y(n_732) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_589), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g626 ( .A(n_589), .Y(n_626) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
AND2x2_ASAP7_75t_L g617 ( .A(n_593), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g662 ( .A(n_595), .Y(n_662) );
AND2x4_ASAP7_75t_L g724 ( .A(n_595), .B(n_693), .Y(n_724) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AOI222xp33_ASAP7_75t_L g675 ( .A1(n_598), .A2(n_664), .B1(n_676), .B2(n_680), .C1(n_682), .C2(n_686), .Y(n_675) );
A2O1A1Ixp33_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B(n_604), .C(n_607), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_601), .B(n_645), .Y(n_668) );
INVx1_ASAP7_75t_L g690 ( .A(n_603), .Y(n_690) );
INVx1_ASAP7_75t_L g624 ( .A(n_605), .Y(n_624) );
OR2x2_ASAP7_75t_L g689 ( .A(n_606), .B(n_690), .Y(n_689) );
OAI21xp33_ASAP7_75t_SL g607 ( .A1(n_608), .A2(n_610), .B(n_614), .Y(n_607) );
NAND3xp33_ASAP7_75t_L g625 ( .A(n_608), .B(n_626), .C(n_627), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_608), .A2(n_645), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_612), .Y(n_665) );
AND2x2_ASAP7_75t_SL g631 ( .A(n_613), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g722 ( .A(n_613), .Y(n_722) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_613), .Y(n_738) );
INVx2_ASAP7_75t_L g696 ( .A(n_614), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_618), .B(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g670 ( .A(n_620), .Y(n_670) );
OAI221xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_624), .B1(n_625), .B2(n_629), .C(n_630), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g703 ( .A(n_624), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_SL g758 ( .A(n_624), .Y(n_758) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g639 ( .A(n_631), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_631), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g697 ( .A(n_631), .B(n_645), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_631), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g730 ( .A(n_631), .B(n_665), .Y(n_730) );
BUFx3_ASAP7_75t_L g693 ( .A(n_632), .Y(n_693) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND5xp2_ASAP7_75t_L g635 ( .A(n_636), .B(n_654), .C(n_675), .D(n_687), .E(n_702), .Y(n_635) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AOI32xp33_ASAP7_75t_L g727 ( .A1(n_639), .A2(n_666), .A3(n_682), .B1(n_728), .B2(n_730), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_641), .B(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_SL g651 ( .A(n_645), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_649), .B1(n_651), .B2(n_652), .Y(n_646) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_661), .B1(n_663), .B2(n_664), .C(n_667), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OR2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g726 ( .A(n_658), .B(n_677), .Y(n_726) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AOI221xp5_ASAP7_75t_L g741 ( .A1(n_663), .A2(n_724), .B1(n_742), .B2(n_747), .C(n_748), .Y(n_741) );
AND2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
INVx2_ASAP7_75t_L g707 ( .A(n_666), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B1(n_671), .B2(n_673), .Y(n_667) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_679), .Y(n_676) );
INVx1_ASAP7_75t_L g685 ( .A(n_677), .Y(n_685) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OR2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
AOI222xp33_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_691), .B1(n_695), .B2(n_696), .C1(n_697), .C2(n_698), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_694), .Y(n_691) );
INVxp67_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
OAI22xp33_ASAP7_75t_L g742 ( .A1(n_696), .A2(n_743), .B1(n_745), .B2(n_746), .Y(n_742) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_705), .B(n_708), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AOI21xp33_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_713), .B(n_715), .Y(n_708) );
INVx2_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g756 ( .A(n_711), .Y(n_756) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
A2O1A1Ixp33_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_723), .B(n_725), .C(n_727), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
AOI211xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_733), .B(n_735), .C(n_760), .Y(n_731) );
CKINVDCx16_ASAP7_75t_R g736 ( .A(n_732), .Y(n_736) );
INVxp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OAI211xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_737), .B(n_741), .C(n_753), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
AOI21xp33_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_751), .B(n_752), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_757), .B1(n_758), .B2(n_759), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
AOI21xp33_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_762), .B(n_764), .Y(n_760) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_SL g769 ( .A(n_770), .Y(n_769) );
NAND2xp33_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
INVx1_ASAP7_75t_SL g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_SL g774 ( .A(n_775), .Y(n_774) );
endmodule