module fake_jpeg_27520_n_106 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_106);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_26),
.B(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_0),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_33),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_20),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_32),
.B(n_16),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_4),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_39),
.A2(n_8),
.B(n_9),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_13),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_48),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_12),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_45),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_29),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_22),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_60),
.Y(n_77)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_31),
.C(n_24),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_47),
.C(n_49),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_18),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_59),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_25),
.B1(n_28),
.B2(n_22),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_57),
.A2(n_61),
.B1(n_35),
.B2(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_23),
.Y(n_58)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_11),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_49),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_36),
.A2(n_25),
.B1(n_9),
.B2(n_10),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_51),
.Y(n_79)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

BUFx4f_ASAP7_75t_SL g74 ( 
.A(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_75),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_76),
.A2(n_41),
.B1(n_65),
.B2(n_56),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_54),
.C(n_51),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_79),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_59),
.B1(n_55),
.B2(n_53),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_80),
.A2(n_81),
.B1(n_82),
.B2(n_73),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_76),
.A2(n_35),
.B1(n_61),
.B2(n_41),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_77),
.B(n_67),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_70),
.B(n_74),
.Y(n_91)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_89),
.Y(n_93)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

NAND2xp33_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_81),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_95),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_91),
.A2(n_84),
.B1(n_78),
.B2(n_79),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_87),
.B(n_72),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_99),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_93),
.A2(n_87),
.B(n_69),
.Y(n_99)
);

BUFx24_ASAP7_75t_SL g101 ( 
.A(n_100),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_101),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_103),
.A2(n_96),
.B(n_95),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_104),
.Y(n_106)
);


endmodule