module real_aes_16340_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g109 ( .A(n_0), .B(n_110), .Y(n_109) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_1), .A2(n_4), .B1(n_267), .B2(n_268), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_2), .A2(n_42), .B1(n_168), .B2(n_216), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_3), .A2(n_24), .B1(n_216), .B2(n_250), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_5), .A2(n_16), .B1(n_517), .B2(n_544), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g152 ( .A1(n_6), .A2(n_59), .B1(n_153), .B2(n_154), .Y(n_152) );
AOI22xp5_ASAP7_75t_L g167 ( .A1(n_7), .A2(n_17), .B1(n_168), .B2(n_169), .Y(n_167) );
INVx1_ASAP7_75t_L g110 ( .A(n_8), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_9), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_10), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_11), .A2(n_18), .B1(n_518), .B2(n_562), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g128 ( .A1(n_12), .A2(n_129), .B1(n_793), .B2(n_794), .Y(n_128) );
INVx1_ASAP7_75t_L g793 ( .A(n_12), .Y(n_793) );
BUFx2_ASAP7_75t_L g115 ( .A(n_13), .Y(n_115) );
OR2x2_ASAP7_75t_L g127 ( .A(n_13), .B(n_37), .Y(n_127) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_14), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g546 ( .A(n_15), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_19), .A2(n_96), .B1(n_268), .B2(n_517), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_20), .A2(n_38), .B1(n_146), .B2(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_21), .B(n_144), .Y(n_578) );
OAI21x1_ASAP7_75t_L g158 ( .A1(n_22), .A2(n_57), .B(n_159), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_23), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_25), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_26), .B(n_141), .Y(n_208) );
INVx4_ASAP7_75t_R g192 ( .A(n_27), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_28), .A2(n_46), .B1(n_172), .B2(n_265), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_29), .A2(n_53), .B1(n_172), .B2(n_517), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g512 ( .A(n_30), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_31), .B(n_542), .Y(n_580) );
CKINVDCx5p33_ASAP7_75t_R g523 ( .A(n_32), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_33), .B(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g272 ( .A(n_34), .Y(n_272) );
A2O1A1Ixp33_ASAP7_75t_SL g247 ( .A1(n_35), .A2(n_140), .B(n_168), .C(n_248), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_36), .A2(n_54), .B1(n_168), .B2(n_172), .Y(n_256) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_37), .Y(n_113) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_39), .A2(n_84), .B1(n_168), .B2(n_509), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g808 ( .A1(n_40), .A2(n_809), .B1(n_810), .B2(n_811), .Y(n_808) );
INVx1_ASAP7_75t_L g811 ( .A(n_40), .Y(n_811) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_41), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_43), .A2(n_45), .B1(n_168), .B2(n_169), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_44), .A2(n_58), .B1(n_517), .B2(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g212 ( .A(n_47), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_48), .B(n_168), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_49), .Y(n_226) );
INVx2_ASAP7_75t_L g122 ( .A(n_50), .Y(n_122) );
INVx1_ASAP7_75t_L g105 ( .A(n_51), .Y(n_105) );
BUFx3_ASAP7_75t_L g125 ( .A(n_51), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g818 ( .A(n_52), .Y(n_818) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_55), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g171 ( .A1(n_56), .A2(n_85), .B1(n_168), .B2(n_172), .Y(n_171) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_60), .A2(n_72), .B1(n_265), .B2(n_534), .Y(n_551) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_61), .Y(n_178) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_62), .A2(n_76), .B1(n_168), .B2(n_169), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_63), .A2(n_95), .B1(n_517), .B2(n_518), .Y(n_516) );
INVx1_ASAP7_75t_L g159 ( .A(n_64), .Y(n_159) );
AND2x4_ASAP7_75t_L g162 ( .A(n_65), .B(n_163), .Y(n_162) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_66), .A2(n_87), .B1(n_172), .B2(n_265), .Y(n_264) );
AO22x1_ASAP7_75t_L g142 ( .A1(n_67), .A2(n_74), .B1(n_143), .B2(n_146), .Y(n_142) );
INVx1_ASAP7_75t_L g163 ( .A(n_68), .Y(n_163) );
AND2x2_ASAP7_75t_L g251 ( .A(n_69), .B(n_204), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_70), .B(n_153), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_71), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_73), .A2(n_100), .B1(n_116), .B2(n_825), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_75), .B(n_216), .Y(n_227) );
INVx2_ASAP7_75t_L g141 ( .A(n_77), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_78), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_79), .B(n_204), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_80), .A2(n_94), .B1(n_153), .B2(n_172), .Y(n_510) );
CKINVDCx5p33_ASAP7_75t_R g554 ( .A(n_81), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_82), .B(n_157), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_83), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_86), .B(n_204), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_88), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_89), .B(n_204), .Y(n_223) );
INVx1_ASAP7_75t_L g108 ( .A(n_90), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g801 ( .A(n_90), .B(n_802), .Y(n_801) );
NAND2xp33_ASAP7_75t_L g581 ( .A(n_91), .B(n_144), .Y(n_581) );
A2O1A1Ixp33_ASAP7_75t_L g187 ( .A1(n_92), .A2(n_153), .B(n_174), .C(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g197 ( .A(n_93), .B(n_198), .Y(n_197) );
NAND2xp33_ASAP7_75t_L g231 ( .A(n_97), .B(n_193), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g797 ( .A(n_98), .Y(n_797) );
CKINVDCx11_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
OR2x6_ASAP7_75t_L g101 ( .A(n_102), .B(n_111), .Y(n_101) );
OR2x6_ASAP7_75t_L g825 ( .A(n_102), .B(n_111), .Y(n_825) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
NOR2x1p5_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
AND3x2_ASAP7_75t_L g816 ( .A(n_104), .B(n_107), .C(n_126), .Y(n_816) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g802 ( .A(n_105), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
BUFx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g489 ( .A(n_108), .Y(n_489) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NOR2x1p5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OR2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_803), .Y(n_116) );
OAI21xp33_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_128), .B(n_795), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
BUFx12f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x6_ASAP7_75t_SL g120 ( .A(n_121), .B(n_123), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx3_ASAP7_75t_L g806 ( .A(n_122), .Y(n_806) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_122), .B(n_822), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_126), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
NOR2x1_ASAP7_75t_L g824 ( .A(n_125), .B(n_127), .Y(n_824) );
AND2x6_ASAP7_75t_SL g800 ( .A(n_126), .B(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g794 ( .A(n_129), .Y(n_794) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OAI22x1_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_487), .B1(n_490), .B2(n_792), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_397), .Y(n_131) );
NOR3xp33_ASAP7_75t_L g132 ( .A(n_133), .B(n_326), .C(n_368), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_300), .Y(n_133) );
AOI22xp33_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_199), .B1(n_275), .B2(n_286), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OR2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_180), .Y(n_136) );
AOI21xp33_ASAP7_75t_L g319 ( .A1(n_137), .A2(n_320), .B(n_322), .Y(n_319) );
AOI21xp33_ASAP7_75t_L g392 ( .A1(n_137), .A2(n_393), .B(n_394), .Y(n_392) );
OR2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_164), .Y(n_137) );
INVx2_ASAP7_75t_L g312 ( .A(n_138), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_138), .B(n_165), .Y(n_342) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_142), .B(n_148), .C(n_160), .Y(n_139) );
INVx6_ASAP7_75t_L g170 ( .A(n_140), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_140), .A2(n_231), .B(n_232), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_140), .B(n_142), .Y(n_284) );
O2A1O1Ixp5_ASAP7_75t_L g576 ( .A1(n_140), .A2(n_169), .B(n_577), .C(n_578), .Y(n_576) );
BUFx8_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g151 ( .A(n_141), .Y(n_151) );
INVx1_ASAP7_75t_L g174 ( .A(n_141), .Y(n_174) );
INVx1_ASAP7_75t_L g211 ( .A(n_141), .Y(n_211) );
INVxp67_ASAP7_75t_SL g143 ( .A(n_144), .Y(n_143) );
INVx3_ASAP7_75t_L g517 ( .A(n_144), .Y(n_517) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g147 ( .A(n_145), .Y(n_147) );
INVx1_ASAP7_75t_L g153 ( .A(n_145), .Y(n_153) );
INVx1_ASAP7_75t_L g155 ( .A(n_145), .Y(n_155) );
INVx3_ASAP7_75t_L g168 ( .A(n_145), .Y(n_168) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_145), .Y(n_172) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_145), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_145), .Y(n_194) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_145), .Y(n_216) );
INVx1_ASAP7_75t_L g244 ( .A(n_145), .Y(n_244) );
INVx2_ASAP7_75t_L g250 ( .A(n_145), .Y(n_250) );
OAI21xp33_ASAP7_75t_SL g207 ( .A1(n_146), .A2(n_208), .B(n_209), .Y(n_207) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g283 ( .A(n_148), .Y(n_283) );
OAI21x1_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_152), .B(n_156), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_149), .A2(n_214), .B(n_215), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g254 ( .A1(n_149), .A2(n_170), .B1(n_255), .B2(n_256), .Y(n_254) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g500 ( .A(n_150), .Y(n_500) );
BUFx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g229 ( .A(n_151), .Y(n_229) );
INVx1_ASAP7_75t_L g562 ( .A(n_154), .Y(n_562) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_155), .B(n_189), .Y(n_188) );
OAI21xp33_ASAP7_75t_L g160 ( .A1(n_156), .A2(n_157), .B(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g175 ( .A(n_157), .Y(n_175) );
INVx2_ASAP7_75t_L g179 ( .A(n_157), .Y(n_179) );
INVx2_ASAP7_75t_L g185 ( .A(n_157), .Y(n_185) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_158), .Y(n_205) );
INVx1_ASAP7_75t_L g285 ( .A(n_160), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_161), .A2(n_240), .B(n_247), .Y(n_239) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
BUFx10_ASAP7_75t_L g176 ( .A(n_162), .Y(n_176) );
BUFx10_ASAP7_75t_L g218 ( .A(n_162), .Y(n_218) );
INVx1_ASAP7_75t_L g270 ( .A(n_162), .Y(n_270) );
AND2x2_ASAP7_75t_L g382 ( .A(n_164), .B(n_221), .Y(n_382) );
INVx1_ASAP7_75t_L g415 ( .A(n_164), .Y(n_415) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g277 ( .A(n_165), .B(n_222), .Y(n_277) );
AND2x2_ASAP7_75t_L g308 ( .A(n_165), .B(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g317 ( .A(n_165), .Y(n_317) );
OR2x2_ASAP7_75t_L g336 ( .A(n_165), .B(n_182), .Y(n_336) );
AND2x2_ASAP7_75t_L g351 ( .A(n_165), .B(n_182), .Y(n_351) );
AO31x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_175), .A3(n_176), .B(n_177), .Y(n_165) );
OAI22x1_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_170), .B1(n_171), .B2(n_173), .Y(n_166) );
INVx4_ASAP7_75t_L g169 ( .A(n_168), .Y(n_169) );
INVx1_ASAP7_75t_L g518 ( .A(n_168), .Y(n_518) );
INVx1_ASAP7_75t_L g534 ( .A(n_168), .Y(n_534) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_169), .A2(n_226), .B(n_227), .C(n_228), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g263 ( .A1(n_170), .A2(n_173), .B1(n_264), .B2(n_266), .Y(n_263) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_170), .A2(n_499), .B1(n_500), .B2(n_501), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_170), .A2(n_173), .B1(n_508), .B2(n_510), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_170), .A2(n_516), .B1(n_519), .B2(n_520), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_170), .A2(n_500), .B1(n_532), .B2(n_533), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_170), .A2(n_500), .B1(n_541), .B2(n_543), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_170), .A2(n_500), .B1(n_551), .B2(n_552), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_170), .A2(n_520), .B1(n_561), .B2(n_563), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_170), .A2(n_580), .B(n_581), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_172), .B(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g267 ( .A(n_172), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_173), .B(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_SL g520 ( .A(n_174), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_175), .B(n_536), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_175), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g196 ( .A(n_176), .Y(n_196) );
AO31x2_ASAP7_75t_L g497 ( .A1(n_176), .A2(n_257), .A3(n_498), .B(n_502), .Y(n_497) );
AO31x2_ASAP7_75t_L g539 ( .A1(n_176), .A2(n_506), .A3(n_540), .B(n_545), .Y(n_539) );
AO31x2_ASAP7_75t_L g559 ( .A1(n_176), .A2(n_238), .A3(n_560), .B(n_564), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
INVx2_ASAP7_75t_L g198 ( .A(n_179), .Y(n_198) );
BUFx2_ASAP7_75t_L g238 ( .A(n_179), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_179), .B(n_259), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_179), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_181), .B(n_350), .Y(n_393) );
OR2x2_ASAP7_75t_L g481 ( .A(n_181), .B(n_342), .Y(n_481) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g309 ( .A(n_182), .Y(n_309) );
AND2x2_ASAP7_75t_L g318 ( .A(n_182), .B(n_281), .Y(n_318) );
AND2x2_ASAP7_75t_L g321 ( .A(n_182), .B(n_222), .Y(n_321) );
AND2x2_ASAP7_75t_L g340 ( .A(n_182), .B(n_221), .Y(n_340) );
AND2x4_ASAP7_75t_L g359 ( .A(n_182), .B(n_282), .Y(n_359) );
AO21x2_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_186), .B(n_197), .Y(n_182) );
AO31x2_ASAP7_75t_L g530 ( .A1(n_183), .A2(n_521), .A3(n_531), .B(n_535), .Y(n_530) );
AO31x2_ASAP7_75t_L g549 ( .A1(n_183), .A2(n_269), .A3(n_550), .B(n_553), .Y(n_549) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_185), .B(n_512), .Y(n_511) );
NOR2xp33_ASAP7_75t_SL g564 ( .A(n_185), .B(n_565), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_190), .B(n_196), .Y(n_186) );
OAI22xp33_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B1(n_194), .B2(n_195), .Y(n_191) );
INVx2_ASAP7_75t_L g265 ( .A(n_193), .Y(n_265) );
INVx1_ASAP7_75t_L g542 ( .A(n_193), .Y(n_542) );
INVx1_ASAP7_75t_L g544 ( .A(n_194), .Y(n_544) );
INVx1_ASAP7_75t_L g521 ( .A(n_196), .Y(n_521) );
OAI21xp33_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_219), .B(n_260), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_200), .B(n_354), .Y(n_457) );
CKINVDCx14_ASAP7_75t_R g200 ( .A(n_201), .Y(n_200) );
BUFx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_202), .B(n_274), .Y(n_273) );
INVx3_ASAP7_75t_L g290 ( .A(n_202), .Y(n_290) );
OR2x2_ASAP7_75t_L g298 ( .A(n_202), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_202), .B(n_291), .Y(n_323) );
AND2x2_ASAP7_75t_L g348 ( .A(n_202), .B(n_262), .Y(n_348) );
AND2x2_ASAP7_75t_L g366 ( .A(n_202), .B(n_296), .Y(n_366) );
INVx1_ASAP7_75t_L g405 ( .A(n_202), .Y(n_405) );
AND2x2_ASAP7_75t_L g407 ( .A(n_202), .B(n_408), .Y(n_407) );
NAND2x1p5_ASAP7_75t_SL g426 ( .A(n_202), .B(n_347), .Y(n_426) );
AND2x4_ASAP7_75t_L g202 ( .A(n_203), .B(n_206), .Y(n_202) );
NOR2x1_ASAP7_75t_L g233 ( .A(n_204), .B(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g257 ( .A(n_204), .Y(n_257) );
INVx4_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g217 ( .A(n_205), .B(n_218), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_205), .B(n_503), .Y(n_502) );
BUFx3_ASAP7_75t_L g506 ( .A(n_205), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_205), .B(n_523), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_205), .B(n_546), .Y(n_545) );
INVx2_ASAP7_75t_SL g574 ( .A(n_205), .Y(n_574) );
OAI21xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_213), .B(n_217), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
BUFx4f_ASAP7_75t_L g246 ( .A(n_211), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_216), .B(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g234 ( .A(n_218), .Y(n_234) );
AO31x2_ASAP7_75t_L g253 ( .A1(n_218), .A2(n_254), .A3(n_257), .B(n_258), .Y(n_253) );
OAI32xp33_ASAP7_75t_L g310 ( .A1(n_219), .A2(n_302), .A3(n_311), .B1(n_313), .B2(n_315), .Y(n_310) );
OR2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_235), .Y(n_219) );
INVx1_ASAP7_75t_L g350 ( .A(n_220), .Y(n_350) );
AND2x2_ASAP7_75t_L g358 ( .A(n_220), .B(n_359), .Y(n_358) );
BUFx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g357 ( .A(n_221), .B(n_281), .Y(n_357) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
BUFx3_ASAP7_75t_L g307 ( .A(n_222), .Y(n_307) );
AND2x2_ASAP7_75t_L g316 ( .A(n_222), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g422 ( .A(n_222), .Y(n_422) );
NAND2x1p5_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
OAI21x1_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_230), .B(n_233), .Y(n_224) );
INVx2_ASAP7_75t_SL g228 ( .A(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g292 ( .A(n_235), .Y(n_292) );
OR2x2_ASAP7_75t_L g302 ( .A(n_235), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g424 ( .A(n_235), .Y(n_424) );
OR2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_252), .Y(n_235) );
AND2x2_ASAP7_75t_L g325 ( .A(n_236), .B(n_253), .Y(n_325) );
INVx2_ASAP7_75t_L g347 ( .A(n_236), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_236), .B(n_262), .Y(n_367) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g274 ( .A(n_237), .Y(n_274) );
AOI21x1_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B(n_251), .Y(n_237) );
AO31x2_ASAP7_75t_L g262 ( .A1(n_238), .A2(n_263), .A3(n_269), .B(n_271), .Y(n_262) );
AO31x2_ASAP7_75t_L g514 ( .A1(n_238), .A2(n_515), .A3(n_521), .B(n_522), .Y(n_514) );
OAI21xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_243), .B(n_246), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
INVx2_ASAP7_75t_L g268 ( .A(n_244), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
INVx2_ASAP7_75t_SL g509 ( .A(n_250), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_252), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g356 ( .A(n_252), .Y(n_356) );
INVx2_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
BUFx2_ASAP7_75t_L g296 ( .A(n_253), .Y(n_296) );
OR2x2_ASAP7_75t_L g362 ( .A(n_253), .B(n_262), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_253), .B(n_262), .Y(n_395) );
INVx2_ASAP7_75t_L g343 ( .A(n_260), .Y(n_343) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_273), .Y(n_260) );
OR2x2_ASAP7_75t_L g330 ( .A(n_261), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g408 ( .A(n_261), .Y(n_408) );
INVx1_ASAP7_75t_L g291 ( .A(n_262), .Y(n_291) );
INVx1_ASAP7_75t_L g299 ( .A(n_262), .Y(n_299) );
INVx1_ASAP7_75t_L g314 ( .A(n_262), .Y(n_314) );
AO31x2_ASAP7_75t_L g505 ( .A1(n_269), .A2(n_506), .A3(n_507), .B(n_511), .Y(n_505) );
INVx2_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
INVx2_ASAP7_75t_SL g582 ( .A(n_270), .Y(n_582) );
OR2x2_ASAP7_75t_L g418 ( .A(n_273), .B(n_395), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_274), .B(n_290), .Y(n_331) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_274), .Y(n_333) );
OR2x2_ASAP7_75t_L g432 ( .A(n_274), .B(n_356), .Y(n_432) );
INVxp67_ASAP7_75t_L g456 ( .A(n_274), .Y(n_456) );
INVx2_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
NAND2x1_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_277), .B(n_318), .Y(n_385) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g334 ( .A(n_279), .B(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g447 ( .A(n_280), .Y(n_447) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g476 ( .A(n_281), .B(n_309), .Y(n_476) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g402 ( .A(n_282), .B(n_309), .Y(n_402) );
AOI21x1_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_284), .B(n_285), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_293), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_292), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_289), .B(n_325), .Y(n_439) );
AND2x4_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx2_ASAP7_75t_L g303 ( .A(n_290), .Y(n_303) );
AND2x2_ASAP7_75t_L g353 ( .A(n_290), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_290), .B(n_347), .Y(n_396) );
OR2x2_ASAP7_75t_L g468 ( .A(n_290), .B(n_355), .Y(n_468) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g388 ( .A(n_294), .B(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
INVx2_ASAP7_75t_L g379 ( .A(n_295), .Y(n_379) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g369 ( .A(n_298), .B(n_370), .Y(n_369) );
INVxp67_ASAP7_75t_SL g380 ( .A(n_298), .Y(n_380) );
OR2x2_ASAP7_75t_L g431 ( .A(n_298), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g486 ( .A(n_298), .Y(n_486) );
AOI211xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_304), .B(n_310), .C(n_319), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g375 ( .A(n_303), .B(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_303), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g448 ( .A(n_303), .B(n_325), .Y(n_448) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_306), .B(n_351), .Y(n_373) );
NAND2x1p5_ASAP7_75t_L g390 ( .A(n_306), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g458 ( .A(n_306), .B(n_459), .Y(n_458) );
INVx3_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx2_ASAP7_75t_L g401 ( .A(n_307), .Y(n_401) );
AND2x2_ASAP7_75t_L g429 ( .A(n_308), .B(n_357), .Y(n_429) );
INVx2_ASAP7_75t_L g452 ( .A(n_308), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_308), .B(n_350), .Y(n_484) );
AND2x4_ASAP7_75t_SL g438 ( .A(n_311), .B(n_316), .Y(n_438) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g391 ( .A(n_312), .B(n_317), .Y(n_391) );
OR2x2_ASAP7_75t_L g443 ( .A(n_312), .B(n_336), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_313), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_313), .B(n_325), .Y(n_479) );
BUFx3_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g427 ( .A(n_314), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
INVx1_ASAP7_75t_L g410 ( .A(n_316), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_316), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g460 ( .A(n_317), .Y(n_460) );
BUFx2_ASAP7_75t_L g328 ( .A(n_318), .Y(n_328) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g446 ( .A(n_321), .B(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g370 ( .A(n_325), .Y(n_370) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_325), .Y(n_387) );
NAND3xp33_ASAP7_75t_SL g326 ( .A(n_327), .B(n_337), .C(n_352), .Y(n_326) );
AOI22xp33_ASAP7_75t_SL g327 ( .A1(n_328), .A2(n_329), .B1(n_332), .B2(n_334), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AOI222xp33_ASAP7_75t_L g440 ( .A1(n_334), .A2(n_360), .B1(n_441), .B2(n_444), .C1(n_446), .C2(n_448), .Y(n_440) );
AND2x2_ASAP7_75t_L g472 ( .A(n_335), .B(n_421), .Y(n_472) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g420 ( .A(n_336), .B(n_421), .Y(n_420) );
AOI22xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_343), .B1(n_344), .B2(n_349), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx2_ASAP7_75t_SL g416 ( .A(n_340), .Y(n_416) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_348), .Y(n_344) );
AND2x2_ASAP7_75t_L g403 ( .A(n_345), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g361 ( .A(n_346), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g355 ( .A(n_347), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g470 ( .A(n_348), .Y(n_470) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_351), .B(n_447), .Y(n_466) );
INVx1_ASAP7_75t_L g483 ( .A(n_351), .Y(n_483) );
AOI222xp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_357), .B1(n_358), .B2(n_360), .C1(n_363), .C2(n_364), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_359), .Y(n_363) );
AND2x2_ASAP7_75t_L g381 ( .A(n_359), .B(n_382), .Y(n_381) );
INVx3_ASAP7_75t_L g412 ( .A(n_359), .Y(n_412) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g376 ( .A(n_362), .Y(n_376) );
OR2x2_ASAP7_75t_L g445 ( .A(n_362), .B(n_426), .Y(n_445) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
OAI211xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_371), .B(n_374), .C(n_383), .Y(n_368) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OAI21xp33_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_377), .B(n_381), .Y(n_374) );
AOI221xp5_ASAP7_75t_L g461 ( .A1(n_375), .A2(n_413), .B1(n_462), .B2(n_465), .C(n_467), .Y(n_461) );
AND2x4_ASAP7_75t_L g404 ( .A(n_376), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
INVx1_ASAP7_75t_L g435 ( .A(n_382), .Y(n_435) );
AOI211x1_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_386), .B(n_388), .C(n_392), .Y(n_383) );
INVxp67_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g453 ( .A(n_391), .Y(n_453) );
NAND3xp33_ASAP7_75t_L g441 ( .A(n_394), .B(n_442), .C(n_443), .Y(n_441) );
OR2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx1_ASAP7_75t_L g477 ( .A(n_395), .Y(n_477) );
NOR2x1_ASAP7_75t_L g397 ( .A(n_398), .B(n_449), .Y(n_397) );
NAND4xp25_ASAP7_75t_L g398 ( .A(n_399), .B(n_406), .C(n_428), .D(n_440), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_403), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
AND2x2_ASAP7_75t_L g459 ( .A(n_402), .B(n_460), .Y(n_459) );
AOI221x1_ASAP7_75t_L g428 ( .A1(n_404), .A2(n_429), .B1(n_430), .B2(n_433), .C(n_436), .Y(n_428) );
AND2x2_ASAP7_75t_L g454 ( .A(n_404), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g464 ( .A(n_405), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_409), .B1(n_413), .B2(n_417), .C(n_419), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_411), .B(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_416), .A2(n_420), .B1(n_423), .B2(n_425), .Y(n_419) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g436 ( .A1(n_420), .A2(n_437), .B(n_439), .Y(n_436) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g442 ( .A(n_422), .Y(n_442) );
OR2x2_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVxp67_ASAP7_75t_L g463 ( .A(n_432), .Y(n_463) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OAI22xp33_ASAP7_75t_L g482 ( .A1(n_445), .A2(n_483), .B1(n_484), .B2(n_485), .Y(n_482) );
NAND3xp33_ASAP7_75t_L g449 ( .A(n_450), .B(n_461), .C(n_473), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_454), .B1(n_457), .B2(n_458), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
INVxp67_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g469 ( .A(n_456), .B(n_470), .Y(n_469) );
NAND2x1_ASAP7_75t_L g485 ( .A(n_456), .B(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
INVx2_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B(n_471), .Y(n_467) );
INVx1_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
AOI221xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_477), .B1(n_478), .B2(n_480), .C(n_482), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx3_ASAP7_75t_R g480 ( .A(n_481), .Y(n_480) );
INVx4_ASAP7_75t_L g792 ( .A(n_487), .Y(n_792) );
BUFx12f_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
CKINVDCx5p33_ASAP7_75t_R g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g823 ( .A(n_489), .B(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g810 ( .A(n_490), .Y(n_810) );
NOR2x1p5_ASAP7_75t_L g490 ( .A(n_491), .B(n_702), .Y(n_490) );
NAND4xp75_ASAP7_75t_L g491 ( .A(n_492), .B(n_647), .C(n_667), .D(n_683), .Y(n_491) );
NOR2x1p5_ASAP7_75t_SL g492 ( .A(n_493), .B(n_617), .Y(n_492) );
NAND4xp75_ASAP7_75t_L g493 ( .A(n_494), .B(n_555), .C(n_594), .D(n_603), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_524), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_504), .Y(n_495) );
AND2x4_ASAP7_75t_L g727 ( .A(n_496), .B(n_654), .Y(n_727) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_497), .Y(n_570) );
INVx2_ASAP7_75t_L g588 ( .A(n_497), .Y(n_588) );
AND2x2_ASAP7_75t_L g611 ( .A(n_497), .B(n_573), .Y(n_611) );
OR2x2_ASAP7_75t_L g666 ( .A(n_497), .B(n_505), .Y(n_666) );
AND2x2_ASAP7_75t_L g584 ( .A(n_504), .B(n_585), .Y(n_584) );
AND2x4_ASAP7_75t_L g734 ( .A(n_504), .B(n_611), .Y(n_734) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_513), .Y(n_504) );
OR2x2_ASAP7_75t_L g571 ( .A(n_505), .B(n_572), .Y(n_571) );
BUFx2_ASAP7_75t_L g602 ( .A(n_505), .Y(n_602) );
AND2x2_ASAP7_75t_L g608 ( .A(n_505), .B(n_514), .Y(n_608) );
INVx1_ASAP7_75t_L g626 ( .A(n_505), .Y(n_626) );
INVx2_ASAP7_75t_L g655 ( .A(n_505), .Y(n_655) );
INVx3_ASAP7_75t_L g631 ( .A(n_513), .Y(n_631) );
INVx2_ASAP7_75t_L g636 ( .A(n_513), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_513), .B(n_587), .Y(n_641) );
AND2x2_ASAP7_75t_L g664 ( .A(n_513), .B(n_643), .Y(n_664) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_513), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_513), .B(n_719), .Y(n_718) );
INVx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
BUFx2_ASAP7_75t_L g653 ( .A(n_514), .Y(n_653) );
AND2x2_ASAP7_75t_L g701 ( .A(n_514), .B(n_655), .Y(n_701) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_537), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_526), .B(n_645), .Y(n_692) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
NAND2x1p5_ASAP7_75t_L g689 ( .A(n_527), .B(n_645), .Y(n_689) );
INVx1_ASAP7_75t_L g790 ( .A(n_527), .Y(n_790) );
INVx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g740 ( .A(n_528), .B(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g593 ( .A(n_529), .Y(n_593) );
OR2x2_ASAP7_75t_L g674 ( .A(n_529), .B(n_548), .Y(n_674) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g616 ( .A(n_530), .Y(n_616) );
AND2x4_ASAP7_75t_L g622 ( .A(n_530), .B(n_623), .Y(n_622) );
AOI32xp33_ASAP7_75t_L g760 ( .A1(n_537), .A2(n_663), .A3(n_761), .B1(n_763), .B2(n_764), .Y(n_760) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g709 ( .A(n_538), .B(n_710), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_547), .Y(n_538) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_539), .Y(n_557) );
OR2x2_ASAP7_75t_L g591 ( .A(n_539), .B(n_549), .Y(n_591) );
INVx1_ASAP7_75t_L g606 ( .A(n_539), .Y(n_606) );
AND2x2_ASAP7_75t_L g615 ( .A(n_539), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g621 ( .A(n_539), .Y(n_621) );
INVx2_ASAP7_75t_L g646 ( .A(n_539), .Y(n_646) );
AND2x2_ASAP7_75t_L g765 ( .A(n_539), .B(n_559), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_547), .B(n_598), .Y(n_685) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g558 ( .A(n_549), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g614 ( .A(n_549), .Y(n_614) );
INVx2_ASAP7_75t_L g623 ( .A(n_549), .Y(n_623) );
AND2x4_ASAP7_75t_L g645 ( .A(n_549), .B(n_646), .Y(n_645) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_549), .Y(n_737) );
AOI22x1_ASAP7_75t_SL g555 ( .A1(n_556), .A2(n_566), .B1(n_584), .B2(n_589), .Y(n_555) );
AND2x4_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
NAND4xp25_ASAP7_75t_L g714 ( .A(n_558), .B(n_715), .C(n_716), .D(n_717), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_558), .B(n_615), .Y(n_745) );
INVx4_ASAP7_75t_SL g598 ( .A(n_559), .Y(n_598) );
BUFx2_ASAP7_75t_L g661 ( .A(n_559), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_559), .B(n_606), .Y(n_724) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g686 ( .A(n_568), .B(n_635), .Y(n_686) );
NOR2x1_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x4_ASAP7_75t_L g609 ( .A(n_572), .B(n_587), .Y(n_609) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_573), .B(n_588), .Y(n_633) );
OAI21x1_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_575), .B(n_583), .Y(n_573) );
OAI21x1_ASAP7_75t_L g628 ( .A1(n_574), .A2(n_575), .B(n_583), .Y(n_628) );
OAI21x1_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_579), .B(n_582), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_585), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g651 ( .A(n_585), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g690 ( .A(n_586), .B(n_608), .Y(n_690) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g733 ( .A(n_588), .B(n_643), .Y(n_733) );
AOI221xp5_ASAP7_75t_L g705 ( .A1(n_589), .A2(n_706), .B1(n_708), .B2(n_711), .C(n_713), .Y(n_705) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx2_ASAP7_75t_L g599 ( .A(n_591), .Y(n_599) );
OR2x2_ASAP7_75t_L g699 ( .A(n_591), .B(n_638), .Y(n_699) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_600), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_595), .A2(n_721), .B1(n_725), .B2(n_728), .Y(n_720) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_599), .Y(n_595) );
AND2x4_ASAP7_75t_L g644 ( .A(n_596), .B(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g756 ( .A(n_596), .B(n_674), .Y(n_756) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x4_ASAP7_75t_L g604 ( .A(n_598), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g620 ( .A(n_598), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g679 ( .A(n_598), .B(n_616), .Y(n_679) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_598), .Y(n_696) );
INVx1_ASAP7_75t_L g710 ( .A(n_598), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_598), .B(n_623), .Y(n_753) );
AND2x4_ASAP7_75t_L g660 ( .A(n_599), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g658 ( .A(n_601), .Y(n_658) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_602), .B(n_643), .Y(n_642) );
NAND2x1_ASAP7_75t_L g762 ( .A(n_602), .B(n_664), .Y(n_762) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_607), .B1(n_610), .B2(n_612), .Y(n_603) );
AND2x2_ASAP7_75t_L g629 ( .A(n_604), .B(n_622), .Y(n_629) );
INVx1_ASAP7_75t_L g670 ( .A(n_604), .Y(n_670) );
AND2x2_ASAP7_75t_L g777 ( .A(n_604), .B(n_638), .Y(n_777) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AND2x4_ASAP7_75t_SL g607 ( .A(n_608), .B(n_609), .Y(n_607) );
AND2x2_ASAP7_75t_L g610 ( .A(n_608), .B(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g750 ( .A(n_608), .Y(n_750) );
AND2x2_ASAP7_75t_L g767 ( .A(n_608), .B(n_627), .Y(n_767) );
AND2x2_ASAP7_75t_L g783 ( .A(n_608), .B(n_733), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_609), .B(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g706 ( .A(n_609), .B(n_707), .Y(n_706) );
OAI22xp33_ASAP7_75t_L g713 ( .A1(n_609), .A2(n_699), .B1(n_714), .B2(n_718), .Y(n_713) );
INVx1_ASAP7_75t_L g669 ( .A(n_611), .Y(n_669) );
AND2x2_ASAP7_75t_L g700 ( .A(n_611), .B(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_611), .B(n_707), .Y(n_729) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g735 ( .A(n_615), .B(n_736), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_615), .A2(n_639), .B1(n_744), .B2(n_746), .Y(n_743) );
INVx3_ASAP7_75t_L g638 ( .A(n_616), .Y(n_638) );
AND2x2_ASAP7_75t_L g770 ( .A(n_616), .B(n_623), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_634), .Y(n_617) );
AOI32xp33_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_624), .A3(n_627), .B1(n_629), .B2(n_630), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_621), .Y(n_716) );
INVx1_ASAP7_75t_L g741 ( .A(n_621), .Y(n_741) );
INVx3_ASAP7_75t_L g697 ( .A(n_622), .Y(n_697) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI221xp5_ASAP7_75t_L g772 ( .A1(n_625), .A2(n_773), .B1(n_774), .B2(n_775), .C(n_776), .Y(n_772) );
BUFx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g749 ( .A(n_627), .B(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_L g785 ( .A(n_627), .B(n_746), .Y(n_785) );
BUFx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g643 ( .A(n_628), .Y(n_643) );
NAND2x1p5_ASAP7_75t_L g657 ( .A(n_630), .B(n_658), .Y(n_657) );
AO22x1_ASAP7_75t_L g687 ( .A1(n_630), .A2(n_688), .B1(n_690), .B2(n_691), .Y(n_687) );
NAND2x1p5_ASAP7_75t_L g791 ( .A(n_630), .B(n_658), .Y(n_791) );
AND2x4_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
INVx2_ASAP7_75t_L g707 ( .A(n_631), .Y(n_707) );
INVx1_ASAP7_75t_L g717 ( .A(n_631), .Y(n_717) );
AND2x2_ASAP7_75t_L g637 ( .A(n_632), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVxp67_ASAP7_75t_SL g719 ( .A(n_633), .Y(n_719) );
INVx1_ASAP7_75t_L g759 ( .A(n_633), .Y(n_759) );
A2O1A1Ixp33_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_637), .B(n_639), .C(n_644), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NOR2x1p5_ASAP7_75t_L g746 ( .A(n_636), .B(n_666), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_637), .B(n_696), .Y(n_773) );
AOI31xp33_ASAP7_75t_L g656 ( .A1(n_638), .A2(n_657), .A3(n_659), .B(n_662), .Y(n_656) );
INVx4_ASAP7_75t_L g715 ( .A(n_638), .Y(n_715) );
OR2x2_ASAP7_75t_L g752 ( .A(n_638), .B(n_753), .Y(n_752) );
INVx2_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
AND2x4_ASAP7_75t_L g654 ( .A(n_643), .B(n_655), .Y(n_654) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_645), .Y(n_650) );
AND2x2_ASAP7_75t_L g681 ( .A(n_645), .B(n_679), .Y(n_681) );
NOR2xp67_ASAP7_75t_L g647 ( .A(n_648), .B(n_656), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx1_ASAP7_75t_L g774 ( .A(n_651), .Y(n_774) );
INVx1_ASAP7_75t_L g682 ( .A(n_652), .Y(n_682) );
AND2x4_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx1_ASAP7_75t_L g712 ( .A(n_653), .Y(n_712) );
AND2x2_ASAP7_75t_L g711 ( .A(n_654), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
OAI322xp33_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_670), .A3(n_671), .B1(n_675), .B2(n_678), .C1(n_680), .C2(n_682), .Y(n_668) );
INVxp67_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AOI211x1_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_686), .B(n_687), .C(n_693), .Y(n_683) );
INVx1_ASAP7_75t_L g788 ( .A(n_684), .Y(n_788) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx2_ASAP7_75t_L g742 ( .A(n_686), .Y(n_742) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OA21x2_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_698), .B(n_700), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OR2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
INVx2_ASAP7_75t_L g763 ( .A(n_697), .Y(n_763) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NAND2xp33_ASAP7_75t_L g758 ( .A(n_701), .B(n_759), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_703), .B(n_771), .Y(n_702) );
NOR3xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_738), .C(n_754), .Y(n_703) );
NAND3xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_720), .C(n_730), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_707), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI21xp33_ASAP7_75t_L g766 ( .A1(n_711), .A2(n_767), .B(n_768), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_715), .B(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_715), .B(n_765), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_716), .B(n_790), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_717), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OAI21xp5_ASAP7_75t_L g776 ( .A1(n_727), .A2(n_777), .B(n_778), .Y(n_776) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
OAI21xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_734), .B(n_735), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
OAI211xp5_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_742), .B(n_743), .C(n_747), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_748), .B(n_751), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
AND2x2_ASAP7_75t_SL g757 ( .A(n_749), .B(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_753), .Y(n_775) );
OAI211xp5_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_757), .B(n_760), .C(n_766), .Y(n_754) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_765), .B(n_770), .Y(n_769) );
INVx2_ASAP7_75t_L g786 ( .A(n_765), .Y(n_786) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g782 ( .A(n_770), .Y(n_782) );
NOR3xp33_ASAP7_75t_L g771 ( .A(n_772), .B(n_780), .C(n_787), .Y(n_771) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
AOI21xp33_ASAP7_75t_SL g780 ( .A1(n_781), .A2(n_784), .B(n_786), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_782), .B(n_783), .Y(n_781) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
AOI21xp33_ASAP7_75t_R g787 ( .A1(n_788), .A2(n_789), .B(n_791), .Y(n_787) );
OAI21xp5_ASAP7_75t_L g807 ( .A1(n_795), .A2(n_808), .B(n_812), .Y(n_807) );
INVxp67_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g796 ( .A(n_797), .B(n_798), .Y(n_796) );
BUFx12f_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx4_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
AO21x1_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_807), .B(n_817), .Y(n_803) );
CKINVDCx11_ASAP7_75t_R g804 ( .A(n_805), .Y(n_804) );
BUFx6f_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx2_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx3_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx4_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_818), .B(n_819), .Y(n_817) );
INVx2_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
BUFx10_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
endmodule