module fake_netlist_1_9091_n_11 (n_1, n_2, n_0, n_11);
input n_1;
input n_2;
input n_0;
output n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
BUFx6f_ASAP7_75t_L g3 ( .A(n_0), .Y(n_3) );
OR2x6_ASAP7_75t_L g4 ( .A(n_1), .B(n_0), .Y(n_4) );
AOI21x1_ASAP7_75t_L g5 ( .A1(n_4), .A2(n_0), .B(n_1), .Y(n_5) );
OR2x2_ASAP7_75t_L g6 ( .A(n_3), .B(n_0), .Y(n_6) );
AND2x2_ASAP7_75t_L g7 ( .A(n_6), .B(n_4), .Y(n_7) );
OAI221xp5_ASAP7_75t_L g8 ( .A1(n_7), .A2(n_4), .B1(n_5), .B2(n_3), .C(n_1), .Y(n_8) );
NAND4xp25_ASAP7_75t_L g9 ( .A(n_8), .B(n_7), .C(n_2), .D(n_3), .Y(n_9) );
OAI22x1_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_2), .B1(n_3), .B2(n_5), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_10), .Y(n_11) );
endmodule