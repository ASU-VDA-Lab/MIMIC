module fake_jpeg_16880_n_201 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_201);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_27),
.B(n_29),
.Y(n_54)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_28),
.Y(n_41)
);

HAxp5_ASAP7_75t_SL g29 ( 
.A(n_15),
.B(n_0),
.CON(n_29),
.SN(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_35),
.A2(n_37),
.B1(n_14),
.B2(n_24),
.Y(n_39)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_25),
.B1(n_17),
.B2(n_20),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_38),
.A2(n_40),
.B1(n_49),
.B2(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_25),
.B1(n_14),
.B2(n_21),
.Y(n_40)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_31),
.A2(n_26),
.B1(n_19),
.B2(n_23),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_29),
.A2(n_26),
.B1(n_23),
.B2(n_21),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_33),
.A2(n_24),
.B1(n_22),
.B2(n_13),
.Y(n_53)
);

AND2x6_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_28),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_57),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_56),
.A2(n_69),
.B1(n_28),
.B2(n_48),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_52),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_61),
.Y(n_83)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_37),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_37),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_49),
.Y(n_75)
);

AOI21xp33_ASAP7_75t_L g74 ( 
.A1(n_70),
.A2(n_54),
.B(n_51),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_74),
.A2(n_32),
.B1(n_36),
.B2(n_46),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_75),
.B(n_81),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_54),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_58),
.A2(n_53),
.B1(n_43),
.B2(n_42),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_78),
.A2(n_45),
.B1(n_41),
.B2(n_66),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_58),
.B(n_50),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_35),
.Y(n_82)
);

MAJx2_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_53),
.C(n_34),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_62),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_53),
.B(n_35),
.C(n_30),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_85),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_41),
.B1(n_36),
.B2(n_48),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_67),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_90),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_74),
.B(n_84),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_27),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_61),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_91),
.B(n_92),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_75),
.B(n_27),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_81),
.B(n_30),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_101),
.Y(n_108)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_97),
.B1(n_63),
.B2(n_69),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_76),
.C(n_82),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_32),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_66),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_79),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_109),
.B(n_119),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

AO21x2_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_85),
.B(n_84),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_SL g137 ( 
.A1(n_111),
.A2(n_34),
.B(n_36),
.C(n_24),
.Y(n_137)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_87),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_79),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_115),
.B(n_117),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_100),
.A2(n_85),
.B1(n_78),
.B2(n_77),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_116),
.A2(n_88),
.B1(n_111),
.B2(n_118),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_89),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_34),
.C(n_79),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_99),
.C(n_96),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_88),
.A2(n_0),
.B(n_15),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_120),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_98),
.Y(n_121)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_134),
.C(n_106),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_124),
.B(n_120),
.Y(n_144)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_98),
.Y(n_126)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

BUFx12_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_127),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_93),
.B1(n_92),
.B2(n_94),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_114),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_136),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_111),
.A2(n_117),
.B1(n_109),
.B2(n_119),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_112),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_94),
.C(n_89),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_108),
.B(n_90),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_137),
.A2(n_71),
.B1(n_68),
.B2(n_60),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_111),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_143),
.C(n_151),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_142),
.A2(n_150),
.B(n_152),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_104),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_71),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_113),
.Y(n_147)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_131),
.B(n_126),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_148),
.B(n_149),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_112),
.Y(n_149)
);

FAx1_ASAP7_75t_SL g153 ( 
.A(n_143),
.B(n_128),
.CI(n_134),
.CON(n_153),
.SN(n_153)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_163),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_139),
.A2(n_130),
.B1(n_122),
.B2(n_125),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_157),
.A2(n_137),
.B1(n_0),
.B2(n_4),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_133),
.C(n_135),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_162),
.C(n_142),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_127),
.Y(n_161)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_132),
.C(n_137),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_127),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_165),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_36),
.Y(n_165)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_150),
.C(n_147),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_172),
.Y(n_177)
);

OAI21x1_ASAP7_75t_L g167 ( 
.A1(n_160),
.A2(n_150),
.B(n_145),
.Y(n_167)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_167),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_170),
.C(n_174),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_152),
.C(n_137),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_34),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_156),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_181),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_154),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_182),
.C(n_22),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_155),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_158),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_171),
.A2(n_162),
.B1(n_157),
.B2(n_158),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_183),
.A2(n_169),
.B1(n_170),
.B2(n_22),
.Y(n_185)
);

NOR2x1_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_166),
.Y(n_184)
);

OAI21x1_ASAP7_75t_L g190 ( 
.A1(n_184),
.A2(n_187),
.B(n_180),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_188),
.C(n_189),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_9),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_177),
.A2(n_8),
.B(n_3),
.Y(n_189)
);

AOI322xp5_ASAP7_75t_L g195 ( 
.A1(n_190),
.A2(n_187),
.A3(n_3),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_180),
.C(n_13),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_192),
.B(n_193),
.Y(n_194)
);

FAx1_ASAP7_75t_SL g193 ( 
.A(n_184),
.B(n_8),
.CI(n_3),
.CON(n_193),
.SN(n_193)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_12),
.C(n_0),
.Y(n_198)
);

AOI322xp5_ASAP7_75t_L g196 ( 
.A1(n_190),
.A2(n_5),
.A3(n_6),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_196),
.A2(n_9),
.B(n_10),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_198),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_194),
.B(n_191),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_12),
.Y(n_201)
);


endmodule