module fake_jpeg_30679_n_63 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_63);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_63;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_48;
wire n_35;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx6_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_24),
.B(n_27),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_28),
.B(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_9),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_30),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_25),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_32),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_47)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

AO21x1_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_27),
.B(n_26),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_39),
.B(n_2),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_31),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_22),
.C(n_23),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_23),
.C(n_1),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_48),
.C(n_4),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_20),
.B1(n_17),
.B2(n_16),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_45),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_0),
.Y(n_45)
);

AOI21x1_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_49),
.B(n_3),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_55),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_41),
.B(n_39),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_53),
.C(n_48),
.Y(n_56)
);

MAJx2_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_42),
.C(n_38),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_54),
.A2(n_50),
.B1(n_6),
.B2(n_7),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_56),
.B(n_57),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_37),
.C(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_59),
.B(n_5),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_58),
.C(n_35),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_SL g63 ( 
.A1(n_62),
.A2(n_60),
.B(n_8),
.Y(n_63)
);


endmodule