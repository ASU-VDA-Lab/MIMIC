module fake_jpeg_10351_n_64 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_64);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_64;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_4),
.B(n_3),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_5),
.B(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_20),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_9),
.B(n_0),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_0),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_19),
.C(n_16),
.Y(n_24)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_16),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_22),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_12),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_24),
.C(n_26),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_15),
.B(n_11),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_31),
.A2(n_32),
.B(n_35),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_25),
.A2(n_13),
.B1(n_18),
.B2(n_15),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_11),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_28),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_31),
.B(n_24),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_6),
.C(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_44),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_28),
.B1(n_25),
.B2(n_37),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_21),
.B1(n_28),
.B2(n_13),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_23),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_45),
.C(n_47),
.Y(n_54)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_52),
.A2(n_55),
.B1(n_10),
.B2(n_0),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_49),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_54),
.C(n_50),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_57),
.C(n_51),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_42),
.C(n_29),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_54),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_60),
.C(n_7),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_62),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_63),
.B(n_8),
.Y(n_64)
);


endmodule