module fake_netlist_6_4150_n_1449 (n_52, n_1, n_91, n_326, n_256, n_209, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_350, n_78, n_84, n_142, n_143, n_180, n_62, n_349, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_280, n_287, n_353, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_352, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_348, n_69, n_293, n_31, n_334, n_53, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_361, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1449);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_350;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_280;
input n_287;
input n_353;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_293;
input n_31;
input n_334;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1449;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1415;
wire n_1370;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1393;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_976;
wire n_1445;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_513;
wire n_645;
wire n_1381;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_1033;
wire n_462;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_595;
wire n_627;
wire n_524;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_527;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1372;
wire n_505;
wire n_1339;
wire n_537;
wire n_1427;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_1429;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_1037;
wire n_621;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1443;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_934;
wire n_482;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_1343;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_799;
wire n_1155;
wire n_787;
wire n_1416;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1373;
wire n_1292;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1177;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_191),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_342),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_50),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_184),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_53),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_359),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_221),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_289),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_111),
.Y(n_372)
);

BUFx8_ASAP7_75t_SL g373 ( 
.A(n_296),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_103),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_255),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_136),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_64),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_36),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_151),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_352),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_199),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_271),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_63),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_47),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_233),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_236),
.Y(n_386)
);

INVxp33_ASAP7_75t_L g387 ( 
.A(n_5),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_9),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g389 ( 
.A(n_281),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_253),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_155),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_272),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_78),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_38),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_363),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_128),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_274),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_354),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_339),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_261),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_206),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_282),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_147),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_104),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_57),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_154),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_247),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_49),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_10),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_160),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_263),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_63),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_300),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_360),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_268),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_56),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_222),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_81),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_138),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_55),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_93),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_139),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_57),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_91),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_237),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_0),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_343),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_218),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_50),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_348),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_99),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_198),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_149),
.Y(n_433)
);

BUFx10_ASAP7_75t_L g434 ( 
.A(n_170),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_26),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_106),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_140),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_89),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_186),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_326),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_66),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_318),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_141),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_162),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_252),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_43),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_179),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_183),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_153),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_262),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_46),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_69),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_137),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g454 ( 
.A(n_55),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_73),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_290),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_195),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_113),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_44),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_107),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_1),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_39),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_190),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_43),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_76),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_304),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_301),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_95),
.Y(n_468)
);

BUFx10_ASAP7_75t_L g469 ( 
.A(n_15),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_266),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_291),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_321),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_219),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_356),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_345),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_172),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_59),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_295),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_223),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_313),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_118),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_117),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_112),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_132),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_85),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_142),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_114),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_358),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_311),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_31),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_280),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_244),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_208),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g494 ( 
.A(n_319),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_6),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_88),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_10),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_240),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_350),
.Y(n_499)
);

BUFx8_ASAP7_75t_SL g500 ( 
.A(n_249),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_323),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_264),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_254),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_38),
.Y(n_504)
);

BUFx8_ASAP7_75t_SL g505 ( 
.A(n_307),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_26),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_4),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_346),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_109),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_53),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_41),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_90),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_334),
.Y(n_513)
);

CKINVDCx14_ASAP7_75t_R g514 ( 
.A(n_238),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_65),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_2),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_129),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_220),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_74),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_335),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_232),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_166),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_143),
.Y(n_523)
);

CKINVDCx14_ASAP7_75t_R g524 ( 
.A(n_212),
.Y(n_524)
);

CKINVDCx14_ASAP7_75t_R g525 ( 
.A(n_124),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_303),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_144),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_332),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_260),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_241),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_74),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_66),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_324),
.Y(n_533)
);

BUFx10_ASAP7_75t_L g534 ( 
.A(n_298),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_329),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_51),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_205),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_245),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_33),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_168),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_94),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_351),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_315),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_69),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_333),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_157),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_33),
.Y(n_547)
);

INVx1_ASAP7_75t_SL g548 ( 
.A(n_228),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_173),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_3),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_276),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_130),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_17),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_341),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_27),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_146),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_361),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_267),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_327),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_49),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_242),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_159),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_22),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_349),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_340),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_131),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_331),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_134),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_167),
.Y(n_569)
);

CKINVDCx16_ASAP7_75t_R g570 ( 
.A(n_52),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_52),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_308),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_455),
.Y(n_573)
);

BUFx12f_ASAP7_75t_L g574 ( 
.A(n_469),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_400),
.B(n_0),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_380),
.B(n_1),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_400),
.B(n_2),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_391),
.B(n_3),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_455),
.Y(n_579)
);

INVx5_ASAP7_75t_L g580 ( 
.A(n_427),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_427),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_465),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_391),
.B(n_4),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_383),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_391),
.B(n_5),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_395),
.B(n_6),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_476),
.B(n_7),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_395),
.B(n_7),
.Y(n_588)
);

BUFx8_ASAP7_75t_SL g589 ( 
.A(n_373),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_427),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_SL g591 ( 
.A(n_570),
.B(n_8),
.Y(n_591)
);

BUFx12f_ASAP7_75t_L g592 ( 
.A(n_469),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_522),
.B(n_8),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_394),
.Y(n_594)
);

BUFx12f_ASAP7_75t_L g595 ( 
.A(n_469),
.Y(n_595)
);

BUFx12f_ASAP7_75t_L g596 ( 
.A(n_434),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_405),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_387),
.B(n_9),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_490),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_427),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_387),
.B(n_11),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_499),
.B(n_11),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_499),
.B(n_538),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_426),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_551),
.Y(n_605)
);

INVx5_ASAP7_75t_L g606 ( 
.A(n_551),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_422),
.B(n_12),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_389),
.B(n_12),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_538),
.B(n_13),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_429),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_552),
.B(n_13),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_430),
.B(n_14),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_514),
.B(n_14),
.Y(n_613)
);

CKINVDCx6p67_ASAP7_75t_R g614 ( 
.A(n_434),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_377),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_368),
.Y(n_616)
);

CKINVDCx11_ASAP7_75t_R g617 ( 
.A(n_366),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_446),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_552),
.B(n_572),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_430),
.B(n_15),
.Y(n_620)
);

INVx5_ASAP7_75t_L g621 ( 
.A(n_551),
.Y(n_621)
);

INVx5_ASAP7_75t_L g622 ( 
.A(n_551),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_442),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_376),
.B(n_365),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_572),
.B(n_16),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_368),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_442),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_420),
.B(n_16),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_478),
.Y(n_629)
);

BUFx8_ASAP7_75t_SL g630 ( 
.A(n_373),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_524),
.B(n_17),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_477),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_382),
.B(n_18),
.Y(n_633)
);

NAND2x1p5_ASAP7_75t_L g634 ( 
.A(n_478),
.B(n_80),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_420),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_402),
.B(n_18),
.Y(n_636)
);

INVx5_ASAP7_75t_L g637 ( 
.A(n_434),
.Y(n_637)
);

AND2x6_ASAP7_75t_L g638 ( 
.A(n_517),
.B(n_82),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_495),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_364),
.Y(n_640)
);

INVx5_ASAP7_75t_L g641 ( 
.A(n_534),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_517),
.Y(n_642)
);

BUFx12f_ASAP7_75t_L g643 ( 
.A(n_534),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_547),
.B(n_19),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_369),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_504),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_542),
.B(n_367),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_450),
.B(n_494),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_547),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_542),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_534),
.Y(n_651)
);

BUFx8_ASAP7_75t_SL g652 ( 
.A(n_500),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_375),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_459),
.B(n_19),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_506),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_507),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_511),
.Y(n_657)
);

BUFx2_ASAP7_75t_L g658 ( 
.A(n_378),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_521),
.B(n_20),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_500),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_516),
.B(n_20),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_531),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_379),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_525),
.B(n_454),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_539),
.B(n_21),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_388),
.Y(n_666)
);

XNOR2x2_ASAP7_75t_L g667 ( 
.A(n_555),
.B(n_21),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_571),
.B(n_22),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_393),
.B(n_23),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_408),
.B(n_23),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_409),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_390),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_412),
.B(n_24),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_396),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_397),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_407),
.B(n_24),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_411),
.B(n_25),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_581),
.Y(n_678)
);

OAI22xp33_ASAP7_75t_SL g679 ( 
.A1(n_591),
.A2(n_423),
.B1(n_435),
.B2(n_416),
.Y(n_679)
);

NAND2xp33_ASAP7_75t_SL g680 ( 
.A(n_598),
.B(n_366),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_664),
.B(n_548),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_648),
.A2(n_613),
.B1(n_631),
.B2(n_608),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_637),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_589),
.Y(n_684)
);

OAI22xp33_ASAP7_75t_L g685 ( 
.A1(n_591),
.A2(n_451),
.B1(n_452),
.B2(n_441),
.Y(n_685)
);

NAND3x1_ASAP7_75t_L g686 ( 
.A(n_601),
.B(n_415),
.C(n_413),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_651),
.B(n_371),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_581),
.Y(n_688)
);

OAI22xp33_ASAP7_75t_R g689 ( 
.A1(n_601),
.A2(n_462),
.B1(n_497),
.B2(n_384),
.Y(n_689)
);

OAI22xp33_ASAP7_75t_L g690 ( 
.A1(n_651),
.A2(n_464),
.B1(n_510),
.B2(n_461),
.Y(n_690)
);

OAI22xp33_ASAP7_75t_L g691 ( 
.A1(n_575),
.A2(n_532),
.B1(n_536),
.B2(n_515),
.Y(n_691)
);

AO22x2_ASAP7_75t_L g692 ( 
.A1(n_612),
.A2(n_419),
.B1(n_436),
.B2(n_418),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_576),
.A2(n_401),
.B1(n_406),
.B2(n_370),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_627),
.Y(n_694)
);

OA22x2_ASAP7_75t_L g695 ( 
.A1(n_599),
.A2(n_550),
.B1(n_553),
.B2(n_544),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_593),
.A2(n_401),
.B1(n_406),
.B2(n_370),
.Y(n_696)
);

OAI22xp33_ASAP7_75t_SL g697 ( 
.A1(n_578),
.A2(n_563),
.B1(n_560),
.B2(n_448),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_671),
.B(n_372),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_640),
.B(n_440),
.Y(n_699)
);

OAI22xp33_ASAP7_75t_R g700 ( 
.A1(n_607),
.A2(n_462),
.B1(n_497),
.B2(n_384),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_581),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_627),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_590),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_590),
.Y(n_704)
);

OAI22xp33_ASAP7_75t_L g705 ( 
.A1(n_575),
.A2(n_519),
.B1(n_482),
.B2(n_492),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_582),
.B(n_25),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_624),
.A2(n_519),
.B1(n_482),
.B2(n_492),
.Y(n_707)
);

OAI22xp33_ASAP7_75t_R g708 ( 
.A1(n_624),
.A2(n_460),
.B1(n_463),
.B2(n_456),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_615),
.B(n_27),
.Y(n_709)
);

AND2x4_ASAP7_75t_L g710 ( 
.A(n_671),
.B(n_471),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_587),
.A2(n_520),
.B1(n_443),
.B2(n_381),
.Y(n_711)
);

OAI22xp33_ASAP7_75t_SL g712 ( 
.A1(n_578),
.A2(n_484),
.B1(n_489),
.B2(n_474),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_658),
.B(n_374),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_590),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_627),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_600),
.Y(n_716)
);

INVx1_ASAP7_75t_SL g717 ( 
.A(n_617),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_633),
.A2(n_520),
.B1(n_443),
.B2(n_386),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_629),
.Y(n_719)
);

OAI22xp33_ASAP7_75t_L g720 ( 
.A1(n_577),
.A2(n_523),
.B1(n_528),
.B2(n_512),
.Y(n_720)
);

AO22x2_ASAP7_75t_L g721 ( 
.A1(n_612),
.A2(n_537),
.B1(n_543),
.B2(n_535),
.Y(n_721)
);

OAI22xp33_ASAP7_75t_L g722 ( 
.A1(n_577),
.A2(n_562),
.B1(n_559),
.B2(n_392),
.Y(n_722)
);

BUFx6f_ASAP7_75t_SL g723 ( 
.A(n_660),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_666),
.B(n_385),
.Y(n_724)
);

OAI22xp33_ASAP7_75t_SL g725 ( 
.A1(n_583),
.A2(n_399),
.B1(n_403),
.B2(n_398),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_623),
.B(n_404),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_637),
.B(n_410),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_637),
.B(n_414),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_600),
.Y(n_729)
);

BUFx2_ASAP7_75t_L g730 ( 
.A(n_630),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_600),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_629),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_629),
.Y(n_733)
);

XNOR2xp5_ASAP7_75t_L g734 ( 
.A(n_667),
.B(n_28),
.Y(n_734)
);

AO22x2_ASAP7_75t_L g735 ( 
.A1(n_620),
.A2(n_585),
.B1(n_583),
.B2(n_676),
.Y(n_735)
);

INVx8_ASAP7_75t_L g736 ( 
.A(n_652),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_637),
.B(n_417),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_645),
.B(n_421),
.Y(n_738)
);

OAI22xp33_ASAP7_75t_L g739 ( 
.A1(n_585),
.A2(n_614),
.B1(n_654),
.B2(n_677),
.Y(n_739)
);

OAI22xp33_ASAP7_75t_L g740 ( 
.A1(n_654),
.A2(n_425),
.B1(n_428),
.B2(n_424),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_642),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_642),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_641),
.B(n_647),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_642),
.Y(n_744)
);

NAND3x1_ASAP7_75t_L g745 ( 
.A(n_633),
.B(n_28),
.C(n_29),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_641),
.B(n_647),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_641),
.B(n_431),
.Y(n_747)
);

OAI22xp33_ASAP7_75t_SL g748 ( 
.A1(n_634),
.A2(n_433),
.B1(n_437),
.B2(n_432),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_636),
.A2(n_439),
.B1(n_444),
.B2(n_438),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_641),
.B(n_445),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_636),
.A2(n_659),
.B1(n_670),
.B2(n_669),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_597),
.Y(n_752)
);

OAI22xp33_ASAP7_75t_L g753 ( 
.A1(n_677),
.A2(n_449),
.B1(n_453),
.B2(n_447),
.Y(n_753)
);

AND2x2_ASAP7_75t_SL g754 ( 
.A(n_659),
.B(n_505),
.Y(n_754)
);

OA22x2_ASAP7_75t_L g755 ( 
.A1(n_573),
.A2(n_458),
.B1(n_466),
.B2(n_457),
.Y(n_755)
);

AND2x2_ASAP7_75t_SL g756 ( 
.A(n_620),
.B(n_505),
.Y(n_756)
);

OAI22xp33_ASAP7_75t_L g757 ( 
.A1(n_586),
.A2(n_468),
.B1(n_470),
.B2(n_467),
.Y(n_757)
);

AO22x2_ASAP7_75t_L g758 ( 
.A1(n_676),
.A2(n_586),
.B1(n_602),
.B2(n_588),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_579),
.B(n_472),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_673),
.A2(n_475),
.B1(n_479),
.B2(n_473),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_588),
.A2(n_481),
.B1(n_483),
.B2(n_480),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_596),
.A2(n_486),
.B1(n_487),
.B2(n_485),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_650),
.Y(n_763)
);

OAI22xp33_ASAP7_75t_SL g764 ( 
.A1(n_634),
.A2(n_609),
.B1(n_611),
.B2(n_602),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_699),
.A2(n_619),
.B(n_603),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_678),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_681),
.B(n_650),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_707),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_678),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_701),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_701),
.Y(n_771)
);

INVxp67_ASAP7_75t_SL g772 ( 
.A(n_688),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_729),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_SL g774 ( 
.A(n_756),
.B(n_638),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_SL g775 ( 
.A(n_754),
.B(n_638),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_731),
.Y(n_776)
);

XOR2xp5_ASAP7_75t_L g777 ( 
.A(n_684),
.B(n_488),
.Y(n_777)
);

INVxp33_ASAP7_75t_L g778 ( 
.A(n_693),
.Y(n_778)
);

INVxp33_ASAP7_75t_L g779 ( 
.A(n_696),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_729),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_733),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_743),
.B(n_650),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_688),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_716),
.Y(n_784)
);

CKINVDCx20_ASAP7_75t_R g785 ( 
.A(n_680),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_706),
.B(n_649),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_716),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_SL g788 ( 
.A(n_705),
.B(n_638),
.Y(n_788)
);

XNOR2x1_ASAP7_75t_L g789 ( 
.A(n_734),
.B(n_661),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_759),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_742),
.Y(n_791)
);

INVxp33_ASAP7_75t_L g792 ( 
.A(n_718),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_703),
.Y(n_793)
);

INVxp33_ASAP7_75t_L g794 ( 
.A(n_711),
.Y(n_794)
);

OR2x2_ASAP7_75t_L g795 ( 
.A(n_709),
.B(n_649),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_764),
.B(n_609),
.Y(n_796)
);

XNOR2x2_ASAP7_75t_L g797 ( 
.A(n_689),
.B(n_611),
.Y(n_797)
);

XOR2xp5_ASAP7_75t_L g798 ( 
.A(n_730),
.B(n_491),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_704),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_714),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_731),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_694),
.Y(n_802)
);

INVx1_ASAP7_75t_SL g803 ( 
.A(n_713),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_702),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_715),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_719),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_732),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_741),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_717),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_744),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_763),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_726),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_731),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_682),
.B(n_603),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_752),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_752),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_710),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_751),
.B(n_685),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_710),
.Y(n_819)
);

INVx3_ASAP7_75t_L g820 ( 
.A(n_746),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_687),
.B(n_672),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_738),
.Y(n_822)
);

INVxp33_ASAP7_75t_L g823 ( 
.A(n_695),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_739),
.B(n_625),
.Y(n_824)
);

INVxp33_ASAP7_75t_SL g825 ( 
.A(n_762),
.Y(n_825)
);

INVxp33_ASAP7_75t_L g826 ( 
.A(n_755),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_698),
.B(n_643),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_735),
.A2(n_619),
.B(n_605),
.Y(n_828)
);

XNOR2x2_ASAP7_75t_L g829 ( 
.A(n_689),
.B(n_625),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_735),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_758),
.Y(n_831)
);

INVxp33_ASAP7_75t_L g832 ( 
.A(n_724),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_758),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_692),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_692),
.Y(n_835)
);

AND2x6_ASAP7_75t_L g836 ( 
.A(n_727),
.B(n_628),
.Y(n_836)
);

INVxp67_ASAP7_75t_SL g837 ( 
.A(n_745),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_721),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_721),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_686),
.A2(n_638),
.B(n_675),
.Y(n_840)
);

OAI21xp5_ASAP7_75t_L g841 ( 
.A1(n_760),
.A2(n_638),
.B(n_628),
.Y(n_841)
);

OR2x2_ASAP7_75t_L g842 ( 
.A(n_749),
.B(n_662),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_728),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_737),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_747),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_750),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_712),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_683),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_679),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_761),
.B(n_662),
.Y(n_850)
);

XOR2xp5_ASAP7_75t_L g851 ( 
.A(n_748),
.B(n_493),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_720),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_725),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_690),
.B(n_653),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_697),
.Y(n_855)
);

NOR2xp67_ASAP7_75t_L g856 ( 
.A(n_723),
.B(n_580),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_708),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_814),
.B(n_604),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_814),
.B(n_610),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_767),
.B(n_618),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_815),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_821),
.B(n_655),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_816),
.Y(n_863)
);

HB1xp67_ASAP7_75t_L g864 ( 
.A(n_849),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_820),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_844),
.B(n_656),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_765),
.B(n_757),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_776),
.Y(n_868)
);

AND2x4_ASAP7_75t_SL g869 ( 
.A(n_853),
.B(n_657),
.Y(n_869)
);

AND2x6_ASAP7_75t_L g870 ( 
.A(n_831),
.B(n_644),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_832),
.B(n_740),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_766),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_820),
.B(n_753),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_769),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_770),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_790),
.B(n_584),
.Y(n_876)
);

INVx1_ASAP7_75t_SL g877 ( 
.A(n_795),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_790),
.B(n_594),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_849),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_832),
.B(n_691),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_771),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_833),
.B(n_632),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_803),
.B(n_639),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_836),
.B(n_722),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_836),
.B(n_843),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_836),
.B(n_845),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_836),
.B(n_653),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_836),
.B(n_653),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_818),
.B(n_646),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_773),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_780),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_782),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_818),
.B(n_644),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_776),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_817),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_846),
.B(n_663),
.Y(n_896)
);

INVxp67_ASAP7_75t_SL g897 ( 
.A(n_772),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_772),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_799),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_793),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_824),
.B(n_661),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_819),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_800),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_830),
.B(n_665),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_841),
.B(n_663),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_781),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_796),
.B(n_663),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_791),
.Y(n_908)
);

INVx1_ASAP7_75t_SL g909 ( 
.A(n_786),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_801),
.Y(n_910)
);

BUFx2_ASAP7_75t_L g911 ( 
.A(n_837),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_801),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_813),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_824),
.B(n_850),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_847),
.B(n_665),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_796),
.B(n_674),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_834),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_813),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_783),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_812),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_R g921 ( 
.A(n_809),
.B(n_736),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_835),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_854),
.B(n_674),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_784),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_802),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_854),
.B(n_674),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_852),
.B(n_827),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_787),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_804),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_828),
.A2(n_668),
.B(n_498),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_768),
.B(n_826),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_788),
.B(n_496),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_805),
.Y(n_933)
);

INVxp67_ASAP7_75t_L g934 ( 
.A(n_789),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_806),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_792),
.B(n_574),
.Y(n_936)
);

BUFx4f_ASAP7_75t_L g937 ( 
.A(n_853),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_840),
.B(n_501),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_807),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_808),
.Y(n_940)
);

NOR2xp67_ASAP7_75t_SL g941 ( 
.A(n_853),
.B(n_580),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_855),
.B(n_502),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_768),
.B(n_826),
.Y(n_943)
);

INVxp67_ASAP7_75t_L g944 ( 
.A(n_842),
.Y(n_944)
);

BUFx5_ASAP7_75t_L g945 ( 
.A(n_838),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_792),
.B(n_668),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_774),
.B(n_503),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_853),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_810),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_811),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_775),
.B(n_508),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_839),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_794),
.B(n_616),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_948),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_893),
.B(n_857),
.Y(n_955)
);

BUFx4f_ASAP7_75t_L g956 ( 
.A(n_948),
.Y(n_956)
);

NAND2x1p5_ASAP7_75t_L g957 ( 
.A(n_948),
.B(n_856),
.Y(n_957)
);

INVx4_ASAP7_75t_L g958 ( 
.A(n_868),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_893),
.B(n_778),
.Y(n_959)
);

OR2x6_ASAP7_75t_L g960 ( 
.A(n_948),
.B(n_736),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_948),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_865),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_861),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_883),
.B(n_778),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_892),
.B(n_848),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_883),
.B(n_779),
.Y(n_966)
);

CKINVDCx11_ASAP7_75t_R g967 ( 
.A(n_877),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_901),
.B(n_779),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_861),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_865),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_946),
.B(n_794),
.Y(n_971)
);

OR2x2_ASAP7_75t_L g972 ( 
.A(n_909),
.B(n_797),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_892),
.B(n_837),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_863),
.Y(n_974)
);

CKINVDCx6p67_ASAP7_75t_R g975 ( 
.A(n_920),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_944),
.B(n_946),
.Y(n_976)
);

NAND2x1_ASAP7_75t_SL g977 ( 
.A(n_914),
.B(n_829),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_868),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_953),
.B(n_823),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_953),
.B(n_823),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_921),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_863),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_868),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_901),
.B(n_822),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_920),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_902),
.B(n_785),
.Y(n_986)
);

INVx4_ASAP7_75t_L g987 ( 
.A(n_868),
.Y(n_987)
);

OR2x6_ASAP7_75t_L g988 ( 
.A(n_911),
.B(n_592),
.Y(n_988)
);

AND2x2_ASAP7_75t_SL g989 ( 
.A(n_937),
.B(n_700),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_902),
.B(n_894),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_872),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_858),
.B(n_825),
.Y(n_992)
);

BUFx12f_ASAP7_75t_L g993 ( 
.A(n_931),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_858),
.B(n_851),
.Y(n_994)
);

CKINVDCx8_ASAP7_75t_R g995 ( 
.A(n_911),
.Y(n_995)
);

BUFx4_ASAP7_75t_SL g996 ( 
.A(n_894),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_872),
.Y(n_997)
);

NOR2xp67_ASAP7_75t_L g998 ( 
.A(n_923),
.B(n_83),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_865),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_859),
.B(n_509),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_912),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_868),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_859),
.B(n_513),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_952),
.Y(n_1004)
);

NAND2xp33_ASAP7_75t_L g1005 ( 
.A(n_945),
.B(n_518),
.Y(n_1005)
);

OR2x2_ASAP7_75t_L g1006 ( 
.A(n_934),
.B(n_777),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_889),
.B(n_798),
.Y(n_1007)
);

NAND2x1p5_ASAP7_75t_L g1008 ( 
.A(n_937),
.B(n_580),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_952),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_SL g1010 ( 
.A(n_937),
.B(n_723),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_931),
.Y(n_1011)
);

NAND2x1p5_ASAP7_75t_L g1012 ( 
.A(n_941),
.B(n_580),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_874),
.Y(n_1013)
);

INVx4_ASAP7_75t_L g1014 ( 
.A(n_952),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_889),
.B(n_595),
.Y(n_1015)
);

INVx1_ASAP7_75t_SL g1016 ( 
.A(n_914),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_952),
.Y(n_1017)
);

OR2x2_ASAP7_75t_L g1018 ( 
.A(n_943),
.B(n_616),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_874),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_895),
.B(n_626),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_943),
.B(n_626),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_875),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_890),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_895),
.B(n_635),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_880),
.B(n_526),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_876),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_993),
.Y(n_1027)
);

INVx5_ASAP7_75t_L g1028 ( 
.A(n_954),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_985),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_963),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_1025),
.B(n_915),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_1001),
.Y(n_1032)
);

INVxp33_ASAP7_75t_L g1033 ( 
.A(n_976),
.Y(n_1033)
);

INVx1_ASAP7_75t_SL g1034 ( 
.A(n_967),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_1025),
.B(n_915),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_1001),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_1013),
.Y(n_1037)
);

INVx4_ASAP7_75t_L g1038 ( 
.A(n_954),
.Y(n_1038)
);

OR2x2_ASAP7_75t_L g1039 ( 
.A(n_959),
.B(n_864),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_1014),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_968),
.B(n_1016),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_954),
.Y(n_1042)
);

INVx2_ASAP7_75t_R g1043 ( 
.A(n_969),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_974),
.Y(n_1044)
);

INVx5_ASAP7_75t_SL g1045 ( 
.A(n_960),
.Y(n_1045)
);

INVx6_ASAP7_75t_SL g1046 ( 
.A(n_960),
.Y(n_1046)
);

BUFx4_ASAP7_75t_SL g1047 ( 
.A(n_960),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_990),
.B(n_952),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_1019),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_982),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_1023),
.Y(n_1051)
);

CKINVDCx20_ASAP7_75t_R g1052 ( 
.A(n_981),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_989),
.A2(n_700),
.B1(n_708),
.B2(n_870),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_991),
.Y(n_1054)
);

NAND2x1p5_ASAP7_75t_L g1055 ( 
.A(n_956),
.B(n_941),
.Y(n_1055)
);

INVx1_ASAP7_75t_SL g1056 ( 
.A(n_996),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_997),
.Y(n_1057)
);

OR2x6_ASAP7_75t_L g1058 ( 
.A(n_1026),
.B(n_1014),
.Y(n_1058)
);

INVx2_ASAP7_75t_SL g1059 ( 
.A(n_1004),
.Y(n_1059)
);

BUFx12f_ASAP7_75t_L g1060 ( 
.A(n_988),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1022),
.Y(n_1061)
);

BUFx4f_ASAP7_75t_L g1062 ( 
.A(n_1004),
.Y(n_1062)
);

INVx1_ASAP7_75t_SL g1063 ( 
.A(n_996),
.Y(n_1063)
);

BUFx4f_ASAP7_75t_SL g1064 ( 
.A(n_975),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1011),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_979),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_999),
.Y(n_1067)
);

CKINVDCx16_ASAP7_75t_R g1068 ( 
.A(n_1010),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_980),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_973),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_956),
.Y(n_1071)
);

BUFx5_ASAP7_75t_L g1072 ( 
.A(n_990),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_999),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_973),
.Y(n_1074)
);

INVx2_ASAP7_75t_SL g1075 ( 
.A(n_1004),
.Y(n_1075)
);

INVx3_ASAP7_75t_L g1076 ( 
.A(n_1009),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_1009),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_962),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_SL g1079 ( 
.A(n_986),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_986),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_995),
.Y(n_1081)
);

CKINVDCx20_ASAP7_75t_R g1082 ( 
.A(n_1006),
.Y(n_1082)
);

INVx5_ASAP7_75t_L g1083 ( 
.A(n_1009),
.Y(n_1083)
);

INVx1_ASAP7_75t_SL g1084 ( 
.A(n_984),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_955),
.A2(n_870),
.B1(n_884),
.B2(n_867),
.Y(n_1085)
);

BUFx2_ASAP7_75t_SL g1086 ( 
.A(n_965),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_1029),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_SL g1088 ( 
.A1(n_1068),
.A2(n_1007),
.B1(n_994),
.B2(n_992),
.Y(n_1088)
);

INVx6_ASAP7_75t_L g1089 ( 
.A(n_1029),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1057),
.Y(n_1090)
);

BUFx3_ASAP7_75t_L g1091 ( 
.A(n_1064),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_1031),
.A2(n_992),
.B1(n_959),
.B2(n_968),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_1071),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_SL g1094 ( 
.A1(n_1079),
.A2(n_936),
.B1(n_1010),
.B2(n_966),
.Y(n_1094)
);

INVx1_ASAP7_75t_SL g1095 ( 
.A(n_1081),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1057),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_SL g1097 ( 
.A1(n_1079),
.A2(n_964),
.B1(n_971),
.B2(n_984),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_1071),
.Y(n_1098)
);

INVx6_ASAP7_75t_L g1099 ( 
.A(n_1027),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_1071),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_1053),
.A2(n_871),
.B1(n_879),
.B2(n_976),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1030),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1044),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1050),
.Y(n_1104)
);

OAI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_1035),
.A2(n_972),
.B1(n_955),
.B2(n_1016),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_1065),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1054),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1037),
.Y(n_1108)
);

OAI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1033),
.A2(n_988),
.B1(n_1003),
.B2(n_1000),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1061),
.Y(n_1110)
);

CKINVDCx6p67_ASAP7_75t_R g1111 ( 
.A(n_1081),
.Y(n_1111)
);

INVx6_ASAP7_75t_L g1112 ( 
.A(n_1027),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1053),
.A2(n_927),
.B1(n_1015),
.B2(n_870),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_1071),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_SL g1115 ( 
.A1(n_1082),
.A2(n_988),
.B1(n_965),
.B2(n_922),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1084),
.A2(n_927),
.B1(n_870),
.B2(n_904),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1066),
.Y(n_1117)
);

OAI22xp33_ASAP7_75t_L g1118 ( 
.A1(n_1033),
.A2(n_1000),
.B1(n_1003),
.B2(n_1018),
.Y(n_1118)
);

OAI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_1039),
.A2(n_1021),
.B1(n_873),
.B2(n_942),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1069),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1041),
.B(n_876),
.Y(n_1121)
);

CKINVDCx20_ASAP7_75t_R g1122 ( 
.A(n_1052),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1037),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1070),
.A2(n_870),
.B1(n_904),
.B2(n_878),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1085),
.A2(n_1017),
.B1(n_897),
.B2(n_951),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1085),
.A2(n_1017),
.B1(n_926),
.B2(n_905),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1049),
.Y(n_1127)
);

BUFx12f_ASAP7_75t_L g1128 ( 
.A(n_1060),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1049),
.Y(n_1129)
);

CKINVDCx11_ASAP7_75t_R g1130 ( 
.A(n_1052),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_1042),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1082),
.A2(n_878),
.B1(n_862),
.B2(n_860),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1070),
.A2(n_870),
.B1(n_904),
.B2(n_932),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1048),
.A2(n_1017),
.B1(n_938),
.B2(n_961),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_1080),
.Y(n_1135)
);

OAI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1074),
.A2(n_935),
.B1(n_940),
.B2(n_925),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_L g1137 ( 
.A1(n_1074),
.A2(n_869),
.B1(n_1024),
.B2(n_1020),
.Y(n_1137)
);

BUFx4_ASAP7_75t_SL g1138 ( 
.A(n_1047),
.Y(n_1138)
);

BUFx8_ASAP7_75t_SL g1139 ( 
.A(n_1079),
.Y(n_1139)
);

BUFx10_ASAP7_75t_L g1140 ( 
.A(n_1048),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_1093),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_1135),
.B(n_977),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1097),
.A2(n_869),
.B1(n_935),
.B2(n_925),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1101),
.A2(n_1113),
.B1(n_1121),
.B2(n_1132),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1102),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_1088),
.A2(n_1055),
.B1(n_1045),
.B2(n_1062),
.Y(n_1146)
);

INVx3_ASAP7_75t_L g1147 ( 
.A(n_1140),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_1093),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1094),
.A2(n_1048),
.B1(n_1086),
.B2(n_1045),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1092),
.B(n_862),
.Y(n_1150)
);

OAI21xp33_ASAP7_75t_L g1151 ( 
.A1(n_1116),
.A2(n_860),
.B(n_930),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1109),
.A2(n_1034),
.B1(n_1060),
.B2(n_947),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1137),
.A2(n_1045),
.B1(n_1055),
.B2(n_1058),
.Y(n_1153)
);

AOI22xp33_ASAP7_75t_L g1154 ( 
.A1(n_1105),
.A2(n_950),
.B1(n_940),
.B2(n_885),
.Y(n_1154)
);

OAI222xp33_ASAP7_75t_L g1155 ( 
.A1(n_1124),
.A2(n_1118),
.B1(n_1117),
.B2(n_1120),
.C1(n_1119),
.C2(n_1133),
.Y(n_1155)
);

AOI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_1115),
.A2(n_950),
.B1(n_886),
.B2(n_866),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1106),
.B(n_1020),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_SL g1158 ( 
.A1(n_1128),
.A2(n_1063),
.B1(n_1056),
.B2(n_1072),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1103),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1104),
.A2(n_1062),
.B1(n_1046),
.B2(n_1058),
.Y(n_1160)
);

AOI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1122),
.A2(n_866),
.B1(n_1072),
.B2(n_1024),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_SL g1162 ( 
.A1(n_1095),
.A2(n_1072),
.B1(n_882),
.B2(n_1005),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1136),
.A2(n_882),
.B1(n_929),
.B2(n_949),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1107),
.A2(n_1110),
.B1(n_1058),
.B2(n_1111),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1096),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_1093),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1090),
.A2(n_1062),
.B1(n_1046),
.B2(n_1058),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1108),
.B(n_1072),
.Y(n_1168)
);

AOI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_1125),
.A2(n_929),
.B1(n_949),
.B2(n_939),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_1098),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1129),
.B(n_1072),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_1139),
.A2(n_949),
.B1(n_933),
.B2(n_939),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1129),
.B(n_1072),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1123),
.Y(n_1174)
);

NOR2x1_ASAP7_75t_L g1175 ( 
.A(n_1087),
.B(n_1038),
.Y(n_1175)
);

NAND3xp33_ASAP7_75t_L g1176 ( 
.A(n_1130),
.B(n_896),
.C(n_933),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1126),
.A2(n_916),
.B(n_907),
.Y(n_1177)
);

BUFx12f_ASAP7_75t_L g1178 ( 
.A(n_1089),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1127),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1134),
.A2(n_890),
.B1(n_1072),
.B2(n_881),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1098),
.A2(n_1046),
.B1(n_961),
.B2(n_1083),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1131),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1140),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_L g1184 ( 
.A1(n_1099),
.A2(n_881),
.B1(n_891),
.B2(n_875),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1131),
.Y(n_1185)
);

NOR3xp33_ASAP7_75t_L g1186 ( 
.A(n_1091),
.B(n_903),
.C(n_900),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1131),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1098),
.A2(n_1083),
.B1(n_1028),
.B2(n_898),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1099),
.A2(n_891),
.B1(n_1043),
.B2(n_924),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_1138),
.Y(n_1190)
);

AOI222xp33_ASAP7_75t_L g1191 ( 
.A1(n_1112),
.A2(n_635),
.B1(n_903),
.B2(n_900),
.C1(n_917),
.C2(n_1051),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1100),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1089),
.B(n_945),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1112),
.A2(n_1043),
.B1(n_924),
.B2(n_928),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1100),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1100),
.B(n_922),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1114),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1114),
.Y(n_1198)
);

OA21x2_ASAP7_75t_L g1199 ( 
.A1(n_1177),
.A2(n_888),
.B(n_887),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1144),
.A2(n_1152),
.B1(n_1146),
.B2(n_1142),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1144),
.A2(n_1146),
.B1(n_1150),
.B2(n_1151),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_SL g1202 ( 
.A1(n_1149),
.A2(n_1176),
.B1(n_1153),
.B2(n_1160),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1186),
.A2(n_1051),
.B1(n_998),
.B2(n_1078),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1157),
.B(n_1183),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1143),
.A2(n_998),
.B1(n_928),
.B2(n_919),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1156),
.A2(n_919),
.B1(n_908),
.B2(n_899),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1161),
.A2(n_908),
.B1(n_899),
.B2(n_906),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1191),
.B(n_1114),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1162),
.A2(n_906),
.B1(n_970),
.B2(n_1078),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1191),
.A2(n_1073),
.B1(n_1067),
.B2(n_1032),
.Y(n_1210)
);

AOI221xp5_ASAP7_75t_SL g1211 ( 
.A1(n_1164),
.A2(n_1042),
.B1(n_910),
.B2(n_1067),
.C(n_1073),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1174),
.B(n_1032),
.Y(n_1212)
);

OAI221xp5_ASAP7_75t_SL g1213 ( 
.A1(n_1172),
.A2(n_1036),
.B1(n_910),
.B2(n_1059),
.C(n_1075),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1158),
.A2(n_1036),
.B1(n_529),
.B2(n_530),
.Y(n_1214)
);

OAI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1160),
.A2(n_1040),
.B1(n_1083),
.B2(n_1075),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1154),
.A2(n_533),
.B1(n_540),
.B2(n_527),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1184),
.A2(n_957),
.B1(n_1040),
.B2(n_1008),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1163),
.A2(n_957),
.B1(n_1040),
.B2(n_1008),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1179),
.B(n_1076),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1189),
.A2(n_1083),
.B1(n_1059),
.B2(n_1077),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1194),
.A2(n_1077),
.B1(n_1076),
.B2(n_1028),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1169),
.A2(n_1077),
.B1(n_1076),
.B2(n_1028),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1180),
.A2(n_545),
.B1(n_546),
.B2(n_541),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1145),
.B(n_945),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_SL g1225 ( 
.A1(n_1167),
.A2(n_1188),
.B1(n_1155),
.B2(n_1181),
.Y(n_1225)
);

AOI222xp33_ASAP7_75t_L g1226 ( 
.A1(n_1159),
.A2(n_549),
.B1(n_554),
.B2(n_556),
.C1(n_557),
.C2(n_558),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1165),
.A2(n_1196),
.B1(n_1167),
.B2(n_1178),
.Y(n_1227)
);

AO22x1_ASAP7_75t_L g1228 ( 
.A1(n_1175),
.A2(n_564),
.B1(n_565),
.B2(n_561),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1192),
.B(n_1198),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_SL g1230 ( 
.A1(n_1188),
.A2(n_1028),
.B1(n_945),
.B2(n_567),
.Y(n_1230)
);

AOI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1181),
.A2(n_568),
.B1(n_569),
.B2(n_566),
.Y(n_1231)
);

NOR3xp33_ASAP7_75t_L g1232 ( 
.A(n_1193),
.B(n_1038),
.C(n_987),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1171),
.A2(n_945),
.B1(n_913),
.B2(n_918),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1173),
.A2(n_945),
.B1(n_913),
.B2(n_918),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1168),
.A2(n_945),
.B1(n_987),
.B2(n_958),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1147),
.A2(n_958),
.B1(n_983),
.B2(n_978),
.Y(n_1236)
);

NAND3xp33_ASAP7_75t_L g1237 ( 
.A(n_1182),
.B(n_1042),
.C(n_983),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1147),
.A2(n_1195),
.B1(n_1197),
.B2(n_1185),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1187),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1141),
.A2(n_983),
.B1(n_1002),
.B2(n_978),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1141),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_SL g1242 ( 
.A1(n_1141),
.A2(n_945),
.B1(n_1038),
.B2(n_1042),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1148),
.A2(n_1002),
.B1(n_978),
.B2(n_912),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_SL g1244 ( 
.A1(n_1148),
.A2(n_1012),
.B(n_1002),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1148),
.A2(n_912),
.B1(n_1012),
.B2(n_622),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_SL g1246 ( 
.A1(n_1166),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1166),
.A2(n_1170),
.B1(n_1190),
.B2(n_622),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1166),
.A2(n_1170),
.B1(n_622),
.B2(n_621),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_SL g1249 ( 
.A1(n_1170),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1144),
.A2(n_622),
.B1(n_621),
.B2(n_606),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1144),
.A2(n_621),
.B1(n_606),
.B2(n_605),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_SL g1252 ( 
.A1(n_1144),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1157),
.B(n_84),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1176),
.A2(n_621),
.B1(n_606),
.B2(n_605),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1200),
.B(n_35),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1201),
.B(n_36),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1202),
.B(n_605),
.Y(n_1257)
);

NAND3xp33_ASAP7_75t_L g1258 ( 
.A(n_1226),
.B(n_606),
.C(n_37),
.Y(n_1258)
);

NAND3xp33_ASAP7_75t_L g1259 ( 
.A(n_1252),
.B(n_37),
.C(n_39),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1201),
.B(n_40),
.Y(n_1260)
);

NAND3xp33_ASAP7_75t_L g1261 ( 
.A(n_1246),
.B(n_40),
.C(n_41),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1204),
.B(n_42),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1239),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1212),
.B(n_42),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1229),
.B(n_44),
.Y(n_1265)
);

NAND3xp33_ASAP7_75t_L g1266 ( 
.A(n_1249),
.B(n_1227),
.C(n_1216),
.Y(n_1266)
);

OAI221xp5_ASAP7_75t_SL g1267 ( 
.A1(n_1225),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.C(n_48),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1227),
.B(n_1238),
.Y(n_1268)
);

NAND3xp33_ASAP7_75t_L g1269 ( 
.A(n_1231),
.B(n_45),
.C(n_48),
.Y(n_1269)
);

OA21x2_ASAP7_75t_L g1270 ( 
.A1(n_1211),
.A2(n_51),
.B(n_54),
.Y(n_1270)
);

AND2x2_ASAP7_75t_SL g1271 ( 
.A(n_1232),
.B(n_54),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1219),
.B(n_56),
.Y(n_1272)
);

OAI21xp33_ASAP7_75t_SL g1273 ( 
.A1(n_1208),
.A2(n_58),
.B(n_59),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1213),
.B(n_58),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1253),
.B(n_60),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_SL g1276 ( 
.A1(n_1254),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_SL g1277 ( 
.A1(n_1214),
.A2(n_61),
.B(n_62),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1241),
.B(n_64),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1224),
.B(n_65),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1250),
.B(n_67),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1209),
.B(n_1203),
.Y(n_1281)
);

NAND3xp33_ASAP7_75t_L g1282 ( 
.A(n_1223),
.B(n_67),
.C(n_68),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1215),
.B(n_68),
.Y(n_1283)
);

AOI221xp5_ASAP7_75t_L g1284 ( 
.A1(n_1251),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.C(n_73),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1247),
.B(n_70),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1210),
.B(n_71),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1207),
.B(n_72),
.Y(n_1287)
);

OAI221xp5_ASAP7_75t_SL g1288 ( 
.A1(n_1205),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.C(n_78),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1206),
.A2(n_75),
.B1(n_77),
.B2(n_79),
.Y(n_1289)
);

OAI221xp5_ASAP7_75t_SL g1290 ( 
.A1(n_1203),
.A2(n_79),
.B1(n_86),
.B2(n_87),
.C(n_92),
.Y(n_1290)
);

AOI211xp5_ASAP7_75t_L g1291 ( 
.A1(n_1228),
.A2(n_96),
.B(n_97),
.C(n_98),
.Y(n_1291)
);

NAND3xp33_ASAP7_75t_L g1292 ( 
.A(n_1230),
.B(n_100),
.C(n_101),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1244),
.B(n_102),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1236),
.B(n_362),
.Y(n_1294)
);

NAND4xp25_ASAP7_75t_L g1295 ( 
.A(n_1237),
.B(n_105),
.C(n_108),
.D(n_110),
.Y(n_1295)
);

OAI21xp5_ASAP7_75t_SL g1296 ( 
.A1(n_1242),
.A2(n_1248),
.B(n_1220),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1235),
.B(n_1240),
.Y(n_1297)
);

AO21x2_ASAP7_75t_L g1298 ( 
.A1(n_1257),
.A2(n_1258),
.B(n_1256),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1263),
.B(n_1199),
.Y(n_1299)
);

NAND3xp33_ASAP7_75t_L g1300 ( 
.A(n_1269),
.B(n_1222),
.C(n_1221),
.Y(n_1300)
);

NOR3xp33_ASAP7_75t_L g1301 ( 
.A(n_1267),
.B(n_1217),
.C(n_1218),
.Y(n_1301)
);

NAND3xp33_ASAP7_75t_L g1302 ( 
.A(n_1291),
.B(n_1235),
.C(n_1199),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1270),
.Y(n_1303)
);

AO21x2_ASAP7_75t_L g1304 ( 
.A1(n_1260),
.A2(n_1199),
.B(n_1233),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1266),
.A2(n_1234),
.B1(n_1233),
.B2(n_1245),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1262),
.B(n_1234),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1297),
.B(n_1243),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1279),
.B(n_115),
.Y(n_1308)
);

AOI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1277),
.A2(n_116),
.B1(n_119),
.B2(n_120),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1268),
.B(n_1275),
.Y(n_1310)
);

NAND4xp75_ASAP7_75t_L g1311 ( 
.A(n_1271),
.B(n_121),
.C(n_122),
.D(n_123),
.Y(n_1311)
);

NAND3xp33_ASAP7_75t_L g1312 ( 
.A(n_1282),
.B(n_1255),
.C(n_1290),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1264),
.B(n_125),
.Y(n_1313)
);

OR2x2_ASAP7_75t_L g1314 ( 
.A(n_1265),
.B(n_126),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1271),
.B(n_127),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1270),
.B(n_133),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1272),
.B(n_135),
.Y(n_1317)
);

NOR3xp33_ASAP7_75t_SL g1318 ( 
.A(n_1273),
.B(n_357),
.C(n_148),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1278),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1281),
.B(n_145),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1283),
.B(n_150),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1286),
.Y(n_1322)
);

NAND4xp75_ASAP7_75t_L g1323 ( 
.A(n_1274),
.B(n_152),
.C(n_156),
.D(n_158),
.Y(n_1323)
);

OAI211xp5_ASAP7_75t_SL g1324 ( 
.A1(n_1285),
.A2(n_161),
.B(n_163),
.C(n_164),
.Y(n_1324)
);

INVxp67_ASAP7_75t_L g1325 ( 
.A(n_1319),
.Y(n_1325)
);

INVxp67_ASAP7_75t_SL g1326 ( 
.A(n_1299),
.Y(n_1326)
);

INVx1_ASAP7_75t_SL g1327 ( 
.A(n_1310),
.Y(n_1327)
);

BUFx2_ASAP7_75t_SL g1328 ( 
.A(n_1299),
.Y(n_1328)
);

NAND3xp33_ASAP7_75t_L g1329 ( 
.A(n_1312),
.B(n_1285),
.C(n_1261),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1303),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1310),
.B(n_1293),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1322),
.Y(n_1332)
);

XNOR2xp5_ASAP7_75t_L g1333 ( 
.A(n_1315),
.B(n_1311),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1304),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1304),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_SL g1336 ( 
.A1(n_1298),
.A2(n_1274),
.B1(n_1259),
.B2(n_1283),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1306),
.B(n_1296),
.Y(n_1337)
);

NAND4xp75_ASAP7_75t_SL g1338 ( 
.A(n_1316),
.B(n_1294),
.C(n_1288),
.D(n_1276),
.Y(n_1338)
);

XNOR2xp5_ASAP7_75t_L g1339 ( 
.A(n_1315),
.B(n_1289),
.Y(n_1339)
);

NAND4xp75_ASAP7_75t_SL g1340 ( 
.A(n_1316),
.B(n_1276),
.C(n_1295),
.D(n_1292),
.Y(n_1340)
);

INVx2_ASAP7_75t_SL g1341 ( 
.A(n_1306),
.Y(n_1341)
);

NAND4xp75_ASAP7_75t_SL g1342 ( 
.A(n_1320),
.B(n_1284),
.C(n_1289),
.D(n_1280),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1304),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1337),
.B(n_1314),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1330),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1330),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1332),
.Y(n_1347)
);

XOR2x2_ASAP7_75t_L g1348 ( 
.A(n_1333),
.B(n_1311),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1332),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1341),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1341),
.B(n_1298),
.Y(n_1351)
);

OA22x2_ASAP7_75t_L g1352 ( 
.A1(n_1333),
.A2(n_1309),
.B1(n_1321),
.B2(n_1320),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1325),
.Y(n_1353)
);

XOR2x2_ASAP7_75t_L g1354 ( 
.A(n_1339),
.B(n_1323),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1349),
.Y(n_1355)
);

AOI22xp5_ASAP7_75t_SL g1356 ( 
.A1(n_1352),
.A2(n_1339),
.B1(n_1331),
.B2(n_1328),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1349),
.Y(n_1357)
);

OA22x2_ASAP7_75t_L g1358 ( 
.A1(n_1353),
.A2(n_1327),
.B1(n_1328),
.B2(n_1331),
.Y(n_1358)
);

AOI22x1_ASAP7_75t_L g1359 ( 
.A1(n_1351),
.A2(n_1334),
.B1(n_1343),
.B2(n_1335),
.Y(n_1359)
);

AOI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1348),
.A2(n_1336),
.B1(n_1329),
.B2(n_1301),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1347),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1345),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1350),
.Y(n_1363)
);

OAI22xp33_ASAP7_75t_SL g1364 ( 
.A1(n_1354),
.A2(n_1326),
.B1(n_1314),
.B2(n_1343),
.Y(n_1364)
);

OA22x2_ASAP7_75t_L g1365 ( 
.A1(n_1346),
.A2(n_1321),
.B1(n_1338),
.B2(n_1342),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1345),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1344),
.B(n_1307),
.Y(n_1367)
);

AOI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1354),
.A2(n_1298),
.B1(n_1323),
.B2(n_1300),
.Y(n_1368)
);

AOI322xp5_ASAP7_75t_L g1369 ( 
.A1(n_1360),
.A2(n_1317),
.A3(n_1307),
.B1(n_1318),
.B2(n_1305),
.C1(n_1287),
.C2(n_1308),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1355),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1357),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1358),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1362),
.Y(n_1373)
);

OAI322xp33_ASAP7_75t_L g1374 ( 
.A1(n_1356),
.A2(n_1313),
.A3(n_1302),
.B1(n_1340),
.B2(n_1324),
.C1(n_175),
.C2(n_176),
.Y(n_1374)
);

AOI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1365),
.A2(n_165),
.B1(n_169),
.B2(n_171),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1361),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1366),
.Y(n_1377)
);

NAND4xp25_ASAP7_75t_L g1378 ( 
.A(n_1375),
.B(n_1368),
.C(n_1367),
.D(n_1364),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1370),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1373),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1371),
.Y(n_1381)
);

AOI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1375),
.A2(n_1368),
.B1(n_1363),
.B2(n_1359),
.Y(n_1382)
);

OAI322xp33_ASAP7_75t_L g1383 ( 
.A1(n_1372),
.A2(n_174),
.A3(n_177),
.B1(n_178),
.B2(n_180),
.C1(n_181),
.C2(n_182),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1377),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1380),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1379),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1381),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1382),
.A2(n_1376),
.B1(n_1374),
.B2(n_1369),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1384),
.Y(n_1389)
);

OAI221xp5_ASAP7_75t_L g1390 ( 
.A1(n_1378),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.C(n_189),
.Y(n_1390)
);

OAI22x1_ASAP7_75t_L g1391 ( 
.A1(n_1383),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1385),
.Y(n_1392)
);

AOI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1388),
.A2(n_196),
.B1(n_197),
.B2(n_200),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1386),
.Y(n_1394)
);

AOI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1390),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_1395)
);

INVxp67_ASAP7_75t_SL g1396 ( 
.A(n_1387),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_SL g1397 ( 
.A1(n_1389),
.A2(n_204),
.B1(n_207),
.B2(n_209),
.Y(n_1397)
);

AOI31xp33_ASAP7_75t_L g1398 ( 
.A1(n_1391),
.A2(n_210),
.A3(n_211),
.B(n_213),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1385),
.B(n_214),
.Y(n_1399)
);

AOI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1388),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_1400)
);

OAI211xp5_ASAP7_75t_L g1401 ( 
.A1(n_1393),
.A2(n_224),
.B(n_225),
.C(n_226),
.Y(n_1401)
);

AOI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1400),
.A2(n_1395),
.B1(n_1392),
.B2(n_1396),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1394),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_SL g1404 ( 
.A(n_1398),
.B(n_1399),
.Y(n_1404)
);

NOR2x1_ASAP7_75t_L g1405 ( 
.A(n_1397),
.B(n_227),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1400),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_1406)
);

AOI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1393),
.A2(n_234),
.B1(n_235),
.B2(n_239),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1392),
.B(n_243),
.Y(n_1408)
);

NOR3xp33_ASAP7_75t_L g1409 ( 
.A(n_1404),
.B(n_246),
.C(n_248),
.Y(n_1409)
);

AO22x2_ASAP7_75t_L g1410 ( 
.A1(n_1403),
.A2(n_250),
.B1(n_251),
.B2(n_256),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1408),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1402),
.Y(n_1412)
);

AO22x2_ASAP7_75t_SL g1413 ( 
.A1(n_1405),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1401),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1407),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1406),
.A2(n_265),
.B1(n_269),
.B2(n_270),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1410),
.Y(n_1417)
);

AOI21xp33_ASAP7_75t_L g1418 ( 
.A1(n_1412),
.A2(n_273),
.B(n_275),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1410),
.Y(n_1419)
);

OAI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1414),
.A2(n_355),
.B1(n_278),
.B2(n_279),
.Y(n_1420)
);

INVx3_ASAP7_75t_L g1421 ( 
.A(n_1411),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1413),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1415),
.Y(n_1423)
);

INVxp67_ASAP7_75t_SL g1424 ( 
.A(n_1409),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1417),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1422),
.A2(n_1416),
.B1(n_283),
.B2(n_284),
.Y(n_1426)
);

OAI22x1_ASAP7_75t_L g1427 ( 
.A1(n_1419),
.A2(n_277),
.B1(n_285),
.B2(n_286),
.Y(n_1427)
);

OA22x2_ASAP7_75t_L g1428 ( 
.A1(n_1423),
.A2(n_287),
.B1(n_288),
.B2(n_292),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1421),
.Y(n_1429)
);

AOI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1424),
.A2(n_293),
.B1(n_294),
.B2(n_297),
.Y(n_1430)
);

AO22x2_ASAP7_75t_L g1431 ( 
.A1(n_1421),
.A2(n_353),
.B1(n_302),
.B2(n_305),
.Y(n_1431)
);

AOI22x1_ASAP7_75t_SL g1432 ( 
.A1(n_1420),
.A2(n_299),
.B1(n_306),
.B2(n_309),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1429),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1425),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1428),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1427),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1431),
.Y(n_1437)
);

AOI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1436),
.A2(n_1426),
.B1(n_1432),
.B2(n_1430),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1435),
.A2(n_1418),
.B1(n_312),
.B2(n_314),
.Y(n_1439)
);

OAI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1437),
.A2(n_1418),
.B1(n_316),
.B2(n_317),
.Y(n_1440)
);

AOI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1433),
.A2(n_310),
.B1(n_320),
.B2(n_322),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1438),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1439),
.Y(n_1443)
);

AOI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1442),
.A2(n_1434),
.B1(n_1437),
.B2(n_1440),
.Y(n_1444)
);

AOI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1443),
.A2(n_1441),
.B1(n_328),
.B2(n_330),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1444),
.Y(n_1446)
);

INVx3_ASAP7_75t_L g1447 ( 
.A(n_1445),
.Y(n_1447)
);

AOI221xp5_ASAP7_75t_L g1448 ( 
.A1(n_1446),
.A2(n_325),
.B1(n_336),
.B2(n_337),
.C(n_338),
.Y(n_1448)
);

AOI211xp5_ASAP7_75t_L g1449 ( 
.A1(n_1448),
.A2(n_1447),
.B(n_344),
.C(n_347),
.Y(n_1449)
);


endmodule