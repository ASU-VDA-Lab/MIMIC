module fake_jpeg_6519_n_231 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_231);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_5),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_26),
.Y(n_34)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_27),
.A2(n_28),
.B1(n_31),
.B2(n_19),
.Y(n_44)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_33),
.Y(n_43)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx2_ASAP7_75t_SL g48 ( 
.A(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_15),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_28),
.A2(n_22),
.B1(n_13),
.B2(n_20),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_20),
.B1(n_13),
.B2(n_25),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_27),
.A2(n_24),
.B1(n_19),
.B2(n_22),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_27),
.B1(n_28),
.B2(n_31),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_46),
.B(n_49),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_60),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_42),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_27),
.B1(n_31),
.B2(n_28),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_52),
.B1(n_56),
.B2(n_61),
.Y(n_66)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_36),
.Y(n_63)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_37),
.Y(n_80)
);

OAI22x1_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_55),
.B1(n_50),
.B2(n_48),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_31),
.B1(n_24),
.B2(n_26),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_32),
.B1(n_29),
.B2(n_26),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_24),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_26),
.B1(n_32),
.B2(n_29),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_25),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_57),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_49),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_67),
.Y(n_81)
);

MAJx2_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_43),
.C(n_34),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_68),
.A2(n_47),
.B(n_51),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_75),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_55),
.B(n_50),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_34),
.Y(n_72)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_56),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_36),
.B1(n_35),
.B2(n_44),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_74),
.A2(n_79),
.B1(n_54),
.B2(n_50),
.Y(n_82)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_62),
.B(n_60),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_78),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_35),
.B1(n_45),
.B2(n_39),
.Y(n_79)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_76),
.B1(n_66),
.B2(n_68),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_70),
.B(n_67),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_88),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_92),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_70),
.B(n_72),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_47),
.B1(n_50),
.B2(n_35),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_90),
.B1(n_91),
.B2(n_74),
.Y(n_106)
);

AO21x2_ASAP7_75t_L g91 ( 
.A1(n_71),
.A2(n_48),
.B(n_53),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_97),
.A2(n_77),
.B(n_78),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_103),
.C(n_104),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_64),
.Y(n_100)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_101),
.B(n_112),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_102),
.A2(n_91),
.B1(n_90),
.B2(n_81),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_68),
.B(n_76),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_94),
.B(n_97),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_40),
.B1(n_33),
.B2(n_41),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_84),
.A2(n_76),
.B(n_79),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_109),
.C(n_95),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_91),
.A2(n_73),
.B1(n_75),
.B2(n_66),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_95),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_80),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_58),
.Y(n_110)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

NOR2x1_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_53),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_58),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_33),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_41),
.Y(n_129)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_113),
.Y(n_118)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_98),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_124),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_102),
.B(n_82),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_127),
.C(n_130),
.Y(n_134)
);

A2O1A1O1Ixp25_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_86),
.B(n_91),
.C(n_85),
.D(n_81),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_121),
.B(n_128),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_113),
.Y(n_125)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_93),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_98),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_129),
.A2(n_131),
.B(n_100),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_96),
.C(n_83),
.Y(n_130)
);

A2O1A1O1Ixp25_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_83),
.B(n_37),
.C(n_40),
.D(n_39),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_92),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_33),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_133),
.A2(n_114),
.B1(n_41),
.B2(n_93),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_99),
.C(n_109),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_141),
.C(n_147),
.Y(n_155)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_139),
.A2(n_143),
.B(n_144),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_107),
.C(n_106),
.Y(n_141)
);

OAI22x1_ASAP7_75t_L g142 ( 
.A1(n_121),
.A2(n_114),
.B1(n_108),
.B2(n_112),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_142),
.A2(n_41),
.B1(n_21),
.B2(n_15),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_129),
.A2(n_105),
.B(n_114),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_150),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_130),
.C(n_120),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_116),
.B(n_110),
.Y(n_149)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_15),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_151),
.A2(n_117),
.B(n_21),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_111),
.C(n_93),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_137),
.C(n_147),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_116),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_166),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_117),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_157),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_126),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_159),
.A2(n_21),
.B(n_23),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_111),
.C(n_33),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_161),
.C(n_167),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_125),
.B1(n_118),
.B2(n_111),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_162),
.A2(n_139),
.B1(n_170),
.B2(n_145),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_41),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_165),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_41),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_41),
.C(n_15),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_17),
.C(n_23),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_156),
.C(n_161),
.Y(n_178)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_171),
.B(n_172),
.Y(n_194)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_158),
.A2(n_142),
.B(n_140),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_173),
.A2(n_178),
.B(n_181),
.Y(n_187)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_167),
.A2(n_135),
.B1(n_148),
.B2(n_150),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_177),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_151),
.C(n_17),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_183),
.C(n_155),
.Y(n_186)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_168),
.B(n_9),
.Y(n_182)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_0),
.B(n_1),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_188),
.A2(n_175),
.B1(n_173),
.B2(n_8),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_177),
.B(n_180),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_190),
.B(n_5),
.Y(n_199)
);

AOI32xp33_ASAP7_75t_L g191 ( 
.A1(n_178),
.A2(n_9),
.A3(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_191),
.Y(n_204)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_176),
.Y(n_197)
);

MAJx2_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_21),
.C(n_23),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_195),
.C(n_196),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_17),
.C(n_23),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_17),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_197),
.A2(n_201),
.B(n_202),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_199),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_0),
.C(n_1),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_8),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_203),
.A2(n_205),
.B(n_206),
.Y(n_211)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_0),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_SL g207 ( 
.A(n_204),
.B(n_187),
.C(n_188),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_12),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_196),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_210),
.B(n_214),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_202),
.B(n_195),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_212),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_200),
.A2(n_193),
.B(n_9),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_213),
.A2(n_10),
.B(n_11),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_8),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_218),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_1),
.C(n_2),
.Y(n_217)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_211),
.B(n_10),
.Y(n_218)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_219),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_208),
.B(n_12),
.Y(n_221)
);

OAI211xp5_ASAP7_75t_L g225 ( 
.A1(n_221),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_225)
);

AOI21x1_ASAP7_75t_L g227 ( 
.A1(n_225),
.A2(n_217),
.B(n_3),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_220),
.C(n_215),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_226),
.A2(n_224),
.B(n_223),
.Y(n_228)
);

XNOR2x2_ASAP7_75t_SL g229 ( 
.A(n_227),
.B(n_3),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_228),
.A2(n_229),
.B(n_4),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_4),
.Y(n_231)
);


endmodule