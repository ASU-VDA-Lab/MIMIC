module fake_jpeg_1065_n_60 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_60);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_60;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_24),
.B(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_21),
.Y(n_25)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_22),
.Y(n_29)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_27),
.B(n_26),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_32),
.B(n_20),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_25),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_28),
.Y(n_40)
);

NAND3xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_35),
.C(n_37),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_25),
.B(n_20),
.Y(n_35)
);

AOI32xp33_ASAP7_75t_L g37 ( 
.A1(n_30),
.A2(n_23),
.A3(n_17),
.B1(n_16),
.B2(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_28),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_44),
.B(n_23),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_1),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_2),
.Y(n_52)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_49),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_43),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_52),
.Y(n_55)
);

A2O1A1O1Ixp25_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_12),
.B(n_14),
.C(n_5),
.D(n_6),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_46),
.C(n_4),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_54),
.A2(n_51),
.B(n_50),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_56),
.A2(n_55),
.B1(n_4),
.B2(n_5),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_57),
.B(n_7),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_58),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_3),
.Y(n_60)
);


endmodule