module real_jpeg_4164_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_534;
wire n_181;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_0),
.B(n_61),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_0),
.B(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_0),
.B(n_321),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_0),
.B(n_306),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_0),
.B(n_365),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_0),
.B(n_398),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_0),
.B(n_409),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_1),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_1),
.B(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_1),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_1),
.B(n_104),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_1),
.B(n_344),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_1),
.B(n_358),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_1),
.B(n_425),
.Y(n_424)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_2),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_2),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_2),
.Y(n_327)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_2),
.Y(n_334)
);

BUFx5_ASAP7_75t_L g361 ( 
.A(n_2),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_3),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_3),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_3),
.B(n_149),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_3),
.B(n_90),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_3),
.B(n_107),
.Y(n_222)
);

AND2x2_ASAP7_75t_SL g297 ( 
.A(n_3),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_3),
.B(n_327),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_3),
.B(n_430),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_4),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_4),
.B(n_198),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_4),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_4),
.B(n_61),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_4),
.B(n_303),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_4),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_4),
.B(n_283),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_4),
.B(n_422),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_5),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_5),
.Y(n_177)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_5),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_6),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_6),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_6),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_6),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_6),
.B(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g191 ( 
.A(n_6),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_6),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_6),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_7),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_7),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_7),
.B(n_68),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_7),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_7),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_7),
.B(n_283),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_7),
.B(n_306),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_7),
.B(n_272),
.Y(n_432)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_8),
.Y(n_87)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_8),
.Y(n_147)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_8),
.Y(n_238)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_9),
.Y(n_543)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_10),
.Y(n_116)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_10),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_10),
.Y(n_300)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_11),
.Y(n_71)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_12),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_12),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_12),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_13),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_13),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_13),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_13),
.B(n_326),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_13),
.B(n_342),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_13),
.B(n_114),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_13),
.B(n_392),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_13),
.B(n_419),
.Y(n_418)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_15),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_15),
.B(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_15),
.B(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_15),
.B(n_351),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_15),
.B(n_139),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_15),
.B(n_396),
.Y(n_395)
);

AND2x4_ASAP7_75t_SL g411 ( 
.A(n_15),
.B(n_412),
.Y(n_411)
);

INVxp33_ASAP7_75t_L g547 ( 
.A(n_16),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_40),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_17),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_17),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_17),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_17),
.B(n_170),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_17),
.B(n_207),
.Y(n_206)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_19),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_19),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_19),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_19),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_19),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_19),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_19),
.B(n_139),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_19),
.B(n_270),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_542),
.B(n_544),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_38),
.B(n_76),
.C(n_541),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_43),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_24),
.B(n_43),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.C(n_34),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_26),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_26),
.A2(n_30),
.B1(n_37),
.B2(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_30),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_30),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_30),
.B(n_47),
.C(n_54),
.Y(n_73)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_32),
.Y(n_396)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_33),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_33),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_34),
.B(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_72),
.C(n_74),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_44),
.B(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_58),
.C(n_62),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_45),
.B(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_54),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_47),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_47),
.A2(n_53),
.B1(n_67),
.B2(n_117),
.Y(n_121)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_49),
.Y(n_398)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_51),
.Y(n_139)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_51),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_51),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_63),
.C(n_67),
.Y(n_62)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_57),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_58),
.B(n_62),
.Y(n_124)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_63),
.A2(n_64),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_67),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_67),
.A2(n_110),
.B1(n_111),
.B2(n_117),
.Y(n_513)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_69),
.Y(n_227)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_70),
.Y(n_152)
);

INVx6_ASAP7_75t_L g367 ( 
.A(n_70),
.Y(n_367)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_71),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_71),
.Y(n_304)
);

BUFx5_ASAP7_75t_L g393 ( 
.A(n_71),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

AO21x1_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_128),
.B(n_540),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_125),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_78),
.B(n_125),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_122),
.C(n_123),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_79),
.A2(n_80),
.B1(n_536),
.B2(n_537),
.Y(n_535)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_105),
.C(n_118),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_81),
.A2(n_82),
.B1(n_517),
.B2(n_519),
.Y(n_516)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_92),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_88),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_88),
.C(n_92),
.Y(n_122)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_91),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g204 ( 
.A(n_91),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.C(n_100),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_93),
.B(n_508),
.Y(n_507)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_96),
.A2(n_97),
.B1(n_100),
.B2(n_101),
.Y(n_508)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_105),
.A2(n_118),
.B1(n_119),
.B2(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_105),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.C(n_117),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g512 ( 
.A(n_106),
.B(n_513),
.Y(n_512)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_110),
.A2(n_111),
.B1(n_206),
.B2(n_209),
.Y(n_205)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_111),
.B(n_203),
.C(n_206),
.Y(n_514)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_115),
.Y(n_330)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_116),
.Y(n_423)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g537 ( 
.A(n_122),
.B(n_123),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_534),
.B(n_539),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_501),
.B(n_531),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_309),
.B(n_500),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_255),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_132),
.B(n_255),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_200),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_133),
.B(n_201),
.C(n_230),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_172),
.C(n_182),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_134),
.B(n_258),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_143),
.C(n_156),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_135),
.B(n_486),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_138),
.C(n_140),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.Y(n_137)
);

INVx6_ASAP7_75t_L g287 ( 
.A(n_139),
.Y(n_287)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_143),
.A2(n_144),
.B1(n_156),
.B2(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.C(n_153),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_145),
.B(n_153),
.Y(n_476)
);

INVx6_ASAP7_75t_L g413 ( 
.A(n_146),
.Y(n_413)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_148),
.B(n_476),
.Y(n_475)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx5_ASAP7_75t_L g351 ( 
.A(n_152),
.Y(n_351)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_152),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_155),
.Y(n_214)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_156),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_161),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_157),
.Y(n_241)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_168),
.B2(n_169),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_163),
.B(n_168),
.C(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_166),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_167),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_168),
.A2(n_169),
.B1(n_206),
.B2(n_209),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_168),
.B(n_206),
.C(n_234),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_171),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_172),
.B(n_182),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_181),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_173)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_174),
.Y(n_179)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_178),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_178),
.A2(n_180),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_178),
.B(n_179),
.C(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_178),
.B(n_247),
.C(n_251),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_181),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_193),
.C(n_197),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_183),
.B(n_290),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.C(n_191),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_184),
.B(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_186),
.B(n_191),
.Y(n_267)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g342 ( 
.A(n_190),
.Y(n_342)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_190),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_193),
.B(n_197),
.Y(n_290)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

BUFx5_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_196),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_230),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_210),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_202),
.B(n_211),
.C(n_229),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_206),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_221),
.B1(n_228),
.B2(n_229),
.Y(n_210)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_211),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.C(n_218),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_218),
.Y(n_243)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_222),
.B(n_224),
.C(n_225),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_244),
.B2(n_245),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_231),
.B(n_246),
.C(n_253),
.Y(n_526)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_240),
.C(n_242),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_233),
.B(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_239),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_238),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_242),
.Y(n_261)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_253),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_251),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_259),
.C(n_262),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_257),
.B(n_260),
.Y(n_496)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_262),
.B(n_496),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_288),
.C(n_291),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_264),
.B(n_489),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_268),
.C(n_277),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_265),
.A2(n_266),
.B1(n_467),
.B2(n_468),
.Y(n_466)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_268),
.A2(n_269),
.B(n_273),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_268),
.B(n_277),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_273),
.Y(n_268)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

MAJx2_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_281),
.C(n_285),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_278),
.A2(n_279),
.B1(n_281),
.B2(n_282),
.Y(n_444)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx8_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_285),
.B(n_444),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_286),
.B(n_307),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_288),
.A2(n_289),
.B1(n_291),
.B2(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_291),
.Y(n_490)
);

MAJx2_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_305),
.C(n_308),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_293),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_293),
.B(n_478),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_297),
.C(n_301),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_294),
.B(n_456),
.Y(n_455)
);

INVx6_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_297),
.A2(n_301),
.B1(n_302),
.B2(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_297),
.Y(n_457)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_305),
.B(n_308),
.Y(n_478)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

AOI21x1_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_494),
.B(n_499),
.Y(n_309)
);

OAI21x1_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_481),
.B(n_493),
.Y(n_310)
);

AOI21x1_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_463),
.B(n_480),
.Y(n_311)
);

OAI21x1_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_437),
.B(n_462),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_402),
.B(n_436),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_373),
.B(n_401),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_353),
.B(n_372),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_336),
.B(n_352),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_331),
.B(n_335),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_328),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_319),
.B(n_328),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_325),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_332),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_320),
.B(n_325),
.Y(n_337)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx5_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_324),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_337),
.B(n_338),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_339),
.A2(n_340),
.B1(n_345),
.B2(n_346),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_339),
.B(n_348),
.C(n_349),
.Y(n_371)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_341),
.B(n_343),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_341),
.B(n_343),
.Y(n_362)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_347),
.A2(n_348),
.B1(n_349),
.B2(n_350),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_354),
.B(n_371),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_354),
.B(n_371),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_363),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_362),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_362),
.C(n_375),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_360),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_357),
.B(n_360),
.Y(n_378)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_363),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_368),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_364),
.B(n_388),
.C(n_389),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx8_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_369),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_370),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_376),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_374),
.B(n_376),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_386),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_377),
.B(n_387),
.C(n_390),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_378),
.B(n_380),
.C(n_381),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_382),
.A2(n_383),
.B1(n_384),
.B2(n_385),
.Y(n_381)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_382),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_383),
.B(n_385),
.Y(n_406)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_390),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_394),
.Y(n_390)
);

MAJx2_ASAP7_75t_L g434 ( 
.A(n_391),
.B(n_397),
.C(n_399),
.Y(n_434)
);

INVx5_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_395),
.A2(n_397),
.B1(n_399),
.B2(n_400),
.Y(n_394)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_395),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_397),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_403),
.B(n_435),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_403),
.B(n_435),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_404),
.B(n_415),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_414),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_405),
.B(n_414),
.C(n_461),
.Y(n_460)
);

XNOR2x1_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_406),
.B(n_451),
.C(n_452),
.Y(n_450)
);

XNOR2x1_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_411),
.Y(n_407)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_408),
.Y(n_451)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_411),
.Y(n_452)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_415),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_426),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_416),
.B(n_428),
.C(n_433),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_424),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_421),
.Y(n_417)
);

MAJx2_ASAP7_75t_L g448 ( 
.A(n_418),
.B(n_421),
.C(n_424),
.Y(n_448)
);

INVx6_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx4_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_428),
.B1(n_433),
.B2(n_434),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_432),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_429),
.B(n_432),
.Y(n_447)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_434),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_460),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_438),
.B(n_460),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_449),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_441),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_440),
.B(n_441),
.C(n_449),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_442),
.A2(n_443),
.B1(n_445),
.B2(n_446),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_442),
.B(n_472),
.C(n_473),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_447),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_448),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_450),
.B(n_453),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_450),
.B(n_454),
.C(n_459),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_454),
.A2(n_455),
.B1(n_458),
.B2(n_459),
.Y(n_453)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_454),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_455),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_464),
.B(n_479),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_464),
.B(n_479),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_465),
.B(n_470),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_469),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_466),
.B(n_469),
.C(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_467),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_470),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_471),
.B(n_474),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_471),
.B(n_475),
.C(n_477),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_477),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_482),
.B(n_491),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_482),
.B(n_491),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_484),
.Y(n_482)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_483),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_488),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_485),
.B(n_488),
.C(n_498),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_495),
.B(n_497),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_495),
.B(n_497),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_527),
.Y(n_501)
);

OAI21xp33_ASAP7_75t_L g531 ( 
.A1(n_502),
.A2(n_532),
.B(n_533),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_503),
.B(n_521),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_503),
.B(n_521),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_504),
.A2(n_505),
.B1(n_510),
.B2(n_520),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_504),
.B(n_511),
.C(n_516),
.Y(n_538)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_507),
.C(n_509),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_506),
.B(n_523),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_507),
.B(n_509),
.Y(n_523)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_510),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_516),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_514),
.C(n_515),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_512),
.B(n_525),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_514),
.B(n_515),
.Y(n_525)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_517),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_524),
.C(n_526),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_522),
.B(n_524),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_526),
.B(n_529),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_528),
.B(n_530),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_528),
.B(n_530),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_535),
.B(n_538),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_535),
.B(n_538),
.Y(n_539)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx6_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx13_ASAP7_75t_L g546 ( 
.A(n_543),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_545),
.B(n_547),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);


endmodule