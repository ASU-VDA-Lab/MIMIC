module real_jpeg_27166_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_0),
.A2(n_35),
.B1(n_36),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_0),
.A2(n_43),
.B1(n_50),
.B2(n_51),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_0),
.A2(n_43),
.B1(n_60),
.B2(n_61),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_0),
.A2(n_22),
.B1(n_27),
.B2(n_43),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_SL g111 ( 
.A1(n_0),
.A2(n_51),
.B(n_65),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_0),
.B(n_66),
.Y(n_145)
);

AOI21xp33_ASAP7_75t_SL g153 ( 
.A1(n_0),
.A2(n_36),
.B(n_154),
.Y(n_153)
);

AOI21xp33_ASAP7_75t_L g173 ( 
.A1(n_0),
.A2(n_22),
.B(n_37),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_0),
.B(n_47),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_4),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_4),
.A2(n_28),
.B1(n_35),
.B2(n_36),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_6),
.A2(n_22),
.B1(n_27),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_8),
.A2(n_22),
.B1(n_27),
.B2(n_38),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_9),
.A2(n_41),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_9),
.A2(n_41),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_9),
.A2(n_22),
.B1(n_27),
.B2(n_41),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_10),
.A2(n_50),
.B1(n_51),
.B2(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_11),
.Y(n_23)
);

HAxp5_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_119),
.CON(n_12),
.SN(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_117),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_100),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_15),
.B(n_100),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_81),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_70),
.B2(n_71),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_44),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_20),
.A2(n_32),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_20),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_21),
.B(n_24),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_21),
.A2(n_29),
.B1(n_87),
.B2(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_24),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_22),
.Y(n_27)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_26),
.A2(n_29),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_27),
.B(n_186),
.Y(n_185)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_29),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_29),
.B(n_43),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_30),
.B(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_32),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_32),
.A2(n_104),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_32),
.A2(n_104),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_32),
.B(n_112),
.C(n_177),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_32),
.B(n_159),
.C(n_167),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_33),
.B(n_42),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_33),
.B(n_39),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_39),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_36),
.A2(n_38),
.B(n_43),
.C(n_173),
.Y(n_172)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_39),
.A2(n_73),
.B(n_74),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_39),
.B(n_43),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_42),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_43),
.A2(n_61),
.B(n_64),
.C(n_111),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_43),
.A2(n_48),
.B(n_51),
.C(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_57),
.B1(n_68),
.B2(n_69),
.Y(n_44)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_45),
.B(n_97),
.C(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_45),
.A2(n_68),
.B1(n_127),
.B2(n_128),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_45),
.A2(n_68),
.B1(n_88),
.B2(n_89),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_49),
.B(n_52),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_46),
.A2(n_49),
.B1(n_95),
.B2(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_47),
.B(n_54),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_51),
.B1(n_64),
.B2(n_65),
.Y(n_66)
);

INVx5_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_56),
.Y(n_154)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_57),
.B(n_108),
.C(n_114),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_57),
.A2(n_69),
.B1(n_114),
.B2(n_115),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_62),
.B1(n_66),
.B2(n_67),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_59),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_67),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_68),
.B(n_89),
.C(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_76),
.B1(n_77),
.B2(n_80),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_72),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_90),
.B(n_91),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

INVxp33_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_79),
.B(n_86),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_92),
.C(n_96),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_88),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_83),
.A2(n_88),
.B1(n_89),
.B2(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_83),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_84),
.A2(n_113),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_88),
.A2(n_89),
.B1(n_172),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_89),
.B(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_92),
.A2(n_93),
.B1(n_96),
.B2(n_97),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_96),
.A2(n_97),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.C(n_106),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_101),
.B(n_103),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_106),
.A2(n_107),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_108),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_110),
.B1(n_112),
.B2(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_112),
.A2(n_139),
.B1(n_175),
.B2(n_178),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_112),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_112),
.B(n_188),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_114),
.A2(n_115),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_141),
.C(n_144),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_146),
.B(n_204),
.C(n_209),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_134),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_121),
.B(n_134),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_122),
.B(n_125),
.C(n_132),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_131),
.B2(n_132),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.C(n_140),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_135),
.B(n_201),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_136),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_138),
.B(n_140),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_141),
.A2(n_144),
.B1(n_145),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_141),
.B(n_185),
.Y(n_184)
);

INVx5_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_203),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_198),
.B(n_202),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_168),
.B(n_197),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_158),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_150),
.B(n_158),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_151),
.B(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_152),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_157),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_164),
.B2(n_165),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_161),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_162),
.B(n_181),
.Y(n_190)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_166),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_192),
.B(n_196),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_179),
.B(n_191),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_174),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_172),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_175),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_176),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_183),
.B(n_190),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_187),
.B(n_189),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_194),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_200),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_205),
.B(n_206),
.Y(n_209)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);


endmodule