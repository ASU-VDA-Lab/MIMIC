module fake_jpeg_31168_n_363 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_363);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_363;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_21),
.B(n_9),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_53),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_0),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_35),
.C(n_23),
.Y(n_59)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_21),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_57),
.Y(n_67)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_26),
.B1(n_25),
.B2(n_37),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_58),
.A2(n_70),
.B1(n_73),
.B2(n_49),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_59),
.B(n_83),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_26),
.B1(n_25),
.B2(n_38),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_62),
.A2(n_65),
.B1(n_78),
.B2(n_82),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_26),
.B1(n_38),
.B2(n_34),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_40),
.A2(n_41),
.B1(n_28),
.B2(n_36),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_68),
.A2(n_72),
.B1(n_90),
.B2(n_57),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_51),
.A2(n_39),
.B1(n_37),
.B2(n_23),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_30),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_71),
.B(n_81),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_40),
.A2(n_18),
.B1(n_36),
.B2(n_28),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_39),
.B1(n_37),
.B2(n_23),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_41),
.A2(n_18),
.B1(n_36),
.B2(n_28),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_34),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_31),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_48),
.B(n_29),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_49),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_43),
.A2(n_18),
.B1(n_39),
.B2(n_24),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_86),
.A2(n_88),
.B1(n_42),
.B2(n_50),
.Y(n_130)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_43),
.A2(n_24),
.B1(n_29),
.B2(n_20),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_20),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_89),
.B(n_52),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_50),
.A2(n_20),
.B1(n_10),
.B2(n_17),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_SL g92 ( 
.A1(n_89),
.A2(n_57),
.B(n_49),
.C(n_52),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_92),
.A2(n_102),
.B(n_128),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_65),
.A2(n_63),
.B1(n_88),
.B2(n_67),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_93),
.A2(n_130),
.B1(n_73),
.B2(n_61),
.Y(n_142)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_95),
.B(n_100),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_97),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_71),
.Y(n_100)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_104),
.B(n_106),
.Y(n_153)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_105),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_81),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_77),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_108),
.B(n_118),
.Y(n_160)
);

AND2x4_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_57),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_110),
.B(n_113),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_111),
.B(n_129),
.Y(n_164)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_82),
.A2(n_63),
.B1(n_78),
.B2(n_76),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_114),
.A2(n_134),
.B1(n_87),
.B2(n_79),
.Y(n_152)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_53),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_116),
.B(n_120),
.Y(n_162)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_76),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_64),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_62),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_126),
.Y(n_166)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_125),
.Y(n_138)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_59),
.B(n_53),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_127),
.Y(n_158)
);

O2A1O1Ixp33_ASAP7_75t_SL g128 ( 
.A1(n_86),
.A2(n_52),
.B(n_44),
.C(n_47),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_58),
.A2(n_47),
.B1(n_44),
.B2(n_42),
.Y(n_129)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_131),
.A2(n_64),
.B1(n_87),
.B2(n_69),
.Y(n_139)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_64),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_132),
.Y(n_159)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_133),
.B(n_80),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_85),
.A2(n_43),
.B1(n_42),
.B2(n_54),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_135),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_139),
.A2(n_118),
.B(n_128),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_85),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_108),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_142),
.A2(n_152),
.B1(n_156),
.B2(n_157),
.Y(n_177)
);

OR2x2_ASAP7_75t_SL g146 ( 
.A(n_109),
.B(n_85),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_L g180 ( 
.A1(n_146),
.A2(n_109),
.B(n_92),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_123),
.A2(n_54),
.B1(n_79),
.B2(n_50),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_79),
.B1(n_56),
.B2(n_69),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_133),
.A2(n_56),
.B1(n_24),
.B2(n_22),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_167),
.A2(n_130),
.B1(n_129),
.B2(n_134),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_121),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_170),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_179),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_121),
.C(n_110),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_171),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_172),
.A2(n_150),
.B(n_165),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_173),
.A2(n_186),
.B1(n_188),
.B2(n_193),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_106),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_187),
.Y(n_204)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_175),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_153),
.B(n_104),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_178),
.B(n_157),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_97),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_180),
.A2(n_140),
.B(n_146),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_122),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_182),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_109),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_107),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_185),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_122),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_166),
.A2(n_115),
.B1(n_119),
.B2(n_117),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_160),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_166),
.A2(n_96),
.B1(n_99),
.B2(n_91),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_132),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_191),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_126),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_164),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_160),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_164),
.A2(n_140),
.B(n_160),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_192),
.A2(n_164),
.B(n_140),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_155),
.A2(n_56),
.B1(n_131),
.B2(n_112),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_145),
.Y(n_194)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_135),
.Y(n_196)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_164),
.B(n_120),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_167),
.Y(n_225)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_149),
.Y(n_198)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_155),
.A2(n_125),
.B1(n_101),
.B2(n_94),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_199),
.A2(n_140),
.B1(n_138),
.B2(n_152),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_187),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_179),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_202),
.B(n_205),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_190),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_207),
.B(n_208),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_185),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_229),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_225),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_215),
.B(n_219),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_216),
.A2(n_173),
.B1(n_196),
.B2(n_176),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_168),
.B(n_142),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_223),
.C(n_171),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_170),
.B(n_156),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_192),
.A2(n_138),
.B(n_159),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_224),
.A2(n_226),
.B(n_231),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_181),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_184),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_169),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_191),
.A2(n_159),
.B(n_149),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_234),
.A2(n_245),
.B1(n_214),
.B2(n_225),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_212),
.B(n_178),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_236),
.Y(n_267)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_256),
.Y(n_272)
);

BUFx24_ASAP7_75t_SL g240 ( 
.A(n_229),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_240),
.B(n_243),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_214),
.A2(n_177),
.B1(n_220),
.B2(n_207),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_241),
.A2(n_206),
.B1(n_215),
.B2(n_221),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_213),
.A2(n_182),
.B(n_172),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_242),
.A2(n_244),
.B(n_250),
.Y(n_270)
);

AOI322xp5_ASAP7_75t_SL g243 ( 
.A1(n_204),
.A2(n_193),
.A3(n_199),
.B1(n_188),
.B2(n_186),
.C1(n_10),
.C2(n_12),
.Y(n_243)
);

A2O1A1Ixp33_ASAP7_75t_SL g244 ( 
.A1(n_224),
.A2(n_177),
.B(n_175),
.C(n_137),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_216),
.A2(n_194),
.B1(n_183),
.B2(n_195),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_204),
.B(n_198),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_248),
.B(n_258),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_249),
.B(n_223),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_202),
.A2(n_150),
.B1(n_147),
.B2(n_165),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_200),
.Y(n_251)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_251),
.Y(n_278)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_200),
.Y(n_252)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_203),
.B(n_136),
.C(n_147),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_254),
.C(n_255),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_203),
.B(n_136),
.C(n_103),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_103),
.C(n_161),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_211),
.Y(n_256)
);

AO22x1_ASAP7_75t_L g257 ( 
.A1(n_220),
.A2(n_151),
.B1(n_148),
.B2(n_137),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_227),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_144),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_218),
.B(n_151),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_259),
.B(n_217),
.Y(n_281)
);

OAI22x1_ASAP7_75t_L g263 ( 
.A1(n_244),
.A2(n_257),
.B1(n_226),
.B2(n_237),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_263),
.A2(n_242),
.B1(n_244),
.B2(n_246),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_265),
.A2(n_268),
.B1(n_269),
.B2(n_233),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_266),
.B(n_277),
.C(n_279),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_234),
.A2(n_245),
.B1(n_239),
.B2(n_241),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_237),
.A2(n_221),
.B1(n_210),
.B2(n_201),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_235),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_280),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_273),
.A2(n_274),
.B1(n_282),
.B2(n_276),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_246),
.A2(n_206),
.B1(n_211),
.B2(n_231),
.Y(n_274)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_276),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_219),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_210),
.C(n_217),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_247),
.Y(n_280)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_281),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_246),
.A2(n_227),
.B1(n_228),
.B2(n_209),
.Y(n_282)
);

BUFx5_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_283),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_284),
.A2(n_292),
.B1(n_293),
.B2(n_301),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_285),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_287),
.A2(n_294),
.B1(n_297),
.B2(n_275),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_265),
.A2(n_244),
.B1(n_255),
.B2(n_251),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_288),
.A2(n_290),
.B1(n_299),
.B2(n_284),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_277),
.B(n_232),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_264),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_252),
.Y(n_290)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_290),
.Y(n_307)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_291),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_263),
.A2(n_244),
.B1(n_253),
.B2(n_250),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_273),
.A2(n_256),
.B1(n_232),
.B2(n_228),
.Y(n_293)
);

AOI221xp5_ASAP7_75t_L g294 ( 
.A1(n_269),
.A2(n_209),
.B1(n_137),
.B2(n_148),
.C(n_151),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_278),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_303),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_209),
.B1(n_161),
.B2(n_105),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_270),
.A2(n_274),
.B(n_282),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_299),
.A2(n_288),
.B(n_298),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_270),
.A2(n_161),
.B1(n_148),
.B2(n_11),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_278),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_260),
.C(n_266),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_310),
.C(n_317),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_267),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_306),
.B(n_311),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_316),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_260),
.C(n_279),
.Y(n_310)
);

AO21x1_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_268),
.B(n_261),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_319),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_275),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_313),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_314),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_293),
.B(n_262),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_289),
.B(n_22),
.C(n_24),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_287),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_318),
.B(n_320),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_316),
.B(n_300),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_321),
.B(n_326),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_319),
.A2(n_292),
.B(n_295),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_324),
.A2(n_331),
.B(n_8),
.Y(n_343)
);

NAND3xp33_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_309),
.C(n_303),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_301),
.C(n_22),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_304),
.Y(n_334)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_307),
.Y(n_328)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_328),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_329),
.A2(n_314),
.B1(n_320),
.B2(n_305),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_313),
.A2(n_9),
.B(n_15),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_334),
.B(n_337),
.Y(n_348)
);

NOR2xp67_ASAP7_75t_L g335 ( 
.A(n_322),
.B(n_312),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g351 ( 
.A(n_335),
.B(n_339),
.Y(n_351)
);

NOR2xp67_ASAP7_75t_SL g336 ( 
.A(n_322),
.B(n_311),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_336),
.B(n_341),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_325),
.B(n_327),
.Y(n_337)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_338),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_330),
.B(n_305),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_332),
.A2(n_317),
.B(n_8),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_343),
.B(n_329),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_340),
.A2(n_323),
.B(n_333),
.Y(n_345)
);

NAND3xp33_ASAP7_75t_SL g353 ( 
.A(n_345),
.B(n_346),
.C(n_347),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_339),
.A2(n_328),
.B(n_324),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_338),
.B(n_325),
.C(n_331),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_349),
.B(n_342),
.C(n_11),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_351),
.A2(n_344),
.B1(n_346),
.B2(n_350),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_352),
.B(n_354),
.C(n_1),
.Y(n_359)
);

OAI321xp33_ASAP7_75t_L g355 ( 
.A1(n_348),
.A2(n_7),
.A3(n_14),
.B1(n_13),
.B2(n_12),
.C(n_24),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_355),
.A2(n_7),
.B1(n_3),
.B2(n_4),
.Y(n_357)
);

AOI321xp33_ASAP7_75t_L g356 ( 
.A1(n_351),
.A2(n_7),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_356),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_357),
.B(n_359),
.Y(n_361)
);

AND2x4_ASAP7_75t_L g360 ( 
.A(n_358),
.B(n_353),
.Y(n_360)
);

AOI322xp5_ASAP7_75t_L g362 ( 
.A1(n_360),
.A2(n_3),
.A3(n_4),
.B1(n_6),
.B2(n_22),
.C1(n_345),
.C2(n_353),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_362),
.B(n_361),
.Y(n_363)
);


endmodule