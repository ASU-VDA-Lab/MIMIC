module real_jpeg_11659_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_17;
wire n_43;
wire n_37;
wire n_21;
wire n_38;
wire n_35;
wire n_33;
wire n_29;
wire n_49;
wire n_31;
wire n_24;
wire n_34;
wire n_44;
wire n_28;
wire n_46;
wire n_23;
wire n_47;
wire n_14;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_40;
wire n_36;
wire n_39;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_48;
wire n_27;
wire n_30;
wire n_16;
wire n_15;

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_0),
.B(n_2),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_0),
.B(n_2),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_0),
.B(n_45),
.C(n_49),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_3),
.A2(n_19),
.B1(n_20),
.B2(n_42),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_4),
.A2(n_9),
.B(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_6),
.B(n_40),
.C(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_7),
.B(n_12),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_8),
.B(n_26),
.C(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_9),
.B(n_32),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_11),
.A2(n_31),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_18),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_16),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_38),
.B(n_41),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_36),
.B(n_37),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.B(n_35),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_26),
.Y(n_35)
);

O2A1O1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_29),
.B(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_40),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);


endmodule