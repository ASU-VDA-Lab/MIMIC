module fake_jpeg_16_n_464 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_464);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_464;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

CKINVDCx11_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_55),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_28),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_56),
.B(n_62),
.Y(n_129)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_54),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g116 ( 
.A(n_57),
.Y(n_116)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_58),
.Y(n_127)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_59),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_39),
.Y(n_60)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_54),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_63),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_L g64 ( 
.A1(n_28),
.A2(n_6),
.B(n_15),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_64),
.B(n_67),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_34),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_68),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_69),
.Y(n_178)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_34),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_74),
.B(n_77),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_75),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_50),
.Y(n_76)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_76),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_34),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_78),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_24),
.B(n_31),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_79),
.B(n_80),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_48),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_81),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_48),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_82),
.B(n_85),
.Y(n_171)
);

BUFx6f_ASAP7_75t_SL g83 ( 
.A(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_83),
.Y(n_175)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_48),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_33),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_88),
.B(n_90),
.Y(n_177)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_89),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_33),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_91),
.Y(n_163)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_93),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_94),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_24),
.B(n_7),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_95),
.B(n_98),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_97),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_25),
.B(n_31),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_99),
.Y(n_182)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_100),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_25),
.B(n_7),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_101),
.B(n_109),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_46),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_102),
.B(n_115),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_104),
.Y(n_169)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_22),
.Y(n_105)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_105),
.Y(n_183)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_29),
.Y(n_106)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_106),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_36),
.Y(n_107)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_107),
.Y(n_172)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_32),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_41),
.B(n_42),
.Y(n_109)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_32),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_111),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_20),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_21),
.Y(n_149)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_20),
.Y(n_113)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_113),
.Y(n_190)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_29),
.Y(n_114)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_114),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_41),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_76),
.A2(n_23),
.B1(n_47),
.B2(n_43),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_117),
.A2(n_123),
.B1(n_124),
.B2(n_138),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_65),
.A2(n_23),
.B1(n_53),
.B2(n_51),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_119),
.A2(n_180),
.B1(n_184),
.B2(n_186),
.Y(n_204)
);

NAND2x1_ASAP7_75t_L g120 ( 
.A(n_58),
.B(n_38),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_120),
.B(n_158),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_111),
.A2(n_47),
.B1(n_43),
.B2(n_42),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_60),
.A2(n_40),
.B1(n_38),
.B2(n_30),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_61),
.A2(n_73),
.B1(n_63),
.B2(n_70),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_75),
.B(n_40),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_139),
.B(n_179),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_72),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_140),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_105),
.A2(n_30),
.B1(n_51),
.B2(n_45),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_141),
.A2(n_145),
.B1(n_150),
.B2(n_156),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_55),
.A2(n_53),
.B1(n_45),
.B2(n_21),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_149),
.B(n_86),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_112),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_151),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_108),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_81),
.B(n_5),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_91),
.A2(n_5),
.B1(n_8),
.B2(n_12),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_176),
.A2(n_174),
.B1(n_165),
.B2(n_122),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_75),
.B(n_5),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_94),
.A2(n_1),
.B1(n_4),
.B2(n_15),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_84),
.B(n_15),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_188),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_96),
.A2(n_4),
.B1(n_16),
.B2(n_97),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_92),
.Y(n_185)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_99),
.A2(n_69),
.B1(n_59),
.B2(n_66),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_103),
.Y(n_187)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_86),
.B(n_57),
.Y(n_188)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_134),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_191),
.Y(n_258)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_189),
.Y(n_192)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_192),
.Y(n_256)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_147),
.Y(n_193)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_193),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_194),
.B(n_234),
.Y(n_263)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_121),
.Y(n_196)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_196),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_143),
.A2(n_68),
.B(n_83),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_197),
.A2(n_211),
.B(n_247),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_177),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_198),
.B(n_227),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_154),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_199),
.Y(n_271)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_137),
.Y(n_200)
);

BUFx4f_ASAP7_75t_SL g285 ( 
.A(n_200),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_129),
.B(n_113),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_201),
.B(n_202),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_153),
.B(n_110),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_130),
.B(n_87),
.C(n_104),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_205),
.B(n_209),
.C(n_247),
.Y(n_272)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_206),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_158),
.B(n_120),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_160),
.B(n_87),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_210),
.B(n_216),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_149),
.A2(n_93),
.B(n_100),
.Y(n_211)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_152),
.Y(n_212)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_212),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_148),
.B(n_107),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_213),
.B(n_241),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_157),
.B(n_173),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_127),
.Y(n_217)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_217),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_155),
.B(n_171),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_218),
.B(n_220),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_219),
.A2(n_238),
.B1(n_194),
.B2(n_205),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_116),
.B(n_159),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_128),
.Y(n_221)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_221),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_184),
.A2(n_180),
.B1(n_145),
.B2(n_123),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_222),
.A2(n_233),
.B1(n_230),
.B2(n_213),
.Y(n_278)
);

INVx11_ASAP7_75t_L g223 ( 
.A(n_116),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_223),
.Y(n_276)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_174),
.Y(n_225)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_225),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_134),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_226),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_154),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_183),
.B(n_126),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_236),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_178),
.Y(n_229)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_229),
.Y(n_288)
);

A2O1A1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_119),
.A2(n_146),
.B(n_144),
.C(n_142),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_230),
.B(n_242),
.Y(n_291)
);

AND2x2_ASAP7_75t_SL g231 ( 
.A(n_136),
.B(n_161),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_231),
.Y(n_265)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_175),
.Y(n_232)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_232),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_156),
.A2(n_117),
.B1(n_124),
.B2(n_163),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_118),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_133),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_235),
.B(n_245),
.Y(n_297)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_133),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_131),
.B(n_118),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_237),
.B(n_246),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_186),
.A2(n_178),
.B1(n_169),
.B2(n_172),
.Y(n_238)
);

INVx11_ASAP7_75t_L g239 ( 
.A(n_166),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_239),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_182),
.B(n_163),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_125),
.Y(n_242)
);

OR2x2_ASAP7_75t_SL g243 ( 
.A(n_150),
.B(n_170),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_243),
.Y(n_298)
);

INVx11_ASAP7_75t_L g245 ( 
.A(n_135),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_135),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_132),
.B(n_162),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_182),
.B(n_162),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_249),
.Y(n_270)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_168),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_164),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_250),
.B(n_251),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_168),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_164),
.B(n_167),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_252),
.B(n_199),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_224),
.A2(n_167),
.B(n_244),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_253),
.Y(n_322)
);

MAJx2_ASAP7_75t_L g255 ( 
.A(n_207),
.B(n_209),
.C(n_244),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_255),
.B(n_267),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_222),
.A2(n_233),
.B1(n_204),
.B2(n_194),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_260),
.B(n_195),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_207),
.B(n_197),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_215),
.A2(n_204),
.B1(n_241),
.B2(n_248),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_268),
.A2(n_278),
.B1(n_286),
.B2(n_208),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_275),
.A2(n_245),
.B1(n_203),
.B2(n_239),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_240),
.A2(n_243),
.B(n_211),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_279),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_231),
.B(n_193),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_281),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_231),
.B(n_217),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_293),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_221),
.A2(n_206),
.B1(n_249),
.B2(n_250),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_235),
.B(n_214),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_191),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_200),
.B(n_234),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_294),
.B(n_276),
.Y(n_319)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_289),
.Y(n_302)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_302),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_266),
.B(n_214),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_303),
.B(n_309),
.Y(n_335)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_292),
.Y(n_304)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_304),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_297),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_305),
.Y(n_348)
);

NAND3xp33_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_223),
.C(n_247),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_306),
.B(n_318),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_298),
.A2(n_212),
.B1(n_229),
.B2(n_208),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_307),
.A2(n_333),
.B(n_263),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_308),
.A2(n_321),
.B1(n_272),
.B2(n_263),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_269),
.B(n_232),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_310),
.B(n_319),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_266),
.B(n_226),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_311),
.B(n_312),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_267),
.B(n_195),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_297),
.Y(n_313)
);

INVx13_ASAP7_75t_L g346 ( 
.A(n_313),
.Y(n_346)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_292),
.Y(n_314)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_314),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_315),
.A2(n_328),
.B1(n_329),
.B2(n_334),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_277),
.B(n_203),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_316),
.B(n_317),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_297),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_260),
.A2(n_278),
.B1(n_253),
.B2(n_268),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_270),
.Y(n_323)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_323),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_282),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_324),
.B(n_325),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_290),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_270),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_327),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_255),
.B(n_280),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_287),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_261),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_277),
.B(n_257),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_330),
.B(n_331),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_262),
.B(n_264),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_281),
.B(n_291),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_332),
.B(n_327),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_264),
.B(n_256),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_261),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_308),
.A2(n_265),
.B1(n_279),
.B2(n_283),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_338),
.A2(n_341),
.B1(n_344),
.B2(n_353),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_342),
.B(n_299),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_321),
.A2(n_272),
.B1(n_263),
.B2(n_256),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_345),
.A2(n_307),
.B(n_301),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_333),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_347),
.B(n_352),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_320),
.B(n_274),
.C(n_276),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_351),
.B(n_359),
.C(n_361),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_330),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_323),
.A2(n_287),
.B1(n_258),
.B2(n_254),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_326),
.A2(n_258),
.B1(n_254),
.B2(n_296),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_355),
.A2(n_362),
.B1(n_305),
.B2(n_318),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_320),
.B(n_312),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_301),
.B(n_274),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_315),
.A2(n_259),
.B1(n_296),
.B2(n_284),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_357),
.A2(n_322),
.B1(n_348),
.B2(n_315),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_363),
.A2(n_379),
.B1(n_381),
.B2(n_382),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_347),
.B(n_302),
.Y(n_365)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_365),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_366),
.B(n_342),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_335),
.B(n_356),
.Y(n_367)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_367),
.Y(n_395)
);

XOR2x2_ASAP7_75t_L g368 ( 
.A(n_359),
.B(n_332),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_368),
.B(n_376),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_352),
.B(n_331),
.Y(n_370)
);

INVxp33_ASAP7_75t_L g399 ( 
.A(n_370),
.Y(n_399)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_340),
.Y(n_371)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_371),
.Y(n_402)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_340),
.Y(n_372)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_372),
.Y(n_403)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_350),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_373),
.B(n_375),
.Y(n_388)
);

AOI21x1_ASAP7_75t_SL g396 ( 
.A1(n_374),
.A2(n_357),
.B(n_338),
.Y(n_396)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_350),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_360),
.B(n_300),
.Y(n_376)
);

AOI32xp33_ASAP7_75t_L g377 ( 
.A1(n_336),
.A2(n_324),
.A3(n_325),
.B1(n_316),
.B2(n_313),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_377),
.A2(n_383),
.B(n_345),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_354),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_378),
.Y(n_390)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_353),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_358),
.B(n_310),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_380),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_358),
.B(n_285),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_355),
.Y(n_382)
);

CKINVDCx14_ASAP7_75t_R g383 ( 
.A(n_343),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_384),
.A2(n_349),
.B1(n_311),
.B2(n_300),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_385),
.B(n_351),
.C(n_344),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_386),
.B(n_387),
.C(n_400),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_385),
.B(n_341),
.C(n_361),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_391),
.B(n_370),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_368),
.B(n_360),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_392),
.B(n_376),
.Y(n_408)
);

AOI21x1_ASAP7_75t_SL g412 ( 
.A1(n_393),
.A2(n_396),
.B(n_377),
.Y(n_412)
);

OAI21xp33_ASAP7_75t_L g406 ( 
.A1(n_396),
.A2(n_374),
.B(n_364),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_368),
.B(n_356),
.C(n_339),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_364),
.A2(n_339),
.B1(n_335),
.B2(n_349),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_401),
.A2(n_404),
.B1(n_365),
.B2(n_367),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_406),
.B(n_413),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_386),
.B(n_387),
.C(n_397),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_407),
.B(n_411),
.C(n_417),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_408),
.B(n_416),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_390),
.B(n_378),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_409),
.B(n_414),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_410),
.A2(n_415),
.B1(n_401),
.B2(n_394),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_397),
.B(n_400),
.C(n_392),
.Y(n_411)
);

OAI21x1_ASAP7_75t_L g429 ( 
.A1(n_412),
.A2(n_419),
.B(n_384),
.Y(n_429)
);

AO22x1_ASAP7_75t_L g413 ( 
.A1(n_394),
.A2(n_382),
.B1(n_379),
.B2(n_369),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_393),
.B(n_375),
.C(n_373),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_389),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_398),
.B(n_372),
.C(n_371),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_391),
.B(n_369),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_418),
.B(n_404),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_399),
.B(n_303),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_422),
.B(n_411),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_423),
.A2(n_424),
.B1(n_427),
.B2(n_388),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_415),
.A2(n_406),
.B(n_412),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_405),
.B(n_395),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_426),
.B(n_407),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_413),
.A2(n_395),
.B1(n_402),
.B2(n_403),
.Y(n_427)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_418),
.Y(n_428)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_428),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_429),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_431),
.B(n_432),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_421),
.B(n_422),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_432),
.B(n_436),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_425),
.B(n_426),
.C(n_405),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_433),
.B(n_435),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_430),
.A2(n_388),
.B(n_408),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_434),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_425),
.B(n_403),
.C(n_402),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_439),
.B(n_421),
.C(n_430),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_440),
.B(n_443),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_438),
.A2(n_420),
.B1(n_428),
.B2(n_362),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_433),
.B(n_309),
.C(n_337),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_445),
.B(n_437),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_434),
.A2(n_346),
.B(n_334),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_446),
.A2(n_346),
.B(n_314),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_447),
.B(n_259),
.C(n_328),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_441),
.A2(n_439),
.B(n_431),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_448),
.B(n_449),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_442),
.B(n_304),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_451),
.B(n_442),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_452),
.B(n_329),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_453),
.B(n_447),
.C(n_444),
.Y(n_457)
);

O2A1O1Ixp33_ASAP7_75t_SL g458 ( 
.A1(n_455),
.A2(n_456),
.B(n_450),
.C(n_288),
.Y(n_458)
);

AOI31xp67_ASAP7_75t_SL g459 ( 
.A1(n_457),
.A2(n_285),
.A3(n_271),
.B(n_288),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_458),
.B(n_459),
.Y(n_460)
);

OAI22xp33_ASAP7_75t_SL g461 ( 
.A1(n_460),
.A2(n_455),
.B1(n_454),
.B2(n_273),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_461),
.B(n_271),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_462),
.B(n_273),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_463),
.B(n_285),
.Y(n_464)
);


endmodule