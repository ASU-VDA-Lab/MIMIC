module real_aes_8217_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_404;
wire n_147;
wire n_288;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_0), .B(n_112), .C(n_113), .Y(n_111) );
INVx1_ASAP7_75t_L g458 ( .A(n_0), .Y(n_458) );
INVx1_ASAP7_75t_L g513 ( .A(n_1), .Y(n_513) );
INVx1_ASAP7_75t_L g204 ( .A(n_2), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_3), .A2(n_37), .B1(n_176), .B2(n_522), .Y(n_521) );
AOI21xp33_ASAP7_75t_L g215 ( .A1(n_4), .A2(n_133), .B(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_5), .B(n_163), .Y(n_505) );
AND2x6_ASAP7_75t_L g138 ( .A(n_6), .B(n_139), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_7), .A2(n_184), .B(n_185), .Y(n_183) );
INVx1_ASAP7_75t_L g109 ( .A(n_8), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_8), .B(n_38), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_9), .B(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g221 ( .A(n_10), .Y(n_221) );
INVx1_ASAP7_75t_L g159 ( .A(n_11), .Y(n_159) );
INVx1_ASAP7_75t_L g509 ( .A(n_12), .Y(n_509) );
INVx1_ASAP7_75t_L g192 ( .A(n_13), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_14), .B(n_207), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_15), .B(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_16), .B(n_155), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_17), .A2(n_41), .B1(n_754), .B2(n_755), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_17), .Y(n_755) );
AO32x2_ASAP7_75t_L g519 ( .A1(n_18), .A2(n_154), .A3(n_163), .B1(n_491), .B2(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_19), .B(n_176), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_20), .B(n_149), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_21), .B(n_155), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_22), .A2(n_49), .B1(n_176), .B2(n_522), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g132 ( .A(n_23), .B(n_133), .Y(n_132) );
AOI22xp33_ASAP7_75t_SL g558 ( .A1(n_24), .A2(n_75), .B1(n_176), .B2(n_207), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_25), .B(n_176), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_26), .B(n_214), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g188 ( .A1(n_27), .A2(n_189), .B(n_191), .C(n_193), .Y(n_188) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_28), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_29), .B(n_167), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_30), .B(n_174), .Y(n_205) );
INVx1_ASAP7_75t_L g231 ( .A(n_31), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_32), .B(n_167), .Y(n_535) );
INVx2_ASAP7_75t_L g136 ( .A(n_33), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_34), .B(n_176), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_35), .B(n_167), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g140 ( .A1(n_36), .A2(n_138), .B(n_141), .C(n_144), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_38), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g229 ( .A(n_39), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_40), .B(n_174), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_41), .Y(n_754) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_42), .B(n_176), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_43), .A2(n_86), .B1(n_152), .B2(n_522), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_44), .B(n_176), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_45), .B(n_176), .Y(n_510) );
CKINVDCx16_ASAP7_75t_R g232 ( .A(n_46), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_47), .B(n_489), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_48), .B(n_133), .Y(n_177) );
AOI22xp33_ASAP7_75t_SL g570 ( .A1(n_50), .A2(n_59), .B1(n_176), .B2(n_207), .Y(n_570) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_51), .A2(n_141), .B1(n_207), .B2(n_228), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g161 ( .A(n_52), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_53), .B(n_176), .Y(n_490) );
CKINVDCx16_ASAP7_75t_R g200 ( .A(n_54), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_55), .B(n_176), .Y(n_539) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_56), .A2(n_219), .B(n_220), .C(n_222), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_57), .Y(n_269) );
INVx1_ASAP7_75t_L g217 ( .A(n_58), .Y(n_217) );
INVx1_ASAP7_75t_L g139 ( .A(n_60), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_61), .B(n_176), .Y(n_514) );
INVx1_ASAP7_75t_L g158 ( .A(n_62), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_63), .Y(n_121) );
AO32x2_ASAP7_75t_L g555 ( .A1(n_64), .A2(n_163), .A3(n_166), .B1(n_491), .B2(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g487 ( .A(n_65), .Y(n_487) );
INVx1_ASAP7_75t_L g530 ( .A(n_66), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_SL g239 ( .A1(n_67), .A2(n_149), .B(n_222), .C(n_240), .Y(n_239) );
INVxp67_ASAP7_75t_L g241 ( .A(n_68), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_69), .B(n_207), .Y(n_531) );
INVx1_ASAP7_75t_L g115 ( .A(n_70), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_71), .Y(n_234) );
INVx1_ASAP7_75t_L g262 ( .A(n_72), .Y(n_262) );
OAI321xp33_ASAP7_75t_L g122 ( .A1(n_73), .A2(n_123), .A3(n_453), .B1(n_460), .B2(n_461), .C(n_463), .Y(n_122) );
CKINVDCx16_ASAP7_75t_R g460 ( .A(n_73), .Y(n_460) );
OAI22xp5_ASAP7_75t_SL g450 ( .A1(n_74), .A2(n_88), .B1(n_451), .B2(n_452), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_74), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g263 ( .A1(n_76), .A2(n_138), .B(n_141), .C(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_77), .B(n_522), .Y(n_544) );
OAI22xp5_ASAP7_75t_SL g751 ( .A1(n_78), .A2(n_752), .B1(n_753), .B2(n_756), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_78), .Y(n_756) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_79), .B(n_207), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_80), .B(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g156 ( .A(n_81), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_82), .B(n_149), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_83), .B(n_207), .Y(n_500) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_84), .A2(n_138), .B(n_141), .C(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g112 ( .A(n_85), .Y(n_112) );
OR2x2_ASAP7_75t_L g455 ( .A(n_85), .B(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g471 ( .A(n_85), .B(n_457), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_87), .A2(n_102), .B1(n_207), .B2(n_208), .Y(n_569) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_88), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_89), .B(n_167), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_90), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g169 ( .A1(n_91), .A2(n_138), .B(n_141), .C(n_170), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_92), .Y(n_179) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_93), .A2(n_104), .B1(n_116), .B2(n_764), .Y(n_103) );
INVx1_ASAP7_75t_L g238 ( .A(n_94), .Y(n_238) );
CKINVDCx16_ASAP7_75t_R g186 ( .A(n_95), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_96), .B(n_146), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_97), .B(n_207), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_98), .B(n_163), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_99), .B(n_115), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_100), .A2(n_133), .B(n_237), .Y(n_236) );
AOI222xp33_ASAP7_75t_L g467 ( .A1(n_101), .A2(n_468), .B1(n_750), .B2(n_751), .C1(n_757), .C2(n_760), .Y(n_467) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g764 ( .A(n_106), .Y(n_764) );
AND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g474 ( .A(n_112), .B(n_457), .Y(n_474) );
NOR2x2_ASAP7_75t_L g759 ( .A(n_112), .B(n_456), .Y(n_759) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
OA21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_122), .B(n_466), .Y(n_116) );
BUFx2_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g763 ( .A(n_120), .Y(n_763) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_123), .B(n_462), .Y(n_461) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_124), .A2(n_125), .B1(n_449), .B2(n_450), .Y(n_123) );
OAI22xp5_ASAP7_75t_SL g760 ( .A1(n_124), .A2(n_471), .B1(n_472), .B2(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_125), .A2(n_469), .B1(n_472), .B2(n_475), .Y(n_468) );
AND2x2_ASAP7_75t_SL g125 ( .A(n_126), .B(n_418), .Y(n_125) );
NOR3xp33_ASAP7_75t_L g126 ( .A(n_127), .B(n_311), .C(n_384), .Y(n_126) );
OAI211xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_196), .B(n_243), .C(n_295), .Y(n_127) );
INVxp67_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_164), .Y(n_129) );
AND2x2_ASAP7_75t_L g259 ( .A(n_130), .B(n_260), .Y(n_259) );
INVx3_ASAP7_75t_L g278 ( .A(n_130), .Y(n_278) );
INVx2_ASAP7_75t_L g293 ( .A(n_130), .Y(n_293) );
INVx1_ASAP7_75t_L g323 ( .A(n_130), .Y(n_323) );
AND2x2_ASAP7_75t_L g373 ( .A(n_130), .B(n_294), .Y(n_373) );
AOI32xp33_ASAP7_75t_L g400 ( .A1(n_130), .A2(n_328), .A3(n_401), .B1(n_403), .B2(n_404), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_130), .B(n_249), .Y(n_406) );
AND2x2_ASAP7_75t_L g433 ( .A(n_130), .B(n_276), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_130), .B(n_442), .Y(n_441) );
OR2x6_ASAP7_75t_L g130 ( .A(n_131), .B(n_160), .Y(n_130) );
AOI21xp5_ASAP7_75t_SL g131 ( .A1(n_132), .A2(n_140), .B(n_153), .Y(n_131) );
BUFx2_ASAP7_75t_L g184 ( .A(n_133), .Y(n_184) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_138), .Y(n_133) );
NAND2x1p5_ASAP7_75t_L g201 ( .A(n_134), .B(n_138), .Y(n_201) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
INVx1_ASAP7_75t_L g489 ( .A(n_135), .Y(n_489) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g142 ( .A(n_136), .Y(n_142) );
INVx1_ASAP7_75t_L g208 ( .A(n_136), .Y(n_208) );
INVx1_ASAP7_75t_L g143 ( .A(n_137), .Y(n_143) );
INVx3_ASAP7_75t_L g147 ( .A(n_137), .Y(n_147) );
INVx1_ASAP7_75t_L g149 ( .A(n_137), .Y(n_149) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_137), .Y(n_174) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_137), .Y(n_190) );
INVx4_ASAP7_75t_SL g194 ( .A(n_138), .Y(n_194) );
BUFx3_ASAP7_75t_L g491 ( .A(n_138), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g497 ( .A1(n_138), .A2(n_498), .B(n_501), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_138), .A2(n_508), .B(n_512), .Y(n_507) );
OAI21xp5_ASAP7_75t_L g528 ( .A1(n_138), .A2(n_529), .B(n_532), .Y(n_528) );
OAI21xp5_ASAP7_75t_L g537 ( .A1(n_138), .A2(n_538), .B(n_542), .Y(n_537) );
INVx5_ASAP7_75t_L g187 ( .A(n_141), .Y(n_187) );
AND2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
BUFx3_ASAP7_75t_L g152 ( .A(n_142), .Y(n_152) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_142), .Y(n_176) );
INVx1_ASAP7_75t_L g522 ( .A(n_142), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_148), .B(n_150), .Y(n_144) );
O2A1O1Ixp33_ASAP7_75t_L g203 ( .A1(n_146), .A2(n_204), .B(n_205), .C(n_206), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_146), .A2(n_484), .B(n_485), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_146), .A2(n_499), .B(n_500), .Y(n_498) );
INVx2_ASAP7_75t_L g504 ( .A(n_146), .Y(n_504) );
O2A1O1Ixp5_ASAP7_75t_SL g529 ( .A1(n_146), .A2(n_222), .B(n_530), .C(n_531), .Y(n_529) );
INVx5_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_147), .B(n_221), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_147), .B(n_241), .Y(n_240) );
OAI22xp5_ASAP7_75t_SL g556 ( .A1(n_147), .A2(n_174), .B1(n_557), .B2(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g541 ( .A(n_149), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_150), .A2(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g193 ( .A(n_152), .Y(n_193) );
INVx1_ASAP7_75t_L g267 ( .A(n_153), .Y(n_267) );
OA21x2_ASAP7_75t_L g481 ( .A1(n_153), .A2(n_482), .B(n_492), .Y(n_481) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_153), .A2(n_507), .B(n_515), .Y(n_506) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AO21x2_ASAP7_75t_L g198 ( .A1(n_154), .A2(n_199), .B(n_209), .Y(n_198) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_154), .A2(n_226), .B(n_233), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_154), .B(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_155), .Y(n_163) );
AND2x2_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
AND2x2_ASAP7_75t_SL g167 ( .A(n_156), .B(n_157), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
NOR2xp33_ASAP7_75t_SL g160 ( .A(n_161), .B(n_162), .Y(n_160) );
INVx3_ASAP7_75t_L g214 ( .A(n_162), .Y(n_214) );
AO21x1_ASAP7_75t_L g567 ( .A1(n_162), .A2(n_568), .B(n_571), .Y(n_567) );
NAND3xp33_ASAP7_75t_L g592 ( .A(n_162), .B(n_491), .C(n_568), .Y(n_592) );
INVx4_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
OA21x2_ASAP7_75t_L g235 ( .A1(n_163), .A2(n_236), .B(n_242), .Y(n_235) );
OA21x2_ASAP7_75t_L g496 ( .A1(n_163), .A2(n_497), .B(n_505), .Y(n_496) );
AND2x2_ASAP7_75t_L g322 ( .A(n_164), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g344 ( .A(n_164), .Y(n_344) );
AND2x2_ASAP7_75t_L g429 ( .A(n_164), .B(n_259), .Y(n_429) );
AND2x2_ASAP7_75t_L g432 ( .A(n_164), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g164 ( .A(n_165), .B(n_181), .Y(n_164) );
INVx2_ASAP7_75t_L g251 ( .A(n_165), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_165), .B(n_276), .Y(n_282) );
AND2x2_ASAP7_75t_L g292 ( .A(n_165), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g328 ( .A(n_165), .Y(n_328) );
AO21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_168), .B(n_178), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g180 ( .A(n_167), .Y(n_180) );
OA21x2_ASAP7_75t_L g182 ( .A1(n_167), .A2(n_183), .B(n_195), .Y(n_182) );
OA21x2_ASAP7_75t_L g527 ( .A1(n_167), .A2(n_528), .B(n_535), .Y(n_527) );
OA21x2_ASAP7_75t_L g536 ( .A1(n_167), .A2(n_537), .B(n_545), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_169), .B(n_177), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_175), .Y(n_170) );
INVx4_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g219 ( .A(n_174), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_174), .A2(n_504), .B1(n_521), .B2(n_523), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_174), .A2(n_504), .B1(n_569), .B2(n_570), .Y(n_568) );
HB1xp67_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx3_ASAP7_75t_L g222 ( .A(n_176), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_180), .B(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_180), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g270 ( .A(n_181), .B(n_251), .Y(n_270) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g252 ( .A(n_182), .Y(n_252) );
AND2x2_ASAP7_75t_L g294 ( .A(n_182), .B(n_276), .Y(n_294) );
AND2x2_ASAP7_75t_L g363 ( .A(n_182), .B(n_260), .Y(n_363) );
O2A1O1Ixp33_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_188), .C(n_194), .Y(n_185) );
O2A1O1Ixp33_ASAP7_75t_L g216 ( .A1(n_187), .A2(n_194), .B(n_217), .C(n_218), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_L g237 ( .A1(n_187), .A2(n_194), .B(n_238), .C(n_239), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_189), .B(n_192), .Y(n_191) );
INVx1_ASAP7_75t_L g511 ( .A(n_189), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_189), .A2(n_533), .B(n_534), .Y(n_532) );
INVx4_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
OAI22xp5_ASAP7_75t_SL g228 ( .A1(n_190), .A2(n_229), .B1(n_230), .B2(n_231), .Y(n_228) );
INVx2_ASAP7_75t_L g230 ( .A(n_190), .Y(n_230) );
OAI22xp33_ASAP7_75t_L g226 ( .A1(n_194), .A2(n_201), .B1(n_227), .B2(n_232), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_197), .B(n_211), .Y(n_196) );
OR2x2_ASAP7_75t_L g257 ( .A(n_197), .B(n_225), .Y(n_257) );
INVx1_ASAP7_75t_L g336 ( .A(n_197), .Y(n_336) );
AND2x2_ASAP7_75t_L g350 ( .A(n_197), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_197), .B(n_224), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_197), .B(n_348), .Y(n_402) );
AND2x2_ASAP7_75t_L g410 ( .A(n_197), .B(n_411), .Y(n_410) );
INVx3_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx3_ASAP7_75t_L g247 ( .A(n_198), .Y(n_247) );
AND2x2_ASAP7_75t_L g317 ( .A(n_198), .B(n_225), .Y(n_317) );
OAI21xp5_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B(n_202), .Y(n_199) );
OAI21xp5_ASAP7_75t_L g261 ( .A1(n_201), .A2(n_262), .B(n_263), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_206), .A2(n_509), .B(n_510), .C(n_511), .Y(n_508) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_211), .B(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g444 ( .A(n_211), .Y(n_444) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_224), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_212), .B(n_288), .Y(n_310) );
OR2x2_ASAP7_75t_L g339 ( .A(n_212), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g371 ( .A(n_212), .B(n_351), .Y(n_371) );
INVx1_ASAP7_75t_SL g391 ( .A(n_212), .Y(n_391) );
AND2x2_ASAP7_75t_L g395 ( .A(n_212), .B(n_256), .Y(n_395) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_SL g248 ( .A(n_213), .B(n_224), .Y(n_248) );
AND2x2_ASAP7_75t_L g255 ( .A(n_213), .B(n_235), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_213), .B(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g298 ( .A(n_213), .B(n_280), .Y(n_298) );
INVx1_ASAP7_75t_SL g305 ( .A(n_213), .Y(n_305) );
BUFx2_ASAP7_75t_L g316 ( .A(n_213), .Y(n_316) );
AND2x2_ASAP7_75t_L g332 ( .A(n_213), .B(n_247), .Y(n_332) );
AND2x2_ASAP7_75t_L g347 ( .A(n_213), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g411 ( .A(n_213), .B(n_225), .Y(n_411) );
OA21x2_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_223), .Y(n_213) );
O2A1O1Ixp5_ASAP7_75t_L g486 ( .A1(n_219), .A2(n_487), .B(n_488), .C(n_490), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_219), .A2(n_543), .B(n_544), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_224), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g335 ( .A(n_224), .B(n_336), .Y(n_335) );
AOI221xp5_ASAP7_75t_L g352 ( .A1(n_224), .A2(n_353), .B1(n_356), .B2(n_359), .C(n_364), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_224), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_235), .Y(n_224) );
INVx3_ASAP7_75t_L g280 ( .A(n_225), .Y(n_280) );
BUFx2_ASAP7_75t_L g290 ( .A(n_235), .Y(n_290) );
AND2x2_ASAP7_75t_L g304 ( .A(n_235), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g321 ( .A(n_235), .Y(n_321) );
OR2x2_ASAP7_75t_L g340 ( .A(n_235), .B(n_280), .Y(n_340) );
INVx3_ASAP7_75t_L g348 ( .A(n_235), .Y(n_348) );
AND2x2_ASAP7_75t_L g351 ( .A(n_235), .B(n_280), .Y(n_351) );
AOI221xp5_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_249), .B1(n_253), .B2(n_258), .C(n_271), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_248), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_246), .B(n_320), .Y(n_445) );
OR2x2_ASAP7_75t_L g448 ( .A(n_246), .B(n_279), .Y(n_448) );
INVx1_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
OAI221xp5_ASAP7_75t_SL g271 ( .A1(n_247), .A2(n_272), .B1(n_279), .B2(n_281), .C(n_284), .Y(n_271) );
AND2x2_ASAP7_75t_L g288 ( .A(n_247), .B(n_280), .Y(n_288) );
AND2x2_ASAP7_75t_L g296 ( .A(n_247), .B(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_247), .B(n_304), .Y(n_303) );
NAND2x1_ASAP7_75t_L g346 ( .A(n_247), .B(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g398 ( .A(n_247), .B(n_340), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_249), .A2(n_358), .B1(n_387), .B2(n_389), .Y(n_386) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AOI322xp5_ASAP7_75t_L g295 ( .A1(n_250), .A2(n_259), .A3(n_296), .B1(n_299), .B2(n_302), .C1(n_306), .C2(n_309), .Y(n_295) );
OR2x2_ASAP7_75t_L g307 ( .A(n_250), .B(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_251), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g286 ( .A(n_251), .B(n_260), .Y(n_286) );
INVx1_ASAP7_75t_L g301 ( .A(n_251), .Y(n_301) );
AND2x2_ASAP7_75t_L g367 ( .A(n_251), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g277 ( .A(n_252), .B(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g368 ( .A(n_252), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_252), .B(n_276), .Y(n_442) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_256), .B(n_391), .Y(n_390) );
INVx3_ASAP7_75t_SL g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g342 ( .A(n_257), .B(n_289), .Y(n_342) );
OR2x2_ASAP7_75t_L g439 ( .A(n_257), .B(n_290), .Y(n_439) );
INVx1_ASAP7_75t_L g420 ( .A(n_258), .Y(n_420) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_270), .Y(n_258) );
INVx4_ASAP7_75t_L g308 ( .A(n_259), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_259), .B(n_327), .Y(n_333) );
INVx2_ASAP7_75t_L g276 ( .A(n_260), .Y(n_276) );
AO21x2_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_267), .B(n_268), .Y(n_260) );
INVx1_ASAP7_75t_L g358 ( .A(n_270), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_270), .B(n_330), .Y(n_399) );
AOI21xp33_ASAP7_75t_L g345 ( .A1(n_272), .A2(n_346), .B(n_349), .Y(n_345) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_277), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g330 ( .A(n_276), .Y(n_330) );
INVx1_ASAP7_75t_L g357 ( .A(n_276), .Y(n_357) );
INVx1_ASAP7_75t_L g283 ( .A(n_277), .Y(n_283) );
AND2x2_ASAP7_75t_L g285 ( .A(n_277), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g381 ( .A(n_278), .B(n_367), .Y(n_381) );
AND2x2_ASAP7_75t_L g403 ( .A(n_278), .B(n_363), .Y(n_403) );
BUFx2_ASAP7_75t_L g355 ( .A(n_280), .Y(n_355) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AOI32xp33_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_287), .A3(n_288), .B1(n_289), .B2(n_291), .Y(n_284) );
INVx1_ASAP7_75t_L g365 ( .A(n_285), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_285), .A2(n_413), .B1(n_414), .B2(n_416), .Y(n_412) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_288), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_288), .B(n_347), .Y(n_388) );
AND2x2_ASAP7_75t_L g435 ( .A(n_288), .B(n_320), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_289), .B(n_336), .Y(n_383) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g436 ( .A(n_291), .Y(n_436) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
INVx1_ASAP7_75t_L g361 ( .A(n_292), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_294), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g408 ( .A(n_294), .B(n_328), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_294), .B(n_323), .Y(n_415) );
INVx1_ASAP7_75t_SL g397 ( .A(n_296), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_297), .B(n_348), .Y(n_375) );
NOR4xp25_ASAP7_75t_L g421 ( .A(n_297), .B(n_320), .C(n_422), .D(n_425), .Y(n_421) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_298), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVxp67_ASAP7_75t_L g378 ( .A(n_301), .Y(n_378) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OAI21xp33_ASAP7_75t_L g428 ( .A1(n_304), .A2(n_395), .B(n_429), .Y(n_428) );
AND2x4_ASAP7_75t_L g320 ( .A(n_305), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g369 ( .A(n_308), .Y(n_369) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND4xp25_ASAP7_75t_SL g311 ( .A(n_312), .B(n_337), .C(n_352), .D(n_372), .Y(n_311) );
O2A1O1Ixp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_318), .B(n_322), .C(n_324), .Y(n_312) );
INVx1_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g404 ( .A(n_317), .B(n_347), .Y(n_404) );
AND2x2_ASAP7_75t_L g413 ( .A(n_317), .B(n_391), .Y(n_413) );
INVx3_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_320), .B(n_355), .Y(n_417) );
AND2x2_ASAP7_75t_L g329 ( .A(n_323), .B(n_330), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_331), .B1(n_333), .B2(n_334), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
AND2x2_ASAP7_75t_L g427 ( .A(n_327), .B(n_373), .Y(n_427) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_329), .B(n_378), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_330), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
O2A1O1Ixp33_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_341), .B(n_343), .C(n_345), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g372 ( .A1(n_338), .A2(n_373), .B1(n_374), .B2(n_376), .C(n_379), .Y(n_372) );
INVx1_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OAI221xp5_ASAP7_75t_L g430 ( .A1(n_346), .A2(n_431), .B1(n_434), .B2(n_436), .C(n_437), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_347), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_355), .B(n_424), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
INVx1_ASAP7_75t_L g385 ( .A(n_357), .Y(n_385) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_360), .A2(n_380), .B1(n_382), .B2(n_383), .Y(n_379) );
OR2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AOI21xp33_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_366), .B(n_370), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_369), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_369), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OAI221xp5_ASAP7_75t_L g443 ( .A1(n_380), .A2(n_406), .B1(n_444), .B2(n_445), .C(n_446), .Y(n_443) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g425 ( .A(n_382), .Y(n_425) );
OAI211xp5_ASAP7_75t_SL g384 ( .A1(n_385), .A2(n_386), .B(n_392), .C(n_412), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI211xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_395), .B(n_396), .C(n_405), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
A2O1A1Ixp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B(n_399), .C(n_400), .Y(n_396) );
INVx1_ASAP7_75t_L g424 ( .A(n_402), .Y(n_424) );
OAI21xp5_ASAP7_75t_SL g446 ( .A1(n_403), .A2(n_429), .B(n_447), .Y(n_446) );
AOI21xp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_407), .B(n_409), .Y(n_405) );
INVx1_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVxp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OAI21xp5_ASAP7_75t_SL g438 ( .A1(n_415), .A2(n_439), .B(n_440), .Y(n_438) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NOR3xp33_ASAP7_75t_L g418 ( .A(n_419), .B(n_430), .C(n_443), .Y(n_418) );
OAI211xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B(n_426), .C(n_428), .Y(n_419) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
CKINVDCx14_ASAP7_75t_R g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx2_ASAP7_75t_L g462 ( .A(n_455), .Y(n_462) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_455), .Y(n_465) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
NAND3xp33_ASAP7_75t_L g466 ( .A(n_463), .B(n_467), .C(n_762), .Y(n_466) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g761 ( .A(n_475), .Y(n_761) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OR3x1_ASAP7_75t_L g476 ( .A(n_477), .B(n_678), .C(n_727), .Y(n_476) );
NAND5xp2_ASAP7_75t_L g477 ( .A(n_478), .B(n_593), .C(n_621), .D(n_651), .E(n_665), .Y(n_477) );
AOI221xp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_516), .B1(n_546), .B2(n_551), .C(n_560), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_480), .B(n_493), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_480), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g573 ( .A(n_481), .Y(n_573) );
AND2x2_ASAP7_75t_L g581 ( .A(n_481), .B(n_496), .Y(n_581) );
AND2x2_ASAP7_75t_L g604 ( .A(n_481), .B(n_495), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_481), .B(n_506), .Y(n_619) );
OR2x2_ASAP7_75t_L g628 ( .A(n_481), .B(n_567), .Y(n_628) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_481), .Y(n_631) );
AND2x2_ASAP7_75t_L g739 ( .A(n_481), .B(n_567), .Y(n_739) );
OAI21xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_486), .B(n_491), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g512 ( .A1(n_488), .A2(n_504), .B(n_513), .C(n_514), .Y(n_512) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_493), .B(n_631), .Y(n_687) );
INVx2_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
OAI311xp33_ASAP7_75t_L g629 ( .A1(n_494), .A2(n_630), .A3(n_631), .B1(n_632), .C1(n_647), .Y(n_629) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_506), .Y(n_494) );
AND2x2_ASAP7_75t_L g590 ( .A(n_495), .B(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g597 ( .A(n_495), .Y(n_597) );
AND2x2_ASAP7_75t_L g718 ( .A(n_495), .B(n_550), .Y(n_718) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_496), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g574 ( .A(n_496), .B(n_506), .Y(n_574) );
AND2x2_ASAP7_75t_L g626 ( .A(n_496), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g640 ( .A(n_496), .B(n_573), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_503), .B(n_504), .Y(n_501) );
INVx2_ASAP7_75t_L g550 ( .A(n_506), .Y(n_550) );
AND2x2_ASAP7_75t_L g589 ( .A(n_506), .B(n_573), .Y(n_589) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_524), .Y(n_516) );
OR2x2_ASAP7_75t_L g684 ( .A(n_517), .B(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_517), .B(n_690), .Y(n_701) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_518), .B(n_697), .Y(n_696) );
BUFx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g559 ( .A(n_519), .Y(n_559) );
AND2x2_ASAP7_75t_L g625 ( .A(n_519), .B(n_555), .Y(n_625) );
AND2x2_ASAP7_75t_L g636 ( .A(n_519), .B(n_536), .Y(n_636) );
AND2x2_ASAP7_75t_L g645 ( .A(n_519), .B(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_524), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_524), .B(n_586), .Y(n_630) );
INVx2_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
OR2x2_ASAP7_75t_L g617 ( .A(n_525), .B(n_576), .Y(n_617) );
OR2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_536), .Y(n_525) );
INVx2_ASAP7_75t_L g553 ( .A(n_526), .Y(n_553) );
AND2x2_ASAP7_75t_L g644 ( .A(n_526), .B(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g563 ( .A(n_527), .Y(n_563) );
OR2x2_ASAP7_75t_L g661 ( .A(n_527), .B(n_662), .Y(n_661) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_527), .Y(n_724) );
AND2x2_ASAP7_75t_L g564 ( .A(n_536), .B(n_559), .Y(n_564) );
INVx1_ASAP7_75t_L g584 ( .A(n_536), .Y(n_584) );
AND2x2_ASAP7_75t_L g605 ( .A(n_536), .B(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g646 ( .A(n_536), .Y(n_646) );
INVx1_ASAP7_75t_L g662 ( .A(n_536), .Y(n_662) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_536), .Y(n_737) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_540), .B(n_541), .Y(n_538) );
INVxp67_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_548), .B(n_650), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_548), .A2(n_635), .B1(n_684), .B2(n_694), .Y(n_693) );
INVx1_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
OAI211xp5_ASAP7_75t_SL g727 ( .A1(n_549), .A2(n_728), .B(n_730), .C(n_748), .Y(n_727) );
INVx2_ASAP7_75t_L g580 ( .A(n_550), .Y(n_580) );
AND2x2_ASAP7_75t_L g638 ( .A(n_550), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g649 ( .A(n_550), .B(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_551), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_554), .Y(n_551) );
AND2x2_ASAP7_75t_L g622 ( .A(n_552), .B(n_586), .Y(n_622) );
BUFx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g654 ( .A(n_553), .B(n_645), .Y(n_654) );
AND2x2_ASAP7_75t_L g673 ( .A(n_553), .B(n_587), .Y(n_673) );
AND2x4_ASAP7_75t_L g609 ( .A(n_554), .B(n_583), .Y(n_609) );
AND2x2_ASAP7_75t_L g747 ( .A(n_554), .B(n_723), .Y(n_747) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_559), .Y(n_554) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_555), .Y(n_576) );
INVx1_ASAP7_75t_L g587 ( .A(n_555), .Y(n_587) );
INVx1_ASAP7_75t_L g686 ( .A(n_555), .Y(n_686) );
OR2x2_ASAP7_75t_L g577 ( .A(n_559), .B(n_563), .Y(n_577) );
AND2x2_ASAP7_75t_L g586 ( .A(n_559), .B(n_587), .Y(n_586) );
NOR2xp67_ASAP7_75t_L g606 ( .A(n_559), .B(n_607), .Y(n_606) );
OAI221xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_565), .B1(n_575), .B2(n_578), .C(n_582), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
A2O1A1Ixp33_ASAP7_75t_L g582 ( .A1(n_562), .A2(n_583), .B(n_585), .C(n_588), .Y(n_582) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
INVx1_ASAP7_75t_L g607 ( .A(n_563), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_563), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_SL g690 ( .A(n_563), .B(n_584), .Y(n_690) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_563), .Y(n_697) );
AND2x2_ASAP7_75t_L g615 ( .A(n_564), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g652 ( .A(n_564), .B(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_574), .Y(n_565) );
INVx2_ASAP7_75t_L g643 ( .A(n_566), .Y(n_643) );
AOI222xp33_ASAP7_75t_L g692 ( .A1(n_566), .A2(n_576), .B1(n_693), .B2(n_695), .C1(n_696), .C2(n_698), .Y(n_692) );
AND2x2_ASAP7_75t_L g749 ( .A(n_566), .B(n_718), .Y(n_749) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_573), .Y(n_566) );
INVx1_ASAP7_75t_L g639 ( .A(n_567), .Y(n_639) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x4_ASAP7_75t_L g591 ( .A(n_572), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g677 ( .A(n_574), .B(n_611), .Y(n_677) );
AOI21xp33_ASAP7_75t_L g688 ( .A1(n_575), .A2(n_689), .B(n_691), .Y(n_688) );
OR2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
INVx2_ASAP7_75t_L g616 ( .A(n_576), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_576), .B(n_583), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_576), .B(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
INVx3_ASAP7_75t_L g642 ( .A(n_580), .Y(n_642) );
OR2x2_ASAP7_75t_L g694 ( .A(n_580), .B(n_616), .Y(n_694) );
AND2x2_ASAP7_75t_L g610 ( .A(n_581), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g648 ( .A(n_581), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_581), .B(n_642), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_581), .B(n_638), .Y(n_664) );
AND2x2_ASAP7_75t_L g668 ( .A(n_581), .B(n_650), .Y(n_668) );
INVxp67_ASAP7_75t_L g600 ( .A(n_583), .Y(n_600) );
BUFx3_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_585), .A2(n_658), .B1(n_663), .B2(n_664), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_585), .B(n_690), .Y(n_720) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g706 ( .A(n_586), .B(n_697), .Y(n_706) );
AND2x2_ASAP7_75t_L g735 ( .A(n_586), .B(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g740 ( .A(n_586), .B(n_690), .Y(n_740) );
INVx1_ASAP7_75t_L g653 ( .A(n_587), .Y(n_653) );
BUFx2_ASAP7_75t_L g659 ( .A(n_587), .Y(n_659) );
INVx1_ASAP7_75t_L g744 ( .A(n_588), .Y(n_744) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
NAND2x1p5_ASAP7_75t_L g595 ( .A(n_589), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g620 ( .A(n_590), .Y(n_620) );
NOR2x1_ASAP7_75t_L g596 ( .A(n_591), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g603 ( .A(n_591), .B(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g612 ( .A(n_591), .Y(n_612) );
INVx3_ASAP7_75t_L g650 ( .A(n_591), .Y(n_650) );
OR2x2_ASAP7_75t_L g716 ( .A(n_591), .B(n_717), .Y(n_716) );
AOI211xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_598), .B(n_601), .C(n_613), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g730 ( .A1(n_594), .A2(n_731), .B1(n_738), .B2(n_740), .C(n_741), .Y(n_730) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_602), .B(n_608), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_605), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_604), .B(n_642), .Y(n_656) );
AND2x2_ASAP7_75t_L g698 ( .A(n_604), .B(n_638), .Y(n_698) );
INVx1_ASAP7_75t_SL g711 ( .A(n_605), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_605), .B(n_659), .Y(n_714) );
INVx1_ASAP7_75t_L g732 ( .A(n_606), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_610), .A2(n_700), .B1(n_702), .B2(n_706), .C(n_707), .Y(n_699) );
AND2x2_ASAP7_75t_L g726 ( .A(n_611), .B(n_718), .Y(n_726) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g710 ( .A(n_612), .Y(n_710) );
AOI21xp33_ASAP7_75t_SL g613 ( .A1(n_614), .A2(n_617), .B(n_618), .Y(n_613) );
INVx1_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
OR2x2_ASAP7_75t_L g681 ( .A(n_616), .B(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g667 ( .A(n_617), .Y(n_667) );
INVx1_ASAP7_75t_L g695 ( .A(n_618), .Y(n_695) );
OR2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
O2A1O1Ixp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_623), .B(n_626), .C(n_629), .Y(n_621) );
OAI31xp33_ASAP7_75t_L g748 ( .A1(n_622), .A2(n_660), .A3(n_747), .B(n_749), .Y(n_748) );
INVxp67_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g722 ( .A(n_625), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_SL g743 ( .A(n_625), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_627), .B(n_642), .Y(n_670) );
INVx1_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g745 ( .A(n_628), .B(n_642), .Y(n_745) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_637), .B1(n_641), .B2(n_644), .Y(n_632) );
NAND2xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_636), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g672 ( .A(n_636), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g675 ( .A(n_636), .B(n_659), .Y(n_675) );
AND2x2_ASAP7_75t_L g729 ( .A(n_636), .B(n_724), .Y(n_729) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
INVx1_ASAP7_75t_L g704 ( .A(n_640), .Y(n_704) );
NOR2xp67_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
OAI32xp33_ASAP7_75t_L g707 ( .A1(n_642), .A2(n_676), .A3(n_708), .B1(n_710), .B2(n_711), .Y(n_707) );
INVx1_ASAP7_75t_L g682 ( .A(n_645), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_645), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g705 ( .A(n_649), .Y(n_705) );
O2A1O1Ixp33_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_654), .B(n_655), .C(n_657), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_653), .B(n_690), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_654), .A2(n_666), .B1(n_667), .B2(n_668), .C(n_669), .Y(n_665) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g666 ( .A(n_664), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_671), .B1(n_674), .B2(n_676), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND4xp25_ASAP7_75t_SL g731 ( .A(n_674), .B(n_732), .C(n_733), .D(n_734), .Y(n_731) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
NAND4xp25_ASAP7_75t_SL g678 ( .A(n_679), .B(n_692), .C(n_699), .D(n_712), .Y(n_678) );
O2A1O1Ixp33_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_683), .B(n_687), .C(n_688), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_SL g709 ( .A(n_685), .Y(n_709) );
INVx2_ASAP7_75t_L g733 ( .A(n_690), .Y(n_733) );
OR2x2_ASAP7_75t_L g742 ( .A(n_697), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
OR2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_715), .B(n_719), .Y(n_712) );
INVxp67_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g738 ( .A(n_718), .B(n_739), .Y(n_738) );
AOI21xp33_ASAP7_75t_SL g719 ( .A1(n_720), .A2(n_721), .B(n_725), .Y(n_719) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
CKINVDCx16_ASAP7_75t_R g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_744), .B1(n_745), .B2(n_746), .Y(n_741) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
endmodule