module fake_jpeg_2367_n_221 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_221);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_221;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_1),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_13),
.B(n_19),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_27),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_51),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_5),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_3),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_23),
.B(n_37),
.Y(n_75)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_11),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_84),
.Y(n_94)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_0),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_85),
.B(n_68),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_86),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_79),
.A2(n_74),
.B1(n_69),
.B2(n_63),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_71),
.B1(n_64),
.B2(n_77),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_74),
.B1(n_63),
.B2(n_67),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_90),
.A2(n_63),
.B1(n_77),
.B2(n_78),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_98),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_53),
.B(n_56),
.C(n_72),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_66),
.B(n_58),
.C(n_67),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_65),
.B1(n_57),
.B2(n_61),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_66),
.B1(n_55),
.B2(n_58),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_101),
.Y(n_135)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_112),
.B1(n_114),
.B2(n_94),
.Y(n_121)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_83),
.B1(n_69),
.B2(n_76),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_115),
.B1(n_92),
.B2(n_64),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_54),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_108),
.Y(n_126)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_107),
.A2(n_118),
.B1(n_64),
.B2(n_78),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_57),
.Y(n_108)
);

NOR2x1_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_0),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_89),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_113),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_91),
.A2(n_76),
.B1(n_59),
.B2(n_70),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_89),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_91),
.A2(n_97),
.B1(n_88),
.B2(n_95),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_109),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_100),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_134),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_120),
.A2(n_125),
.B1(n_136),
.B2(n_10),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_SL g162 ( 
.A1(n_121),
.A2(n_133),
.B(n_138),
.Y(n_162)
);

AND2x6_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_24),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_123),
.Y(n_147)
);

AND2x6_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_38),
.Y(n_123)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_124),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_115),
.A2(n_92),
.B1(n_94),
.B2(n_65),
.Y(n_125)
);

XOR2x2_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_61),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_132),
.C(n_101),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_135),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_75),
.C(n_64),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_117),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_4),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_140),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_101),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_6),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_109),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_149),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_155),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_107),
.B1(n_8),
.B2(n_9),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_143),
.A2(n_144),
.B1(n_17),
.B2(n_18),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_129),
.A2(n_139),
.B1(n_135),
.B2(n_131),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_52),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_163),
.C(n_19),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_7),
.B(n_9),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_151),
.B(n_145),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_134),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_130),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_150),
.B(n_154),
.Y(n_174)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_49),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_157),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_124),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_131),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_123),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_L g182 ( 
.A1(n_158),
.A2(n_159),
.B(n_20),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_12),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

FAx1_ASAP7_75t_SL g161 ( 
.A(n_119),
.B(n_14),
.CI(n_15),
.CON(n_161),
.SN(n_161)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_16),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_26),
.C(n_43),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_149),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_168),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_167),
.A2(n_182),
.B(n_146),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_156),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_141),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_169),
.B(n_178),
.Y(n_190)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_173),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_181),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_33),
.C(n_42),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_163),
.C(n_153),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_152),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

HAxp5_ASAP7_75t_SL g184 ( 
.A(n_165),
.B(n_161),
.CON(n_184),
.SN(n_184)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_193),
.Y(n_196)
);

AND2x2_ASAP7_75t_SL g191 ( 
.A(n_171),
.B(n_162),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_191),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_147),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_179),
.Y(n_201)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_192),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_195),
.B(n_198),
.Y(n_205)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_186),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_189),
.A2(n_165),
.B1(n_170),
.B2(n_167),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_200),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_188),
.A2(n_172),
.B1(n_174),
.B2(n_176),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_166),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_188),
.A2(n_173),
.B1(n_171),
.B2(n_180),
.Y(n_203)
);

OAI321xp33_ASAP7_75t_L g206 ( 
.A1(n_203),
.A2(n_191),
.A3(n_190),
.B1(n_172),
.B2(n_183),
.C(n_194),
.Y(n_206)
);

A2O1A1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_202),
.A2(n_184),
.B(n_191),
.C(n_185),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_197),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_206),
.A2(n_197),
.B1(n_203),
.B2(n_161),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_193),
.C(n_178),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_208),
.C(n_201),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_211),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_204),
.C(n_209),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_214),
.A2(n_212),
.B(n_205),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_215),
.A2(n_213),
.B(n_34),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_32),
.Y(n_217)
);

AOI322xp5_ASAP7_75t_L g218 ( 
.A1(n_217),
.A2(n_25),
.A3(n_45),
.B1(n_40),
.B2(n_36),
.C1(n_157),
.C2(n_22),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_20),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_21),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_21),
.Y(n_221)
);


endmodule