module fake_ariane_2229_n_1876 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1876);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1876;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_604;
wire n_439;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_106),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_80),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_152),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_13),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_66),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_107),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_30),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_93),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_6),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_69),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_25),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_165),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_96),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_22),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_15),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_19),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_132),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_137),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_5),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_73),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_43),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_26),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_50),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_64),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_99),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_65),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_122),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_23),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_117),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_87),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_92),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_102),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_28),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_155),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_101),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_149),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_35),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_109),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_163),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_118),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_108),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_60),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_110),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_81),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_34),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_60),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_11),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_136),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_66),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_50),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_140),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_148),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_54),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_166),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_95),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_5),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_39),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_159),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_131),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_168),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_76),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_104),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_39),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_34),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_133),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_30),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_170),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_28),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_115),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_126),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_6),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_55),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_150),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_121),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_1),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_164),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_68),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_63),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_83),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_74),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_20),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_82),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_145),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_49),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_20),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_120),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_26),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_29),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_157),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_57),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_97),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_38),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_127),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_61),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_7),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_10),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_141),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_139),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_19),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_3),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_33),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_18),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_169),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_45),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_54),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_23),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_32),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_144),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_63),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_113),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_143),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_160),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_103),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_9),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_128),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_94),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_72),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_162),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_0),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_146),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_1),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_13),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_114),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_125),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_130),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_11),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_58),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_112),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_25),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_37),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_70),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_27),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_22),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_55),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_42),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_85),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_138),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_129),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_119),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_147),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_135),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_14),
.Y(n_312)
);

BUFx2_ASAP7_75t_SL g313 ( 
.A(n_61),
.Y(n_313)
);

BUFx5_ASAP7_75t_L g314 ( 
.A(n_36),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_88),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_111),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_49),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_18),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_40),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_58),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_142),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_56),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_77),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_46),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_79),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_16),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_56),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_37),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_84),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_4),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_86),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_98),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_90),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_31),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_47),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_32),
.Y(n_336)
);

BUFx10_ASAP7_75t_L g337 ( 
.A(n_15),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_2),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_153),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_62),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_184),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_277),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_171),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_184),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_225),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_214),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_268),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_280),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_184),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_184),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_184),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_184),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_184),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_192),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_219),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_220),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_184),
.B(n_314),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_314),
.B(n_0),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_226),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_314),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_314),
.Y(n_361)
);

NAND2xp33_ASAP7_75t_R g362 ( 
.A(n_183),
.B(n_123),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_198),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_227),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_242),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_257),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_314),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_203),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_320),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_314),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_314),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_206),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_206),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_314),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_255),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_174),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_262),
.Y(n_377)
);

NOR2xp67_ASAP7_75t_L g378 ( 
.A(n_245),
.B(n_2),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_337),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_175),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_213),
.B(n_3),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_174),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_337),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_276),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_175),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_175),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_175),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_301),
.B(n_245),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_175),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_337),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_177),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_181),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_181),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_181),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_181),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_181),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_233),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_233),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_233),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_233),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g401 ( 
.A(n_179),
.B(n_4),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_177),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_301),
.B(n_7),
.Y(n_403)
);

NOR2xp67_ASAP7_75t_L g404 ( 
.A(n_301),
.B(n_8),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_191),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_233),
.Y(n_406)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_276),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_238),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_191),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_238),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_238),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_193),
.Y(n_412)
);

INVxp33_ASAP7_75t_L g413 ( 
.A(n_185),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_193),
.Y(n_414)
);

INVxp33_ASAP7_75t_SL g415 ( 
.A(n_264),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_264),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_238),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_238),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_172),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_R g420 ( 
.A(n_221),
.B(n_167),
.Y(n_420)
);

NOR2xp67_ASAP7_75t_L g421 ( 
.A(n_217),
.B(n_8),
.Y(n_421)
);

NOR2xp67_ASAP7_75t_L g422 ( 
.A(n_179),
.B(n_9),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_300),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_347),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_357),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_344),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_388),
.B(n_187),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_344),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_419),
.B(n_340),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_344),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_354),
.A2(n_284),
.B1(n_266),
.B2(n_271),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_384),
.B(n_283),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_341),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_419),
.B(n_195),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_419),
.B(n_189),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_413),
.B(n_189),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_350),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_350),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_350),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_341),
.B(n_200),
.Y(n_440)
);

OAI21x1_ASAP7_75t_L g441 ( 
.A1(n_367),
.A2(n_273),
.B(n_190),
.Y(n_441)
);

INVx6_ASAP7_75t_L g442 ( 
.A(n_401),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_367),
.Y(n_443)
);

NOR2x1_ASAP7_75t_L g444 ( 
.A(n_381),
.B(n_230),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_349),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_349),
.B(n_205),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_351),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_404),
.B(n_196),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_351),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_367),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_402),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_352),
.B(n_208),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_394),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_352),
.Y(n_454)
);

OA21x2_ASAP7_75t_L g455 ( 
.A1(n_358),
.A2(n_273),
.B(n_190),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_353),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_407),
.B(n_196),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_353),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_360),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_360),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_361),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_361),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_343),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_370),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_404),
.B(n_216),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_370),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_345),
.B(n_216),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_345),
.B(n_270),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_371),
.Y(n_469)
);

CKINVDCx6p67_ASAP7_75t_R g470 ( 
.A(n_379),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_371),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_374),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_374),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_380),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_394),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_405),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_394),
.Y(n_477)
);

BUFx8_ASAP7_75t_L g478 ( 
.A(n_401),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_395),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_377),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_395),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_395),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_380),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_385),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_403),
.B(n_385),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_363),
.B(n_266),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_386),
.Y(n_487)
);

BUFx8_ASAP7_75t_L g488 ( 
.A(n_379),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_396),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_386),
.B(n_211),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_376),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_387),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_387),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_389),
.B(n_392),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_375),
.B(n_340),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_389),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_422),
.B(n_270),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_392),
.B(n_296),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_393),
.B(n_237),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_428),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_458),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_456),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_436),
.B(n_382),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_442),
.B(n_415),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_478),
.A2(n_378),
.B1(n_422),
.B2(n_391),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_428),
.Y(n_506)
);

AND2x6_ASAP7_75t_L g507 ( 
.A(n_425),
.B(n_315),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_444),
.B(n_355),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_442),
.B(n_356),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_428),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_425),
.B(n_359),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_430),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_433),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_444),
.B(n_364),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_432),
.B(n_365),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_430),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_436),
.B(n_412),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_463),
.Y(n_518)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_426),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_458),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_442),
.B(n_366),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_467),
.B(n_369),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_432),
.B(n_416),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_426),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_458),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_458),
.Y(n_526)
);

NAND2xp33_ASAP7_75t_SL g527 ( 
.A(n_491),
.B(n_362),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_480),
.B(n_342),
.Y(n_528)
);

AO21x2_ASAP7_75t_L g529 ( 
.A1(n_441),
.A2(n_243),
.B(n_240),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_436),
.B(n_378),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_430),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_426),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_460),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_460),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_443),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_456),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_478),
.A2(n_448),
.B1(n_465),
.B2(n_442),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_443),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_467),
.B(n_468),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_443),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_438),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_460),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_460),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_467),
.B(n_372),
.Y(n_544)
);

NOR3xp33_ASAP7_75t_L g545 ( 
.A(n_431),
.B(n_421),
.C(n_269),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_478),
.A2(n_421),
.B1(n_373),
.B2(n_296),
.Y(n_546)
);

BUFx4f_ASAP7_75t_L g547 ( 
.A(n_455),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_456),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_438),
.Y(n_549)
);

OAI22xp33_ASAP7_75t_SL g550 ( 
.A1(n_442),
.A2(n_299),
.B1(n_275),
.B2(n_274),
.Y(n_550)
);

NAND2xp33_ASAP7_75t_R g551 ( 
.A(n_424),
.B(n_346),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_442),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_438),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_478),
.A2(n_251),
.B1(n_194),
.B2(n_248),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_468),
.B(n_173),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_438),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_426),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_427),
.B(n_393),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_470),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_474),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_427),
.B(n_398),
.Y(n_561)
);

OR2x6_ASAP7_75t_L g562 ( 
.A(n_448),
.B(n_313),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_488),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_468),
.B(n_409),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_478),
.B(n_173),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_426),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_474),
.Y(n_567)
);

AND2x2_ASAP7_75t_SL g568 ( 
.A(n_455),
.B(n_315),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_456),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_485),
.B(n_398),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_491),
.B(n_176),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_483),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_483),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_448),
.B(n_176),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_485),
.B(n_399),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_431),
.A2(n_414),
.B1(n_284),
.B2(n_299),
.Y(n_576)
);

INVx5_ASAP7_75t_L g577 ( 
.A(n_461),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_426),
.Y(n_578)
);

BUFx4f_ASAP7_75t_L g579 ( 
.A(n_455),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_448),
.B(n_178),
.Y(n_580)
);

INVx4_ASAP7_75t_L g581 ( 
.A(n_461),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_457),
.Y(n_582)
);

INVx6_ASAP7_75t_L g583 ( 
.A(n_461),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_434),
.B(n_383),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_433),
.B(n_445),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_451),
.Y(n_586)
);

INVx4_ASAP7_75t_L g587 ( 
.A(n_461),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_470),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_448),
.B(n_178),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_457),
.B(n_429),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_484),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_434),
.B(n_445),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_465),
.B(n_180),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_465),
.A2(n_215),
.B1(n_212),
.B2(n_223),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_480),
.B(n_271),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_484),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_487),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_487),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_456),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_461),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_492),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_426),
.Y(n_602)
);

NAND3xp33_ASAP7_75t_L g603 ( 
.A(n_447),
.B(n_300),
.C(n_423),
.Y(n_603)
);

BUFx10_ASAP7_75t_L g604 ( 
.A(n_465),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_426),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_492),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_465),
.B(n_457),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_461),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_493),
.Y(n_609)
);

BUFx10_ASAP7_75t_L g610 ( 
.A(n_429),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_461),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_488),
.B(n_180),
.Y(n_612)
);

OR2x6_ASAP7_75t_L g613 ( 
.A(n_497),
.B(n_283),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_447),
.B(n_399),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_493),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_449),
.B(n_390),
.Y(n_616)
);

AND2x6_ASAP7_75t_L g617 ( 
.A(n_429),
.B(n_222),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_488),
.Y(n_618)
);

NAND2xp33_ASAP7_75t_R g619 ( 
.A(n_451),
.B(n_348),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_449),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_461),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_454),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_429),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_429),
.B(n_186),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_454),
.B(n_400),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_459),
.B(n_400),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_459),
.B(n_406),
.Y(n_627)
);

AND2x6_ASAP7_75t_L g628 ( 
.A(n_435),
.B(n_222),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_462),
.B(n_406),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_462),
.B(n_408),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_488),
.B(n_182),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_437),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_437),
.Y(n_633)
);

NAND3xp33_ASAP7_75t_L g634 ( 
.A(n_464),
.B(n_300),
.C(n_423),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_437),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_496),
.Y(n_636)
);

AND2x6_ASAP7_75t_L g637 ( 
.A(n_435),
.B(n_222),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_435),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_496),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_464),
.B(n_408),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_466),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_435),
.B(n_207),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_437),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_437),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_466),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_497),
.A2(n_326),
.B1(n_234),
.B2(n_236),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_437),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_471),
.B(n_410),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_471),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_435),
.B(n_241),
.Y(n_650)
);

INVx1_ASAP7_75t_SL g651 ( 
.A(n_451),
.Y(n_651)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_476),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_509),
.B(n_488),
.Y(n_653)
);

INVx5_ASAP7_75t_L g654 ( 
.A(n_524),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_521),
.B(n_473),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_504),
.B(n_473),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_513),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_584),
.B(n_470),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_500),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_592),
.B(n_497),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_500),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_506),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_641),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_519),
.A2(n_446),
.B(n_440),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_527),
.B(n_476),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_607),
.A2(n_497),
.B1(n_455),
.B2(n_452),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_530),
.B(n_497),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_515),
.B(n_476),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_506),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_511),
.B(n_440),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_523),
.B(n_446),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_530),
.B(n_452),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_641),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_552),
.B(n_182),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_510),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_616),
.B(n_368),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_582),
.B(n_498),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_552),
.B(n_188),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_582),
.B(n_498),
.Y(n_679)
);

INVxp67_ASAP7_75t_L g680 ( 
.A(n_564),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_SL g681 ( 
.A(n_563),
.B(n_495),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_604),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_503),
.B(n_188),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_645),
.Y(n_684)
);

OAI22xp5_ASAP7_75t_L g685 ( 
.A1(n_513),
.A2(n_272),
.B1(n_304),
.B2(n_302),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_503),
.B(n_197),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_522),
.B(n_495),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_607),
.B(n_498),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_607),
.A2(n_455),
.B1(n_495),
.B2(n_490),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_528),
.B(n_486),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_607),
.B(n_455),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_604),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_623),
.B(n_469),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_623),
.B(n_469),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_645),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_517),
.B(n_197),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_528),
.B(n_486),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_510),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_638),
.B(n_469),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_517),
.B(n_199),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_508),
.B(n_486),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_649),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_514),
.B(n_272),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_638),
.B(n_469),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_590),
.B(n_469),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_604),
.B(n_199),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_649),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_590),
.B(n_469),
.Y(n_708)
);

INVxp67_ASAP7_75t_SL g709 ( 
.A(n_620),
.Y(n_709)
);

NOR3xp33_ASAP7_75t_L g710 ( 
.A(n_571),
.B(n_258),
.C(n_254),
.Y(n_710)
);

INVxp67_ASAP7_75t_R g711 ( 
.A(n_652),
.Y(n_711)
);

NOR2xp67_ASAP7_75t_L g712 ( 
.A(n_502),
.B(n_490),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_620),
.B(n_469),
.Y(n_713)
);

NOR3xp33_ASAP7_75t_L g714 ( 
.A(n_550),
.B(n_265),
.C(n_260),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_560),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_560),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_622),
.B(n_469),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_567),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_507),
.A2(n_274),
.B1(n_336),
.B2(n_334),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_622),
.B(n_472),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_512),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_567),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_502),
.B(n_472),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_512),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_604),
.B(n_201),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_610),
.B(n_201),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_524),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_651),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_507),
.A2(n_275),
.B1(n_336),
.B2(n_334),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_516),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_568),
.A2(n_499),
.B1(n_300),
.B2(n_450),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_SL g732 ( 
.A1(n_518),
.A2(n_327),
.B1(n_289),
.B2(n_317),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_572),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_572),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_573),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_524),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_610),
.B(n_202),
.Y(n_737)
);

NAND2xp33_ASAP7_75t_L g738 ( 
.A(n_507),
.B(n_472),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_539),
.B(n_289),
.Y(n_739)
);

NOR3xp33_ASAP7_75t_L g740 ( 
.A(n_550),
.B(n_291),
.C(n_279),
.Y(n_740)
);

INVx2_ASAP7_75t_SL g741 ( 
.A(n_610),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_544),
.B(n_555),
.Y(n_742)
);

AOI221xp5_ASAP7_75t_L g743 ( 
.A1(n_576),
.A2(n_302),
.B1(n_292),
.B2(n_312),
.C(n_317),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_502),
.B(n_472),
.Y(n_744)
);

O2A1O1Ixp5_ASAP7_75t_L g745 ( 
.A1(n_547),
.A2(n_499),
.B(n_249),
.C(n_316),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_574),
.B(n_292),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_536),
.B(n_472),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_610),
.B(n_202),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_536),
.B(n_472),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_516),
.Y(n_750)
);

OR2x2_ASAP7_75t_L g751 ( 
.A(n_651),
.B(n_304),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_562),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_531),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_536),
.B(n_472),
.Y(n_754)
);

AND2x4_ASAP7_75t_SL g755 ( 
.A(n_559),
.B(n_297),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_531),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_580),
.B(n_312),
.Y(n_757)
);

A2O1A1Ixp33_ASAP7_75t_L g758 ( 
.A1(n_548),
.A2(n_441),
.B(n_303),
.C(n_305),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_535),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_537),
.B(n_505),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_535),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_548),
.B(n_472),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_538),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_573),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_591),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_554),
.B(n_204),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_589),
.B(n_327),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_538),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_548),
.B(n_437),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_569),
.B(n_437),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_569),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_524),
.Y(n_772)
);

O2A1O1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_585),
.A2(n_338),
.B(n_319),
.C(n_322),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_546),
.B(n_204),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_569),
.B(n_599),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_599),
.B(n_439),
.Y(n_776)
);

NOR3xp33_ASAP7_75t_L g777 ( 
.A(n_576),
.B(n_335),
.C(n_328),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_540),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_593),
.B(n_253),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_618),
.B(n_209),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_540),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_599),
.B(n_439),
.Y(n_782)
);

AND2x6_ASAP7_75t_SL g783 ( 
.A(n_562),
.B(n_318),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_558),
.B(n_561),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_501),
.B(n_439),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_541),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_524),
.Y(n_787)
);

NOR3xp33_ASAP7_75t_L g788 ( 
.A(n_545),
.B(n_330),
.C(n_324),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_501),
.B(n_439),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_541),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_568),
.A2(n_300),
.B1(n_439),
.B2(n_450),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_591),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_596),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_596),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_520),
.B(n_439),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_568),
.A2(n_450),
.B1(n_439),
.B2(n_331),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_520),
.B(n_525),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_525),
.B(n_439),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_562),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_526),
.B(n_533),
.Y(n_800)
);

AND2x6_ASAP7_75t_SL g801 ( 
.A(n_562),
.B(n_642),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_562),
.Y(n_802)
);

AND2x4_ASAP7_75t_SL g803 ( 
.A(n_588),
.B(n_481),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_526),
.B(n_450),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_533),
.B(n_450),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_597),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_597),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_507),
.A2(n_450),
.B1(n_281),
.B2(n_308),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_570),
.A2(n_450),
.B(n_441),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_549),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_534),
.B(n_450),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_534),
.B(n_481),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_549),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_542),
.B(n_481),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_507),
.A2(n_247),
.B1(n_261),
.B2(n_278),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_618),
.B(n_563),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_598),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_553),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_595),
.B(n_209),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_598),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_565),
.B(n_210),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_542),
.B(n_481),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_553),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_595),
.B(n_210),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_655),
.A2(n_547),
.B1(n_579),
.B2(n_615),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_769),
.A2(n_776),
.B(n_770),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_672),
.B(n_642),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_782),
.A2(n_579),
.B(n_547),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_723),
.A2(n_579),
.B(n_566),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_658),
.B(n_642),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_660),
.B(n_642),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_656),
.B(n_624),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_823),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_667),
.B(n_624),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_670),
.B(n_671),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_727),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_680),
.A2(n_612),
.B1(n_631),
.B2(n_613),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_663),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_744),
.A2(n_566),
.B(n_557),
.Y(n_839)
);

NAND2x1_ASAP7_75t_L g840 ( 
.A(n_823),
.B(n_657),
.Y(n_840)
);

NOR2x1p5_ASAP7_75t_L g841 ( 
.A(n_751),
.B(n_551),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_747),
.A2(n_578),
.B(n_557),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_663),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_819),
.B(n_650),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_749),
.A2(n_762),
.B(n_754),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_803),
.B(n_752),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_664),
.A2(n_605),
.B(n_578),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_777),
.A2(n_613),
.B1(n_507),
.B2(n_586),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_784),
.B(n_650),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_785),
.A2(n_633),
.B(n_605),
.Y(n_850)
);

NAND2x1p5_ASAP7_75t_L g851 ( 
.A(n_752),
.B(n_601),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_673),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_789),
.A2(n_635),
.B(n_633),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_795),
.A2(n_643),
.B(n_635),
.Y(n_854)
);

NOR2x1_ASAP7_75t_L g855 ( 
.A(n_816),
.B(n_613),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_709),
.B(n_613),
.Y(n_856)
);

NAND3xp33_ASAP7_75t_L g857 ( 
.A(n_743),
.B(n_619),
.C(n_606),
.Y(n_857)
);

OAI21x1_ASAP7_75t_L g858 ( 
.A1(n_809),
.A2(n_644),
.B(n_643),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_728),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_687),
.B(n_613),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_681),
.B(n_575),
.Y(n_861)
);

NAND2xp33_ASAP7_75t_L g862 ( 
.A(n_727),
.B(n_507),
.Y(n_862)
);

NAND3xp33_ASAP7_75t_SL g863 ( 
.A(n_676),
.B(n_420),
.C(n_594),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_803),
.B(n_601),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_742),
.B(n_581),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_688),
.B(n_646),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_677),
.B(n_543),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_691),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_665),
.B(n_824),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_741),
.B(n_532),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_798),
.A2(n_647),
.B(n_644),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_804),
.A2(n_647),
.B(n_587),
.Y(n_872)
);

INVx4_ASAP7_75t_L g873 ( 
.A(n_801),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_779),
.A2(n_609),
.B1(n_639),
.B2(n_606),
.Y(n_874)
);

NAND2xp33_ASAP7_75t_SL g875 ( 
.A(n_741),
.B(n_609),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_682),
.B(n_532),
.Y(n_876)
);

NAND2xp33_ASAP7_75t_L g877 ( 
.A(n_727),
.B(n_736),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_683),
.B(n_581),
.Y(n_878)
);

A2O1A1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_684),
.A2(n_543),
.B(n_615),
.C(n_639),
.Y(n_879)
);

O2A1O1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_705),
.A2(n_636),
.B(n_640),
.C(n_626),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_679),
.B(n_556),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_823),
.Y(n_882)
);

A2O1A1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_684),
.A2(n_636),
.B(n_556),
.C(n_608),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_805),
.A2(n_621),
.B(n_587),
.Y(n_884)
);

BUFx12f_ASAP7_75t_L g885 ( 
.A(n_783),
.Y(n_885)
);

BUFx2_ASAP7_75t_L g886 ( 
.A(n_783),
.Y(n_886)
);

O2A1O1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_708),
.A2(n_625),
.B(n_614),
.C(n_630),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_695),
.A2(n_583),
.B1(n_600),
.B2(n_608),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_755),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_811),
.A2(n_621),
.B(n_587),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_657),
.B(n_581),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_682),
.B(n_532),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_727),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_751),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_657),
.B(n_581),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_775),
.A2(n_587),
.B(n_621),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_713),
.A2(n_621),
.B(n_600),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_717),
.A2(n_611),
.B(n_608),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_711),
.B(n_617),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_799),
.B(n_617),
.Y(n_900)
);

AO21x1_ASAP7_75t_L g901 ( 
.A1(n_653),
.A2(n_648),
.B(n_627),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_727),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_720),
.A2(n_611),
.B(n_600),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_695),
.B(n_702),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_692),
.B(n_532),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_758),
.A2(n_611),
.B(n_629),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_797),
.A2(n_602),
.B(n_532),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_702),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_736),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_707),
.B(n_602),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_715),
.B(n_602),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_736),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_715),
.Y(n_913)
);

NAND2xp33_ASAP7_75t_L g914 ( 
.A(n_736),
.B(n_602),
.Y(n_914)
);

INVx1_ASAP7_75t_SL g915 ( 
.A(n_755),
.Y(n_915)
);

O2A1O1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_716),
.A2(n_494),
.B(n_290),
.C(n_293),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_771),
.Y(n_917)
);

NAND2xp33_ASAP7_75t_L g918 ( 
.A(n_736),
.B(n_602),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_800),
.A2(n_632),
.B(n_577),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_716),
.B(n_632),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_718),
.B(n_632),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_693),
.A2(n_632),
.B(n_577),
.Y(n_922)
);

BUFx4f_ASAP7_75t_L g923 ( 
.A(n_799),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_694),
.A2(n_632),
.B(n_577),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_692),
.B(n_577),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_718),
.B(n_617),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_686),
.B(n_583),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_699),
.A2(n_577),
.B(n_529),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_722),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_722),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_733),
.B(n_577),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_704),
.A2(n_529),
.B(n_583),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_696),
.B(n_583),
.Y(n_933)
);

INVxp67_ASAP7_75t_L g934 ( 
.A(n_739),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_786),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_719),
.A2(n_637),
.B1(n_628),
.B2(n_617),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_733),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_719),
.B(n_218),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_734),
.B(n_617),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_712),
.A2(n_529),
.B(n_634),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_802),
.B(n_617),
.Y(n_941)
);

NOR2x1_ASAP7_75t_L g942 ( 
.A(n_780),
.B(n_603),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_729),
.B(n_218),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_734),
.B(n_735),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_729),
.B(n_256),
.Y(n_945)
);

O2A1O1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_735),
.A2(n_494),
.B(n_306),
.C(n_311),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_712),
.A2(n_603),
.B(n_634),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_764),
.B(n_617),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_771),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_764),
.B(n_628),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_700),
.B(n_256),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_812),
.A2(n_307),
.B(n_263),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_765),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_668),
.B(n_263),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_691),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_765),
.B(n_628),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_814),
.A2(n_309),
.B(n_267),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_711),
.B(n_628),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_745),
.A2(n_637),
.B(n_628),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_822),
.A2(n_309),
.B(n_267),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_792),
.B(n_628),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_792),
.B(n_628),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_793),
.A2(n_637),
.B(n_329),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_793),
.A2(n_307),
.B(n_285),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_794),
.B(n_806),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_794),
.A2(n_298),
.B(n_285),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_806),
.A2(n_286),
.B(n_287),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_807),
.B(n_637),
.Y(n_968)
);

OAI21xp5_ASAP7_75t_L g969 ( 
.A1(n_807),
.A2(n_637),
.B(n_333),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_817),
.A2(n_282),
.B(n_325),
.C(n_332),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_817),
.A2(n_820),
.B(n_771),
.Y(n_971)
);

BUFx12f_ASAP7_75t_L g972 ( 
.A(n_801),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_732),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_760),
.B(n_286),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_786),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_820),
.A2(n_298),
.B(n_287),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_772),
.A2(n_787),
.B(n_790),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_772),
.A2(n_288),
.B(n_294),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_689),
.B(n_637),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_746),
.B(n_637),
.Y(n_980)
);

AO21x1_ASAP7_75t_L g981 ( 
.A1(n_815),
.A2(n_411),
.B(n_410),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_772),
.A2(n_295),
.B(n_294),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_802),
.B(n_288),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_690),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_788),
.B(n_710),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_757),
.B(n_295),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_685),
.A2(n_481),
.B(n_417),
.C(n_411),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_659),
.Y(n_988)
);

OAI21xp5_ASAP7_75t_L g989 ( 
.A1(n_790),
.A2(n_479),
.B(n_482),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_772),
.A2(n_339),
.B(n_224),
.Y(n_990)
);

O2A1O1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_706),
.A2(n_417),
.B(n_418),
.C(n_479),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_767),
.B(n_339),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_772),
.A2(n_259),
.B(n_228),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_725),
.A2(n_418),
.B(n_479),
.C(n_482),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_703),
.B(n_10),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_810),
.Y(n_996)
);

AO21x1_ASAP7_75t_L g997 ( 
.A1(n_815),
.A2(n_479),
.B(n_396),
.Y(n_997)
);

AOI21xp33_ASAP7_75t_L g998 ( 
.A1(n_701),
.A2(n_766),
.B(n_774),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_810),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_659),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_654),
.B(n_229),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_654),
.B(n_231),
.Y(n_1002)
);

OAI21x1_ASAP7_75t_L g1003 ( 
.A1(n_813),
.A2(n_489),
.B(n_482),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_787),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_697),
.B(n_489),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_813),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_666),
.B(n_489),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_787),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_661),
.Y(n_1009)
);

NAND2x1p5_ASAP7_75t_L g1010 ( 
.A(n_654),
.B(n_787),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_787),
.A2(n_252),
.B(n_246),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_726),
.A2(n_475),
.B(n_453),
.C(n_397),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_737),
.A2(n_310),
.B1(n_232),
.B2(n_235),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_818),
.B(n_475),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_654),
.B(n_791),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_838),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_914),
.A2(n_738),
.B(n_654),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_849),
.A2(n_731),
.B1(n_796),
.B2(n_808),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_918),
.A2(n_738),
.B(n_748),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_995),
.A2(n_714),
.B(n_740),
.C(n_773),
.Y(n_1020)
);

A2O1A1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_995),
.A2(n_821),
.B(n_674),
.C(n_678),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_843),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_860),
.B(n_818),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_984),
.B(n_661),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_935),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_825),
.A2(n_781),
.B(n_778),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_828),
.A2(n_698),
.B(n_778),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_832),
.A2(n_781),
.B1(n_768),
.B2(n_763),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_904),
.A2(n_768),
.B1(n_763),
.B2(n_761),
.Y(n_1029)
);

AOI21x1_ASAP7_75t_L g1030 ( 
.A1(n_901),
.A2(n_761),
.B(n_759),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_R g1031 ( 
.A(n_973),
.B(n_662),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_826),
.A2(n_865),
.B(n_845),
.Y(n_1032)
);

BUFx8_ASAP7_75t_L g1033 ( 
.A(n_894),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_984),
.A2(n_759),
.B1(n_756),
.B2(n_753),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_860),
.B(n_756),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_934),
.B(n_662),
.Y(n_1036)
);

AOI21xp33_ASAP7_75t_L g1037 ( 
.A1(n_974),
.A2(n_753),
.B(n_750),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_852),
.Y(n_1038)
);

OAI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_971),
.A2(n_750),
.B(n_730),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_944),
.A2(n_730),
.B1(n_724),
.B2(n_721),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_830),
.B(n_724),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_844),
.A2(n_721),
.B1(n_698),
.B2(n_675),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_864),
.B(n_675),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_934),
.B(n_1005),
.Y(n_1044)
);

NOR3xp33_ASAP7_75t_SL g1045 ( 
.A(n_951),
.B(n_323),
.C(n_250),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_R g1046 ( 
.A(n_859),
.B(n_669),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_861),
.B(n_669),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_861),
.A2(n_475),
.B(n_453),
.C(n_396),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_827),
.B(n_453),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_889),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_975),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_858),
.A2(n_397),
.B(n_477),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_865),
.A2(n_244),
.B(n_239),
.Y(n_1053)
);

NOR3xp33_ASAP7_75t_SL g1054 ( 
.A(n_951),
.B(n_12),
.C(n_14),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_908),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_841),
.B(n_397),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_986),
.A2(n_12),
.B(n_16),
.C(n_17),
.Y(n_1057)
);

AOI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_863),
.A2(n_477),
.B1(n_321),
.B2(n_222),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_864),
.B(n_17),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_877),
.A2(n_321),
.B(n_222),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_866),
.B(n_21),
.Y(n_1061)
);

AOI22xp33_ASAP7_75t_SL g1062 ( 
.A1(n_857),
.A2(n_321),
.B1(n_477),
.B2(n_27),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_996),
.Y(n_1063)
);

NAND3xp33_ASAP7_75t_SL g1064 ( 
.A(n_992),
.B(n_21),
.C(n_24),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_837),
.B(n_477),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_848),
.B(n_24),
.Y(n_1066)
);

NOR2xp67_ASAP7_75t_L g1067 ( 
.A(n_873),
.B(n_161),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_907),
.A2(n_321),
.B(n_477),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_886),
.B(n_29),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_913),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_915),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_910),
.A2(n_321),
.B(n_477),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_911),
.A2(n_477),
.B(n_158),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_836),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_929),
.Y(n_1075)
);

AOI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_863),
.A2(n_477),
.B1(n_33),
.B2(n_35),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_930),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_998),
.B(n_31),
.Y(n_1078)
);

NOR3xp33_ASAP7_75t_SL g1079 ( 
.A(n_964),
.B(n_36),
.C(n_38),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_985),
.B(n_40),
.Y(n_1080)
);

BUFx12f_ASAP7_75t_L g1081 ( 
.A(n_885),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_869),
.B(n_985),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_836),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_874),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_1084)
);

NAND2x1p5_ASAP7_75t_L g1085 ( 
.A(n_923),
.B(n_156),
.Y(n_1085)
);

INVx4_ASAP7_75t_L g1086 ( 
.A(n_846),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_937),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_974),
.A2(n_41),
.B(n_44),
.C(n_45),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_900),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_900),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_920),
.A2(n_154),
.B(n_151),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_999),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_836),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_953),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1006),
.Y(n_1095)
);

BUFx8_ASAP7_75t_L g1096 ( 
.A(n_972),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_836),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_835),
.B(n_44),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_831),
.B(n_46),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_868),
.A2(n_955),
.B1(n_834),
.B2(n_867),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_869),
.B(n_47),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_921),
.A2(n_71),
.B(n_124),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_954),
.B(n_48),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_988),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1000),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_893),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_829),
.A2(n_134),
.B(n_116),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1009),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_847),
.A2(n_105),
.B(n_100),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_846),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_868),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_1111)
);

NAND3xp33_ASAP7_75t_SL g1112 ( 
.A(n_954),
.B(n_51),
.C(n_52),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_888),
.A2(n_91),
.B(n_89),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_965),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_872),
.A2(n_78),
.B(n_75),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_955),
.B(n_67),
.Y(n_1116)
);

HB1xp67_ASAP7_75t_L g1117 ( 
.A(n_899),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_884),
.A2(n_53),
.B(n_57),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_856),
.B(n_53),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_833),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_916),
.A2(n_59),
.B(n_62),
.C(n_64),
.Y(n_1121)
);

NAND3xp33_ASAP7_75t_SL g1122 ( 
.A(n_946),
.B(n_59),
.C(n_65),
.Y(n_1122)
);

NOR3xp33_ASAP7_75t_SL g1123 ( 
.A(n_966),
.B(n_67),
.C(n_967),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_890),
.A2(n_896),
.B(n_919),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_850),
.A2(n_853),
.B(n_854),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_882),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_958),
.B(n_923),
.Y(n_1127)
);

INVx1_ASAP7_75t_SL g1128 ( 
.A(n_941),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_873),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_965),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_855),
.B(n_851),
.Y(n_1131)
);

INVx1_ASAP7_75t_SL g1132 ( 
.A(n_941),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_881),
.A2(n_879),
.B1(n_943),
.B2(n_945),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_L g1134 ( 
.A1(n_938),
.A2(n_979),
.B1(n_983),
.B2(n_933),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_917),
.B(n_949),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_936),
.A2(n_851),
.B1(n_969),
.B2(n_963),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_917),
.B(n_949),
.Y(n_1137)
);

AOI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_878),
.A2(n_927),
.B1(n_933),
.B2(n_862),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_SL g1139 ( 
.A(n_1010),
.B(n_980),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1014),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_878),
.B(n_1004),
.Y(n_1141)
);

INVx5_ASAP7_75t_L g1142 ( 
.A(n_893),
.Y(n_1142)
);

O2A1O1Ixp33_ASAP7_75t_SL g1143 ( 
.A1(n_931),
.A2(n_883),
.B(n_925),
.C(n_840),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1004),
.B(n_927),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_970),
.B(n_976),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_931),
.B(n_1013),
.Y(n_1146)
);

INVx5_ASAP7_75t_L g1147 ( 
.A(n_893),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_893),
.B(n_909),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_902),
.B(n_912),
.Y(n_1149)
);

O2A1O1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_880),
.A2(n_987),
.B(n_887),
.C(n_906),
.Y(n_1150)
);

NOR2x1_ASAP7_75t_L g1151 ( 
.A(n_942),
.B(n_1001),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1012),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_994),
.Y(n_1153)
);

AND2x4_ASAP7_75t_L g1154 ( 
.A(n_902),
.B(n_912),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_SL g1155 ( 
.A(n_1010),
.B(n_909),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_926),
.A2(n_948),
.B1(n_968),
.B2(n_962),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_939),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_871),
.A2(n_839),
.B(n_842),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_902),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_981),
.A2(n_1015),
.B1(n_1007),
.B2(n_950),
.Y(n_1160)
);

NAND2x1_ASAP7_75t_L g1161 ( 
.A(n_902),
.B(n_909),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_956),
.Y(n_1162)
);

AOI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_875),
.A2(n_1015),
.B1(n_961),
.B2(n_925),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_940),
.A2(n_947),
.B(n_959),
.C(n_957),
.Y(n_1164)
);

INVx2_ASAP7_75t_SL g1165 ( 
.A(n_909),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_912),
.B(n_1008),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_912),
.B(n_1008),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_SL g1168 ( 
.A(n_1008),
.B(n_977),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_1008),
.B(n_870),
.Y(n_1169)
);

INVxp67_ASAP7_75t_L g1170 ( 
.A(n_978),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_982),
.B(n_990),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_997),
.A2(n_960),
.B1(n_952),
.B2(n_1002),
.Y(n_1172)
);

NAND2x1p5_ASAP7_75t_L g1173 ( 
.A(n_876),
.B(n_892),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_1050),
.Y(n_1174)
);

INVx3_ASAP7_75t_L g1175 ( 
.A(n_1142),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1044),
.B(n_1011),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1016),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1022),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_1031),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1024),
.B(n_993),
.Y(n_1180)
);

O2A1O1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_1103),
.A2(n_1020),
.B(n_1080),
.C(n_1021),
.Y(n_1181)
);

AO21x1_ASAP7_75t_L g1182 ( 
.A1(n_1100),
.A2(n_932),
.B(n_928),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1023),
.B(n_891),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1052),
.A2(n_1003),
.B(n_898),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1082),
.B(n_989),
.Y(n_1185)
);

AOI221x1_ASAP7_75t_L g1186 ( 
.A1(n_1084),
.A2(n_903),
.B1(n_897),
.B2(n_922),
.C(n_924),
.Y(n_1186)
);

INVxp67_ASAP7_75t_SL g1187 ( 
.A(n_1035),
.Y(n_1187)
);

OR2x2_ASAP7_75t_L g1188 ( 
.A(n_1101),
.B(n_895),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1032),
.A2(n_905),
.B(n_991),
.Y(n_1189)
);

AOI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1078),
.A2(n_1112),
.B1(n_1033),
.B2(n_1122),
.Y(n_1190)
);

OAI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1150),
.A2(n_1164),
.B(n_1061),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1100),
.B(n_1128),
.Y(n_1192)
);

AO31x2_ASAP7_75t_L g1193 ( 
.A1(n_1042),
.A2(n_1028),
.A3(n_1029),
.B(n_1040),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1104),
.Y(n_1194)
);

O2A1O1Ixp5_ASAP7_75t_L g1195 ( 
.A1(n_1133),
.A2(n_1119),
.B(n_1019),
.C(n_1171),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1128),
.B(n_1132),
.Y(n_1196)
);

OAI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1133),
.A2(n_1026),
.B(n_1027),
.Y(n_1197)
);

AO32x2_ASAP7_75t_L g1198 ( 
.A1(n_1111),
.A2(n_1042),
.A3(n_1028),
.B1(n_1040),
.B2(n_1029),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1038),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1124),
.A2(n_1017),
.B(n_1158),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1125),
.A2(n_1027),
.B(n_1030),
.Y(n_1201)
);

A2O1A1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1146),
.A2(n_1076),
.B(n_1123),
.C(n_1066),
.Y(n_1202)
);

O2A1O1Ixp5_ASAP7_75t_L g1203 ( 
.A1(n_1113),
.A2(n_1073),
.B(n_1068),
.C(n_1072),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1098),
.A2(n_1099),
.B(n_1156),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1156),
.A2(n_1138),
.B(n_1163),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1055),
.Y(n_1206)
);

AO31x2_ASAP7_75t_L g1207 ( 
.A1(n_1136),
.A2(n_1018),
.A3(n_1162),
.B(n_1157),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1039),
.A2(n_1109),
.B(n_1107),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1136),
.A2(n_1139),
.B(n_1143),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1086),
.B(n_1142),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1139),
.A2(n_1141),
.B(n_1168),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1105),
.Y(n_1212)
);

A2O1A1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_1145),
.A2(n_1045),
.B(n_1057),
.C(n_1088),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1168),
.A2(n_1115),
.B(n_1039),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1060),
.A2(n_1144),
.B(n_1160),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1148),
.A2(n_1149),
.B(n_1018),
.Y(n_1216)
);

INVx3_ASAP7_75t_SL g1217 ( 
.A(n_1129),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1043),
.A2(n_1025),
.B1(n_1095),
.B2(n_1092),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1155),
.A2(n_1166),
.B(n_1091),
.Y(n_1219)
);

O2A1O1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1121),
.A2(n_1064),
.B(n_1111),
.C(n_1054),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1116),
.A2(n_1094),
.B1(n_1070),
.B2(n_1075),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1132),
.B(n_1077),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1155),
.A2(n_1102),
.B(n_1041),
.Y(n_1223)
);

BUFx2_ASAP7_75t_R g1224 ( 
.A(n_1127),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1161),
.A2(n_1135),
.B(n_1137),
.Y(n_1225)
);

INVx4_ASAP7_75t_SL g1226 ( 
.A(n_1154),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1087),
.B(n_1089),
.Y(n_1227)
);

BUFx10_ASAP7_75t_L g1228 ( 
.A(n_1154),
.Y(n_1228)
);

INVxp67_ASAP7_75t_L g1229 ( 
.A(n_1033),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1108),
.Y(n_1230)
);

AOI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1065),
.A2(n_1047),
.B(n_1131),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_1046),
.Y(n_1232)
);

OA21x2_ASAP7_75t_L g1233 ( 
.A1(n_1037),
.A2(n_1152),
.B(n_1048),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1173),
.A2(n_1114),
.B(n_1130),
.Y(n_1234)
);

O2A1O1Ixp33_ASAP7_75t_SL g1235 ( 
.A1(n_1170),
.A2(n_1118),
.B(n_1036),
.C(n_1165),
.Y(n_1235)
);

O2A1O1Ixp33_ASAP7_75t_SL g1236 ( 
.A1(n_1153),
.A2(n_1059),
.B(n_1053),
.C(n_1049),
.Y(n_1236)
);

AO21x1_ASAP7_75t_L g1237 ( 
.A1(n_1173),
.A2(n_1085),
.B(n_1034),
.Y(n_1237)
);

A2O1A1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1058),
.A2(n_1062),
.B(n_1079),
.C(n_1151),
.Y(n_1238)
);

OR2x6_ASAP7_75t_L g1239 ( 
.A(n_1086),
.B(n_1110),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1089),
.B(n_1090),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1172),
.A2(n_1134),
.B(n_1140),
.Y(n_1241)
);

INVxp67_ASAP7_75t_L g1242 ( 
.A(n_1071),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1167),
.A2(n_1147),
.B(n_1142),
.Y(n_1243)
);

AO21x1_ASAP7_75t_L g1244 ( 
.A1(n_1085),
.A2(n_1169),
.B(n_1056),
.Y(n_1244)
);

BUFx8_ASAP7_75t_L g1245 ( 
.A(n_1081),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1167),
.A2(n_1142),
.B(n_1147),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1090),
.B(n_1043),
.Y(n_1247)
);

OAI22x1_ASAP7_75t_L g1248 ( 
.A1(n_1069),
.A2(n_1117),
.B1(n_1126),
.B2(n_1120),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1051),
.A2(n_1063),
.B(n_1067),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1169),
.Y(n_1250)
);

O2A1O1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1147),
.A2(n_1096),
.B(n_1083),
.C(n_1093),
.Y(n_1251)
);

O2A1O1Ixp5_ASAP7_75t_L g1252 ( 
.A1(n_1147),
.A2(n_1074),
.B(n_1083),
.C(n_1093),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1159),
.B(n_1074),
.Y(n_1253)
);

BUFx3_ASAP7_75t_L g1254 ( 
.A(n_1096),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1074),
.A2(n_1083),
.B(n_1093),
.Y(n_1255)
);

A2O1A1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1097),
.A2(n_1103),
.B(n_995),
.C(n_658),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1097),
.B(n_1106),
.Y(n_1257)
);

BUFx12f_ASAP7_75t_L g1258 ( 
.A(n_1106),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1106),
.A2(n_1103),
.B1(n_995),
.B2(n_860),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1159),
.A2(n_995),
.B(n_1150),
.Y(n_1260)
);

AOI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1159),
.A2(n_1032),
.B(n_1124),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1023),
.B(n_1035),
.Y(n_1262)
);

AOI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1032),
.A2(n_1124),
.B(n_1158),
.Y(n_1263)
);

AOI221xp5_ASAP7_75t_L g1264 ( 
.A1(n_1103),
.A2(n_676),
.B1(n_743),
.B2(n_680),
.C(n_777),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1044),
.B(n_680),
.Y(n_1265)
);

A2O1A1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1103),
.A2(n_995),
.B(n_658),
.C(n_934),
.Y(n_1266)
);

AO32x2_ASAP7_75t_L g1267 ( 
.A1(n_1100),
.A2(n_1111),
.A3(n_1084),
.B1(n_1042),
.B2(n_1133),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_1142),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1082),
.B(n_984),
.Y(n_1269)
);

O2A1O1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1103),
.A2(n_680),
.B(n_995),
.C(n_934),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1150),
.A2(n_995),
.B(n_1103),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1103),
.A2(n_676),
.B1(n_697),
.B2(n_690),
.Y(n_1272)
);

OAI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1150),
.A2(n_995),
.B(n_1103),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1032),
.A2(n_918),
.B(n_914),
.Y(n_1274)
);

AND2x4_ASAP7_75t_SL g1275 ( 
.A(n_1086),
.B(n_518),
.Y(n_1275)
);

BUFx24_ASAP7_75t_L g1276 ( 
.A(n_1154),
.Y(n_1276)
);

AOI221x1_ASAP7_75t_L g1277 ( 
.A1(n_1103),
.A2(n_995),
.B1(n_1084),
.B2(n_1088),
.C(n_1020),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1104),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1052),
.A2(n_858),
.B(n_1124),
.Y(n_1279)
);

AOI221xp5_ASAP7_75t_L g1280 ( 
.A1(n_1103),
.A2(n_676),
.B1(n_743),
.B2(n_680),
.C(n_777),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_1046),
.Y(n_1281)
);

NOR2xp67_ASAP7_75t_SL g1282 ( 
.A(n_1081),
.B(n_652),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1150),
.A2(n_995),
.B(n_1103),
.Y(n_1283)
);

NOR2xp67_ASAP7_75t_L g1284 ( 
.A(n_1082),
.B(n_728),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1016),
.Y(n_1285)
);

INVx4_ASAP7_75t_L g1286 ( 
.A(n_1050),
.Y(n_1286)
);

AO31x2_ASAP7_75t_L g1287 ( 
.A1(n_1164),
.A2(n_825),
.A3(n_901),
.B(n_1042),
.Y(n_1287)
);

O2A1O1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1103),
.A2(n_680),
.B(n_995),
.C(n_934),
.Y(n_1288)
);

NAND3xp33_ASAP7_75t_L g1289 ( 
.A(n_1103),
.B(n_995),
.C(n_1078),
.Y(n_1289)
);

O2A1O1Ixp33_ASAP7_75t_SL g1290 ( 
.A1(n_1021),
.A2(n_1088),
.B(n_995),
.C(n_1103),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1104),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1032),
.A2(n_918),
.B(n_914),
.Y(n_1292)
);

BUFx2_ASAP7_75t_L g1293 ( 
.A(n_1033),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1082),
.B(n_984),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_SL g1295 ( 
.A1(n_1023),
.A2(n_1035),
.B(n_830),
.Y(n_1295)
);

AO21x1_ASAP7_75t_L g1296 ( 
.A1(n_1103),
.A2(n_995),
.B(n_1100),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1023),
.B(n_1035),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1032),
.A2(n_918),
.B(n_914),
.Y(n_1298)
);

O2A1O1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1103),
.A2(n_680),
.B(n_995),
.C(n_934),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1052),
.A2(n_858),
.B(n_1124),
.Y(n_1300)
);

AO31x2_ASAP7_75t_L g1301 ( 
.A1(n_1164),
.A2(n_825),
.A3(n_901),
.B(n_1042),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1103),
.A2(n_995),
.B1(n_860),
.B2(n_849),
.Y(n_1302)
);

INVxp67_ASAP7_75t_L g1303 ( 
.A(n_1033),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1082),
.B(n_984),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1032),
.A2(n_918),
.B(n_914),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1103),
.A2(n_995),
.B1(n_860),
.B2(n_849),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1032),
.A2(n_918),
.B(n_914),
.Y(n_1307)
);

NAND3xp33_ASAP7_75t_SL g1308 ( 
.A(n_1103),
.B(n_676),
.C(n_424),
.Y(n_1308)
);

OAI22x1_ASAP7_75t_L g1309 ( 
.A1(n_1103),
.A2(n_576),
.B1(n_486),
.B2(n_676),
.Y(n_1309)
);

NAND2x1p5_ASAP7_75t_L g1310 ( 
.A(n_1086),
.B(n_1142),
.Y(n_1310)
);

INVx5_ASAP7_75t_L g1311 ( 
.A(n_1142),
.Y(n_1311)
);

BUFx2_ASAP7_75t_L g1312 ( 
.A(n_1033),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1033),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1044),
.B(n_680),
.Y(n_1314)
);

BUFx6f_ASAP7_75t_L g1315 ( 
.A(n_1142),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1086),
.B(n_1089),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1044),
.B(n_680),
.Y(n_1317)
);

BUFx6f_ASAP7_75t_L g1318 ( 
.A(n_1142),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1032),
.A2(n_918),
.B(n_914),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1103),
.A2(n_676),
.B1(n_697),
.B2(n_690),
.Y(n_1320)
);

AOI221xp5_ASAP7_75t_L g1321 ( 
.A1(n_1103),
.A2(n_676),
.B1(n_743),
.B2(n_680),
.C(n_777),
.Y(n_1321)
);

AOI221xp5_ASAP7_75t_L g1322 ( 
.A1(n_1103),
.A2(n_676),
.B1(n_743),
.B2(n_680),
.C(n_777),
.Y(n_1322)
);

AO32x2_ASAP7_75t_L g1323 ( 
.A1(n_1100),
.A2(n_1111),
.A3(n_1084),
.B1(n_1042),
.B2(n_1133),
.Y(n_1323)
);

INVxp67_ASAP7_75t_SL g1324 ( 
.A(n_1024),
.Y(n_1324)
);

AO31x2_ASAP7_75t_L g1325 ( 
.A1(n_1164),
.A2(n_825),
.A3(n_901),
.B(n_1042),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1023),
.B(n_1035),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1052),
.A2(n_858),
.B(n_1124),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1032),
.A2(n_918),
.B(n_914),
.Y(n_1328)
);

AO31x2_ASAP7_75t_L g1329 ( 
.A1(n_1164),
.A2(n_825),
.A3(n_901),
.B(n_1042),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1150),
.A2(n_995),
.B(n_1103),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1044),
.B(n_680),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1104),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1104),
.Y(n_1333)
);

BUFx6f_ASAP7_75t_L g1334 ( 
.A(n_1142),
.Y(n_1334)
);

AOI21xp33_ASAP7_75t_L g1335 ( 
.A1(n_1289),
.A2(n_1273),
.B(n_1271),
.Y(n_1335)
);

OAI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1289),
.A2(n_1309),
.B1(n_1271),
.B2(n_1283),
.Y(n_1336)
);

CKINVDCx14_ASAP7_75t_R g1337 ( 
.A(n_1254),
.Y(n_1337)
);

INVx1_ASAP7_75t_SL g1338 ( 
.A(n_1275),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1177),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_SL g1340 ( 
.A1(n_1302),
.A2(n_1306),
.B1(n_1330),
.B2(n_1273),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_SL g1341 ( 
.A1(n_1302),
.A2(n_1306),
.B1(n_1283),
.B2(n_1330),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1232),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1266),
.A2(n_1320),
.B1(n_1272),
.B2(n_1288),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1264),
.A2(n_1280),
.B1(n_1321),
.B2(n_1322),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_SL g1345 ( 
.A1(n_1259),
.A2(n_1205),
.B1(n_1221),
.B2(n_1192),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_1245),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1296),
.A2(n_1308),
.B1(n_1259),
.B2(n_1248),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1258),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1174),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1270),
.A2(n_1299),
.B1(n_1256),
.B2(n_1190),
.Y(n_1350)
);

CKINVDCx11_ASAP7_75t_R g1351 ( 
.A(n_1293),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1205),
.A2(n_1324),
.B1(n_1212),
.B2(n_1291),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1269),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1181),
.A2(n_1202),
.B1(n_1213),
.B2(n_1317),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1178),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1194),
.A2(n_1278),
.B1(n_1333),
.B2(n_1332),
.Y(n_1356)
);

OAI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1277),
.A2(n_1331),
.B1(n_1314),
.B2(n_1265),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1185),
.A2(n_1192),
.B1(n_1187),
.B2(n_1221),
.Y(n_1358)
);

CKINVDCx14_ASAP7_75t_R g1359 ( 
.A(n_1312),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_1245),
.Y(n_1360)
);

OAI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1284),
.A2(n_1179),
.B1(n_1260),
.B2(n_1304),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_SL g1362 ( 
.A1(n_1260),
.A2(n_1204),
.B1(n_1191),
.B2(n_1294),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1222),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_1313),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_SL g1365 ( 
.A1(n_1204),
.A2(n_1191),
.B1(n_1290),
.B2(n_1209),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1311),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1199),
.Y(n_1367)
);

CKINVDCx11_ASAP7_75t_R g1368 ( 
.A(n_1217),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1206),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1234),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1250),
.A2(n_1218),
.B1(n_1176),
.B2(n_1180),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1239),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1220),
.A2(n_1238),
.B1(n_1188),
.B2(n_1297),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_1229),
.Y(n_1374)
);

BUFx2_ASAP7_75t_L g1375 ( 
.A(n_1315),
.Y(n_1375)
);

INVx1_ASAP7_75t_SL g1376 ( 
.A(n_1281),
.Y(n_1376)
);

OAI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1303),
.A2(n_1297),
.B1(n_1326),
.B2(n_1262),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_1315),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_1286),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_SL g1380 ( 
.A1(n_1197),
.A2(n_1326),
.B1(n_1262),
.B2(n_1222),
.Y(n_1380)
);

INVx6_ASAP7_75t_L g1381 ( 
.A(n_1228),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_SL g1382 ( 
.A1(n_1197),
.A2(n_1267),
.B1(n_1323),
.B2(n_1247),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1244),
.A2(n_1196),
.B1(n_1230),
.B2(n_1247),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1196),
.A2(n_1285),
.B1(n_1237),
.B2(n_1282),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_SL g1385 ( 
.A1(n_1286),
.A2(n_1242),
.B1(n_1316),
.B2(n_1227),
.Y(n_1385)
);

INVx6_ASAP7_75t_L g1386 ( 
.A(n_1226),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_SL g1387 ( 
.A1(n_1267),
.A2(n_1323),
.B1(n_1276),
.B2(n_1241),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1227),
.Y(n_1388)
);

CKINVDCx20_ASAP7_75t_R g1389 ( 
.A(n_1226),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1240),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1183),
.A2(n_1249),
.B1(n_1182),
.B2(n_1233),
.Y(n_1391)
);

CKINVDCx11_ASAP7_75t_R g1392 ( 
.A(n_1318),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_SL g1393 ( 
.A1(n_1267),
.A2(n_1323),
.B1(n_1233),
.B2(n_1183),
.Y(n_1393)
);

INVxp67_ASAP7_75t_L g1394 ( 
.A(n_1253),
.Y(n_1394)
);

BUFx3_ASAP7_75t_L g1395 ( 
.A(n_1318),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1240),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1316),
.A2(n_1216),
.B1(n_1226),
.B2(n_1211),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1224),
.B(n_1310),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1253),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_SL g1400 ( 
.A1(n_1214),
.A2(n_1215),
.B1(n_1198),
.B2(n_1219),
.Y(n_1400)
);

CKINVDCx11_ASAP7_75t_R g1401 ( 
.A(n_1318),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1231),
.Y(n_1402)
);

INVx1_ASAP7_75t_SL g1403 ( 
.A(n_1257),
.Y(n_1403)
);

INVx1_ASAP7_75t_SL g1404 ( 
.A(n_1334),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1210),
.A2(n_1223),
.B1(n_1225),
.B2(n_1334),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1207),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_1175),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1295),
.A2(n_1305),
.B1(n_1328),
.B2(n_1319),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1195),
.A2(n_1236),
.B(n_1189),
.Y(n_1409)
);

BUFx4f_ASAP7_75t_L g1410 ( 
.A(n_1310),
.Y(n_1410)
);

CKINVDCx10_ASAP7_75t_R g1411 ( 
.A(n_1251),
.Y(n_1411)
);

OAI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1175),
.A2(n_1268),
.B1(n_1246),
.B2(n_1243),
.Y(n_1412)
);

INVx5_ASAP7_75t_L g1413 ( 
.A(n_1268),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1208),
.A2(n_1292),
.B1(n_1274),
.B2(n_1298),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1307),
.A2(n_1255),
.B1(n_1201),
.B2(n_1198),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1198),
.A2(n_1200),
.B1(n_1184),
.B2(n_1327),
.Y(n_1416)
);

OAI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1186),
.A2(n_1261),
.B1(n_1325),
.B2(n_1301),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1263),
.A2(n_1235),
.B1(n_1329),
.B2(n_1287),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1279),
.A2(n_1300),
.B1(n_1193),
.B2(n_1287),
.Y(n_1419)
);

CKINVDCx11_ASAP7_75t_R g1420 ( 
.A(n_1252),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1193),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1287),
.A2(n_1301),
.B1(n_1325),
.B2(n_1329),
.Y(n_1422)
);

BUFx4_ASAP7_75t_R g1423 ( 
.A(n_1301),
.Y(n_1423)
);

CKINVDCx6p67_ASAP7_75t_R g1424 ( 
.A(n_1325),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1329),
.A2(n_1309),
.B1(n_1320),
.B2(n_1272),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1203),
.A2(n_1309),
.B1(n_1320),
.B2(n_1272),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_1258),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1289),
.A2(n_676),
.B1(n_1306),
.B2(n_1302),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1177),
.Y(n_1429)
);

BUFx2_ASAP7_75t_SL g1430 ( 
.A(n_1174),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1177),
.Y(n_1431)
);

CKINVDCx11_ASAP7_75t_R g1432 ( 
.A(n_1254),
.Y(n_1432)
);

OAI21xp5_ASAP7_75t_SL g1433 ( 
.A1(n_1271),
.A2(n_1283),
.B(n_1273),
.Y(n_1433)
);

INVx6_ASAP7_75t_L g1434 ( 
.A(n_1311),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1309),
.A2(n_1320),
.B1(n_1272),
.B2(n_676),
.Y(n_1435)
);

OAI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1289),
.A2(n_576),
.B1(n_1309),
.B2(n_1273),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1269),
.Y(n_1437)
);

INVx3_ASAP7_75t_L g1438 ( 
.A(n_1234),
.Y(n_1438)
);

BUFx4f_ASAP7_75t_L g1439 ( 
.A(n_1275),
.Y(n_1439)
);

BUFx12f_ASAP7_75t_L g1440 ( 
.A(n_1245),
.Y(n_1440)
);

CKINVDCx6p67_ASAP7_75t_R g1441 ( 
.A(n_1254),
.Y(n_1441)
);

INVx6_ASAP7_75t_L g1442 ( 
.A(n_1311),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1289),
.A2(n_1283),
.B(n_1271),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_SL g1444 ( 
.A1(n_1289),
.A2(n_676),
.B1(n_1306),
.B2(n_1302),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_SL g1445 ( 
.A1(n_1289),
.A2(n_676),
.B1(n_1306),
.B2(n_1302),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1177),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1177),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1289),
.A2(n_1266),
.B1(n_1320),
.B2(n_1272),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1309),
.A2(n_1320),
.B1(n_1272),
.B2(n_676),
.Y(n_1449)
);

CKINVDCx6p67_ASAP7_75t_R g1450 ( 
.A(n_1254),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1177),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1289),
.A2(n_1266),
.B1(n_1320),
.B2(n_1272),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1289),
.A2(n_1266),
.B1(n_1320),
.B2(n_1272),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1234),
.Y(n_1454)
);

BUFx8_ASAP7_75t_L g1455 ( 
.A(n_1293),
.Y(n_1455)
);

INVx6_ASAP7_75t_L g1456 ( 
.A(n_1311),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_1245),
.Y(n_1457)
);

CKINVDCx11_ASAP7_75t_R g1458 ( 
.A(n_1254),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1177),
.Y(n_1459)
);

BUFx10_ASAP7_75t_L g1460 ( 
.A(n_1275),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1177),
.Y(n_1461)
);

CKINVDCx20_ASAP7_75t_R g1462 ( 
.A(n_1245),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1258),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1289),
.A2(n_1266),
.B1(n_1320),
.B2(n_1272),
.Y(n_1464)
);

AOI22x1_ASAP7_75t_SL g1465 ( 
.A1(n_1179),
.A2(n_518),
.B1(n_973),
.B2(n_192),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1234),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1309),
.A2(n_1320),
.B1(n_1272),
.B2(n_676),
.Y(n_1467)
);

AND2x4_ASAP7_75t_L g1468 ( 
.A(n_1438),
.B(n_1370),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1409),
.A2(n_1408),
.B(n_1414),
.Y(n_1469)
);

BUFx2_ASAP7_75t_SL g1470 ( 
.A(n_1389),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1421),
.Y(n_1471)
);

INVx1_ASAP7_75t_SL g1472 ( 
.A(n_1420),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1382),
.B(n_1353),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1402),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1437),
.B(n_1345),
.Y(n_1475)
);

AOI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1418),
.A2(n_1350),
.B(n_1448),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1394),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_1424),
.Y(n_1478)
);

INVx4_ASAP7_75t_L g1479 ( 
.A(n_1413),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1416),
.A2(n_1419),
.B(n_1391),
.Y(n_1480)
);

INVxp67_ASAP7_75t_L g1481 ( 
.A(n_1342),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1388),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1390),
.Y(n_1483)
);

NAND3xp33_ASAP7_75t_L g1484 ( 
.A(n_1344),
.B(n_1444),
.C(n_1428),
.Y(n_1484)
);

INVx3_ASAP7_75t_L g1485 ( 
.A(n_1424),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1339),
.B(n_1355),
.Y(n_1486)
);

AOI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1433),
.A2(n_1340),
.B(n_1341),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1396),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1380),
.B(n_1358),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1406),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1363),
.B(n_1443),
.Y(n_1491)
);

INVxp33_ASAP7_75t_L g1492 ( 
.A(n_1368),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1367),
.B(n_1369),
.Y(n_1493)
);

AOI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1452),
.A2(n_1453),
.B(n_1464),
.Y(n_1494)
);

OAI21x1_ASAP7_75t_L g1495 ( 
.A1(n_1415),
.A2(n_1454),
.B(n_1466),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1377),
.B(n_1362),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_SL g1497 ( 
.A(n_1445),
.B(n_1357),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1434),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1429),
.B(n_1431),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_1440),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1440),
.Y(n_1501)
);

OA21x2_ASAP7_75t_L g1502 ( 
.A1(n_1422),
.A2(n_1335),
.B(n_1466),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1457),
.Y(n_1503)
);

INVxp67_ASAP7_75t_L g1504 ( 
.A(n_1403),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1399),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1446),
.Y(n_1506)
);

AO21x2_ASAP7_75t_L g1507 ( 
.A1(n_1417),
.A2(n_1336),
.B(n_1436),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1393),
.B(n_1373),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1365),
.B(n_1447),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1451),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1459),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1461),
.B(n_1387),
.Y(n_1512)
);

BUFx3_ASAP7_75t_L g1513 ( 
.A(n_1372),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1423),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1343),
.A2(n_1426),
.B1(n_1354),
.B2(n_1449),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1425),
.B(n_1352),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1400),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1371),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1435),
.A2(n_1467),
.B1(n_1383),
.B2(n_1347),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1405),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1397),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1356),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1412),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1407),
.B(n_1378),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1378),
.B(n_1384),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1385),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1361),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1366),
.Y(n_1528)
);

OAI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1410),
.A2(n_1439),
.B(n_1366),
.Y(n_1529)
);

OA21x2_ASAP7_75t_L g1530 ( 
.A1(n_1375),
.A2(n_1404),
.B(n_1398),
.Y(n_1530)
);

INVxp67_ASAP7_75t_R g1531 ( 
.A(n_1439),
.Y(n_1531)
);

OA21x2_ASAP7_75t_L g1532 ( 
.A1(n_1420),
.A2(n_1379),
.B(n_1376),
.Y(n_1532)
);

BUFx2_ASAP7_75t_L g1533 ( 
.A(n_1395),
.Y(n_1533)
);

AOI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1348),
.A2(n_1463),
.B(n_1442),
.Y(n_1534)
);

INVx5_ASAP7_75t_L g1535 ( 
.A(n_1386),
.Y(n_1535)
);

INVx2_ASAP7_75t_SL g1536 ( 
.A(n_1456),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1389),
.B(n_1349),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1349),
.B(n_1359),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1386),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1386),
.Y(n_1540)
);

OAI21x1_ASAP7_75t_L g1541 ( 
.A1(n_1392),
.A2(n_1401),
.B(n_1381),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1359),
.B(n_1430),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1338),
.A2(n_1364),
.B1(n_1337),
.B2(n_1379),
.Y(n_1543)
);

AO32x2_ASAP7_75t_L g1544 ( 
.A1(n_1515),
.A2(n_1536),
.A3(n_1498),
.B1(n_1543),
.B2(n_1479),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1485),
.B(n_1427),
.Y(n_1545)
);

NAND2xp33_ASAP7_75t_L g1546 ( 
.A(n_1484),
.B(n_1457),
.Y(n_1546)
);

NAND3xp33_ASAP7_75t_L g1547 ( 
.A(n_1487),
.B(n_1455),
.C(n_1401),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1477),
.B(n_1364),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1537),
.B(n_1337),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1537),
.B(n_1351),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1471),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1511),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1484),
.A2(n_1374),
.B1(n_1450),
.B2(n_1441),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1485),
.B(n_1427),
.Y(n_1554)
);

A2O1A1Ixp33_ASAP7_75t_L g1555 ( 
.A1(n_1515),
.A2(n_1411),
.B(n_1392),
.C(n_1465),
.Y(n_1555)
);

A2O1A1Ixp33_ASAP7_75t_L g1556 ( 
.A1(n_1496),
.A2(n_1374),
.B(n_1460),
.C(n_1360),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1537),
.B(n_1351),
.Y(n_1557)
);

AO32x2_ASAP7_75t_L g1558 ( 
.A1(n_1498),
.A2(n_1455),
.A3(n_1368),
.B1(n_1441),
.B2(n_1450),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_1500),
.Y(n_1559)
);

OR2x6_ASAP7_75t_L g1560 ( 
.A(n_1478),
.B(n_1381),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1538),
.B(n_1460),
.Y(n_1561)
);

INVx4_ASAP7_75t_L g1562 ( 
.A(n_1479),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1491),
.B(n_1455),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1496),
.A2(n_1462),
.B1(n_1360),
.B2(n_1346),
.Y(n_1564)
);

AND2x4_ASAP7_75t_L g1565 ( 
.A(n_1485),
.B(n_1346),
.Y(n_1565)
);

OA21x2_ASAP7_75t_L g1566 ( 
.A1(n_1469),
.A2(n_1432),
.B(n_1458),
.Y(n_1566)
);

NOR4xp25_ASAP7_75t_SL g1567 ( 
.A(n_1497),
.B(n_1462),
.C(n_1432),
.D(n_1458),
.Y(n_1567)
);

AO21x2_ASAP7_75t_L g1568 ( 
.A1(n_1507),
.A2(n_1517),
.B(n_1520),
.Y(n_1568)
);

AOI221xp5_ASAP7_75t_L g1569 ( 
.A1(n_1508),
.A2(n_1489),
.B1(n_1519),
.B2(n_1517),
.C(n_1509),
.Y(n_1569)
);

AOI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1508),
.A2(n_1507),
.B1(n_1489),
.B2(n_1526),
.Y(n_1570)
);

INVx1_ASAP7_75t_SL g1571 ( 
.A(n_1542),
.Y(n_1571)
);

BUFx4f_ASAP7_75t_SL g1572 ( 
.A(n_1542),
.Y(n_1572)
);

NAND3xp33_ASAP7_75t_L g1573 ( 
.A(n_1527),
.B(n_1520),
.C(n_1509),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1470),
.B(n_1486),
.Y(n_1574)
);

INVxp67_ASAP7_75t_L g1575 ( 
.A(n_1491),
.Y(n_1575)
);

OA21x2_ASAP7_75t_L g1576 ( 
.A1(n_1469),
.A2(n_1480),
.B(n_1495),
.Y(n_1576)
);

O2A1O1Ixp33_ASAP7_75t_L g1577 ( 
.A1(n_1507),
.A2(n_1527),
.B(n_1481),
.C(n_1523),
.Y(n_1577)
);

OAI21xp33_ASAP7_75t_L g1578 ( 
.A1(n_1494),
.A2(n_1476),
.B(n_1475),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1533),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1505),
.B(n_1475),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1516),
.A2(n_1518),
.B1(n_1507),
.B2(n_1473),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1493),
.B(n_1499),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1483),
.B(n_1488),
.Y(n_1583)
);

A2O1A1Ixp33_ASAP7_75t_L g1584 ( 
.A1(n_1521),
.A2(n_1516),
.B(n_1473),
.C(n_1512),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1493),
.B(n_1499),
.Y(n_1585)
);

AO32x2_ASAP7_75t_L g1586 ( 
.A1(n_1536),
.A2(n_1543),
.A3(n_1479),
.B1(n_1530),
.B2(n_1494),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_L g1587 ( 
.A(n_1476),
.B(n_1523),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1512),
.A2(n_1532),
.B1(n_1518),
.B2(n_1472),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1468),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1513),
.B(n_1524),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1513),
.B(n_1524),
.Y(n_1591)
);

INVx4_ASAP7_75t_L g1592 ( 
.A(n_1535),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1521),
.A2(n_1472),
.B1(n_1532),
.B2(n_1522),
.Y(n_1593)
);

AO32x1_ASAP7_75t_L g1594 ( 
.A1(n_1490),
.A2(n_1528),
.A3(n_1525),
.B1(n_1506),
.B2(n_1510),
.Y(n_1594)
);

AO32x2_ASAP7_75t_L g1595 ( 
.A1(n_1530),
.A2(n_1504),
.A3(n_1506),
.B1(n_1510),
.B2(n_1488),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1551),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1582),
.B(n_1480),
.Y(n_1597)
);

BUFx2_ASAP7_75t_L g1598 ( 
.A(n_1544),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1585),
.B(n_1589),
.Y(n_1599)
);

OAI221xp5_ASAP7_75t_L g1600 ( 
.A1(n_1570),
.A2(n_1532),
.B1(n_1529),
.B2(n_1525),
.C(n_1482),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1544),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1595),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1595),
.Y(n_1603)
);

NAND2x1p5_ASAP7_75t_L g1604 ( 
.A(n_1592),
.B(n_1535),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1595),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1595),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1590),
.B(n_1502),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1591),
.B(n_1502),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_SL g1609 ( 
.A1(n_1573),
.A2(n_1532),
.B1(n_1514),
.B2(n_1530),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1544),
.B(n_1502),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1563),
.B(n_1492),
.Y(n_1611)
);

CKINVDCx20_ASAP7_75t_R g1612 ( 
.A(n_1559),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1544),
.B(n_1502),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1569),
.A2(n_1522),
.B1(n_1490),
.B2(n_1530),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1575),
.B(n_1580),
.Y(n_1615)
);

BUFx6f_ASAP7_75t_L g1616 ( 
.A(n_1576),
.Y(n_1616)
);

INVx2_ASAP7_75t_SL g1617 ( 
.A(n_1560),
.Y(n_1617)
);

OAI222xp33_ASAP7_75t_L g1618 ( 
.A1(n_1581),
.A2(n_1534),
.B1(n_1474),
.B2(n_1540),
.C1(n_1539),
.C2(n_1535),
.Y(n_1618)
);

BUFx2_ASAP7_75t_SL g1619 ( 
.A(n_1592),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1594),
.Y(n_1620)
);

NOR2xp67_ASAP7_75t_L g1621 ( 
.A(n_1587),
.B(n_1562),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1598),
.B(n_1575),
.Y(n_1622)
);

INVxp67_ASAP7_75t_SL g1623 ( 
.A(n_1616),
.Y(n_1623)
);

BUFx3_ASAP7_75t_L g1624 ( 
.A(n_1604),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1607),
.B(n_1586),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1616),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1607),
.B(n_1586),
.Y(n_1627)
);

INVxp67_ASAP7_75t_SL g1628 ( 
.A(n_1616),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1607),
.B(n_1586),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1596),
.Y(n_1630)
);

NAND3xp33_ASAP7_75t_L g1631 ( 
.A(n_1598),
.B(n_1546),
.C(n_1578),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1607),
.B(n_1586),
.Y(n_1632)
);

NOR2x1_ASAP7_75t_SL g1633 ( 
.A(n_1619),
.B(n_1560),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1608),
.B(n_1574),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1598),
.B(n_1552),
.Y(n_1635)
);

OA21x2_ASAP7_75t_L g1636 ( 
.A1(n_1620),
.A2(n_1584),
.B(n_1581),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1601),
.B(n_1587),
.Y(n_1637)
);

NAND4xp25_ASAP7_75t_SL g1638 ( 
.A(n_1612),
.B(n_1556),
.C(n_1555),
.D(n_1547),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1600),
.A2(n_1568),
.B1(n_1546),
.B2(n_1588),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1602),
.Y(n_1640)
);

INVx1_ASAP7_75t_SL g1641 ( 
.A(n_1615),
.Y(n_1641)
);

AO21x2_ASAP7_75t_L g1642 ( 
.A1(n_1620),
.A2(n_1577),
.B(n_1568),
.Y(n_1642)
);

INVx4_ASAP7_75t_L g1643 ( 
.A(n_1604),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1601),
.B(n_1583),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1620),
.Y(n_1645)
);

BUFx3_ASAP7_75t_L g1646 ( 
.A(n_1612),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1601),
.B(n_1579),
.Y(n_1647)
);

INVx3_ASAP7_75t_L g1648 ( 
.A(n_1616),
.Y(n_1648)
);

OAI221xp5_ASAP7_75t_L g1649 ( 
.A1(n_1600),
.A2(n_1555),
.B1(n_1584),
.B2(n_1588),
.C(n_1556),
.Y(n_1649)
);

AOI211xp5_ASAP7_75t_L g1650 ( 
.A1(n_1610),
.A2(n_1553),
.B(n_1564),
.C(n_1531),
.Y(n_1650)
);

INVxp67_ASAP7_75t_SL g1651 ( 
.A(n_1616),
.Y(n_1651)
);

AOI33xp33_ASAP7_75t_L g1652 ( 
.A1(n_1620),
.A2(n_1567),
.A3(n_1593),
.B1(n_1571),
.B2(n_1557),
.B3(n_1550),
.Y(n_1652)
);

BUFx3_ASAP7_75t_L g1653 ( 
.A(n_1617),
.Y(n_1653)
);

NAND3xp33_ASAP7_75t_L g1654 ( 
.A(n_1610),
.B(n_1566),
.C(n_1593),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1624),
.B(n_1621),
.Y(n_1655)
);

NOR2x1_ASAP7_75t_L g1656 ( 
.A(n_1638),
.B(n_1565),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1626),
.Y(n_1657)
);

NAND4xp25_ASAP7_75t_L g1658 ( 
.A(n_1650),
.B(n_1548),
.C(n_1610),
.D(n_1613),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1622),
.B(n_1602),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1640),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1622),
.B(n_1602),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1626),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1625),
.B(n_1608),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1640),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1626),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1625),
.B(n_1608),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1648),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1622),
.B(n_1602),
.Y(n_1668)
);

INVx3_ASAP7_75t_L g1669 ( 
.A(n_1643),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1635),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1635),
.Y(n_1671)
);

INVx1_ASAP7_75t_SL g1672 ( 
.A(n_1646),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1648),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1641),
.B(n_1603),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_SL g1675 ( 
.A(n_1652),
.B(n_1621),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1645),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1635),
.Y(n_1677)
);

NAND2x1p5_ASAP7_75t_L g1678 ( 
.A(n_1643),
.B(n_1566),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1630),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1641),
.B(n_1603),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1645),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1625),
.B(n_1627),
.Y(n_1682)
);

NAND4xp25_ASAP7_75t_L g1683 ( 
.A(n_1650),
.B(n_1610),
.C(n_1613),
.D(n_1611),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1644),
.B(n_1603),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1627),
.B(n_1599),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1646),
.B(n_1501),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1627),
.B(n_1599),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1630),
.Y(n_1688)
);

INVx2_ASAP7_75t_SL g1689 ( 
.A(n_1653),
.Y(n_1689)
);

INVx3_ASAP7_75t_L g1690 ( 
.A(n_1643),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1629),
.B(n_1599),
.Y(n_1691)
);

INVx4_ASAP7_75t_L g1692 ( 
.A(n_1646),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1624),
.B(n_1621),
.Y(n_1693)
);

INVx1_ASAP7_75t_SL g1694 ( 
.A(n_1645),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1676),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1672),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1682),
.B(n_1637),
.Y(n_1697)
);

NAND2x1p5_ASAP7_75t_L g1698 ( 
.A(n_1656),
.B(n_1692),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1676),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1681),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1681),
.Y(n_1701)
);

NAND3xp33_ASAP7_75t_L g1702 ( 
.A(n_1683),
.B(n_1631),
.C(n_1652),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1679),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_SL g1704 ( 
.A(n_1656),
.B(n_1631),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1694),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1682),
.B(n_1637),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1679),
.Y(n_1707)
);

AND2x4_ASAP7_75t_L g1708 ( 
.A(n_1692),
.B(n_1643),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1694),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1688),
.Y(n_1710)
);

OAI211xp5_ASAP7_75t_L g1711 ( 
.A1(n_1658),
.A2(n_1649),
.B(n_1639),
.C(n_1654),
.Y(n_1711)
);

INVx3_ASAP7_75t_SL g1712 ( 
.A(n_1692),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1672),
.B(n_1692),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1692),
.B(n_1629),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1688),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1670),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1682),
.B(n_1629),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1670),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1683),
.B(n_1644),
.Y(n_1719)
);

NAND2x1_ASAP7_75t_L g1720 ( 
.A(n_1689),
.B(n_1632),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1685),
.B(n_1632),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1685),
.B(n_1632),
.Y(n_1722)
);

NAND2xp67_ASAP7_75t_L g1723 ( 
.A(n_1674),
.B(n_1680),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1685),
.B(n_1597),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1671),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1671),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1663),
.B(n_1647),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1677),
.Y(n_1728)
);

AND3x2_ASAP7_75t_L g1729 ( 
.A(n_1686),
.B(n_1638),
.C(n_1565),
.Y(n_1729)
);

NAND2x1p5_ASAP7_75t_L g1730 ( 
.A(n_1669),
.B(n_1565),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1677),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1663),
.B(n_1647),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1660),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1663),
.B(n_1647),
.Y(n_1734)
);

INVx1_ASAP7_75t_SL g1735 ( 
.A(n_1675),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1687),
.B(n_1643),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1687),
.B(n_1597),
.Y(n_1737)
);

NAND2xp67_ASAP7_75t_L g1738 ( 
.A(n_1709),
.B(n_1666),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1703),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1698),
.B(n_1687),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1723),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1698),
.B(n_1691),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1717),
.B(n_1691),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1717),
.B(n_1730),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1707),
.Y(n_1745)
);

INVx3_ASAP7_75t_SL g1746 ( 
.A(n_1712),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1710),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1697),
.B(n_1658),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1730),
.B(n_1691),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1696),
.B(n_1666),
.Y(n_1750)
);

INVx1_ASAP7_75t_SL g1751 ( 
.A(n_1735),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1699),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1696),
.B(n_1666),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1721),
.B(n_1689),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1715),
.Y(n_1755)
);

OR2x6_ASAP7_75t_L g1756 ( 
.A(n_1704),
.B(n_1541),
.Y(n_1756)
);

NAND4xp25_ASAP7_75t_L g1757 ( 
.A(n_1702),
.B(n_1690),
.C(n_1669),
.D(n_1649),
.Y(n_1757)
);

INVx4_ASAP7_75t_L g1758 ( 
.A(n_1729),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1712),
.B(n_1559),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1721),
.B(n_1689),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1733),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1713),
.B(n_1503),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1706),
.B(n_1674),
.Y(n_1763)
);

AND3x2_ASAP7_75t_L g1764 ( 
.A(n_1705),
.B(n_1549),
.C(n_1611),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1722),
.B(n_1704),
.Y(n_1765)
);

NOR2xp67_ASAP7_75t_SL g1766 ( 
.A(n_1711),
.B(n_1654),
.Y(n_1766)
);

NOR2x1_ASAP7_75t_L g1767 ( 
.A(n_1709),
.B(n_1669),
.Y(n_1767)
);

NAND2x1_ASAP7_75t_SL g1768 ( 
.A(n_1705),
.B(n_1669),
.Y(n_1768)
);

INVx1_ASAP7_75t_SL g1769 ( 
.A(n_1729),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1722),
.B(n_1669),
.Y(n_1770)
);

NAND3xp33_ASAP7_75t_L g1771 ( 
.A(n_1719),
.B(n_1664),
.C(n_1660),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1716),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1708),
.B(n_1690),
.Y(n_1773)
);

AND2x4_ASAP7_75t_SL g1774 ( 
.A(n_1759),
.B(n_1561),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1765),
.B(n_1708),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1766),
.B(n_1714),
.Y(n_1776)
);

AOI222xp33_ASAP7_75t_L g1777 ( 
.A1(n_1766),
.A2(n_1613),
.B1(n_1603),
.B2(n_1606),
.C1(n_1605),
.C2(n_1639),
.Y(n_1777)
);

AOI221xp5_ASAP7_75t_L g1778 ( 
.A1(n_1771),
.A2(n_1684),
.B1(n_1606),
.B2(n_1605),
.C(n_1680),
.Y(n_1778)
);

NAND3xp33_ASAP7_75t_SL g1779 ( 
.A(n_1769),
.B(n_1720),
.C(n_1699),
.Y(n_1779)
);

NAND2xp33_ASAP7_75t_R g1780 ( 
.A(n_1764),
.B(n_1708),
.Y(n_1780)
);

AO22x1_ASAP7_75t_L g1781 ( 
.A1(n_1758),
.A2(n_1695),
.B1(n_1700),
.B2(n_1701),
.Y(n_1781)
);

NOR2xp67_ASAP7_75t_L g1782 ( 
.A(n_1758),
.B(n_1736),
.Y(n_1782)
);

OAI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1756),
.A2(n_1636),
.B1(n_1605),
.B2(n_1606),
.Y(n_1783)
);

NOR2xp33_ASAP7_75t_L g1784 ( 
.A(n_1751),
.B(n_1736),
.Y(n_1784)
);

OAI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1758),
.A2(n_1727),
.B1(n_1734),
.B2(n_1732),
.Y(n_1785)
);

OAI21xp33_ASAP7_75t_SL g1786 ( 
.A1(n_1768),
.A2(n_1765),
.B(n_1757),
.Y(n_1786)
);

A2O1A1Ixp33_ASAP7_75t_L g1787 ( 
.A1(n_1748),
.A2(n_1606),
.B(n_1605),
.C(n_1613),
.Y(n_1787)
);

AOI222xp33_ASAP7_75t_L g1788 ( 
.A1(n_1771),
.A2(n_1684),
.B1(n_1614),
.B2(n_1664),
.C1(n_1616),
.C2(n_1618),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1746),
.B(n_1736),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1750),
.B(n_1753),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1748),
.B(n_1718),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1758),
.A2(n_1636),
.B1(n_1642),
.B2(n_1609),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1768),
.Y(n_1793)
);

AOI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1756),
.A2(n_1636),
.B1(n_1642),
.B2(n_1609),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_L g1795 ( 
.A1(n_1756),
.A2(n_1636),
.B1(n_1642),
.B2(n_1616),
.Y(n_1795)
);

OAI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1767),
.A2(n_1726),
.B(n_1725),
.Y(n_1796)
);

AOI21xp33_ASAP7_75t_L g1797 ( 
.A1(n_1741),
.A2(n_1731),
.B(n_1728),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1739),
.Y(n_1798)
);

OR2x6_ASAP7_75t_L g1799 ( 
.A(n_1752),
.B(n_1541),
.Y(n_1799)
);

OAI32xp33_ASAP7_75t_L g1800 ( 
.A1(n_1786),
.A2(n_1741),
.A3(n_1763),
.B1(n_1740),
.B2(n_1742),
.Y(n_1800)
);

AOI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1777),
.A2(n_1756),
.B1(n_1636),
.B2(n_1642),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1798),
.Y(n_1802)
);

OAI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1776),
.A2(n_1756),
.B1(n_1767),
.B2(n_1741),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1775),
.B(n_1754),
.Y(n_1804)
);

AOI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1788),
.A2(n_1642),
.B1(n_1740),
.B2(n_1742),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1781),
.A2(n_1752),
.B(n_1761),
.Y(n_1806)
);

BUFx3_ASAP7_75t_L g1807 ( 
.A(n_1784),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1785),
.Y(n_1808)
);

A2O1A1Ixp33_ASAP7_75t_L g1809 ( 
.A1(n_1794),
.A2(n_1668),
.B(n_1661),
.C(n_1659),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1774),
.B(n_1746),
.Y(n_1810)
);

OAI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1779),
.A2(n_1752),
.B(n_1761),
.Y(n_1811)
);

INVxp67_ASAP7_75t_L g1812 ( 
.A(n_1789),
.Y(n_1812)
);

AOI322xp5_ASAP7_75t_L g1813 ( 
.A1(n_1783),
.A2(n_1743),
.A3(n_1772),
.B1(n_1744),
.B2(n_1724),
.C1(n_1737),
.C2(n_1749),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1793),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1799),
.Y(n_1815)
);

AOI221xp5_ASAP7_75t_L g1816 ( 
.A1(n_1778),
.A2(n_1772),
.B1(n_1747),
.B2(n_1739),
.C(n_1745),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1791),
.B(n_1763),
.Y(n_1817)
);

OAI322xp33_ASAP7_75t_L g1818 ( 
.A1(n_1790),
.A2(n_1792),
.A3(n_1780),
.B1(n_1755),
.B2(n_1747),
.C1(n_1745),
.C2(n_1661),
.Y(n_1818)
);

AOI211xp5_ASAP7_75t_L g1819 ( 
.A1(n_1782),
.A2(n_1746),
.B(n_1755),
.C(n_1744),
.Y(n_1819)
);

OAI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1808),
.A2(n_1787),
.B1(n_1795),
.B2(n_1796),
.Y(n_1820)
);

AOI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1805),
.A2(n_1797),
.B1(n_1799),
.B2(n_1754),
.Y(n_1821)
);

NAND3xp33_ASAP7_75t_L g1822 ( 
.A(n_1811),
.B(n_1760),
.C(n_1799),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1817),
.Y(n_1823)
);

AOI322xp5_ASAP7_75t_L g1824 ( 
.A1(n_1801),
.A2(n_1743),
.A3(n_1760),
.B1(n_1749),
.B2(n_1738),
.C1(n_1770),
.C2(n_1614),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1802),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1804),
.B(n_1770),
.Y(n_1826)
);

AND2x4_ASAP7_75t_L g1827 ( 
.A(n_1807),
.B(n_1773),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1814),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_SL g1829 ( 
.A(n_1819),
.B(n_1773),
.Y(n_1829)
);

AOI22xp33_ASAP7_75t_L g1830 ( 
.A1(n_1818),
.A2(n_1616),
.B1(n_1566),
.B2(n_1661),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1806),
.Y(n_1831)
);

AOI22xp5_ASAP7_75t_L g1832 ( 
.A1(n_1820),
.A2(n_1815),
.B1(n_1811),
.B2(n_1816),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1823),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1827),
.Y(n_1834)
);

NOR2xp33_ASAP7_75t_L g1835 ( 
.A(n_1827),
.B(n_1812),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1828),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1831),
.B(n_1813),
.Y(n_1837)
);

AND3x1_ASAP7_75t_L g1838 ( 
.A(n_1825),
.B(n_1810),
.C(n_1762),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1826),
.B(n_1738),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1829),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1822),
.Y(n_1841)
);

INVxp67_ASAP7_75t_L g1842 ( 
.A(n_1821),
.Y(n_1842)
);

O2A1O1Ixp33_ASAP7_75t_L g1843 ( 
.A1(n_1837),
.A2(n_1800),
.B(n_1803),
.C(n_1809),
.Y(n_1843)
);

OAI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1837),
.A2(n_1830),
.B1(n_1803),
.B2(n_1821),
.Y(n_1844)
);

OAI211xp5_ASAP7_75t_L g1845 ( 
.A1(n_1840),
.A2(n_1824),
.B(n_1690),
.C(n_1623),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1832),
.A2(n_1668),
.B(n_1659),
.Y(n_1846)
);

OAI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1841),
.A2(n_1668),
.B1(n_1659),
.B2(n_1678),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1834),
.B(n_1634),
.Y(n_1848)
);

AOI211xp5_ASAP7_75t_SL g1849 ( 
.A1(n_1845),
.A2(n_1835),
.B(n_1833),
.C(n_1836),
.Y(n_1849)
);

OAI221xp5_ASAP7_75t_SL g1850 ( 
.A1(n_1843),
.A2(n_1842),
.B1(n_1839),
.B2(n_1838),
.C(n_1690),
.Y(n_1850)
);

XOR2xp5_ASAP7_75t_L g1851 ( 
.A(n_1844),
.B(n_1531),
.Y(n_1851)
);

AOI221xp5_ASAP7_75t_L g1852 ( 
.A1(n_1846),
.A2(n_1651),
.B1(n_1628),
.B2(n_1623),
.C(n_1616),
.Y(n_1852)
);

INVx1_ASAP7_75t_SL g1853 ( 
.A(n_1848),
.Y(n_1853)
);

HB1xp67_ASAP7_75t_L g1854 ( 
.A(n_1847),
.Y(n_1854)
);

BUFx2_ASAP7_75t_SL g1855 ( 
.A(n_1848),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_L g1856 ( 
.A(n_1850),
.B(n_1690),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1855),
.B(n_1628),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1853),
.A2(n_1678),
.B1(n_1657),
.B2(n_1662),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1849),
.B(n_1634),
.Y(n_1859)
);

XOR2xp5_ASAP7_75t_SL g1860 ( 
.A(n_1854),
.B(n_1558),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1859),
.B(n_1851),
.Y(n_1861)
);

OAI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1857),
.A2(n_1852),
.B1(n_1678),
.B2(n_1665),
.Y(n_1862)
);

OAI221xp5_ASAP7_75t_L g1863 ( 
.A1(n_1856),
.A2(n_1858),
.B1(n_1860),
.B2(n_1678),
.C(n_1651),
.Y(n_1863)
);

NOR2xp33_ASAP7_75t_SL g1864 ( 
.A(n_1861),
.B(n_1572),
.Y(n_1864)
);

OA22x2_ASAP7_75t_L g1865 ( 
.A1(n_1864),
.A2(n_1862),
.B1(n_1863),
.B2(n_1673),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1865),
.Y(n_1866)
);

XOR2x1_ASAP7_75t_L g1867 ( 
.A(n_1865),
.B(n_1655),
.Y(n_1867)
);

OAI322xp33_ASAP7_75t_L g1868 ( 
.A1(n_1866),
.A2(n_1867),
.A3(n_1657),
.B1(n_1662),
.B2(n_1665),
.C1(n_1667),
.C2(n_1673),
.Y(n_1868)
);

OAI31xp33_ASAP7_75t_L g1869 ( 
.A1(n_1867),
.A2(n_1665),
.A3(n_1662),
.B(n_1657),
.Y(n_1869)
);

OAI22xp33_ASAP7_75t_L g1870 ( 
.A1(n_1869),
.A2(n_1673),
.B1(n_1667),
.B2(n_1572),
.Y(n_1870)
);

AO21x2_ASAP7_75t_L g1871 ( 
.A1(n_1868),
.A2(n_1667),
.B(n_1633),
.Y(n_1871)
);

AOI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1870),
.A2(n_1693),
.B(n_1655),
.Y(n_1872)
);

OAI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1872),
.A2(n_1871),
.B(n_1693),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_SL g1874 ( 
.A1(n_1873),
.A2(n_1558),
.B1(n_1693),
.B2(n_1655),
.Y(n_1874)
);

OAI221xp5_ASAP7_75t_L g1875 ( 
.A1(n_1874),
.A2(n_1558),
.B1(n_1529),
.B2(n_1648),
.C(n_1653),
.Y(n_1875)
);

AOI211xp5_ASAP7_75t_L g1876 ( 
.A1(n_1875),
.A2(n_1558),
.B(n_1545),
.C(n_1554),
.Y(n_1876)
);


endmodule