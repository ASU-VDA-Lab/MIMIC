module fake_netlist_1_11595_n_29 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_29);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
INVx1_ASAP7_75t_L g13 ( .A(n_7), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_8), .B(n_2), .Y(n_14) );
OA21x2_ASAP7_75t_L g15 ( .A1(n_5), .A2(n_9), .B(n_2), .Y(n_15) );
NOR2xp33_ASAP7_75t_R g16 ( .A(n_4), .B(n_1), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_12), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_4), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_13), .B(n_0), .Y(n_19) );
NAND2xp33_ASAP7_75t_SL g20 ( .A(n_16), .B(n_0), .Y(n_20) );
AOI22xp33_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_18), .B1(n_14), .B2(n_15), .Y(n_21) );
AND2x4_ASAP7_75t_L g22 ( .A(n_19), .B(n_18), .Y(n_22) );
OAI22xp5_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_18), .B1(n_13), .B2(n_14), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_23), .B(n_22), .Y(n_24) );
OAI22xp5_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_22), .B1(n_17), .B2(n_15), .Y(n_25) );
OAI211xp5_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_15), .B(n_22), .C(n_1), .Y(n_26) );
NOR2x1p5_ASAP7_75t_L g27 ( .A(n_26), .B(n_3), .Y(n_27) );
BUFx2_ASAP7_75t_SL g28 ( .A(n_27), .Y(n_28) );
AOI322xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_3), .A3(n_6), .B1(n_10), .B2(n_11), .C1(n_15), .C2(n_20), .Y(n_29) );
endmodule