module fake_jpeg_27070_n_5 (n_0, n_1, n_5);

input n_0;
input n_1;

output n_5;

wire n_3;
wire n_2;
wire n_4;

AND2x2_ASAP7_75t_L g2 ( 
.A(n_1),
.B(n_0),
.Y(n_2)
);

AND2x2_ASAP7_75t_L g3 ( 
.A(n_2),
.B(n_0),
.Y(n_3)
);

CKINVDCx16_ASAP7_75t_R g4 ( 
.A(n_3),
.Y(n_4)
);

NOR3xp33_ASAP7_75t_L g5 ( 
.A(n_4),
.B(n_2),
.C(n_1),
.Y(n_5)
);


endmodule