module real_aes_6858_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_449;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g105 ( .A(n_0), .Y(n_105) );
INVx1_ASAP7_75t_L g455 ( .A(n_1), .Y(n_455) );
INVx1_ASAP7_75t_L g258 ( .A(n_2), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_3), .A2(n_36), .B1(n_208), .B2(n_494), .Y(n_530) );
AOI21xp33_ASAP7_75t_L g219 ( .A1(n_4), .A2(n_141), .B(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_5), .B(n_163), .Y(n_480) );
AND2x6_ASAP7_75t_L g146 ( .A(n_6), .B(n_147), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_7), .A2(n_140), .B(n_148), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_8), .B(n_111), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g122 ( .A(n_8), .B(n_37), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_9), .B(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g225 ( .A(n_10), .Y(n_225) );
INVx1_ASAP7_75t_L g138 ( .A(n_11), .Y(n_138) );
INVx1_ASAP7_75t_L g449 ( .A(n_12), .Y(n_449) );
INVx1_ASAP7_75t_L g158 ( .A(n_13), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_14), .B(n_232), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_15), .B(n_164), .Y(n_482) );
AO32x2_ASAP7_75t_L g528 ( .A1(n_16), .A2(n_163), .A3(n_179), .B1(n_468), .B2(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_17), .B(n_208), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_18), .B(n_175), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_19), .B(n_164), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_20), .A2(n_48), .B1(n_208), .B2(n_494), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_21), .B(n_141), .Y(n_168) );
AOI22xp33_ASAP7_75t_SL g495 ( .A1(n_22), .A2(n_73), .B1(n_208), .B2(n_232), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_23), .B(n_208), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_24), .B(n_218), .Y(n_248) );
A2O1A1Ixp33_ASAP7_75t_L g154 ( .A1(n_25), .A2(n_155), .B(n_157), .C(n_159), .Y(n_154) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_26), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_27), .B(n_134), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_28), .B(n_190), .Y(n_259) );
AOI222xp33_ASAP7_75t_SL g124 ( .A1(n_29), .A2(n_88), .B1(n_125), .B2(n_714), .C1(n_715), .C2(n_718), .Y(n_124) );
INVx1_ASAP7_75t_L g714 ( .A(n_29), .Y(n_714) );
INVx1_ASAP7_75t_L g237 ( .A(n_30), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_31), .B(n_134), .Y(n_506) );
INVx2_ASAP7_75t_L g144 ( .A(n_32), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_33), .B(n_208), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_34), .B(n_134), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g169 ( .A1(n_35), .A2(n_146), .B(n_151), .C(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g111 ( .A(n_37), .Y(n_111) );
INVx1_ASAP7_75t_L g235 ( .A(n_38), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_39), .B(n_190), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_40), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_41), .B(n_208), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_42), .A2(n_84), .B1(n_160), .B2(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_43), .B(n_208), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_44), .B(n_208), .Y(n_450) );
CKINVDCx16_ASAP7_75t_R g238 ( .A(n_45), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_46), .B(n_454), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_47), .B(n_141), .Y(n_209) );
AOI22xp33_ASAP7_75t_SL g486 ( .A1(n_49), .A2(n_58), .B1(n_208), .B2(n_232), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_50), .A2(n_151), .B1(n_232), .B2(n_234), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_51), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_52), .B(n_208), .Y(n_467) );
CKINVDCx16_ASAP7_75t_R g255 ( .A(n_53), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_54), .B(n_208), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_55), .A2(n_223), .B(n_224), .C(n_226), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_56), .Y(n_194) );
INVx1_ASAP7_75t_L g221 ( .A(n_57), .Y(n_221) );
INVx1_ASAP7_75t_L g147 ( .A(n_59), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_60), .B(n_208), .Y(n_456) );
INVx1_ASAP7_75t_L g137 ( .A(n_61), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_62), .Y(n_116) );
AO32x2_ASAP7_75t_L g491 ( .A1(n_63), .A2(n_163), .A3(n_200), .B1(n_468), .B2(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g466 ( .A(n_64), .Y(n_466) );
INVx1_ASAP7_75t_L g501 ( .A(n_65), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_SL g245 ( .A1(n_66), .A2(n_175), .B(n_226), .C(n_246), .Y(n_245) );
INVxp67_ASAP7_75t_L g247 ( .A(n_67), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_68), .B(n_232), .Y(n_502) );
INVx1_ASAP7_75t_L g108 ( .A(n_69), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_70), .Y(n_240) );
INVx1_ASAP7_75t_L g185 ( .A(n_71), .Y(n_185) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_72), .A2(n_127), .B1(n_716), .B2(n_726), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_72), .Y(n_726) );
A2O1A1Ixp33_ASAP7_75t_L g187 ( .A1(n_74), .A2(n_146), .B(n_151), .C(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_75), .B(n_494), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_76), .B(n_232), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_77), .A2(n_100), .B1(n_112), .B2(n_729), .Y(n_99) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_78), .B(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g135 ( .A(n_79), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_80), .B(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_81), .B(n_232), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_82), .A2(n_146), .B(n_151), .C(n_257), .Y(n_256) );
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_83), .B(n_105), .C(n_106), .Y(n_104) );
OR2x2_ASAP7_75t_L g119 ( .A(n_83), .B(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g126 ( .A(n_83), .B(n_121), .Y(n_126) );
INVx2_ASAP7_75t_L g438 ( .A(n_83), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_85), .A2(n_98), .B1(n_232), .B2(n_233), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_86), .B(n_134), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g262 ( .A(n_87), .Y(n_262) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_89), .A2(n_146), .B(n_151), .C(n_203), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_90), .Y(n_211) );
INVx1_ASAP7_75t_L g244 ( .A(n_91), .Y(n_244) );
CKINVDCx16_ASAP7_75t_R g149 ( .A(n_92), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_93), .B(n_172), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_94), .B(n_232), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_95), .B(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_96), .B(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_97), .A2(n_141), .B(n_243), .Y(n_242) );
INVx1_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx2_ASAP7_75t_SL g731 ( .A(n_102), .Y(n_731) );
AND2x2_ASAP7_75t_SL g102 ( .A(n_103), .B(n_109), .Y(n_102) );
CKINVDCx16_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_L g121 ( .A(n_105), .B(n_122), .Y(n_121) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVxp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AOI22x1_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_124), .B1(n_721), .B2(n_724), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_117), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g723 ( .A(n_116), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g724 ( .A1(n_117), .A2(n_725), .B(n_727), .Y(n_724) );
NOR2xp33_ASAP7_75t_SL g117 ( .A(n_118), .B(n_123), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g728 ( .A(n_119), .Y(n_728) );
NOR2x2_ASAP7_75t_L g720 ( .A(n_120), .B(n_438), .Y(n_720) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g437 ( .A(n_121), .B(n_438), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_127), .B1(n_435), .B2(n_439), .Y(n_125) );
OAI22xp5_ASAP7_75t_SL g715 ( .A1(n_126), .A2(n_437), .B1(n_716), .B2(n_717), .Y(n_715) );
INVx2_ASAP7_75t_SL g716 ( .A(n_127), .Y(n_716) );
OR4x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_331), .C(n_390), .D(n_417), .Y(n_127) );
NAND3xp33_ASAP7_75t_SL g128 ( .A(n_129), .B(n_273), .C(n_298), .Y(n_128) );
O2A1O1Ixp33_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_196), .B(n_216), .C(n_249), .Y(n_129) );
AOI211xp5_ASAP7_75t_SL g421 ( .A1(n_130), .A2(n_422), .B(n_424), .C(n_427), .Y(n_421) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_165), .Y(n_130) );
INVx1_ASAP7_75t_L g296 ( .A(n_131), .Y(n_296) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OR2x2_ASAP7_75t_L g271 ( .A(n_132), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g303 ( .A(n_132), .Y(n_303) );
AND2x2_ASAP7_75t_L g358 ( .A(n_132), .B(n_327), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_132), .B(n_214), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_132), .B(n_215), .Y(n_416) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g277 ( .A(n_133), .Y(n_277) );
AND2x2_ASAP7_75t_L g320 ( .A(n_133), .B(n_183), .Y(n_320) );
AND2x2_ASAP7_75t_L g338 ( .A(n_133), .B(n_215), .Y(n_338) );
OA21x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_139), .B(n_162), .Y(n_133) );
INVx1_ASAP7_75t_L g195 ( .A(n_134), .Y(n_195) );
INVx2_ASAP7_75t_L g200 ( .A(n_134), .Y(n_200) );
OA21x2_ASAP7_75t_L g498 ( .A1(n_134), .A2(n_499), .B(n_506), .Y(n_498) );
OA21x2_ASAP7_75t_L g507 ( .A1(n_134), .A2(n_508), .B(n_516), .Y(n_507) );
AND2x2_ASAP7_75t_SL g134 ( .A(n_135), .B(n_136), .Y(n_134) );
AND2x2_ASAP7_75t_L g164 ( .A(n_135), .B(n_136), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
BUFx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_146), .Y(n_141) );
NAND2x1p5_ASAP7_75t_L g186 ( .A(n_142), .B(n_146), .Y(n_186) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_145), .Y(n_142) );
INVx1_ASAP7_75t_L g454 ( .A(n_143), .Y(n_454) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g152 ( .A(n_144), .Y(n_152) );
INVx1_ASAP7_75t_L g233 ( .A(n_144), .Y(n_233) );
INVx1_ASAP7_75t_L g153 ( .A(n_145), .Y(n_153) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_145), .Y(n_156) );
INVx3_ASAP7_75t_L g173 ( .A(n_145), .Y(n_173) );
INVx1_ASAP7_75t_L g175 ( .A(n_145), .Y(n_175) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_145), .Y(n_190) );
INVx4_ASAP7_75t_SL g161 ( .A(n_146), .Y(n_161) );
OAI21xp5_ASAP7_75t_L g447 ( .A1(n_146), .A2(n_448), .B(n_452), .Y(n_447) );
BUFx3_ASAP7_75t_L g468 ( .A(n_146), .Y(n_468) );
OAI21xp5_ASAP7_75t_L g473 ( .A1(n_146), .A2(n_474), .B(n_477), .Y(n_473) );
OAI21xp5_ASAP7_75t_L g499 ( .A1(n_146), .A2(n_500), .B(n_503), .Y(n_499) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_146), .A2(n_509), .B(n_513), .Y(n_508) );
O2A1O1Ixp33_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B(n_154), .C(n_161), .Y(n_148) );
O2A1O1Ixp33_ASAP7_75t_L g220 ( .A1(n_150), .A2(n_161), .B(n_221), .C(n_222), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_150), .A2(n_161), .B(n_244), .C(n_245), .Y(n_243) );
INVx5_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x6_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
BUFx3_ASAP7_75t_L g160 ( .A(n_152), .Y(n_160) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_152), .Y(n_208) );
INVx1_ASAP7_75t_L g494 ( .A(n_152), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_155), .B(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g451 ( .A(n_155), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_155), .A2(n_504), .B(n_505), .Y(n_503) );
INVx4_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
OAI22xp5_ASAP7_75t_SL g234 ( .A1(n_156), .A2(n_235), .B1(n_236), .B2(n_237), .Y(n_234) );
INVx2_ASAP7_75t_L g236 ( .A(n_156), .Y(n_236) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g177 ( .A(n_160), .Y(n_177) );
OAI22xp33_ASAP7_75t_L g230 ( .A1(n_161), .A2(n_186), .B1(n_231), .B2(n_238), .Y(n_230) );
INVx4_ASAP7_75t_L g182 ( .A(n_163), .Y(n_182) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_163), .A2(n_242), .B(n_248), .Y(n_241) );
OA21x2_ASAP7_75t_L g472 ( .A1(n_163), .A2(n_473), .B(n_480), .Y(n_472) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g179 ( .A(n_164), .Y(n_179) );
INVx4_ASAP7_75t_L g270 ( .A(n_165), .Y(n_270) );
OAI21xp5_ASAP7_75t_L g325 ( .A1(n_165), .A2(n_326), .B(n_328), .Y(n_325) );
AND2x2_ASAP7_75t_L g406 ( .A(n_165), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_183), .Y(n_165) );
INVx1_ASAP7_75t_L g213 ( .A(n_166), .Y(n_213) );
AND2x2_ASAP7_75t_L g275 ( .A(n_166), .B(n_215), .Y(n_275) );
OR2x2_ASAP7_75t_L g304 ( .A(n_166), .B(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g318 ( .A(n_166), .Y(n_318) );
INVx3_ASAP7_75t_L g327 ( .A(n_166), .Y(n_327) );
AND2x2_ASAP7_75t_L g337 ( .A(n_166), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g370 ( .A(n_166), .B(n_276), .Y(n_370) );
AND2x2_ASAP7_75t_L g394 ( .A(n_166), .B(n_350), .Y(n_394) );
OR2x6_ASAP7_75t_L g166 ( .A(n_167), .B(n_180), .Y(n_166) );
AOI21xp5_ASAP7_75t_SL g167 ( .A1(n_168), .A2(n_169), .B(n_178), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_174), .B(n_176), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_L g257 ( .A1(n_172), .A2(n_258), .B(n_259), .C(n_260), .Y(n_257) );
INVx2_ASAP7_75t_L g457 ( .A(n_172), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_172), .A2(n_463), .B(n_464), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_172), .A2(n_475), .B(n_476), .Y(n_474) );
O2A1O1Ixp5_ASAP7_75t_SL g500 ( .A1(n_172), .A2(n_226), .B(n_501), .C(n_502), .Y(n_500) );
INVx5_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_173), .B(n_225), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_173), .B(n_247), .Y(n_246) );
OAI22xp5_ASAP7_75t_SL g492 ( .A1(n_173), .A2(n_190), .B1(n_493), .B2(n_495), .Y(n_492) );
INVx1_ASAP7_75t_L g512 ( .A(n_175), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_176), .A2(n_189), .B(n_191), .Y(n_188) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g192 ( .A(n_178), .Y(n_192) );
OA21x2_ASAP7_75t_L g446 ( .A1(n_178), .A2(n_447), .B(n_458), .Y(n_446) );
OA21x2_ASAP7_75t_L g460 ( .A1(n_178), .A2(n_461), .B(n_469), .Y(n_460) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_179), .A2(n_230), .B(n_239), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_179), .B(n_240), .Y(n_239) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_179), .A2(n_254), .B(n_261), .Y(n_253) );
NOR2xp33_ASAP7_75t_SL g180 ( .A(n_181), .B(n_182), .Y(n_180) );
INVx3_ASAP7_75t_L g218 ( .A(n_182), .Y(n_218) );
NAND3xp33_ASAP7_75t_L g483 ( .A(n_182), .B(n_468), .C(n_484), .Y(n_483) );
AO21x1_ASAP7_75t_L g562 ( .A1(n_182), .A2(n_484), .B(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g215 ( .A(n_183), .Y(n_215) );
AND2x2_ASAP7_75t_L g430 ( .A(n_183), .B(n_272), .Y(n_430) );
AO21x2_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_192), .B(n_193), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_187), .Y(n_184) );
OAI21xp5_ASAP7_75t_L g254 ( .A1(n_186), .A2(n_255), .B(n_256), .Y(n_254) );
INVx4_ASAP7_75t_L g206 ( .A(n_190), .Y(n_206) );
INVx2_ASAP7_75t_L g223 ( .A(n_190), .Y(n_223) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_190), .A2(n_457), .B1(n_485), .B2(n_486), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_190), .A2(n_457), .B1(n_530), .B2(n_531), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_195), .B(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_195), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_212), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_198), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g350 ( .A(n_198), .B(n_338), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_198), .B(n_327), .Y(n_412) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g272 ( .A(n_199), .Y(n_272) );
AND2x2_ASAP7_75t_L g276 ( .A(n_199), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g317 ( .A(n_199), .B(n_318), .Y(n_317) );
AO21x2_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B(n_210), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_202), .B(n_209), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_207), .Y(n_203) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx3_ASAP7_75t_L g226 ( .A(n_208), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_212), .B(n_313), .Y(n_335) );
INVx1_ASAP7_75t_L g374 ( .A(n_212), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_212), .B(n_301), .Y(n_418) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
AND2x2_ASAP7_75t_L g281 ( .A(n_213), .B(n_276), .Y(n_281) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_215), .B(n_272), .Y(n_305) );
INVx1_ASAP7_75t_L g384 ( .A(n_215), .Y(n_384) );
AOI322xp5_ASAP7_75t_L g408 ( .A1(n_216), .A2(n_323), .A3(n_383), .B1(n_409), .B2(n_411), .C1(n_413), .C2(n_415), .Y(n_408) );
AND2x2_ASAP7_75t_SL g216 ( .A(n_217), .B(n_228), .Y(n_216) );
AND2x2_ASAP7_75t_L g263 ( .A(n_217), .B(n_241), .Y(n_263) );
INVx1_ASAP7_75t_SL g266 ( .A(n_217), .Y(n_266) );
AND2x2_ASAP7_75t_L g268 ( .A(n_217), .B(n_229), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_217), .B(n_285), .Y(n_291) );
INVx2_ASAP7_75t_L g310 ( .A(n_217), .Y(n_310) );
AND2x2_ASAP7_75t_L g323 ( .A(n_217), .B(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g361 ( .A(n_217), .B(n_285), .Y(n_361) );
BUFx2_ASAP7_75t_L g378 ( .A(n_217), .Y(n_378) );
AND2x2_ASAP7_75t_L g392 ( .A(n_217), .B(n_252), .Y(n_392) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_227), .Y(n_217) );
O2A1O1Ixp5_ASAP7_75t_L g465 ( .A1(n_223), .A2(n_453), .B(n_466), .C(n_467), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_223), .A2(n_514), .B(n_515), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_228), .B(n_280), .Y(n_307) );
AND2x2_ASAP7_75t_L g434 ( .A(n_228), .B(n_310), .Y(n_434) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_241), .Y(n_228) );
OR2x2_ASAP7_75t_L g279 ( .A(n_229), .B(n_280), .Y(n_279) );
INVx3_ASAP7_75t_L g285 ( .A(n_229), .Y(n_285) );
AND2x2_ASAP7_75t_L g330 ( .A(n_229), .B(n_253), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_229), .B(n_378), .Y(n_377) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_229), .Y(n_414) );
INVx2_ASAP7_75t_L g260 ( .A(n_232), .Y(n_260) );
INVx3_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g265 ( .A(n_241), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g287 ( .A(n_241), .Y(n_287) );
BUFx2_ASAP7_75t_L g293 ( .A(n_241), .Y(n_293) );
AND2x2_ASAP7_75t_L g312 ( .A(n_241), .B(n_285), .Y(n_312) );
INVx3_ASAP7_75t_L g324 ( .A(n_241), .Y(n_324) );
OR2x2_ASAP7_75t_L g334 ( .A(n_241), .B(n_285), .Y(n_334) );
AOI31xp33_ASAP7_75t_SL g249 ( .A1(n_250), .A2(n_264), .A3(n_267), .B(n_269), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_263), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_251), .B(n_286), .Y(n_297) );
OR2x2_ASAP7_75t_L g321 ( .A(n_251), .B(n_291), .Y(n_321) );
INVx1_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_252), .B(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g342 ( .A(n_252), .B(n_334), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_252), .B(n_324), .Y(n_352) );
AND2x2_ASAP7_75t_L g359 ( .A(n_252), .B(n_360), .Y(n_359) );
NAND2x1_ASAP7_75t_L g387 ( .A(n_252), .B(n_323), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_252), .B(n_378), .Y(n_388) );
AND2x2_ASAP7_75t_L g400 ( .A(n_252), .B(n_285), .Y(n_400) );
INVx3_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx3_ASAP7_75t_L g280 ( .A(n_253), .Y(n_280) );
O2A1O1Ixp33_ASAP7_75t_L g448 ( .A1(n_260), .A2(n_449), .B(n_450), .C(n_451), .Y(n_448) );
INVx1_ASAP7_75t_L g346 ( .A(n_263), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_263), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_265), .B(n_341), .Y(n_375) );
AND2x4_ASAP7_75t_L g286 ( .A(n_266), .B(n_287), .Y(n_286) );
CKINVDCx16_ASAP7_75t_R g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx2_ASAP7_75t_L g365 ( .A(n_271), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_271), .B(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g313 ( .A(n_272), .B(n_303), .Y(n_313) );
AND2x2_ASAP7_75t_L g407 ( .A(n_272), .B(n_277), .Y(n_407) );
INVx1_ASAP7_75t_L g432 ( .A(n_272), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_278), .B1(n_281), .B2(n_282), .C(n_288), .Y(n_273) );
CKINVDCx14_ASAP7_75t_R g294 ( .A(n_274), .Y(n_294) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_275), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_278), .B(n_329), .Y(n_348) );
INVx3_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g397 ( .A(n_279), .B(n_293), .Y(n_397) );
AND2x2_ASAP7_75t_L g311 ( .A(n_280), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g341 ( .A(n_280), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_280), .B(n_324), .Y(n_369) );
NOR3xp33_ASAP7_75t_L g411 ( .A(n_280), .B(n_381), .C(n_412), .Y(n_411) );
AOI211xp5_ASAP7_75t_SL g344 ( .A1(n_281), .A2(n_345), .B(n_347), .C(n_355), .Y(n_344) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OAI22xp33_ASAP7_75t_L g333 ( .A1(n_283), .A2(n_334), .B1(n_335), .B2(n_336), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_284), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_284), .B(n_368), .Y(n_367) );
BUFx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g426 ( .A(n_286), .B(n_400), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_294), .B1(n_295), .B2(n_297), .Y(n_288) );
NOR2xp33_ASAP7_75t_SL g289 ( .A(n_290), .B(n_292), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_292), .B(n_341), .Y(n_372) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_295), .A2(n_387), .B1(n_418), .B2(n_425), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_306), .B1(n_308), .B2(n_313), .C(n_314), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_304), .Y(n_300) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVxp67_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OAI221xp5_ASAP7_75t_L g314 ( .A1(n_304), .A2(n_315), .B1(n_321), .B2(n_322), .C(n_325), .Y(n_314) );
INVx1_ASAP7_75t_L g357 ( .A(n_305), .Y(n_357) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_SL g329 ( .A(n_310), .Y(n_329) );
OR2x2_ASAP7_75t_L g402 ( .A(n_310), .B(n_334), .Y(n_402) );
AND2x2_ASAP7_75t_L g404 ( .A(n_310), .B(n_312), .Y(n_404) );
INVx1_ASAP7_75t_L g343 ( .A(n_313), .Y(n_343) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_319), .Y(n_315) );
AOI21xp33_ASAP7_75t_SL g373 ( .A1(n_316), .A2(n_374), .B(n_375), .Y(n_373) );
OR2x2_ASAP7_75t_L g380 ( .A(n_316), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g354 ( .A(n_317), .B(n_338), .Y(n_354) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp33_ASAP7_75t_SL g371 ( .A(n_322), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_323), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_324), .B(n_360), .Y(n_423) );
O2A1O1Ixp33_ASAP7_75t_L g339 ( .A1(n_327), .A2(n_340), .B(n_342), .C(n_343), .Y(n_339) );
NAND2x1_ASAP7_75t_SL g364 ( .A(n_327), .B(n_365), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_328), .A2(n_377), .B1(n_379), .B2(n_382), .Y(n_376) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_330), .B(n_420), .Y(n_419) );
NAND5xp2_ASAP7_75t_L g331 ( .A(n_332), .B(n_344), .C(n_362), .D(n_376), .E(n_385), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_333), .B(n_339), .Y(n_332) );
INVx1_ASAP7_75t_L g389 ( .A(n_335), .Y(n_389) );
INVx1_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g395 ( .A1(n_337), .A2(n_356), .B1(n_396), .B2(n_398), .C(n_401), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_338), .B(n_432), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_341), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_341), .B(n_407), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_349), .B1(n_351), .B2(n_353), .Y(n_347) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_359), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
AND2x2_ASAP7_75t_L g429 ( .A(n_358), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_366), .B1(n_370), .B2(n_371), .C(n_373), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g413 ( .A(n_368), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_SL g420 ( .A(n_378), .Y(n_420) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OAI21xp5_ASAP7_75t_SL g385 ( .A1(n_386), .A2(n_388), .B(n_389), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI211xp5_ASAP7_75t_SL g390 ( .A1(n_391), .A2(n_393), .B(n_395), .C(n_408), .Y(n_390) );
INVx1_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
A2O1A1Ixp33_ASAP7_75t_L g417 ( .A1(n_393), .A2(n_418), .B(n_419), .C(n_421), .Y(n_417) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_397), .B(n_399), .Y(n_398) );
AOI21xp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B(n_405), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AOI21xp33_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_431), .B(n_433), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g717 ( .A(n_439), .Y(n_717) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OR5x1_ASAP7_75t_L g441 ( .A(n_442), .B(n_605), .C(n_663), .D(n_699), .E(n_706), .Y(n_441) );
NAND3xp33_ASAP7_75t_SL g442 ( .A(n_443), .B(n_551), .C(n_575), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_487), .B1(n_517), .B2(n_522), .C(n_532), .Y(n_443) );
OAI21xp5_ASAP7_75t_SL g685 ( .A1(n_444), .A2(n_686), .B(n_688), .Y(n_685) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_470), .Y(n_444) );
NAND2x1p5_ASAP7_75t_L g675 ( .A(n_445), .B(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_459), .Y(n_445) );
INVx2_ASAP7_75t_L g521 ( .A(n_446), .Y(n_521) );
AND2x2_ASAP7_75t_L g534 ( .A(n_446), .B(n_472), .Y(n_534) );
AND2x2_ASAP7_75t_L g588 ( .A(n_446), .B(n_471), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_446), .B(n_460), .Y(n_603) );
O2A1O1Ixp33_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_455), .B(n_456), .C(n_457), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_457), .A2(n_478), .B(n_479), .Y(n_477) );
AND2x2_ASAP7_75t_L g621 ( .A(n_459), .B(n_562), .Y(n_621) );
AND2x2_ASAP7_75t_L g654 ( .A(n_459), .B(n_472), .Y(n_654) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OR2x2_ASAP7_75t_L g561 ( .A(n_460), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g574 ( .A(n_460), .B(n_472), .Y(n_574) );
AND2x2_ASAP7_75t_L g581 ( .A(n_460), .B(n_562), .Y(n_581) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_460), .Y(n_590) );
AND2x2_ASAP7_75t_L g597 ( .A(n_460), .B(n_471), .Y(n_597) );
INVx1_ASAP7_75t_L g628 ( .A(n_460), .Y(n_628) );
OAI21xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_465), .B(n_468), .Y(n_461) );
INVx1_ASAP7_75t_L g604 ( .A(n_470), .Y(n_604) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_481), .Y(n_470) );
INVx2_ASAP7_75t_L g560 ( .A(n_471), .Y(n_560) );
AND2x2_ASAP7_75t_L g582 ( .A(n_471), .B(n_521), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_471), .B(n_628), .Y(n_633) );
INVx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_472), .B(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g705 ( .A(n_472), .B(n_669), .Y(n_705) );
INVx2_ASAP7_75t_L g519 ( .A(n_481), .Y(n_519) );
INVx3_ASAP7_75t_L g620 ( .A(n_481), .Y(n_620) );
OR2x2_ASAP7_75t_L g650 ( .A(n_481), .B(n_651), .Y(n_650) );
NOR2x1_ASAP7_75t_L g676 ( .A(n_481), .B(n_560), .Y(n_676) );
AND2x4_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
INVx1_ASAP7_75t_L g563 ( .A(n_482), .Y(n_563) );
AOI33xp33_ASAP7_75t_L g696 ( .A1(n_487), .A2(n_534), .A3(n_548), .B1(n_620), .B2(n_697), .B3(n_698), .Y(n_696) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_496), .Y(n_488) );
OR2x2_ASAP7_75t_L g549 ( .A(n_489), .B(n_550), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_489), .B(n_546), .Y(n_608) );
OR2x2_ASAP7_75t_L g661 ( .A(n_489), .B(n_662), .Y(n_661) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g587 ( .A(n_490), .B(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g612 ( .A(n_490), .B(n_496), .Y(n_612) );
AND2x2_ASAP7_75t_L g679 ( .A(n_490), .B(n_524), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g704 ( .A1(n_490), .A2(n_579), .B(n_705), .Y(n_704) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g526 ( .A(n_491), .Y(n_526) );
INVx1_ASAP7_75t_L g539 ( .A(n_491), .Y(n_539) );
AND2x2_ASAP7_75t_L g558 ( .A(n_491), .B(n_528), .Y(n_558) );
AND2x2_ASAP7_75t_L g607 ( .A(n_491), .B(n_527), .Y(n_607) );
INVx2_ASAP7_75t_SL g649 ( .A(n_496), .Y(n_649) );
OR2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_507), .Y(n_496) );
INVx2_ASAP7_75t_L g569 ( .A(n_497), .Y(n_569) );
INVx1_ASAP7_75t_L g700 ( .A(n_497), .Y(n_700) );
AND2x2_ASAP7_75t_L g713 ( .A(n_497), .B(n_594), .Y(n_713) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g540 ( .A(n_498), .Y(n_540) );
OR2x2_ASAP7_75t_L g546 ( .A(n_498), .B(n_547), .Y(n_546) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_498), .Y(n_557) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_507), .Y(n_524) );
AND2x2_ASAP7_75t_L g541 ( .A(n_507), .B(n_527), .Y(n_541) );
INVx1_ASAP7_75t_L g547 ( .A(n_507), .Y(n_547) );
INVx1_ASAP7_75t_L g554 ( .A(n_507), .Y(n_554) );
AND2x2_ASAP7_75t_L g579 ( .A(n_507), .B(n_528), .Y(n_579) );
INVx2_ASAP7_75t_L g595 ( .A(n_507), .Y(n_595) );
AND2x2_ASAP7_75t_L g688 ( .A(n_507), .B(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_507), .B(n_569), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_511), .B(n_512), .Y(n_509) );
INVx1_ASAP7_75t_SL g517 ( .A(n_518), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
INVx2_ASAP7_75t_L g543 ( .A(n_519), .Y(n_543) );
INVx1_ASAP7_75t_L g572 ( .A(n_519), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_519), .B(n_603), .Y(n_669) );
INVx1_ASAP7_75t_SL g629 ( .A(n_520), .Y(n_629) );
INVx2_ASAP7_75t_L g550 ( .A(n_521), .Y(n_550) );
AND2x2_ASAP7_75t_L g619 ( .A(n_521), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g635 ( .A(n_521), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_525), .Y(n_522) );
INVx1_ASAP7_75t_L g697 ( .A(n_523), .Y(n_697) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g552 ( .A(n_525), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g655 ( .A(n_525), .B(n_645), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_525), .A2(n_666), .B(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
AND2x2_ASAP7_75t_L g568 ( .A(n_526), .B(n_569), .Y(n_568) );
BUFx2_ASAP7_75t_L g593 ( .A(n_526), .Y(n_593) );
INVx1_ASAP7_75t_L g617 ( .A(n_526), .Y(n_617) );
OR2x2_ASAP7_75t_L g681 ( .A(n_527), .B(n_540), .Y(n_681) );
NOR2xp67_ASAP7_75t_L g689 ( .A(n_527), .B(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g594 ( .A(n_528), .B(n_595), .Y(n_594) );
BUFx2_ASAP7_75t_L g601 ( .A(n_528), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_535), .B1(n_542), .B2(n_544), .Y(n_532) );
OR2x2_ASAP7_75t_L g611 ( .A(n_533), .B(n_561), .Y(n_611) );
INVx1_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
AOI222xp33_ASAP7_75t_L g652 ( .A1(n_534), .A2(n_653), .B1(n_655), .B2(n_656), .C1(n_657), .C2(n_660), .Y(n_652) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_541), .Y(n_536) );
INVx1_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g599 ( .A(n_538), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
AND2x2_ASAP7_75t_SL g553 ( .A(n_540), .B(n_554), .Y(n_553) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_540), .Y(n_624) );
AND2x2_ASAP7_75t_L g672 ( .A(n_540), .B(n_541), .Y(n_672) );
INVx1_ASAP7_75t_L g690 ( .A(n_540), .Y(n_690) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g656 ( .A(n_543), .B(n_582), .Y(n_656) );
AND2x2_ASAP7_75t_L g698 ( .A(n_543), .B(n_574), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_548), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_545), .B(n_593), .Y(n_680) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_546), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g573 ( .A(n_550), .B(n_574), .Y(n_573) );
INVx3_ASAP7_75t_L g641 ( .A(n_550), .Y(n_641) );
O2A1O1Ixp33_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_555), .B(n_559), .C(n_564), .Y(n_551) );
INVxp67_ASAP7_75t_L g565 ( .A(n_552), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_553), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_553), .B(n_600), .Y(n_695) );
BUFx3_ASAP7_75t_L g659 ( .A(n_554), .Y(n_659) );
INVx1_ASAP7_75t_L g566 ( .A(n_555), .Y(n_566) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g585 ( .A(n_557), .B(n_579), .Y(n_585) );
INVx1_ASAP7_75t_SL g625 ( .A(n_558), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
INVx1_ASAP7_75t_L g615 ( .A(n_560), .Y(n_615) );
AND2x2_ASAP7_75t_L g638 ( .A(n_560), .B(n_621), .Y(n_638) );
INVx1_ASAP7_75t_SL g609 ( .A(n_561), .Y(n_609) );
INVx1_ASAP7_75t_L g636 ( .A(n_562), .Y(n_636) );
AOI31xp33_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_566), .A3(n_567), .B(n_570), .Y(n_564) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g657 ( .A(n_568), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g631 ( .A(n_569), .Y(n_631) );
BUFx2_ASAP7_75t_L g645 ( .A(n_569), .Y(n_645) );
AND2x2_ASAP7_75t_L g673 ( .A(n_569), .B(n_594), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_SL g646 ( .A(n_573), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_574), .B(n_641), .Y(n_687) );
AND2x2_ASAP7_75t_L g694 ( .A(n_574), .B(n_620), .Y(n_694) );
AOI211xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_580), .B(n_583), .C(n_598), .Y(n_575) );
INVxp67_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AOI221xp5_ASAP7_75t_L g606 ( .A1(n_580), .A2(n_607), .B1(n_608), .B2(n_609), .C(n_610), .Y(n_606) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
AND2x2_ASAP7_75t_L g614 ( .A(n_581), .B(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g651 ( .A(n_582), .Y(n_651) );
OAI32xp33_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_586), .A3(n_589), .B1(n_591), .B2(n_596), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
O2A1O1Ixp33_ASAP7_75t_L g637 ( .A1(n_585), .A2(n_638), .B(n_639), .C(n_642), .Y(n_637) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
OAI21xp5_ASAP7_75t_SL g701 ( .A1(n_593), .A2(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_L g662 ( .A(n_594), .Y(n_662) );
INVxp67_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_599), .B(n_602), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_600), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g648 ( .A(n_600), .B(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g665 ( .A(n_602), .Y(n_665) );
OR2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
NAND4xp25_ASAP7_75t_SL g605 ( .A(n_606), .B(n_618), .C(n_637), .D(n_652), .Y(n_605) );
AND2x2_ASAP7_75t_L g644 ( .A(n_607), .B(n_645), .Y(n_644) );
AND2x4_ASAP7_75t_L g666 ( .A(n_607), .B(n_659), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_609), .B(n_641), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_612), .B1(n_613), .B2(n_616), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_611), .A2(n_662), .B1(n_693), .B2(n_695), .Y(n_692) );
O2A1O1Ixp33_ASAP7_75t_L g699 ( .A1(n_611), .A2(n_700), .B(n_701), .C(n_704), .Y(n_699) );
INVx2_ASAP7_75t_L g670 ( .A(n_612), .Y(n_670) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AOI222xp33_ASAP7_75t_L g664 ( .A1(n_614), .A2(n_648), .B1(n_665), .B2(n_666), .C1(n_667), .C2(n_670), .Y(n_664) );
O2A1O1Ixp33_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_621), .B(n_622), .C(n_626), .Y(n_618) );
INVx1_ASAP7_75t_L g684 ( .A(n_619), .Y(n_684) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OAI22xp33_ASAP7_75t_L g626 ( .A1(n_623), .A2(n_627), .B1(n_630), .B2(n_632), .Y(n_626) );
OR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
OR2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g653 ( .A(n_635), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g711 ( .A(n_638), .Y(n_711) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI22xp33_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_646), .B1(n_647), .B2(n_650), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_645), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g702 ( .A(n_650), .Y(n_702) );
INVx1_ASAP7_75t_L g683 ( .A(n_654), .Y(n_683) );
CKINVDCx16_ASAP7_75t_R g710 ( .A(n_656), .Y(n_710) );
INVxp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND5xp2_ASAP7_75t_L g663 ( .A(n_664), .B(n_671), .C(n_685), .D(n_691), .E(n_696), .Y(n_663) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
O2A1O1Ixp33_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .B(n_674), .C(n_677), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AOI31xp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_680), .A3(n_681), .B(n_682), .Y(n_677) );
INVx1_ASAP7_75t_L g703 ( .A(n_679), .Y(n_703) );
OR2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OAI222xp33_ASAP7_75t_L g706 ( .A1(n_693), .A2(n_695), .B1(n_707), .B2(n_710), .C1(n_711), .C2(n_712), .Y(n_706) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
BUFx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
endmodule