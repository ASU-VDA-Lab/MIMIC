module real_jpeg_13320_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_308, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_308;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_215;
wire n_221;
wire n_176;
wire n_249;
wire n_292;
wire n_288;
wire n_300;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_184;
wire n_164;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_305;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_285;
wire n_45;
wire n_172;
wire n_304;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_225;
wire n_103;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_295;
wire n_213;
wire n_202;
wire n_167;
wire n_179;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g110 ( 
.A(n_0),
.Y(n_110)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_30),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_3),
.A2(n_30),
.B1(n_48),
.B2(n_49),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_3),
.A2(n_30),
.B1(n_42),
.B2(n_46),
.Y(n_235)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_6),
.A2(n_42),
.B1(n_46),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_6),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_54),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_54),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_6),
.A2(n_48),
.B1(n_49),
.B2(n_54),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_6),
.B(n_60),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_6),
.B(n_45),
.C(n_49),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_6),
.B(n_109),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_6),
.B(n_47),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_6),
.A2(n_24),
.B(n_62),
.C(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_6),
.B(n_20),
.Y(n_188)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_9),
.A2(n_48),
.B1(n_49),
.B2(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_9),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_9),
.A2(n_42),
.B1(n_46),
.B2(n_115),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_115),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_115),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_35),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_10),
.A2(n_35),
.B1(n_42),
.B2(n_46),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_10),
.A2(n_35),
.B1(n_48),
.B2(n_49),
.Y(n_146)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_94),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_92),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_84),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_15),
.B(n_84),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_70),
.C(n_76),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_16),
.A2(n_17),
.B1(n_70),
.B2(n_78),
.Y(n_302)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_36),
.B1(n_37),
.B2(n_69),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_18),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_25),
.B(n_31),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_19),
.A2(n_74),
.B(n_75),
.Y(n_279)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_20),
.B(n_34),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_20),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_20),
.B(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_21),
.A2(n_22),
.B1(n_26),
.B2(n_27),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_21),
.B(n_24),
.C(n_54),
.Y(n_200)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_23),
.A2(n_24),
.B1(n_62),
.B2(n_63),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_25),
.A2(n_71),
.B(n_74),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_26),
.B(n_200),
.Y(n_199)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_31),
.B(n_208),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_32),
.B(n_209),
.Y(n_219)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_55),
.B1(n_56),
.B2(n_68),
.Y(n_37)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_38),
.B(n_78),
.C(n_79),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_38),
.B(n_56),
.C(n_69),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_38),
.A2(n_68),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_38),
.A2(n_68),
.B1(n_79),
.B2(n_296),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_52),
.B(n_53),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_39),
.A2(n_119),
.B(n_235),
.Y(n_265)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_40),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_40),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_40),
.B(n_120),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_47),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_41)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_46),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_42),
.B(n_130),
.Y(n_129)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AO22x1_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_45),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_46),
.A2(n_54),
.B(n_63),
.Y(n_171)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_47),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_47),
.B(n_122),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_47),
.B(n_134),
.Y(n_178)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_49),
.B(n_110),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_49),
.B(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_52),
.A2(n_166),
.B(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_53),
.Y(n_134)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_64),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_58),
.B(n_221),
.Y(n_220)
);

NAND2x1_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_59),
.A2(n_60),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_59),
.B(n_87),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_60),
.B(n_163),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_60),
.A2(n_64),
.B(n_81),
.Y(n_283)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_61),
.B(n_67),
.Y(n_83)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_64),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_65),
.A2(n_80),
.B(n_82),
.Y(n_79)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_65),
.B(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_68),
.B(n_206),
.C(n_212),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_70),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_70),
.A2(n_78),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_71),
.B(n_219),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_73),
.B(n_207),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_75),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_76),
.A2(n_77),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_79),
.Y(n_296)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_83),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_83),
.B(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_91),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_86),
.A2(n_90),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_86),
.B(n_225),
.C(n_231),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_286),
.B(n_303),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_269),
.B(n_285),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_248),
.B(n_268),
.Y(n_97)
);

AOI321xp33_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_215),
.A3(n_241),
.B1(n_246),
.B2(n_247),
.C(n_308),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_191),
.B(n_214),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_174),
.B(n_190),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_157),
.B(n_173),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_135),
.B(n_156),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_127),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_104),
.B(n_127),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_116),
.B1(n_117),
.B2(n_126),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_105),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_111),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_106),
.B(n_153),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_113),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_108),
.A2(n_110),
.B(n_113),
.Y(n_169)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_114),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_110),
.A2(n_153),
.B(n_202),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_146),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_113),
.A2(n_202),
.B(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_117)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_119),
.B(n_133),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_121),
.B(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_124),
.C(n_126),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_131),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_128),
.A2(n_129),
.B1(n_131),
.B2(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_149),
.B(n_155),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_143),
.B(n_148),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_142),
.B(n_145),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_147),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_145),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_152),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_159),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_167),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_165),
.C(n_167),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_162),
.Y(n_213)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

INVxp33_ASAP7_75t_L g262 ( 
.A(n_164),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_166),
.B(n_178),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_170),
.B2(n_172),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_168),
.A2(n_169),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_168),
.A2(n_169),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_170),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_169),
.B(n_265),
.Y(n_276)
);

AOI21xp33_ASAP7_75t_L g290 ( 
.A1(n_169),
.A2(n_276),
.B(n_278),
.Y(n_290)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_170),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_189),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_189),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_182),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_176)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_177),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_179),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_180),
.C(n_182),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_187),
.C(n_188),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_184),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_193),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_204),
.B2(n_205),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_196),
.B(n_197),
.C(n_204),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_201),
.B2(n_203),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_203),
.Y(n_222)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_210),
.Y(n_205)
);

INVxp33_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_236),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_236),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_223),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_224),
.C(n_232),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.C(n_222),
.Y(n_217)
);

FAx1_ASAP7_75t_SL g238 ( 
.A(n_218),
.B(n_220),
.CI(n_222),
.CON(n_238),
.SN(n_238)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_219),
.B(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_232),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_229),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_228),
.Y(n_239)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_230),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_234),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_239),
.C(n_240),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_237),
.A2(n_238),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx24_ASAP7_75t_SL g306 ( 
.A(n_238),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_240),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_245),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_245),
.Y(n_246)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_250),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_267),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_263),
.B2(n_264),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_264),
.C(n_267),
.Y(n_270)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_256),
.C(n_261),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_260),
.B2(n_261),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_265),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_271),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_274),
.C(n_281),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_280),
.B2(n_281),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_283),
.B(n_284),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_282),
.B(n_283),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_284),
.A2(n_292),
.B1(n_293),
.B2(n_297),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_284),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_290),
.C(n_292),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_298),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_289),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_298),
.A2(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_300),
.Y(n_305)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);


endmodule