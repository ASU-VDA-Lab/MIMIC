module fake_jpeg_5450_n_337 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_46),
.Y(n_63)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_25),
.B1(n_24),
.B2(n_35),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_19),
.B1(n_34),
.B2(n_31),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_50),
.A2(n_71),
.B1(n_32),
.B2(n_20),
.Y(n_95)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_28),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_54),
.B(n_64),
.Y(n_92)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_57),
.Y(n_74)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_25),
.B1(n_24),
.B2(n_19),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_59),
.A2(n_22),
.B1(n_1),
.B2(n_2),
.Y(n_87)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_61),
.Y(n_73)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_62),
.B(n_0),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_65),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_68),
.Y(n_79)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_70),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_45),
.A2(n_23),
.B1(n_34),
.B2(n_31),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_48),
.A2(n_47),
.B1(n_45),
.B2(n_35),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_57),
.A2(n_47),
.B1(n_29),
.B2(n_27),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_80),
.A2(n_81),
.B1(n_98),
.B2(n_62),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_48),
.A2(n_27),
.B1(n_22),
.B2(n_29),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_60),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_82),
.Y(n_113)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_86),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_43),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_68),
.C(n_49),
.Y(n_107)
);

AO22x2_ASAP7_75t_L g85 ( 
.A1(n_72),
.A2(n_43),
.B1(n_40),
.B2(n_32),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_85),
.A2(n_58),
.B1(n_66),
.B2(n_67),
.Y(n_117)
);

INVxp33_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_99),
.B1(n_54),
.B2(n_51),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_52),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_89),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_63),
.Y(n_89)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_30),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_91),
.B(n_54),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_95),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_55),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_100),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_61),
.A2(n_43),
.B1(n_40),
.B2(n_32),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_49),
.A2(n_70),
.B1(n_69),
.B2(n_64),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_108),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_125),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_102),
.Y(n_108)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_111),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_92),
.B1(n_82),
.B2(n_86),
.Y(n_140)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_115),
.Y(n_157)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g137 ( 
.A(n_116),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_96),
.B1(n_88),
.B2(n_78),
.Y(n_146)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_118),
.B(n_119),
.Y(n_150)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

NOR2x1_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_67),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_94),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_79),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_121),
.B(n_77),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_66),
.B1(n_67),
.B2(n_32),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_122),
.A2(n_101),
.B1(n_73),
.B2(n_79),
.Y(n_135)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

INVxp33_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

INVx3_ASAP7_75t_SL g126 ( 
.A(n_75),
.Y(n_126)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_131),
.Y(n_158)
);

BUFx24_ASAP7_75t_SL g130 ( 
.A(n_74),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_130),
.Y(n_134)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_135),
.A2(n_140),
.B1(n_148),
.B2(n_116),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

INVx6_ASAP7_75t_SL g194 ( 
.A(n_136),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_74),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_138),
.A2(n_149),
.B(n_161),
.Y(n_193)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_142),
.Y(n_173)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_144),
.Y(n_185)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_146),
.A2(n_154),
.B1(n_104),
.B2(n_18),
.Y(n_179)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_147),
.B(n_151),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_106),
.A2(n_94),
.B1(n_97),
.B2(n_77),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_125),
.A2(n_100),
.B(n_97),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_114),
.A2(n_96),
.B1(n_93),
.B2(n_66),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_152),
.A2(n_155),
.B1(n_159),
.B2(n_131),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_20),
.B1(n_18),
.B2(n_17),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_119),
.A2(n_20),
.B1(n_18),
.B2(n_17),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_160),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_103),
.A2(n_30),
.B(n_20),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_163),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_142),
.B(n_113),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_164),
.B(n_167),
.Y(n_217)
);

NOR2x1p5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_120),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_165),
.A2(n_191),
.B(n_0),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_103),
.B(n_128),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_166),
.A2(n_176),
.B(n_178),
.Y(n_224)
);

BUFx24_ASAP7_75t_SL g167 ( 
.A(n_134),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_151),
.A2(n_144),
.B1(n_157),
.B2(n_110),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_168),
.Y(n_201)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_135),
.A2(n_115),
.B1(n_122),
.B2(n_105),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_170),
.A2(n_136),
.B1(n_17),
.B2(n_30),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_105),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_182),
.Y(n_205)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_172),
.Y(n_209)
);

BUFx12_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_174),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_137),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_175),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_153),
.A2(n_158),
.B(n_149),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_132),
.Y(n_177)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_158),
.A2(n_30),
.B(n_18),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_SL g197 ( 
.A1(n_179),
.A2(n_189),
.B(n_190),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_145),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_180),
.Y(n_225)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

O2A1O1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_155),
.A2(n_17),
.B(n_30),
.C(n_127),
.Y(n_183)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_183),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_152),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_186),
.Y(n_210)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_187),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_138),
.B(n_30),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_0),
.Y(n_206)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_141),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_133),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_192),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_139),
.C(n_143),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_199),
.C(n_202),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_139),
.C(n_133),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_147),
.C(n_160),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_204),
.A2(n_218),
.B1(n_183),
.B2(n_163),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_168),
.Y(n_234)
);

OAI22x1_ASAP7_75t_L g207 ( 
.A1(n_165),
.A2(n_194),
.B1(n_166),
.B2(n_189),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_207),
.A2(n_182),
.B1(n_186),
.B2(n_169),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_134),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_215),
.C(n_174),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_181),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_162),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_165),
.A2(n_162),
.B(n_3),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_220),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_170),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_196),
.A2(n_3),
.B(n_4),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_223),
.B(n_174),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_221),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_226),
.B(n_232),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_228),
.A2(n_235),
.B(n_237),
.Y(n_265)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_229),
.B(n_234),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_230),
.A2(n_220),
.B1(n_203),
.B2(n_206),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_231),
.A2(n_239),
.B(n_241),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_213),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_178),
.Y(n_233)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_233),
.Y(n_259)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

NOR3xp33_ASAP7_75t_SL g236 ( 
.A(n_207),
.B(n_185),
.C(n_187),
.Y(n_236)
);

A2O1A1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_236),
.A2(n_224),
.B(n_216),
.C(n_211),
.Y(n_252)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_225),
.Y(n_238)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_191),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

INVx11_ASAP7_75t_L g269 ( 
.A(n_240),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_190),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_209),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_201),
.A2(n_195),
.B1(n_173),
.B2(n_192),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_243),
.A2(n_200),
.B1(n_204),
.B2(n_202),
.Y(n_255)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_244),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_251),
.C(n_208),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_246),
.A2(n_247),
.B1(n_249),
.B2(n_223),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_172),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_4),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_199),
.B(n_16),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_8),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_198),
.B(n_5),
.C(n_6),
.Y(n_251)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_254),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_256),
.B(n_271),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_240),
.A2(n_219),
.B1(n_197),
.B2(n_224),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_257),
.A2(n_260),
.B1(n_228),
.B2(n_243),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_234),
.B(n_245),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_263),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_209),
.C(n_203),
.Y(n_263)
);

MAJx2_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_6),
.C(n_7),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_268),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_8),
.C(n_9),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_9),
.Y(n_272)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_264),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_281),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_270),
.A2(n_230),
.B1(n_241),
.B2(n_233),
.Y(n_279)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_279),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_269),
.A2(n_239),
.B1(n_231),
.B2(n_236),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_280),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_253),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_264),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_284),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_257),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_265),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_261),
.B(n_248),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_263),
.C(n_256),
.Y(n_295)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_255),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_289),
.Y(n_293)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_282),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_292),
.A2(n_295),
.B(n_301),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_273),
.B(n_266),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_296),
.B(n_297),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_286),
.B(n_248),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_258),
.C(n_268),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_299),
.A2(n_302),
.B(n_303),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_292),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_262),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_275),
.B(n_272),
.C(n_271),
.Y(n_302)
);

XNOR2x1_ASAP7_75t_L g303 ( 
.A(n_276),
.B(n_267),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_304),
.A2(n_305),
.B(n_306),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_269),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_274),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_290),
.B(n_288),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_309),
.B(n_311),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_280),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_310),
.B(n_312),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_291),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_303),
.B(n_276),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_300),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_313),
.B(n_287),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_299),
.A2(n_283),
.B1(n_252),
.B2(n_287),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_315),
.A2(n_11),
.B(n_13),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_316),
.A2(n_317),
.B(n_323),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_251),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_302),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_320),
.B(n_14),
.Y(n_327)
);

OAI21x1_ASAP7_75t_L g321 ( 
.A1(n_307),
.A2(n_277),
.B(n_12),
.Y(n_321)
);

AOI21x1_ASAP7_75t_SL g326 ( 
.A1(n_321),
.A2(n_11),
.B(n_13),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_311),
.A2(n_11),
.B(n_13),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_14),
.C(n_15),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_315),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_326),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_328),
.C(n_329),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_15),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_330),
.A2(n_318),
.B(n_319),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_332),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_333),
.Y(n_337)
);


endmodule