module fake_jpeg_22711_n_191 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_191);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_191;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_5),
.B(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_0),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_39),
.B(n_29),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_0),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_15),
.B(n_1),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_44),
.B(n_14),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_26),
.C(n_19),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_31),
.Y(n_89)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_32),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_54),
.B(n_4),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_22),
.Y(n_55)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_22),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_57),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_28),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_28),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_36),
.A2(n_43),
.B1(n_42),
.B2(n_34),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_64),
.B1(n_67),
.B2(n_69),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_20),
.B1(n_21),
.B2(n_17),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_29),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_23),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_34),
.A2(n_20),
.B1(n_21),
.B2(n_26),
.Y(n_67)
);

AO22x1_ASAP7_75t_SL g69 ( 
.A1(n_43),
.A2(n_26),
.B1(n_19),
.B2(n_23),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_37),
.A2(n_21),
.B1(n_30),
.B2(n_25),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_73),
.B1(n_67),
.B2(n_69),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_33),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_31),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_37),
.A2(n_30),
.B1(n_25),
.B2(n_15),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_35),
.B(n_1),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_1),
.B(n_3),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_69),
.A2(n_40),
.B1(n_41),
.B2(n_16),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_82),
.Y(n_114)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_100),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_23),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_45),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_85),
.Y(n_118)
);

OR2x4_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_97),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_45),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_45),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_63),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_33),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_46),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_64),
.C(n_62),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_51),
.A2(n_41),
.B1(n_40),
.B2(n_5),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_31),
.B1(n_4),
.B2(n_6),
.Y(n_91)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_31),
.Y(n_93)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_3),
.Y(n_95)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_6),
.Y(n_98)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_89),
.C(n_88),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_10),
.C(n_11),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_115),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_99),
.Y(n_107)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_49),
.Y(n_111)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_91),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_112),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_49),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_113),
.B(n_97),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_80),
.A2(n_60),
.B1(n_51),
.B2(n_46),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_87),
.Y(n_123)
);

AO22x1_ASAP7_75t_SL g117 ( 
.A1(n_80),
.A2(n_72),
.B1(n_52),
.B2(n_63),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_117),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_72),
.B(n_52),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_119),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_86),
.A2(n_10),
.B1(n_13),
.B2(n_7),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_121),
.Y(n_130)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_7),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_136),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_139),
.C(n_104),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_78),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_128),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_82),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_132),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_106),
.B(n_94),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_133),
.C(n_101),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_75),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_96),
.Y(n_137)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_75),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_113),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_140),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_141),
.A2(n_119),
.B(n_122),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_154),
.C(n_146),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_148),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_134),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_117),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_141),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_117),
.B1(n_109),
.B2(n_115),
.Y(n_151)
);

O2A1O1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_151),
.A2(n_125),
.B(n_141),
.C(n_128),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_127),
.A2(n_103),
.B(n_101),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_SL g166 ( 
.A1(n_152),
.A2(n_153),
.B(n_110),
.C(n_106),
.Y(n_166)
);

HAxp5_ASAP7_75t_SL g153 ( 
.A(n_127),
.B(n_103),
.CON(n_153),
.SN(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_123),
.C(n_126),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_120),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_145),
.B(n_137),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_163),
.Y(n_167)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_165),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_159),
.C(n_164),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_108),
.C(n_129),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_160),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_162),
.A2(n_153),
.B1(n_152),
.B2(n_149),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_136),
.C(n_139),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_166),
.A2(n_160),
.B1(n_144),
.B2(n_161),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_168),
.A2(n_173),
.B1(n_167),
.B2(n_171),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_145),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_173),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_172),
.A2(n_174),
.B(n_79),
.Y(n_176)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_166),
.A2(n_79),
.B(n_100),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_175),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_167),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_178),
.B(n_121),
.Y(n_183)
);

AOI21xp33_ASAP7_75t_L g179 ( 
.A1(n_169),
.A2(n_146),
.B(n_150),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_180),
.B(n_172),
.Y(n_182)
);

OAI21x1_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_150),
.B(n_96),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_181),
.B(n_175),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_182),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_183),
.A2(n_185),
.B1(n_13),
.B2(n_7),
.Y(n_188)
);

AOI21x1_ASAP7_75t_L g186 ( 
.A1(n_184),
.A2(n_181),
.B(n_177),
.Y(n_186)
);

OAI21x1_ASAP7_75t_L g189 ( 
.A1(n_186),
.A2(n_187),
.B(n_184),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_188),
.B(n_9),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_190),
.Y(n_191)
);


endmodule