module fake_ariane_2537_n_1996 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1996);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1996;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_851;
wire n_212;
wire n_444;
wire n_355;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_604;
wire n_439;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_1126;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_97),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_65),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_126),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_174),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_123),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_127),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_103),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_85),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_48),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_106),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_44),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_7),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_13),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_170),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_186),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_163),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g226 ( 
.A(n_91),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_55),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_15),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_112),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_70),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_86),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_168),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_69),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_77),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g235 ( 
.A(n_102),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_120),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_195),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_153),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_142),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_10),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_88),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_99),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_63),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_156),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_162),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_41),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_208),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_7),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_176),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_25),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_24),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_134),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_200),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_132),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_137),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_104),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_42),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_30),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_50),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_36),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_164),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_17),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_136),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_28),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_76),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_69),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_89),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_40),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_1),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_179),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_205),
.Y(n_271)
);

BUFx5_ASAP7_75t_L g272 ( 
.A(n_52),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_32),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_82),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_95),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_116),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_6),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_207),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_161),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_139),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_125),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_56),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_167),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_47),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_147),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_148),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_70),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_26),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_118),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_56),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_55),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_37),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_140),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_35),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_40),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_93),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_143),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_202),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_0),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_100),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_191),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_37),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_204),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_62),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_181),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_8),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_71),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_17),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_10),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_92),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_146),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_185),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_44),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_113),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_20),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_180),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_203),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_16),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_0),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_47),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_67),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_52),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_157),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_34),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_63),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_184),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_133),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_22),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_49),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_21),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_135),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_38),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_60),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_178),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_187),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_39),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_192),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_151),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_183),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_188),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_114),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_34),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_62),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_26),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_14),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_43),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_11),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_145),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_58),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_165),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_61),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_175),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_42),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_21),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_149),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_194),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_129),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_25),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_80),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_159),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_206),
.Y(n_361)
);

CKINVDCx14_ASAP7_75t_R g362 ( 
.A(n_152),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_201),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_66),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_198),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_177),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_65),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_150),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_31),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_11),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_39),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_28),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_20),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_51),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_68),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_79),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_101),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_197),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_23),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_173),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_67),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_96),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_75),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_109),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_14),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_12),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_169),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_59),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_60),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_111),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_36),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_193),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_141),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_130),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_105),
.Y(n_395)
);

BUFx10_ASAP7_75t_L g396 ( 
.A(n_122),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_166),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_57),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_84),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_117),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_23),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_121),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_19),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_16),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_1),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_8),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_45),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_155),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_46),
.Y(n_409)
);

BUFx10_ASAP7_75t_L g410 ( 
.A(n_172),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_196),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_74),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_4),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_6),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_107),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_333),
.Y(n_416)
);

INVxp33_ASAP7_75t_SL g417 ( 
.A(n_354),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_342),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_272),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_272),
.B(n_359),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_287),
.Y(n_421)
);

INVxp33_ASAP7_75t_SL g422 ( 
.A(n_210),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_288),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_272),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_329),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_272),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_237),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_272),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_247),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_272),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_271),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_272),
.Y(n_432)
);

INVxp33_ASAP7_75t_SL g433 ( 
.A(n_210),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_272),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_213),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_278),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_224),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_228),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_297),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_228),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_409),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_326),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_360),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_409),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_368),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_222),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_L g447 ( 
.A(n_217),
.B(n_2),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_222),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_376),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_397),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_415),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_259),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_230),
.B(n_2),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_223),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_262),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_223),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_258),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_345),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_264),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_245),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_269),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_398),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_245),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_273),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_277),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_282),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_284),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_249),
.Y(n_468)
);

INVxp67_ASAP7_75t_SL g469 ( 
.A(n_264),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_211),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_244),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_291),
.Y(n_472)
);

INVxp33_ASAP7_75t_SL g473 ( 
.A(n_217),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_230),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_256),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_383),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_249),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_292),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_294),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_289),
.Y(n_480)
);

NOR2xp67_ASAP7_75t_L g481 ( 
.A(n_220),
.B(n_3),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_289),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_302),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_293),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_293),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_261),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g487 ( 
.A(n_266),
.Y(n_487)
);

INVxp33_ASAP7_75t_L g488 ( 
.A(n_219),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_304),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_306),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_300),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_338),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_230),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_300),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_392),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_339),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_308),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_315),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_392),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_318),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_400),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_320),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_362),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_325),
.Y(n_504)
);

INVxp67_ASAP7_75t_SL g505 ( 
.A(n_266),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_328),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_400),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_220),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_226),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_257),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_229),
.B(n_3),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_336),
.Y(n_512)
);

INVxp67_ASAP7_75t_SL g513 ( 
.A(n_299),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_260),
.Y(n_514)
);

NOR2xp67_ASAP7_75t_L g515 ( 
.A(n_221),
.B(n_4),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_343),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_236),
.Y(n_517)
);

INVxp67_ASAP7_75t_SL g518 ( 
.A(n_299),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_268),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_241),
.B(n_5),
.Y(n_520)
);

NAND2x1_ASAP7_75t_L g521 ( 
.A(n_453),
.B(n_234),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_419),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_419),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_487),
.B(n_226),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_424),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_487),
.B(n_226),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_420),
.B(n_234),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_459),
.B(n_253),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_469),
.B(n_505),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_435),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_435),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_424),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_513),
.B(n_254),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_426),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_417),
.A2(n_386),
.B1(n_351),
.B2(n_251),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_508),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_518),
.B(n_276),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_435),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_488),
.B(n_235),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_426),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_422),
.B(n_279),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_428),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_470),
.B(n_517),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_435),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_428),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_421),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_430),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_430),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_435),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_432),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_432),
.Y(n_551)
);

AND3x2_ASAP7_75t_L g552 ( 
.A(n_453),
.B(n_322),
.C(n_307),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_470),
.B(n_323),
.Y(n_553)
);

AND2x6_ASAP7_75t_L g554 ( 
.A(n_434),
.B(n_213),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_434),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_446),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_446),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_517),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_448),
.B(n_335),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_448),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_454),
.B(n_279),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_454),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_456),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_456),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_460),
.B(n_463),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_460),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_463),
.B(n_337),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_468),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_468),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_423),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_477),
.B(n_340),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_477),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_480),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_480),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_482),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_482),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_484),
.B(n_341),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_484),
.B(n_485),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_485),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_491),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_452),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_471),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_491),
.B(n_352),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_494),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_494),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_495),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_495),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_499),
.B(n_357),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_499),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_501),
.B(n_290),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_501),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_507),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_507),
.B(n_363),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_438),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g595 ( 
.A(n_455),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_510),
.B(n_295),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_438),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_440),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_461),
.B(n_366),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_433),
.B(n_377),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_440),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_441),
.Y(n_602)
);

AND2x6_ASAP7_75t_L g603 ( 
.A(n_520),
.B(n_213),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_603),
.A2(n_561),
.B1(n_527),
.B2(n_590),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_550),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_550),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_554),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_522),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_539),
.B(n_437),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_581),
.B(n_541),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_522),
.Y(n_611)
);

INVx1_ASAP7_75t_SL g612 ( 
.A(n_539),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_523),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_529),
.B(n_437),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_523),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_601),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_556),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_525),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_582),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_525),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_532),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_524),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_556),
.Y(n_623)
);

INVx4_ASAP7_75t_L g624 ( 
.A(n_554),
.Y(n_624)
);

NAND2xp33_ASAP7_75t_SL g625 ( 
.A(n_581),
.B(n_464),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_532),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_534),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_534),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_540),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_540),
.Y(n_630)
);

OR2x6_ASAP7_75t_L g631 ( 
.A(n_521),
.B(n_511),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_600),
.B(n_465),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_526),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_556),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_536),
.B(n_418),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_596),
.B(n_474),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_542),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_542),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_526),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_599),
.B(n_466),
.Y(n_640)
);

BUFx10_ASAP7_75t_L g641 ( 
.A(n_595),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_556),
.Y(n_642)
);

BUFx2_ASAP7_75t_L g643 ( 
.A(n_546),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_590),
.B(n_596),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_545),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_545),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_603),
.A2(n_561),
.B1(n_590),
.B2(n_596),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_547),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_535),
.B(n_467),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_547),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_601),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_548),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_548),
.B(n_472),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_551),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_570),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_535),
.B(n_478),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_603),
.A2(n_561),
.B1(n_590),
.B2(n_596),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_551),
.Y(n_658)
);

INVx5_ASAP7_75t_L g659 ( 
.A(n_554),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_555),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_555),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_521),
.B(n_479),
.Y(n_662)
);

AND2x6_ASAP7_75t_L g663 ( 
.A(n_561),
.B(n_213),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_528),
.B(n_483),
.Y(n_664)
);

INVx6_ASAP7_75t_L g665 ( 
.A(n_556),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_560),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_560),
.Y(n_667)
);

INVx4_ASAP7_75t_L g668 ( 
.A(n_554),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_533),
.B(n_489),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_537),
.B(n_490),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_560),
.Y(n_671)
);

INVx5_ASAP7_75t_L g672 ( 
.A(n_554),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_560),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_558),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_582),
.B(n_416),
.Y(n_675)
);

AND2x6_ASAP7_75t_L g676 ( 
.A(n_563),
.B(n_213),
.Y(n_676)
);

XOR2xp5_ASAP7_75t_L g677 ( 
.A(n_543),
.B(n_427),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_552),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_563),
.B(n_497),
.Y(n_679)
);

OR2x6_ASAP7_75t_L g680 ( 
.A(n_565),
.B(n_514),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_560),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_560),
.Y(n_682)
);

NAND2x1p5_ASAP7_75t_L g683 ( 
.A(n_563),
.B(n_382),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_575),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_575),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_575),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_558),
.B(n_514),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_563),
.B(n_498),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_575),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_575),
.Y(n_690)
);

INVx6_ASAP7_75t_L g691 ( 
.A(n_575),
.Y(n_691)
);

BUFx4f_ASAP7_75t_L g692 ( 
.A(n_603),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_589),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_558),
.B(n_500),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_589),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_558),
.B(n_502),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_557),
.B(n_473),
.Y(n_697)
);

NOR2x1p5_ASAP7_75t_L g698 ( 
.A(n_597),
.B(n_504),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_589),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_589),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_589),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_589),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_566),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_566),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_566),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_568),
.Y(n_706)
);

OR2x6_ASAP7_75t_L g707 ( 
.A(n_578),
.B(n_519),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_557),
.B(n_506),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_568),
.Y(n_709)
);

AND2x6_ASAP7_75t_L g710 ( 
.A(n_562),
.B(n_242),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_568),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_562),
.B(n_512),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_569),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_597),
.B(n_493),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_564),
.B(n_516),
.Y(n_715)
);

AO22x1_ASAP7_75t_L g716 ( 
.A1(n_603),
.A2(n_227),
.B1(n_233),
.B2(n_221),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_603),
.A2(n_372),
.B1(n_344),
.B2(n_332),
.Y(n_717)
);

AND3x2_ASAP7_75t_L g718 ( 
.A(n_564),
.B(n_313),
.C(n_309),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_601),
.B(n_486),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_597),
.B(n_447),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_603),
.A2(n_481),
.B1(n_515),
.B2(n_381),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_572),
.B(n_573),
.Y(n_722)
);

INVx5_ASAP7_75t_L g723 ( 
.A(n_554),
.Y(n_723)
);

INVxp67_ASAP7_75t_SL g724 ( 
.A(n_553),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_597),
.Y(n_725)
);

AND2x6_ASAP7_75t_L g726 ( 
.A(n_572),
.B(n_242),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_569),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_L g728 ( 
.A1(n_573),
.A2(n_248),
.B1(n_373),
.B2(n_374),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_574),
.Y(n_729)
);

BUFx2_ASAP7_75t_L g730 ( 
.A(n_574),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_576),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_601),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_601),
.A2(n_379),
.B1(n_364),
.B2(n_319),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_569),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_576),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_579),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_601),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_602),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_602),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_602),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_602),
.A2(n_371),
.B1(n_404),
.B2(n_349),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_579),
.Y(n_742)
);

INVx6_ASAP7_75t_L g743 ( 
.A(n_602),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_580),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_602),
.Y(n_745)
);

CKINVDCx6p67_ASAP7_75t_R g746 ( 
.A(n_554),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_580),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_594),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_584),
.A2(n_321),
.B1(n_330),
.B2(n_324),
.Y(n_749)
);

INVx4_ASAP7_75t_L g750 ( 
.A(n_530),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_584),
.B(n_519),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_585),
.B(n_586),
.Y(n_752)
);

INVx1_ASAP7_75t_SL g753 ( 
.A(n_559),
.Y(n_753)
);

INVxp33_ASAP7_75t_L g754 ( 
.A(n_567),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_674),
.Y(n_755)
);

OAI221xp5_ASAP7_75t_L g756 ( 
.A1(n_749),
.A2(n_414),
.B1(n_251),
.B2(n_385),
.C(n_391),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_L g757 ( 
.A1(n_632),
.A2(n_604),
.B1(n_731),
.B2(n_657),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_753),
.B(n_492),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_724),
.B(n_496),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_692),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_643),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_712),
.B(n_503),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_658),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_622),
.A2(n_475),
.B1(n_476),
.B2(n_442),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_754),
.B(n_585),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_643),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_674),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_731),
.B(n_586),
.Y(n_768)
);

INVxp67_ASAP7_75t_L g769 ( 
.A(n_655),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_669),
.B(n_571),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_611),
.Y(n_771)
);

INVxp33_ASAP7_75t_L g772 ( 
.A(n_635),
.Y(n_772)
);

O2A1O1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_608),
.A2(n_620),
.B(n_621),
.C(n_613),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_658),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_692),
.B(n_209),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_660),
.Y(n_776)
);

AOI22x1_ASAP7_75t_L g777 ( 
.A1(n_611),
.A2(n_587),
.B1(n_591),
.B2(n_592),
.Y(n_777)
);

NAND2xp33_ASAP7_75t_L g778 ( 
.A(n_683),
.B(n_653),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_612),
.B(n_577),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_622),
.B(n_583),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_730),
.B(n_592),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_635),
.B(n_431),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_660),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_692),
.B(n_209),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_683),
.B(n_647),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_730),
.B(n_697),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_633),
.B(n_588),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_729),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_R g789 ( 
.A(n_625),
.B(n_436),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_655),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_633),
.B(n_593),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_729),
.B(n_509),
.Y(n_792)
);

INVxp67_ASAP7_75t_SL g793 ( 
.A(n_683),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_605),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_735),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_610),
.A2(n_391),
.B1(n_389),
.B2(n_388),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_639),
.B(n_425),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_735),
.B(n_598),
.Y(n_798)
);

OR2x2_ASAP7_75t_L g799 ( 
.A(n_675),
.B(n_439),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_747),
.B(n_598),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_747),
.Y(n_801)
);

INVxp67_ASAP7_75t_L g802 ( 
.A(n_675),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_615),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_639),
.A2(n_680),
.B1(n_707),
.B2(n_609),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_725),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_641),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_644),
.B(n_594),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_618),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_618),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_608),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_613),
.B(n_212),
.Y(n_811)
);

NAND3xp33_ASAP7_75t_L g812 ( 
.A(n_609),
.B(n_445),
.C(n_443),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_620),
.B(n_212),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_645),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_645),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_644),
.B(n_594),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_680),
.A2(n_449),
.B1(n_450),
.B2(n_451),
.Y(n_817)
);

NAND2xp33_ASAP7_75t_L g818 ( 
.A(n_679),
.B(n_214),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_650),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_621),
.B(n_214),
.Y(n_820)
);

NOR3xp33_ASAP7_75t_L g821 ( 
.A(n_640),
.B(n_233),
.C(n_227),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_725),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_680),
.B(n_232),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_626),
.Y(n_824)
);

O2A1O1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_626),
.A2(n_441),
.B(n_444),
.C(n_411),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_680),
.B(n_274),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_614),
.B(n_346),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_614),
.B(n_347),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_680),
.B(n_283),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_707),
.B(n_285),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_627),
.B(n_215),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_L g832 ( 
.A1(n_707),
.A2(n_250),
.B1(n_385),
.B2(n_248),
.Y(n_832)
);

NAND2xp33_ASAP7_75t_SL g833 ( 
.A(n_698),
.B(n_240),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_636),
.B(n_429),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_627),
.B(n_215),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_677),
.Y(n_836)
);

NAND3xp33_ASAP7_75t_SL g837 ( 
.A(n_619),
.B(n_243),
.C(n_240),
.Y(n_837)
);

AO221x1_ASAP7_75t_L g838 ( 
.A1(n_728),
.A2(n_716),
.B1(n_634),
.B2(n_682),
.C(n_740),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_707),
.B(n_310),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_628),
.B(n_216),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_636),
.B(n_457),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_707),
.B(n_395),
.Y(n_842)
);

BUFx5_ASAP7_75t_L g843 ( 
.A(n_676),
.Y(n_843)
);

BUFx3_ASAP7_75t_L g844 ( 
.A(n_700),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_650),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_636),
.B(n_458),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_736),
.A2(n_235),
.B1(n_270),
.B2(n_396),
.Y(n_847)
);

OAI22xp33_ASAP7_75t_L g848 ( 
.A1(n_721),
.A2(n_246),
.B1(n_243),
.B2(n_250),
.Y(n_848)
);

OAI22xp5_ASAP7_75t_L g849 ( 
.A1(n_688),
.A2(n_246),
.B1(n_388),
.B2(n_389),
.Y(n_849)
);

A2O1A1Ixp33_ASAP7_75t_L g850 ( 
.A1(n_736),
.A2(n_405),
.B(n_375),
.C(n_374),
.Y(n_850)
);

OR2x2_ASAP7_75t_L g851 ( 
.A(n_619),
.B(n_462),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_714),
.B(n_216),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_636),
.B(n_641),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_628),
.B(n_218),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_661),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_700),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_708),
.B(n_353),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_629),
.B(n_218),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_714),
.B(n_225),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_661),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_665),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_714),
.B(n_225),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_714),
.B(n_231),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_706),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_715),
.B(n_358),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_706),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_631),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_630),
.B(n_231),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_720),
.B(n_238),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_720),
.B(n_238),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_720),
.B(n_751),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_641),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_720),
.B(n_239),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_637),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_638),
.Y(n_875)
);

INVxp67_ASAP7_75t_SL g876 ( 
.A(n_739),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_638),
.B(n_239),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_646),
.B(n_252),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_646),
.B(n_648),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_641),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_709),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_677),
.B(n_444),
.Y(n_882)
);

BUFx3_ASAP7_75t_L g883 ( 
.A(n_665),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_648),
.B(n_652),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_751),
.B(n_687),
.Y(n_885)
);

AND2x6_ASAP7_75t_L g886 ( 
.A(n_721),
.B(n_242),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_687),
.B(n_252),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_652),
.Y(n_888)
);

NAND2x1_ASAP7_75t_L g889 ( 
.A(n_624),
.B(n_530),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_665),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_654),
.B(n_378),
.Y(n_891)
);

NAND3xp33_ASAP7_75t_L g892 ( 
.A(n_649),
.B(n_375),
.C(n_403),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_654),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_631),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_698),
.A2(n_380),
.B1(n_402),
.B2(n_387),
.Y(n_895)
);

BUFx5_ASAP7_75t_L g896 ( 
.A(n_676),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_616),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_742),
.A2(n_235),
.B1(n_396),
.B2(n_270),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_656),
.A2(n_631),
.B1(n_664),
.B2(n_670),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_744),
.B(n_380),
.Y(n_900)
);

AND2x6_ASAP7_75t_SL g901 ( 
.A(n_662),
.B(n_373),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_694),
.B(n_367),
.Y(n_902)
);

AND2x6_ASAP7_75t_L g903 ( 
.A(n_744),
.B(n_703),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_722),
.A2(n_384),
.B(n_390),
.C(n_538),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_631),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_678),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_752),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_709),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_703),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_704),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_606),
.B(n_387),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_606),
.B(n_394),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_704),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_705),
.B(n_394),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_631),
.A2(n_401),
.B1(n_403),
.B2(n_381),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_716),
.A2(n_399),
.B1(n_402),
.B2(n_408),
.Y(n_916)
);

O2A1O1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_696),
.A2(n_544),
.B(n_538),
.C(n_549),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_705),
.B(n_399),
.Y(n_918)
);

NOR3xp33_ASAP7_75t_L g919 ( 
.A(n_762),
.B(n_719),
.C(n_370),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_770),
.A2(n_713),
.B(n_748),
.C(n_727),
.Y(n_920)
);

NAND3xp33_ASAP7_75t_L g921 ( 
.A(n_786),
.B(n_717),
.C(n_713),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_760),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_778),
.A2(n_623),
.B(n_617),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_871),
.A2(n_682),
.B(n_737),
.C(n_740),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_770),
.B(n_711),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_805),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_779),
.B(n_711),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_879),
.A2(n_623),
.B(n_617),
.Y(n_928)
);

BUFx2_ASAP7_75t_L g929 ( 
.A(n_761),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_810),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_824),
.Y(n_931)
);

INVx4_ASAP7_75t_L g932 ( 
.A(n_903),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_757),
.A2(n_737),
.B(n_740),
.C(n_732),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_779),
.B(n_727),
.Y(n_934)
);

INVx1_ASAP7_75t_SL g935 ( 
.A(n_766),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_879),
.A2(n_623),
.B(n_617),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_760),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_780),
.B(n_734),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_884),
.A2(n_642),
.B(n_634),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_780),
.B(n_734),
.Y(n_940)
);

AOI22xp5_ASAP7_75t_L g941 ( 
.A1(n_857),
.A2(n_678),
.B1(n_663),
.B2(n_691),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_874),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_760),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_884),
.A2(n_642),
.B(n_634),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_773),
.A2(n_667),
.B(n_666),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_807),
.A2(n_667),
.B(n_666),
.Y(n_946)
);

CKINVDCx6p67_ASAP7_75t_R g947 ( 
.A(n_851),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_768),
.A2(n_682),
.B(n_642),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_775),
.A2(n_732),
.B(n_699),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_775),
.A2(n_732),
.B(n_699),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_R g951 ( 
.A(n_806),
.B(n_746),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_857),
.A2(n_663),
.B1(n_691),
.B2(n_743),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_794),
.Y(n_953)
);

NOR3xp33_ASAP7_75t_L g954 ( 
.A(n_782),
.B(n_369),
.C(n_401),
.Y(n_954)
);

O2A1O1Ixp5_ASAP7_75t_L g955 ( 
.A1(n_784),
.A2(n_902),
.B(n_865),
.C(n_813),
.Y(n_955)
);

NOR2x1_ASAP7_75t_R g956 ( 
.A(n_834),
.B(n_405),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_787),
.B(n_748),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_865),
.A2(n_663),
.B1(n_691),
.B2(n_743),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_784),
.A2(n_737),
.B(n_699),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_875),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_907),
.A2(n_673),
.B(n_671),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_769),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_787),
.B(n_791),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_791),
.B(n_663),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_790),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_802),
.B(n_733),
.Y(n_966)
);

CKINVDCx10_ASAP7_75t_R g967 ( 
.A(n_772),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_864),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_760),
.B(n_616),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_885),
.B(n_663),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_793),
.A2(n_673),
.B(n_671),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_902),
.B(n_663),
.Y(n_972)
);

OAI21xp33_ASAP7_75t_L g973 ( 
.A1(n_827),
.A2(n_828),
.B(n_916),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_827),
.B(n_663),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_804),
.B(n_616),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_816),
.A2(n_695),
.B(n_689),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_828),
.B(n_741),
.Y(n_977)
);

AOI22xp5_ASAP7_75t_L g978 ( 
.A1(n_853),
.A2(n_665),
.B1(n_691),
.B2(n_743),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_781),
.B(n_689),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_909),
.A2(n_695),
.B(n_701),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_910),
.A2(n_701),
.B(n_745),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_866),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_913),
.A2(n_690),
.B(n_745),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_888),
.Y(n_984)
);

BUFx4f_ASAP7_75t_L g985 ( 
.A(n_841),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_771),
.A2(n_686),
.B(n_738),
.Y(n_986)
);

AOI22xp5_ASAP7_75t_L g987 ( 
.A1(n_848),
.A2(n_743),
.B1(n_681),
.B2(n_684),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_893),
.A2(n_690),
.B(n_738),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_798),
.A2(n_684),
.B(n_681),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_765),
.B(n_887),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_800),
.A2(n_702),
.B(n_693),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_889),
.A2(n_702),
.B(n_693),
.Y(n_992)
);

OAI21xp33_ASAP7_75t_L g993 ( 
.A1(n_832),
.A2(n_859),
.B(n_852),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_899),
.A2(n_686),
.B(n_685),
.C(n_413),
.Y(n_994)
);

BUFx2_ASAP7_75t_SL g995 ( 
.A(n_906),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_867),
.B(n_616),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_867),
.B(n_616),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_914),
.A2(n_685),
.B(n_651),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_846),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_918),
.A2(n_651),
.B(n_750),
.Y(n_1000)
);

O2A1O1Ixp5_ASAP7_75t_L g1001 ( 
.A1(n_811),
.A2(n_750),
.B(n_607),
.C(n_624),
.Y(n_1001)
);

O2A1O1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_848),
.A2(n_538),
.B(n_544),
.C(n_549),
.Y(n_1002)
);

OAI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_803),
.A2(n_750),
.B(n_668),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_755),
.A2(n_651),
.B(n_750),
.Y(n_1004)
);

AO21x1_ASAP7_75t_L g1005 ( 
.A1(n_785),
.A2(n_624),
.B(n_668),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_767),
.A2(n_651),
.B(n_624),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_805),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_881),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_789),
.Y(n_1009)
);

NAND2x1p5_ASAP7_75t_L g1010 ( 
.A(n_822),
.B(n_668),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_759),
.B(n_607),
.Y(n_1011)
);

BUFx3_ASAP7_75t_L g1012 ( 
.A(n_822),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_850),
.A2(n_915),
.B(n_849),
.C(n_796),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_823),
.B(n_826),
.Y(n_1014)
);

NOR3xp33_ASAP7_75t_L g1015 ( 
.A(n_837),
.B(n_892),
.C(n_797),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_829),
.B(n_607),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_882),
.B(n_406),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_799),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_900),
.A2(n_723),
.B(n_672),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_818),
.A2(n_723),
.B(n_672),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_808),
.A2(n_723),
.B(n_672),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_908),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_894),
.B(n_659),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_830),
.B(n_839),
.Y(n_1024)
);

BUFx4f_ASAP7_75t_L g1025 ( 
.A(n_872),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_844),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_809),
.Y(n_1027)
);

HB1xp67_ASAP7_75t_L g1028 ( 
.A(n_894),
.Y(n_1028)
);

NAND2xp33_ASAP7_75t_L g1029 ( 
.A(n_903),
.B(n_897),
.Y(n_1029)
);

NAND2xp33_ASAP7_75t_L g1030 ( 
.A(n_903),
.B(n_897),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_758),
.B(n_406),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_792),
.B(n_718),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_814),
.A2(n_723),
.B(n_672),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_842),
.B(n_746),
.Y(n_1034)
);

INVx2_ASAP7_75t_SL g1035 ( 
.A(n_880),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_897),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_763),
.B(n_407),
.Y(n_1037)
);

AOI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_886),
.A2(n_270),
.B1(n_410),
.B2(n_396),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_815),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_850),
.A2(n_544),
.B(n_549),
.C(n_531),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_774),
.B(n_407),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_819),
.Y(n_1042)
);

OR2x6_ASAP7_75t_L g1043 ( 
.A(n_812),
.B(n_242),
.Y(n_1043)
);

AO21x1_ASAP7_75t_L g1044 ( 
.A1(n_785),
.A2(n_531),
.B(n_410),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_845),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_776),
.B(n_783),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_855),
.A2(n_723),
.B(n_659),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_788),
.B(n_413),
.Y(n_1048)
);

O2A1O1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_811),
.A2(n_5),
.B(n_9),
.C(n_12),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_860),
.A2(n_676),
.B(n_723),
.Y(n_1050)
);

OAI21xp33_ASAP7_75t_L g1051 ( 
.A1(n_862),
.A2(n_412),
.B(n_408),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_795),
.B(n_412),
.Y(n_1052)
);

OAI21xp33_ASAP7_75t_L g1053 ( 
.A1(n_863),
.A2(n_275),
.B(n_267),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_797),
.B(n_410),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_911),
.A2(n_659),
.B(n_672),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_912),
.A2(n_659),
.B(n_672),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_869),
.A2(n_873),
.B(n_870),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_825),
.A2(n_393),
.B(n_301),
.C(n_242),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_813),
.A2(n_877),
.B(n_835),
.C(n_854),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_820),
.A2(n_659),
.B(n_255),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_756),
.A2(n_393),
.B(n_301),
.C(n_280),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_801),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_876),
.B(n_676),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_847),
.B(n_676),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_897),
.B(n_659),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_847),
.B(n_676),
.Y(n_1066)
);

OAI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_777),
.A2(n_676),
.B(n_726),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_820),
.A2(n_316),
.B(n_265),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_831),
.A2(n_317),
.B(n_281),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_844),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_898),
.B(n_263),
.Y(n_1071)
);

AOI22x1_ASAP7_75t_L g1072 ( 
.A1(n_905),
.A2(n_838),
.B1(n_903),
.B2(n_917),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_831),
.A2(n_331),
.B(n_296),
.Y(n_1073)
);

AO21x1_ASAP7_75t_L g1074 ( 
.A1(n_835),
.A2(n_726),
.B(n_710),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_861),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_840),
.A2(n_334),
.B(n_298),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_898),
.B(n_286),
.Y(n_1077)
);

AO21x1_ASAP7_75t_L g1078 ( 
.A1(n_840),
.A2(n_726),
.B(n_710),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_764),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_854),
.A2(n_726),
.B(n_710),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_858),
.A2(n_348),
.B(n_303),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_858),
.B(n_305),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_856),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_868),
.B(n_311),
.Y(n_1084)
);

BUFx12f_ASAP7_75t_L g1085 ( 
.A(n_901),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_868),
.A2(n_355),
.B(n_312),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_856),
.B(n_301),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_861),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_883),
.Y(n_1089)
);

NAND2x1p5_ASAP7_75t_L g1090 ( 
.A(n_883),
.B(n_301),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_877),
.A2(n_878),
.B(n_891),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_878),
.A2(n_356),
.B(n_314),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_891),
.B(n_9),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_890),
.A2(n_361),
.B(n_327),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_890),
.B(n_393),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_903),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_843),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_821),
.A2(n_13),
.B(n_15),
.C(n_18),
.Y(n_1098)
);

INVx2_ASAP7_75t_SL g1099 ( 
.A(n_789),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_895),
.B(n_365),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_843),
.Y(n_1101)
);

NOR3xp33_ASAP7_75t_L g1102 ( 
.A(n_833),
.B(n_350),
.C(n_19),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_935),
.B(n_817),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_1036),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_930),
.Y(n_1105)
);

AO21x2_ASAP7_75t_L g1106 ( 
.A1(n_1044),
.A2(n_904),
.B(n_886),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_973),
.A2(n_886),
.B(n_836),
.C(n_393),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_955),
.A2(n_886),
.B(n_393),
.C(n_301),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_1093),
.A2(n_886),
.B(n_896),
.C(n_843),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_963),
.A2(n_896),
.B(n_843),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_1093),
.A2(n_896),
.B(n_843),
.C(n_726),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_925),
.A2(n_18),
.B1(n_22),
.B2(n_24),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_SL g1113 ( 
.A(n_932),
.B(n_896),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_1036),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_931),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_938),
.A2(n_896),
.B(n_843),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_1036),
.Y(n_1117)
);

AOI22xp33_ASAP7_75t_L g1118 ( 
.A1(n_1079),
.A2(n_896),
.B1(n_726),
.B2(n_710),
.Y(n_1118)
);

OR2x6_ASAP7_75t_L g1119 ( 
.A(n_1099),
.B(n_726),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_1018),
.B(n_27),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_1013),
.A2(n_710),
.B(n_29),
.C(n_30),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_990),
.B(n_27),
.Y(n_1122)
);

NAND3xp33_ASAP7_75t_L g1123 ( 
.A(n_954),
.B(n_29),
.C(n_31),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_927),
.B(n_32),
.Y(n_1124)
);

NOR2xp67_ASAP7_75t_SL g1125 ( 
.A(n_1018),
.B(n_33),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_934),
.B(n_33),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_929),
.B(n_710),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_965),
.B(n_710),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_940),
.A2(n_81),
.B(n_190),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_957),
.A2(n_78),
.B(n_182),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_942),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_R g1132 ( 
.A(n_1009),
.B(n_73),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_962),
.B(n_35),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1014),
.B(n_38),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_960),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1029),
.A2(n_83),
.B(n_171),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1024),
.B(n_41),
.Y(n_1137)
);

OR2x2_ASAP7_75t_L g1138 ( 
.A(n_1017),
.B(n_43),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1030),
.A2(n_87),
.B(n_160),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_966),
.B(n_45),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_947),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_R g1142 ( 
.A(n_967),
.B(n_90),
.Y(n_1142)
);

INVx4_ASAP7_75t_L g1143 ( 
.A(n_932),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_985),
.Y(n_1144)
);

INVx5_ASAP7_75t_L g1145 ( 
.A(n_1036),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_972),
.A2(n_72),
.B(n_158),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_962),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1054),
.B(n_46),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_985),
.Y(n_1149)
);

INVxp67_ASAP7_75t_L g1150 ( 
.A(n_999),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_999),
.B(n_1031),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_1028),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1028),
.B(n_48),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_926),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_956),
.B(n_49),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1057),
.A2(n_98),
.B(n_154),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_977),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_984),
.B(n_53),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1011),
.B(n_54),
.Y(n_1159)
);

NAND2x1p5_ASAP7_75t_L g1160 ( 
.A(n_926),
.B(n_108),
.Y(n_1160)
);

CKINVDCx8_ASAP7_75t_R g1161 ( 
.A(n_995),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_954),
.B(n_54),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_1098),
.A2(n_57),
.B(n_58),
.C(n_59),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_979),
.A2(n_61),
.B1(n_64),
.B2(n_66),
.Y(n_1164)
);

AO32x1_ASAP7_75t_L g1165 ( 
.A1(n_1039),
.A2(n_64),
.A3(n_68),
.B1(n_94),
.B2(n_110),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_1011),
.B(n_115),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1032),
.B(n_119),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_1059),
.A2(n_124),
.B(n_128),
.C(n_131),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_993),
.A2(n_138),
.B(n_144),
.C(n_199),
.Y(n_1169)
);

BUFx12f_ASAP7_75t_L g1170 ( 
.A(n_1085),
.Y(n_1170)
);

AO21x1_ASAP7_75t_L g1171 ( 
.A1(n_1091),
.A2(n_975),
.B(n_974),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_998),
.A2(n_923),
.B(n_1000),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_964),
.A2(n_1025),
.B1(n_1096),
.B2(n_941),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_988),
.A2(n_920),
.B(n_976),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_1007),
.Y(n_1175)
);

OR2x6_ASAP7_75t_L g1176 ( 
.A(n_1096),
.B(n_1007),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1012),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1012),
.Y(n_1178)
);

AND2x6_ASAP7_75t_L g1179 ( 
.A(n_943),
.B(n_922),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1025),
.B(n_951),
.Y(n_1180)
);

BUFx8_ASAP7_75t_L g1181 ( 
.A(n_1035),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_951),
.B(n_919),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_1032),
.B(n_1062),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1070),
.Y(n_1184)
);

INVxp67_ASAP7_75t_L g1185 ( 
.A(n_1037),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1015),
.A2(n_1102),
.B(n_1049),
.C(n_1052),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_921),
.A2(n_970),
.B1(n_1100),
.B2(n_1038),
.Y(n_1187)
);

NAND2x1p5_ASAP7_75t_L g1188 ( 
.A(n_1026),
.B(n_1089),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_919),
.B(n_1015),
.Y(n_1189)
);

INVx2_ASAP7_75t_SL g1190 ( 
.A(n_1083),
.Y(n_1190)
);

O2A1O1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1102),
.A2(n_1082),
.B(n_1084),
.C(n_1048),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_953),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1071),
.B(n_1077),
.Y(n_1193)
);

INVx1_ASAP7_75t_SL g1194 ( 
.A(n_1026),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_943),
.B(n_1089),
.Y(n_1195)
);

INVxp67_ASAP7_75t_L g1196 ( 
.A(n_1037),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_1010),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_1043),
.Y(n_1198)
);

NOR3xp33_ASAP7_75t_SL g1199 ( 
.A(n_1041),
.B(n_1051),
.C(n_1076),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_SL g1200 ( 
.A1(n_920),
.A2(n_969),
.B(n_1061),
.C(n_933),
.Y(n_1200)
);

AO21x1_ASAP7_75t_L g1201 ( 
.A1(n_975),
.A2(n_946),
.B(n_924),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1043),
.B(n_1042),
.Y(n_1202)
);

INVxp67_ASAP7_75t_L g1203 ( 
.A(n_1043),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_943),
.B(n_922),
.Y(n_1204)
);

NAND3xp33_ASAP7_75t_L g1205 ( 
.A(n_1061),
.B(n_994),
.C(n_1038),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_943),
.B(n_1034),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_981),
.A2(n_983),
.B(n_961),
.Y(n_1207)
);

AO32x1_ASAP7_75t_L g1208 ( 
.A1(n_968),
.A2(n_982),
.A3(n_1008),
.B1(n_1045),
.B2(n_1027),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1046),
.B(n_1053),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1075),
.B(n_1088),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_994),
.A2(n_1001),
.B(n_945),
.C(n_1040),
.Y(n_1211)
);

OR2x2_ASAP7_75t_L g1212 ( 
.A(n_1022),
.B(n_1008),
.Y(n_1212)
);

OAI22x1_ASAP7_75t_L g1213 ( 
.A1(n_1072),
.A2(n_996),
.B1(n_997),
.B2(n_987),
.Y(n_1213)
);

BUFx4f_ASAP7_75t_L g1214 ( 
.A(n_937),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_937),
.B(n_978),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1064),
.B(n_1066),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_949),
.A2(n_950),
.B(n_959),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_996),
.Y(n_1218)
);

INVx1_ASAP7_75t_SL g1219 ( 
.A(n_997),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1016),
.B(n_1023),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_948),
.A2(n_928),
.B(n_936),
.Y(n_1221)
);

BUFx3_ASAP7_75t_L g1222 ( 
.A(n_1010),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1023),
.B(n_1097),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_986),
.Y(n_1224)
);

AOI21x1_ASAP7_75t_L g1225 ( 
.A1(n_969),
.A2(n_1087),
.B(n_991),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1068),
.B(n_1081),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1090),
.Y(n_1227)
);

BUFx10_ASAP7_75t_L g1228 ( 
.A(n_1069),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1097),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1090),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_939),
.A2(n_944),
.B(n_992),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_980),
.A2(n_989),
.B(n_1004),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1002),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_952),
.A2(n_958),
.B1(n_1063),
.B2(n_1058),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1073),
.B(n_1092),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1086),
.A2(n_1005),
.B1(n_1003),
.B2(n_1074),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1087),
.B(n_1094),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_971),
.B(n_1095),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1006),
.A2(n_1101),
.B1(n_1060),
.B2(n_1065),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1065),
.A2(n_1058),
.B1(n_1067),
.B2(n_1080),
.Y(n_1240)
);

OAI22x1_ASAP7_75t_L g1241 ( 
.A1(n_1095),
.A2(n_1078),
.B1(n_1050),
.B2(n_1021),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1033),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1019),
.B(n_1055),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1056),
.B(n_1020),
.Y(n_1244)
);

INVx4_ASAP7_75t_L g1245 ( 
.A(n_1047),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_963),
.B(n_786),
.Y(n_1246)
);

INVx1_ASAP7_75t_SL g1247 ( 
.A(n_935),
.Y(n_1247)
);

HB1xp67_ASAP7_75t_L g1248 ( 
.A(n_929),
.Y(n_1248)
);

HB1xp67_ASAP7_75t_L g1249 ( 
.A(n_929),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_973),
.A2(n_955),
.B(n_1093),
.C(n_1013),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_963),
.A2(n_925),
.B(n_778),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_963),
.A2(n_925),
.B(n_778),
.Y(n_1252)
);

NOR2xp67_ASAP7_75t_L g1253 ( 
.A(n_932),
.B(n_1026),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_929),
.Y(n_1254)
);

AO31x2_ASAP7_75t_L g1255 ( 
.A1(n_1171),
.A2(n_1201),
.A3(n_1250),
.B(n_1241),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1232),
.A2(n_1231),
.B(n_1172),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1246),
.B(n_1220),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_1181),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1212),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1185),
.A2(n_1196),
.B1(n_1189),
.B2(n_1122),
.Y(n_1260)
);

AO32x2_ASAP7_75t_L g1261 ( 
.A1(n_1112),
.A2(n_1164),
.A3(n_1187),
.B1(n_1157),
.B2(n_1234),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1221),
.A2(n_1217),
.B(n_1207),
.Y(n_1262)
);

AO31x2_ASAP7_75t_L g1263 ( 
.A1(n_1213),
.A2(n_1108),
.A3(n_1240),
.B(n_1211),
.Y(n_1263)
);

INVx6_ASAP7_75t_L g1264 ( 
.A(n_1181),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_SL g1265 ( 
.A1(n_1191),
.A2(n_1186),
.B(n_1168),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1105),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1225),
.A2(n_1243),
.B(n_1174),
.Y(n_1267)
);

NOR4xp25_ASAP7_75t_L g1268 ( 
.A(n_1112),
.B(n_1123),
.C(n_1163),
.D(n_1164),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1166),
.A2(n_1110),
.B(n_1200),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1115),
.Y(n_1270)
);

BUFx10_ASAP7_75t_L g1271 ( 
.A(n_1120),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1239),
.A2(n_1244),
.B(n_1216),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1242),
.A2(n_1238),
.B(n_1116),
.Y(n_1273)
);

O2A1O1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1148),
.A2(n_1162),
.B(n_1159),
.C(n_1121),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1236),
.A2(n_1156),
.B(n_1234),
.Y(n_1275)
);

AOI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1151),
.A2(n_1123),
.B1(n_1140),
.B2(n_1133),
.Y(n_1276)
);

AO31x2_ASAP7_75t_L g1277 ( 
.A1(n_1107),
.A2(n_1224),
.A3(n_1109),
.B(n_1111),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1146),
.A2(n_1235),
.B(n_1206),
.Y(n_1278)
);

AO31x2_ASAP7_75t_L g1279 ( 
.A1(n_1169),
.A2(n_1226),
.A3(n_1173),
.B(n_1193),
.Y(n_1279)
);

A2O1A1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_1209),
.A2(n_1205),
.B(n_1167),
.C(n_1134),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1113),
.A2(n_1126),
.B(n_1124),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_1144),
.B(n_1149),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1237),
.A2(n_1136),
.B(n_1139),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1141),
.Y(n_1284)
);

NOR2xp67_ASAP7_75t_L g1285 ( 
.A(n_1180),
.B(n_1248),
.Y(n_1285)
);

NAND3xp33_ASAP7_75t_L g1286 ( 
.A(n_1199),
.B(n_1125),
.C(n_1205),
.Y(n_1286)
);

OR2x2_ASAP7_75t_L g1287 ( 
.A(n_1247),
.B(n_1152),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1137),
.A2(n_1138),
.B1(n_1158),
.B2(n_1153),
.Y(n_1288)
);

A2O1A1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1183),
.A2(n_1210),
.B(n_1218),
.C(n_1182),
.Y(n_1289)
);

AOI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1233),
.A2(n_1215),
.B(n_1128),
.Y(n_1290)
);

A2O1A1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_1219),
.A2(n_1214),
.B(n_1155),
.C(n_1253),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1113),
.A2(n_1130),
.B(n_1129),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1229),
.A2(n_1197),
.B(n_1160),
.Y(n_1293)
);

AOI31xp67_ASAP7_75t_L g1294 ( 
.A1(n_1227),
.A2(n_1223),
.A3(n_1195),
.B(n_1127),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1131),
.B(n_1135),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1150),
.A2(n_1194),
.B1(n_1103),
.B2(n_1143),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1194),
.B(n_1223),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1253),
.A2(n_1245),
.B(n_1219),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_1249),
.Y(n_1299)
);

AOI21xp33_ASAP7_75t_L g1300 ( 
.A1(n_1203),
.A2(n_1198),
.B(n_1106),
.Y(n_1300)
);

AO21x1_ASAP7_75t_L g1301 ( 
.A1(n_1160),
.A2(n_1202),
.B(n_1188),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1229),
.A2(n_1165),
.B(n_1143),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1165),
.A2(n_1145),
.B(n_1188),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1214),
.A2(n_1176),
.B1(n_1254),
.B2(n_1161),
.Y(n_1304)
);

INVx1_ASAP7_75t_SL g1305 ( 
.A(n_1247),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1184),
.B(n_1178),
.Y(n_1306)
);

AO31x2_ASAP7_75t_L g1307 ( 
.A1(n_1208),
.A2(n_1192),
.A3(n_1165),
.B(n_1228),
.Y(n_1307)
);

AO31x2_ASAP7_75t_L g1308 ( 
.A1(n_1208),
.A2(n_1228),
.A3(n_1176),
.B(n_1118),
.Y(n_1308)
);

O2A1O1Ixp33_ASAP7_75t_SL g1309 ( 
.A1(n_1197),
.A2(n_1190),
.B(n_1145),
.C(n_1179),
.Y(n_1309)
);

OR2x2_ASAP7_75t_L g1310 ( 
.A(n_1154),
.B(n_1175),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1154),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1175),
.B(n_1178),
.Y(n_1312)
);

O2A1O1Ixp5_ASAP7_75t_L g1313 ( 
.A1(n_1204),
.A2(n_1179),
.B(n_1145),
.C(n_1117),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1177),
.Y(n_1314)
);

AO31x2_ASAP7_75t_L g1315 ( 
.A1(n_1208),
.A2(n_1230),
.A3(n_1179),
.B(n_1222),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1177),
.A2(n_1178),
.B1(n_1119),
.B2(n_1117),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1230),
.A2(n_1104),
.B(n_1114),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1230),
.A2(n_1104),
.B(n_1114),
.Y(n_1318)
);

BUFx8_ASAP7_75t_L g1319 ( 
.A(n_1170),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1104),
.A2(n_1114),
.B(n_1117),
.Y(n_1320)
);

CKINVDCx11_ASAP7_75t_R g1321 ( 
.A(n_1177),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1204),
.Y(n_1322)
);

NAND3xp33_ASAP7_75t_L g1323 ( 
.A(n_1119),
.B(n_1132),
.C(n_1142),
.Y(n_1323)
);

A2O1A1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1119),
.A2(n_973),
.B(n_1193),
.C(n_955),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1246),
.B(n_963),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1105),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1246),
.B(n_963),
.Y(n_1327)
);

AOI221xp5_ASAP7_75t_SL g1328 ( 
.A1(n_1112),
.A2(n_1164),
.B1(n_973),
.B2(n_1013),
.C(n_1157),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1185),
.B(n_851),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1212),
.Y(n_1330)
);

AOI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1185),
.A2(n_973),
.B1(n_1093),
.B2(n_1018),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1212),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1232),
.A2(n_1231),
.B(n_1172),
.Y(n_1333)
);

OAI221xp5_ASAP7_75t_L g1334 ( 
.A1(n_1185),
.A2(n_973),
.B1(n_954),
.B2(n_632),
.C(n_762),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1232),
.A2(n_1231),
.B(n_1172),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1232),
.A2(n_1231),
.B(n_1172),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1144),
.B(n_1149),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1105),
.Y(n_1338)
);

BUFx3_ASAP7_75t_L g1339 ( 
.A(n_1181),
.Y(n_1339)
);

BUFx8_ASAP7_75t_L g1340 ( 
.A(n_1170),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1246),
.B(n_963),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1246),
.B(n_963),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1105),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1147),
.B(n_1018),
.Y(n_1344)
);

AOI221x1_ASAP7_75t_L g1345 ( 
.A1(n_1250),
.A2(n_973),
.B1(n_1205),
.B2(n_1123),
.C(n_1112),
.Y(n_1345)
);

AO31x2_ASAP7_75t_L g1346 ( 
.A1(n_1171),
.A2(n_1044),
.A3(n_1201),
.B(n_1250),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1212),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1105),
.Y(n_1348)
);

AOI221x1_ASAP7_75t_L g1349 ( 
.A1(n_1250),
.A2(n_973),
.B1(n_1205),
.B2(n_1123),
.C(n_1112),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1232),
.A2(n_1231),
.B(n_1172),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1232),
.A2(n_1231),
.B(n_1172),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1105),
.Y(n_1352)
);

AO31x2_ASAP7_75t_L g1353 ( 
.A1(n_1171),
.A2(n_1044),
.A3(n_1201),
.B(n_1250),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1246),
.A2(n_963),
.B1(n_973),
.B2(n_1185),
.Y(n_1354)
);

AOI221x1_ASAP7_75t_L g1355 ( 
.A1(n_1250),
.A2(n_973),
.B1(n_1205),
.B2(n_1123),
.C(n_1112),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1105),
.Y(n_1356)
);

O2A1O1Ixp33_ASAP7_75t_SL g1357 ( 
.A1(n_1246),
.A2(n_963),
.B(n_1250),
.C(n_973),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1185),
.B(n_851),
.Y(n_1358)
);

O2A1O1Ixp33_ASAP7_75t_SL g1359 ( 
.A1(n_1246),
.A2(n_963),
.B(n_1250),
.C(n_973),
.Y(n_1359)
);

INVx3_ASAP7_75t_L g1360 ( 
.A(n_1143),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1105),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1143),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1232),
.A2(n_1231),
.B(n_1172),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1232),
.A2(n_1231),
.B(n_1172),
.Y(n_1364)
);

OA21x2_ASAP7_75t_L g1365 ( 
.A1(n_1172),
.A2(n_1221),
.B(n_1217),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1246),
.B(n_963),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1246),
.B(n_963),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_1185),
.B(n_963),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1212),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1246),
.B(n_963),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1212),
.Y(n_1371)
);

A2O1A1Ixp33_ASAP7_75t_L g1372 ( 
.A1(n_1193),
.A2(n_973),
.B(n_955),
.C(n_1191),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1151),
.B(n_1017),
.Y(n_1373)
);

O2A1O1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1185),
.A2(n_973),
.B(n_632),
.C(n_1196),
.Y(n_1374)
);

O2A1O1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1185),
.A2(n_973),
.B(n_632),
.C(n_1196),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1232),
.A2(n_1231),
.B(n_1172),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1232),
.A2(n_1231),
.B(n_1172),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1105),
.Y(n_1378)
);

AOI221xp5_ASAP7_75t_L g1379 ( 
.A1(n_1185),
.A2(n_954),
.B1(n_973),
.B2(n_827),
.C(n_828),
.Y(n_1379)
);

AO31x2_ASAP7_75t_L g1380 ( 
.A1(n_1171),
.A2(n_1044),
.A3(n_1201),
.B(n_1250),
.Y(n_1380)
);

INVx1_ASAP7_75t_SL g1381 ( 
.A(n_1247),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1246),
.B(n_963),
.Y(n_1382)
);

AOI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1243),
.A2(n_1231),
.B(n_1172),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1147),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1185),
.B(n_851),
.Y(n_1385)
);

OAI21xp5_ASAP7_75t_SL g1386 ( 
.A1(n_1162),
.A2(n_973),
.B(n_1123),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1212),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1181),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1144),
.B(n_1149),
.Y(n_1389)
);

AO31x2_ASAP7_75t_L g1390 ( 
.A1(n_1171),
.A2(n_1044),
.A3(n_1201),
.B(n_1250),
.Y(n_1390)
);

A2O1A1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1193),
.A2(n_973),
.B(n_955),
.C(n_1191),
.Y(n_1391)
);

INVx3_ASAP7_75t_L g1392 ( 
.A(n_1143),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1232),
.A2(n_1231),
.B(n_1172),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1246),
.A2(n_963),
.B1(n_973),
.B2(n_1185),
.Y(n_1394)
);

A2O1A1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1193),
.A2(n_973),
.B(n_955),
.C(n_1191),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1105),
.Y(n_1396)
);

OA21x2_ASAP7_75t_L g1397 ( 
.A1(n_1172),
.A2(n_1221),
.B(n_1217),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1147),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1251),
.A2(n_1252),
.B(n_1030),
.Y(n_1399)
);

AND2x4_ASAP7_75t_L g1400 ( 
.A(n_1144),
.B(n_1149),
.Y(n_1400)
);

OAI22x1_ASAP7_75t_L g1401 ( 
.A1(n_1162),
.A2(n_1123),
.B1(n_817),
.B2(n_1079),
.Y(n_1401)
);

A2O1A1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1193),
.A2(n_973),
.B(n_955),
.C(n_1191),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_SL g1403 ( 
.A1(n_1107),
.A2(n_932),
.B(n_925),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1246),
.B(n_963),
.Y(n_1404)
);

BUFx6f_ASAP7_75t_L g1405 ( 
.A(n_1154),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1151),
.B(n_1017),
.Y(n_1406)
);

O2A1O1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1185),
.A2(n_973),
.B(n_632),
.C(n_1196),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_1319),
.Y(n_1408)
);

CKINVDCx16_ASAP7_75t_R g1409 ( 
.A(n_1258),
.Y(n_1409)
);

BUFx12f_ASAP7_75t_L g1410 ( 
.A(n_1319),
.Y(n_1410)
);

BUFx6f_ASAP7_75t_L g1411 ( 
.A(n_1321),
.Y(n_1411)
);

BUFx2_ASAP7_75t_L g1412 ( 
.A(n_1344),
.Y(n_1412)
);

INVx1_ASAP7_75t_SL g1413 ( 
.A(n_1287),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1379),
.A2(n_1401),
.B1(n_1334),
.B2(n_1260),
.Y(n_1414)
);

BUFx12f_ASAP7_75t_L g1415 ( 
.A(n_1340),
.Y(n_1415)
);

INVx1_ASAP7_75t_SL g1416 ( 
.A(n_1305),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1260),
.A2(n_1276),
.B1(n_1288),
.B2(n_1354),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1272),
.Y(n_1418)
);

OAI22x1_ASAP7_75t_L g1419 ( 
.A1(n_1276),
.A2(n_1331),
.B1(n_1286),
.B2(n_1323),
.Y(n_1419)
);

BUFx12f_ASAP7_75t_L g1420 ( 
.A(n_1264),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1331),
.A2(n_1386),
.B1(n_1354),
.B2(n_1394),
.Y(n_1421)
);

INVx4_ASAP7_75t_L g1422 ( 
.A(n_1339),
.Y(n_1422)
);

CKINVDCx6p67_ASAP7_75t_R g1423 ( 
.A(n_1388),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1373),
.A2(n_1406),
.B1(n_1288),
.B2(n_1385),
.Y(n_1424)
);

CKINVDCx11_ASAP7_75t_R g1425 ( 
.A(n_1284),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1295),
.Y(n_1426)
);

CKINVDCx11_ASAP7_75t_R g1427 ( 
.A(n_1271),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1394),
.A2(n_1286),
.B1(n_1271),
.B2(n_1341),
.Y(n_1428)
);

CKINVDCx11_ASAP7_75t_R g1429 ( 
.A(n_1299),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1386),
.A2(n_1280),
.B1(n_1325),
.B2(n_1382),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1322),
.B(n_1310),
.Y(n_1431)
);

INVx4_ASAP7_75t_L g1432 ( 
.A(n_1282),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1266),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1306),
.Y(n_1434)
);

INVx4_ASAP7_75t_L g1435 ( 
.A(n_1282),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_SL g1436 ( 
.A1(n_1257),
.A2(n_1265),
.B1(n_1296),
.B2(n_1323),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1270),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1327),
.A2(n_1341),
.B1(n_1404),
.B2(n_1366),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1327),
.A2(n_1342),
.B1(n_1404),
.B2(n_1367),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1384),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_SL g1441 ( 
.A1(n_1257),
.A2(n_1296),
.B1(n_1304),
.B2(n_1367),
.Y(n_1441)
);

BUFx3_ASAP7_75t_L g1442 ( 
.A(n_1398),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1329),
.A2(n_1358),
.B1(n_1347),
.B2(n_1259),
.Y(n_1443)
);

NAND2x1p5_ASAP7_75t_L g1444 ( 
.A(n_1381),
.B(n_1312),
.Y(n_1444)
);

NAND2x1p5_ASAP7_75t_L g1445 ( 
.A(n_1293),
.B(n_1285),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_SL g1446 ( 
.A1(n_1304),
.A2(n_1370),
.B1(n_1268),
.B2(n_1261),
.Y(n_1446)
);

OAI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1345),
.A2(n_1355),
.B1(n_1349),
.B2(n_1368),
.Y(n_1447)
);

INVx8_ASAP7_75t_L g1448 ( 
.A(n_1337),
.Y(n_1448)
);

CKINVDCx11_ASAP7_75t_R g1449 ( 
.A(n_1389),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_1311),
.Y(n_1450)
);

BUFx4f_ASAP7_75t_L g1451 ( 
.A(n_1389),
.Y(n_1451)
);

CKINVDCx20_ASAP7_75t_R g1452 ( 
.A(n_1314),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1400),
.Y(n_1453)
);

BUFx4f_ASAP7_75t_SL g1454 ( 
.A(n_1400),
.Y(n_1454)
);

INVx6_ASAP7_75t_L g1455 ( 
.A(n_1313),
.Y(n_1455)
);

BUFx10_ASAP7_75t_L g1456 ( 
.A(n_1326),
.Y(n_1456)
);

OAI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1297),
.A2(n_1352),
.B1(n_1348),
.B2(n_1378),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1330),
.A2(n_1332),
.B1(n_1369),
.B2(n_1371),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1374),
.A2(n_1407),
.B1(n_1375),
.B2(n_1391),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1289),
.B(n_1387),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1338),
.B(n_1343),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1356),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_SL g1463 ( 
.A1(n_1268),
.A2(n_1261),
.B1(n_1328),
.B2(n_1275),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_SL g1464 ( 
.A1(n_1261),
.A2(n_1328),
.B1(n_1361),
.B2(n_1396),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_SL g1465 ( 
.A1(n_1316),
.A2(n_1297),
.B1(n_1274),
.B2(n_1281),
.Y(n_1465)
);

BUFx2_ASAP7_75t_L g1466 ( 
.A(n_1320),
.Y(n_1466)
);

BUFx12f_ASAP7_75t_L g1467 ( 
.A(n_1291),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1255),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1372),
.B(n_1395),
.Y(n_1469)
);

INVx2_ASAP7_75t_SL g1470 ( 
.A(n_1317),
.Y(n_1470)
);

INVx1_ASAP7_75t_SL g1471 ( 
.A(n_1316),
.Y(n_1471)
);

INVx6_ASAP7_75t_L g1472 ( 
.A(n_1309),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1301),
.A2(n_1300),
.B1(n_1298),
.B2(n_1269),
.Y(n_1473)
);

OAI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1298),
.A2(n_1290),
.B1(n_1357),
.B2(n_1359),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1402),
.B(n_1324),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1300),
.A2(n_1292),
.B1(n_1303),
.B2(n_1302),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1283),
.A2(n_1392),
.B1(n_1362),
.B2(n_1360),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1318),
.Y(n_1478)
);

CKINVDCx11_ASAP7_75t_R g1479 ( 
.A(n_1294),
.Y(n_1479)
);

INVx3_ASAP7_75t_SL g1480 ( 
.A(n_1362),
.Y(n_1480)
);

BUFx3_ASAP7_75t_L g1481 ( 
.A(n_1392),
.Y(n_1481)
);

INVx4_ASAP7_75t_L g1482 ( 
.A(n_1365),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1399),
.A2(n_1279),
.B1(n_1278),
.B2(n_1267),
.Y(n_1483)
);

OAI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1263),
.A2(n_1279),
.B1(n_1403),
.B2(n_1255),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1279),
.A2(n_1273),
.B1(n_1397),
.B2(n_1365),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1315),
.Y(n_1486)
);

BUFx10_ASAP7_75t_L g1487 ( 
.A(n_1346),
.Y(n_1487)
);

BUFx8_ASAP7_75t_SL g1488 ( 
.A(n_1383),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1397),
.A2(n_1263),
.B1(n_1262),
.B2(n_1256),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_SL g1490 ( 
.A1(n_1353),
.A2(n_1390),
.B1(n_1380),
.B2(n_1277),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1308),
.Y(n_1491)
);

OAI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1277),
.A2(n_1307),
.B1(n_1333),
.B2(n_1335),
.Y(n_1492)
);

OAI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1277),
.A2(n_1336),
.B1(n_1350),
.B2(n_1351),
.Y(n_1493)
);

INVx3_ASAP7_75t_SL g1494 ( 
.A(n_1363),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1364),
.Y(n_1495)
);

INVx6_ASAP7_75t_L g1496 ( 
.A(n_1376),
.Y(n_1496)
);

CKINVDCx11_ASAP7_75t_R g1497 ( 
.A(n_1377),
.Y(n_1497)
);

INVx1_ASAP7_75t_SL g1498 ( 
.A(n_1393),
.Y(n_1498)
);

INVx5_ASAP7_75t_L g1499 ( 
.A(n_1405),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1379),
.A2(n_973),
.B1(n_1401),
.B2(n_1334),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_SL g1501 ( 
.A1(n_1334),
.A2(n_1155),
.B1(n_1196),
.B2(n_1185),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1295),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1295),
.Y(n_1503)
);

OAI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1379),
.A2(n_1334),
.B1(n_963),
.B2(n_973),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1379),
.A2(n_973),
.B1(n_1401),
.B2(n_1334),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1379),
.A2(n_1334),
.B1(n_963),
.B2(n_973),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1319),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1344),
.Y(n_1508)
);

CKINVDCx11_ASAP7_75t_R g1509 ( 
.A(n_1321),
.Y(n_1509)
);

INVx6_ASAP7_75t_L g1510 ( 
.A(n_1405),
.Y(n_1510)
);

INVx5_ASAP7_75t_L g1511 ( 
.A(n_1405),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_SL g1512 ( 
.A1(n_1288),
.A2(n_1162),
.B1(n_429),
.B2(n_427),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1288),
.A2(n_1162),
.B1(n_429),
.B2(n_427),
.Y(n_1513)
);

INVx4_ASAP7_75t_L g1514 ( 
.A(n_1321),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_SL g1515 ( 
.A1(n_1288),
.A2(n_1162),
.B1(n_429),
.B2(n_427),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1379),
.A2(n_1334),
.B1(n_963),
.B2(n_973),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1295),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1284),
.Y(n_1518)
);

CKINVDCx11_ASAP7_75t_R g1519 ( 
.A(n_1321),
.Y(n_1519)
);

BUFx2_ASAP7_75t_L g1520 ( 
.A(n_1344),
.Y(n_1520)
);

INVxp67_ASAP7_75t_L g1521 ( 
.A(n_1384),
.Y(n_1521)
);

CKINVDCx11_ASAP7_75t_R g1522 ( 
.A(n_1321),
.Y(n_1522)
);

BUFx8_ASAP7_75t_SL g1523 ( 
.A(n_1258),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1295),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1379),
.A2(n_973),
.B1(n_1401),
.B2(n_1334),
.Y(n_1525)
);

CKINVDCx6p67_ASAP7_75t_R g1526 ( 
.A(n_1321),
.Y(n_1526)
);

OAI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1280),
.A2(n_973),
.B(n_1379),
.Y(n_1527)
);

BUFx12f_ASAP7_75t_L g1528 ( 
.A(n_1319),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1272),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1379),
.A2(n_973),
.B1(n_1079),
.B2(n_882),
.Y(n_1530)
);

OAI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1331),
.A2(n_1386),
.B1(n_1276),
.B2(n_1349),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1379),
.A2(n_973),
.B1(n_1401),
.B2(n_1334),
.Y(n_1532)
);

BUFx3_ASAP7_75t_L g1533 ( 
.A(n_1284),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1379),
.A2(n_973),
.B1(n_1401),
.B2(n_1334),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1295),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1379),
.A2(n_973),
.B1(n_1401),
.B2(n_1334),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1421),
.B(n_1412),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1488),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1466),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1468),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1468),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1508),
.B(n_1520),
.Y(n_1542)
);

AO21x1_ASAP7_75t_SL g1543 ( 
.A1(n_1417),
.A2(n_1475),
.B(n_1527),
.Y(n_1543)
);

AOI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1459),
.A2(n_1495),
.B(n_1419),
.Y(n_1544)
);

OAI21x1_ASAP7_75t_L g1545 ( 
.A1(n_1485),
.A2(n_1489),
.B(n_1483),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1418),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1456),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1418),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1529),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1529),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1433),
.Y(n_1551)
);

INVx1_ASAP7_75t_SL g1552 ( 
.A(n_1449),
.Y(n_1552)
);

INVx2_ASAP7_75t_SL g1553 ( 
.A(n_1456),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1494),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1437),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1512),
.A2(n_1515),
.B1(n_1513),
.B2(n_1530),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1429),
.B(n_1432),
.Y(n_1557)
);

BUFx2_ASAP7_75t_SL g1558 ( 
.A(n_1499),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1482),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1427),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_L g1561 ( 
.A(n_1472),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1521),
.Y(n_1562)
);

BUFx2_ASAP7_75t_L g1563 ( 
.A(n_1494),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1491),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1457),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1438),
.B(n_1439),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1457),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1518),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1426),
.Y(n_1569)
);

OA21x2_ASAP7_75t_L g1570 ( 
.A1(n_1476),
.A2(n_1473),
.B(n_1486),
.Y(n_1570)
);

HB1xp67_ASAP7_75t_L g1571 ( 
.A(n_1462),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1440),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1442),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1482),
.Y(n_1574)
);

NAND2x1p5_ASAP7_75t_L g1575 ( 
.A(n_1471),
.B(n_1478),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1469),
.B(n_1463),
.Y(n_1576)
);

INVx3_ASAP7_75t_L g1577 ( 
.A(n_1496),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1502),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1503),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1517),
.Y(n_1580)
);

INVxp67_ASAP7_75t_L g1581 ( 
.A(n_1434),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1444),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_SL g1583 ( 
.A1(n_1504),
.A2(n_1506),
.B1(n_1516),
.B2(n_1430),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1417),
.B(n_1413),
.Y(n_1584)
);

INVx5_ASAP7_75t_L g1585 ( 
.A(n_1472),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1463),
.B(n_1464),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1464),
.B(n_1446),
.Y(n_1587)
);

AOI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1470),
.A2(n_1460),
.B(n_1461),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1524),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1535),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1487),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1416),
.Y(n_1592)
);

AND3x1_ASAP7_75t_L g1593 ( 
.A(n_1414),
.B(n_1428),
.C(n_1500),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1487),
.Y(n_1594)
);

CKINVDCx6p67_ASAP7_75t_R g1595 ( 
.A(n_1410),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1490),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1490),
.Y(n_1597)
);

OAI21x1_ASAP7_75t_L g1598 ( 
.A1(n_1477),
.A2(n_1476),
.B(n_1473),
.Y(n_1598)
);

BUFx12f_ASAP7_75t_L g1599 ( 
.A(n_1509),
.Y(n_1599)
);

AOI21x1_ASAP7_75t_L g1600 ( 
.A1(n_1431),
.A2(n_1493),
.B(n_1497),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1484),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1492),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1450),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1492),
.Y(n_1604)
);

OAI21x1_ASAP7_75t_L g1605 ( 
.A1(n_1445),
.A2(n_1536),
.B(n_1534),
.Y(n_1605)
);

INVx11_ASAP7_75t_L g1606 ( 
.A(n_1415),
.Y(n_1606)
);

AO21x2_ASAP7_75t_L g1607 ( 
.A1(n_1531),
.A2(n_1493),
.B(n_1474),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1498),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1446),
.B(n_1441),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1465),
.Y(n_1610)
);

O2A1O1Ixp5_ASAP7_75t_L g1611 ( 
.A1(n_1531),
.A2(n_1447),
.B(n_1474),
.C(n_1451),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1479),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1455),
.Y(n_1613)
);

BUFx3_ASAP7_75t_L g1614 ( 
.A(n_1455),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1465),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1455),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1447),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1441),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1436),
.B(n_1467),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1424),
.B(n_1436),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1500),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1505),
.Y(n_1622)
);

NAND2x1p5_ASAP7_75t_L g1623 ( 
.A(n_1499),
.B(n_1511),
.Y(n_1623)
);

CKINVDCx6p67_ASAP7_75t_R g1624 ( 
.A(n_1528),
.Y(n_1624)
);

INVx3_ASAP7_75t_L g1625 ( 
.A(n_1481),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1525),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_1408),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1532),
.Y(n_1628)
);

INVx2_ASAP7_75t_SL g1629 ( 
.A(n_1448),
.Y(n_1629)
);

BUFx3_ASAP7_75t_L g1630 ( 
.A(n_1448),
.Y(n_1630)
);

NAND2x1p5_ASAP7_75t_L g1631 ( 
.A(n_1511),
.B(n_1451),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1443),
.B(n_1432),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1571),
.B(n_1411),
.Y(n_1633)
);

OAI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1583),
.A2(n_1515),
.B(n_1513),
.Y(n_1634)
);

A2O1A1Ixp33_ASAP7_75t_L g1635 ( 
.A1(n_1611),
.A2(n_1512),
.B(n_1448),
.C(n_1501),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1603),
.B(n_1411),
.Y(n_1636)
);

OAI21xp5_ASAP7_75t_L g1637 ( 
.A1(n_1593),
.A2(n_1435),
.B(n_1453),
.Y(n_1637)
);

OA21x2_ASAP7_75t_L g1638 ( 
.A1(n_1598),
.A2(n_1458),
.B(n_1480),
.Y(n_1638)
);

INVxp67_ASAP7_75t_L g1639 ( 
.A(n_1539),
.Y(n_1639)
);

O2A1O1Ixp33_ASAP7_75t_L g1640 ( 
.A1(n_1609),
.A2(n_1480),
.B(n_1533),
.C(n_1452),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1551),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1573),
.B(n_1514),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1618),
.A2(n_1454),
.B1(n_1526),
.B2(n_1409),
.Y(n_1643)
);

AOI221xp5_ASAP7_75t_SL g1644 ( 
.A1(n_1576),
.A2(n_1522),
.B1(n_1519),
.B2(n_1423),
.C(n_1425),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1572),
.B(n_1422),
.Y(n_1645)
);

A2O1A1Ixp33_ASAP7_75t_L g1646 ( 
.A1(n_1620),
.A2(n_1587),
.B(n_1610),
.C(n_1615),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1537),
.B(n_1510),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1562),
.B(n_1510),
.Y(n_1648)
);

O2A1O1Ixp33_ASAP7_75t_SL g1649 ( 
.A1(n_1619),
.A2(n_1523),
.B(n_1507),
.C(n_1420),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1555),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1555),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_1606),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1542),
.B(n_1537),
.Y(n_1653)
);

AOI221xp5_ASAP7_75t_L g1654 ( 
.A1(n_1617),
.A2(n_1587),
.B1(n_1586),
.B2(n_1621),
.C(n_1622),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1542),
.B(n_1592),
.Y(n_1655)
);

A2O1A1Ixp33_ASAP7_75t_L g1656 ( 
.A1(n_1615),
.A2(n_1605),
.B(n_1586),
.C(n_1566),
.Y(n_1656)
);

OR2x6_ASAP7_75t_L g1657 ( 
.A(n_1600),
.B(n_1613),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1612),
.B(n_1581),
.Y(n_1658)
);

AOI21x1_ASAP7_75t_L g1659 ( 
.A1(n_1617),
.A2(n_1544),
.B(n_1588),
.Y(n_1659)
);

A2O1A1Ixp33_ASAP7_75t_L g1660 ( 
.A1(n_1605),
.A2(n_1622),
.B(n_1621),
.C(n_1626),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1538),
.B(n_1625),
.Y(n_1661)
);

AOI221xp5_ASAP7_75t_L g1662 ( 
.A1(n_1626),
.A2(n_1628),
.B1(n_1556),
.B2(n_1565),
.C(n_1567),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1569),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1538),
.B(n_1625),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1538),
.B(n_1625),
.Y(n_1665)
);

NOR3xp33_ASAP7_75t_SL g1666 ( 
.A(n_1627),
.B(n_1557),
.C(n_1599),
.Y(n_1666)
);

AO32x2_ASAP7_75t_L g1667 ( 
.A1(n_1547),
.A2(n_1553),
.A3(n_1629),
.B1(n_1596),
.B2(n_1597),
.Y(n_1667)
);

INVx1_ASAP7_75t_SL g1668 ( 
.A(n_1568),
.Y(n_1668)
);

A2O1A1Ixp33_ASAP7_75t_L g1669 ( 
.A1(n_1628),
.A2(n_1565),
.B(n_1567),
.C(n_1598),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1607),
.A2(n_1616),
.B1(n_1613),
.B2(n_1597),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1606),
.Y(n_1671)
);

O2A1O1Ixp33_ASAP7_75t_SL g1672 ( 
.A1(n_1560),
.A2(n_1553),
.B(n_1552),
.C(n_1629),
.Y(n_1672)
);

A2O1A1Ixp33_ASAP7_75t_L g1673 ( 
.A1(n_1584),
.A2(n_1601),
.B(n_1543),
.C(n_1596),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1578),
.B(n_1579),
.Y(n_1674)
);

AND2x4_ASAP7_75t_L g1675 ( 
.A(n_1582),
.B(n_1614),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_1595),
.Y(n_1676)
);

A2O1A1Ixp33_ASAP7_75t_L g1677 ( 
.A1(n_1601),
.A2(n_1543),
.B(n_1614),
.C(n_1602),
.Y(n_1677)
);

OAI21x1_ASAP7_75t_L g1678 ( 
.A1(n_1545),
.A2(n_1575),
.B(n_1623),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_1595),
.Y(n_1679)
);

O2A1O1Ixp33_ASAP7_75t_L g1680 ( 
.A1(n_1607),
.A2(n_1602),
.B(n_1604),
.C(n_1632),
.Y(n_1680)
);

OA21x2_ASAP7_75t_L g1681 ( 
.A1(n_1604),
.A2(n_1549),
.B(n_1546),
.Y(n_1681)
);

OR2x6_ASAP7_75t_L g1682 ( 
.A(n_1575),
.B(n_1558),
.Y(n_1682)
);

O2A1O1Ixp5_ASAP7_75t_L g1683 ( 
.A1(n_1540),
.A2(n_1541),
.B(n_1591),
.C(n_1594),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1548),
.Y(n_1684)
);

A2O1A1Ixp33_ASAP7_75t_L g1685 ( 
.A1(n_1585),
.A2(n_1561),
.B(n_1540),
.C(n_1541),
.Y(n_1685)
);

AOI21x1_ASAP7_75t_L g1686 ( 
.A1(n_1554),
.A2(n_1563),
.B(n_1591),
.Y(n_1686)
);

AO32x2_ASAP7_75t_L g1687 ( 
.A1(n_1570),
.A2(n_1578),
.A3(n_1590),
.B1(n_1579),
.B2(n_1580),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1653),
.B(n_1559),
.Y(n_1688)
);

BUFx3_ASAP7_75t_L g1689 ( 
.A(n_1678),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1687),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1687),
.Y(n_1691)
);

BUFx12f_ASAP7_75t_L g1692 ( 
.A(n_1676),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1681),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1687),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1667),
.B(n_1559),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1667),
.B(n_1574),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1667),
.B(n_1574),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1687),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1667),
.B(n_1574),
.Y(n_1699)
);

BUFx2_ASAP7_75t_L g1700 ( 
.A(n_1639),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1684),
.B(n_1549),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1641),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1655),
.B(n_1570),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1634),
.A2(n_1654),
.B1(n_1662),
.B2(n_1670),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1681),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1650),
.B(n_1651),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1681),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1663),
.Y(n_1708)
);

HB1xp67_ASAP7_75t_L g1709 ( 
.A(n_1686),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1674),
.Y(n_1710)
);

INVx4_ASAP7_75t_L g1711 ( 
.A(n_1682),
.Y(n_1711)
);

OAI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1646),
.A2(n_1630),
.B1(n_1589),
.B2(n_1631),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1669),
.B(n_1550),
.Y(n_1713)
);

AND2x4_ASAP7_75t_L g1714 ( 
.A(n_1685),
.B(n_1577),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1683),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1683),
.Y(n_1716)
);

INVxp67_ASAP7_75t_SL g1717 ( 
.A(n_1680),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1659),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1693),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1695),
.B(n_1638),
.Y(n_1720)
);

CKINVDCx20_ASAP7_75t_R g1721 ( 
.A(n_1692),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1689),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1695),
.B(n_1638),
.Y(n_1723)
);

OR2x6_ASAP7_75t_L g1724 ( 
.A(n_1714),
.B(n_1657),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1710),
.B(n_1680),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1696),
.B(n_1661),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1690),
.B(n_1648),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1696),
.B(n_1664),
.Y(n_1728)
);

AND2x2_ASAP7_75t_SL g1729 ( 
.A(n_1714),
.B(n_1675),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1690),
.B(n_1656),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1696),
.B(n_1697),
.Y(n_1731)
);

INVxp67_ASAP7_75t_L g1732 ( 
.A(n_1715),
.Y(n_1732)
);

INVx3_ASAP7_75t_L g1733 ( 
.A(n_1689),
.Y(n_1733)
);

INVx4_ASAP7_75t_L g1734 ( 
.A(n_1692),
.Y(n_1734)
);

AOI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1704),
.A2(n_1635),
.B1(n_1646),
.B2(n_1673),
.Y(n_1735)
);

INVx1_ASAP7_75t_SL g1736 ( 
.A(n_1700),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1708),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1708),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1690),
.B(n_1656),
.Y(n_1739)
);

NOR3xp33_ASAP7_75t_L g1740 ( 
.A(n_1717),
.B(n_1635),
.C(n_1715),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1696),
.B(n_1665),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1701),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1697),
.B(n_1685),
.Y(n_1743)
);

INVx3_ASAP7_75t_L g1744 ( 
.A(n_1689),
.Y(n_1744)
);

INVx1_ASAP7_75t_SL g1745 ( 
.A(n_1700),
.Y(n_1745)
);

OAI221xp5_ASAP7_75t_L g1746 ( 
.A1(n_1704),
.A2(n_1673),
.B1(n_1677),
.B2(n_1640),
.C(n_1660),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1710),
.B(n_1647),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1693),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1691),
.Y(n_1749)
);

INVx1_ASAP7_75t_SL g1750 ( 
.A(n_1700),
.Y(n_1750)
);

BUFx3_ASAP7_75t_L g1751 ( 
.A(n_1714),
.Y(n_1751)
);

INVx4_ASAP7_75t_L g1752 ( 
.A(n_1692),
.Y(n_1752)
);

AO21x2_ASAP7_75t_L g1753 ( 
.A1(n_1717),
.A2(n_1660),
.B(n_1608),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1715),
.B(n_1716),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_1692),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1716),
.B(n_1608),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1702),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1699),
.B(n_1658),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1716),
.B(n_1564),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1757),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1757),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1748),
.Y(n_1762)
);

BUFx2_ASAP7_75t_SL g1763 ( 
.A(n_1721),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1732),
.B(n_1694),
.Y(n_1764)
);

AOI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1735),
.A2(n_1740),
.B1(n_1746),
.B2(n_1712),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1731),
.B(n_1699),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1737),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1754),
.B(n_1694),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1731),
.B(n_1699),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1731),
.B(n_1703),
.Y(n_1770)
);

AOI21xp33_ASAP7_75t_L g1771 ( 
.A1(n_1732),
.A2(n_1709),
.B(n_1713),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1743),
.B(n_1703),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1749),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1749),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1754),
.B(n_1694),
.Y(n_1775)
);

AO21x2_ASAP7_75t_L g1776 ( 
.A1(n_1740),
.A2(n_1718),
.B(n_1705),
.Y(n_1776)
);

INVxp67_ASAP7_75t_SL g1777 ( 
.A(n_1756),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1743),
.B(n_1703),
.Y(n_1778)
);

AND2x4_ASAP7_75t_L g1779 ( 
.A(n_1751),
.B(n_1689),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1759),
.B(n_1756),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1743),
.B(n_1703),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1727),
.B(n_1698),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1729),
.B(n_1714),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1759),
.B(n_1698),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1726),
.B(n_1688),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1725),
.B(n_1706),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1742),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1748),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1737),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1738),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1738),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1748),
.Y(n_1792)
);

NAND2x1p5_ASAP7_75t_L g1793 ( 
.A(n_1729),
.B(n_1711),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1748),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1719),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1726),
.B(n_1688),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1728),
.B(n_1741),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1719),
.Y(n_1798)
);

BUFx3_ASAP7_75t_L g1799 ( 
.A(n_1721),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1719),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1742),
.Y(n_1801)
);

HB1xp67_ASAP7_75t_L g1802 ( 
.A(n_1727),
.Y(n_1802)
);

NAND2x1_ASAP7_75t_L g1803 ( 
.A(n_1779),
.B(n_1722),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1760),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1797),
.B(n_1758),
.Y(n_1805)
);

OR2x2_ASAP7_75t_L g1806 ( 
.A(n_1786),
.B(n_1730),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1776),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1776),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1776),
.Y(n_1809)
);

OAI22xp33_ASAP7_75t_SL g1810 ( 
.A1(n_1765),
.A2(n_1730),
.B1(n_1739),
.B2(n_1735),
.Y(n_1810)
);

AND2x2_ASAP7_75t_SL g1811 ( 
.A(n_1765),
.B(n_1729),
.Y(n_1811)
);

NAND3xp33_ASAP7_75t_L g1812 ( 
.A(n_1771),
.B(n_1746),
.C(n_1725),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1760),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1761),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1797),
.B(n_1758),
.Y(n_1815)
);

AND2x4_ASAP7_75t_L g1816 ( 
.A(n_1783),
.B(n_1751),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1797),
.B(n_1758),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1761),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1776),
.Y(n_1819)
);

AND2x4_ASAP7_75t_L g1820 ( 
.A(n_1783),
.B(n_1751),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1767),
.Y(n_1821)
);

INVx1_ASAP7_75t_SL g1822 ( 
.A(n_1763),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1776),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1767),
.Y(n_1824)
);

INVxp33_ASAP7_75t_L g1825 ( 
.A(n_1799),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1789),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1789),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1790),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1786),
.B(n_1730),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1780),
.B(n_1739),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1777),
.B(n_1747),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1790),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1791),
.Y(n_1833)
);

INVx2_ASAP7_75t_SL g1834 ( 
.A(n_1799),
.Y(n_1834)
);

INVxp67_ASAP7_75t_SL g1835 ( 
.A(n_1799),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1791),
.Y(n_1836)
);

NAND2x1p5_ASAP7_75t_L g1837 ( 
.A(n_1799),
.B(n_1734),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1777),
.B(n_1747),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1773),
.Y(n_1839)
);

OAI211xp5_ASAP7_75t_L g1840 ( 
.A1(n_1771),
.A2(n_1709),
.B(n_1722),
.C(n_1733),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_SL g1841 ( 
.A(n_1793),
.B(n_1729),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1785),
.B(n_1796),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1773),
.Y(n_1843)
);

INVx2_ASAP7_75t_SL g1844 ( 
.A(n_1793),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1780),
.B(n_1736),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1774),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1772),
.B(n_1736),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1763),
.B(n_1734),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1818),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1835),
.B(n_1772),
.Y(n_1850)
);

BUFx3_ASAP7_75t_L g1851 ( 
.A(n_1834),
.Y(n_1851)
);

AOI211x1_ASAP7_75t_L g1852 ( 
.A1(n_1812),
.A2(n_1772),
.B(n_1781),
.C(n_1778),
.Y(n_1852)
);

NAND4xp25_ASAP7_75t_L g1853 ( 
.A(n_1822),
.B(n_1644),
.C(n_1734),
.D(n_1752),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1830),
.B(n_1778),
.Y(n_1854)
);

NAND3xp33_ASAP7_75t_L g1855 ( 
.A(n_1840),
.B(n_1774),
.C(n_1764),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1818),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1830),
.B(n_1778),
.Y(n_1857)
);

OR2x6_ASAP7_75t_L g1858 ( 
.A(n_1837),
.B(n_1834),
.Y(n_1858)
);

INVx2_ASAP7_75t_SL g1859 ( 
.A(n_1837),
.Y(n_1859)
);

NOR2xp33_ASAP7_75t_L g1860 ( 
.A(n_1825),
.B(n_1763),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1826),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1810),
.B(n_1781),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1806),
.B(n_1781),
.Y(n_1863)
);

NAND4xp25_ASAP7_75t_L g1864 ( 
.A(n_1848),
.B(n_1752),
.C(n_1734),
.D(n_1774),
.Y(n_1864)
);

NOR2xp67_ASAP7_75t_L g1865 ( 
.A(n_1841),
.B(n_1751),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1825),
.B(n_1734),
.Y(n_1866)
);

INVx1_ASAP7_75t_SL g1867 ( 
.A(n_1811),
.Y(n_1867)
);

INVx5_ASAP7_75t_L g1868 ( 
.A(n_1807),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1816),
.B(n_1770),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1806),
.B(n_1802),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1837),
.B(n_1811),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1807),
.Y(n_1872)
);

AOI22xp33_ASAP7_75t_L g1873 ( 
.A1(n_1808),
.A2(n_1753),
.B1(n_1739),
.B2(n_1720),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1829),
.B(n_1802),
.Y(n_1874)
);

INVxp67_ASAP7_75t_SL g1875 ( 
.A(n_1808),
.Y(n_1875)
);

OAI21xp33_ASAP7_75t_L g1876 ( 
.A1(n_1831),
.A2(n_1764),
.B(n_1779),
.Y(n_1876)
);

HB1xp67_ASAP7_75t_L g1877 ( 
.A(n_1839),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1829),
.B(n_1785),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_L g1879 ( 
.A(n_1816),
.B(n_1752),
.Y(n_1879)
);

NOR3xp33_ASAP7_75t_L g1880 ( 
.A(n_1809),
.B(n_1733),
.C(n_1722),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_L g1881 ( 
.A(n_1816),
.B(n_1752),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1843),
.B(n_1796),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1838),
.B(n_1796),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1820),
.B(n_1752),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1826),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1854),
.B(n_1845),
.Y(n_1886)
);

OAI221xp5_ASAP7_75t_L g1887 ( 
.A1(n_1873),
.A2(n_1809),
.B1(n_1819),
.B2(n_1823),
.C(n_1744),
.Y(n_1887)
);

HB1xp67_ASAP7_75t_L g1888 ( 
.A(n_1851),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1871),
.B(n_1842),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1868),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1849),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1860),
.B(n_1755),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1856),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1861),
.Y(n_1894)
);

INVx2_ASAP7_75t_SL g1895 ( 
.A(n_1858),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1858),
.B(n_1842),
.Y(n_1896)
);

NOR2xp33_ASAP7_75t_L g1897 ( 
.A(n_1860),
.B(n_1624),
.Y(n_1897)
);

INVxp67_ASAP7_75t_L g1898 ( 
.A(n_1851),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1885),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1877),
.Y(n_1900)
);

AOI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1867),
.A2(n_1753),
.B1(n_1723),
.B2(n_1720),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1870),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1874),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1858),
.B(n_1805),
.Y(n_1904)
);

OAI22xp33_ASAP7_75t_L g1905 ( 
.A1(n_1862),
.A2(n_1724),
.B1(n_1865),
.B2(n_1863),
.Y(n_1905)
);

INVx1_ASAP7_75t_SL g1906 ( 
.A(n_1866),
.Y(n_1906)
);

AOI22xp33_ASAP7_75t_L g1907 ( 
.A1(n_1873),
.A2(n_1753),
.B1(n_1823),
.B2(n_1819),
.Y(n_1907)
);

AOI221x1_ASAP7_75t_L g1908 ( 
.A1(n_1864),
.A2(n_1846),
.B1(n_1828),
.B2(n_1821),
.C(n_1836),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1868),
.Y(n_1909)
);

INVxp67_ASAP7_75t_SL g1910 ( 
.A(n_1859),
.Y(n_1910)
);

AOI22xp5_ASAP7_75t_L g1911 ( 
.A1(n_1857),
.A2(n_1753),
.B1(n_1720),
.B2(n_1723),
.Y(n_1911)
);

OAI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1855),
.A2(n_1841),
.B(n_1820),
.Y(n_1912)
);

OAI211xp5_ASAP7_75t_L g1913 ( 
.A1(n_1908),
.A2(n_1852),
.B(n_1876),
.C(n_1853),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1888),
.B(n_1850),
.Y(n_1914)
);

INVx1_ASAP7_75t_SL g1915 ( 
.A(n_1906),
.Y(n_1915)
);

OAI22xp33_ASAP7_75t_L g1916 ( 
.A1(n_1911),
.A2(n_1782),
.B1(n_1724),
.B2(n_1793),
.Y(n_1916)
);

OAI21xp33_ASAP7_75t_L g1917 ( 
.A1(n_1912),
.A2(n_1881),
.B(n_1879),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1896),
.Y(n_1918)
);

NAND3xp33_ASAP7_75t_SL g1919 ( 
.A(n_1901),
.B(n_1881),
.C(n_1879),
.Y(n_1919)
);

OAI221xp5_ASAP7_75t_L g1920 ( 
.A1(n_1907),
.A2(n_1858),
.B1(n_1844),
.B2(n_1859),
.C(n_1733),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1889),
.B(n_1884),
.Y(n_1921)
);

AOI22xp5_ASAP7_75t_L g1922 ( 
.A1(n_1905),
.A2(n_1753),
.B1(n_1723),
.B2(n_1779),
.Y(n_1922)
);

OR2x2_ASAP7_75t_L g1923 ( 
.A(n_1886),
.B(n_1878),
.Y(n_1923)
);

AOI222xp33_ASAP7_75t_L g1924 ( 
.A1(n_1887),
.A2(n_1875),
.B1(n_1872),
.B2(n_1868),
.C1(n_1705),
.C2(n_1707),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1898),
.B(n_1883),
.Y(n_1925)
);

A2O1A1Ixp33_ASAP7_75t_L g1926 ( 
.A1(n_1895),
.A2(n_1722),
.B(n_1744),
.C(n_1733),
.Y(n_1926)
);

AOI21xp33_ASAP7_75t_L g1927 ( 
.A1(n_1890),
.A2(n_1872),
.B(n_1846),
.Y(n_1927)
);

OAI21xp33_ASAP7_75t_L g1928 ( 
.A1(n_1889),
.A2(n_1882),
.B(n_1869),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1891),
.Y(n_1929)
);

OAI22xp5_ASAP7_75t_L g1930 ( 
.A1(n_1896),
.A2(n_1820),
.B1(n_1793),
.B2(n_1869),
.Y(n_1930)
);

OAI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1908),
.A2(n_1895),
.B(n_1904),
.Y(n_1931)
);

AOI221xp5_ASAP7_75t_L g1932 ( 
.A1(n_1902),
.A2(n_1880),
.B1(n_1868),
.B2(n_1722),
.C(n_1733),
.Y(n_1932)
);

AOI221xp5_ASAP7_75t_L g1933 ( 
.A1(n_1903),
.A2(n_1868),
.B1(n_1744),
.B2(n_1784),
.C(n_1794),
.Y(n_1933)
);

OAI322xp33_ASAP7_75t_L g1934 ( 
.A1(n_1915),
.A2(n_1900),
.A3(n_1891),
.B1(n_1899),
.B2(n_1893),
.C1(n_1894),
.C2(n_1910),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1915),
.B(n_1893),
.Y(n_1935)
);

AOI22xp5_ASAP7_75t_L g1936 ( 
.A1(n_1913),
.A2(n_1904),
.B1(n_1897),
.B2(n_1890),
.Y(n_1936)
);

NOR2xp33_ASAP7_75t_L g1937 ( 
.A(n_1921),
.B(n_1892),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1929),
.Y(n_1938)
);

AOI32xp33_ASAP7_75t_L g1939 ( 
.A1(n_1916),
.A2(n_1920),
.A3(n_1933),
.B1(n_1918),
.B2(n_1909),
.Y(n_1939)
);

BUFx2_ASAP7_75t_L g1940 ( 
.A(n_1931),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1923),
.Y(n_1941)
);

OAI21xp33_ASAP7_75t_SL g1942 ( 
.A1(n_1927),
.A2(n_1909),
.B(n_1899),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1928),
.B(n_1886),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1914),
.B(n_1894),
.Y(n_1944)
);

NOR2xp33_ASAP7_75t_L g1945 ( 
.A(n_1917),
.B(n_1925),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1930),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1935),
.Y(n_1947)
);

NOR2x1_ASAP7_75t_L g1948 ( 
.A(n_1940),
.B(n_1919),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1941),
.B(n_1924),
.Y(n_1949)
);

OAI221xp5_ASAP7_75t_L g1950 ( 
.A1(n_1942),
.A2(n_1922),
.B1(n_1932),
.B2(n_1926),
.C(n_1844),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1945),
.B(n_1935),
.Y(n_1951)
);

AOI211xp5_ASAP7_75t_SL g1952 ( 
.A1(n_1934),
.A2(n_1649),
.B(n_1672),
.C(n_1847),
.Y(n_1952)
);

AOI211xp5_ASAP7_75t_L g1953 ( 
.A1(n_1946),
.A2(n_1649),
.B(n_1672),
.C(n_1643),
.Y(n_1953)
);

O2A1O1Ixp5_ASAP7_75t_L g1954 ( 
.A1(n_1937),
.A2(n_1803),
.B(n_1779),
.C(n_1832),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1944),
.B(n_1805),
.Y(n_1955)
);

AOI221xp5_ASAP7_75t_L g1956 ( 
.A1(n_1939),
.A2(n_1744),
.B1(n_1833),
.B2(n_1827),
.C(n_1824),
.Y(n_1956)
);

OAI221xp5_ASAP7_75t_L g1957 ( 
.A1(n_1936),
.A2(n_1744),
.B1(n_1803),
.B2(n_1782),
.C(n_1775),
.Y(n_1957)
);

NAND3xp33_ASAP7_75t_L g1958 ( 
.A(n_1938),
.B(n_1813),
.C(n_1804),
.Y(n_1958)
);

A2O1A1Ixp33_ASAP7_75t_L g1959 ( 
.A1(n_1948),
.A2(n_1943),
.B(n_1779),
.C(n_1666),
.Y(n_1959)
);

AOI31xp33_ASAP7_75t_L g1960 ( 
.A1(n_1951),
.A2(n_1679),
.A3(n_1652),
.B(n_1671),
.Y(n_1960)
);

OAI21xp5_ASAP7_75t_L g1961 ( 
.A1(n_1956),
.A2(n_1779),
.B(n_1815),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1954),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1947),
.B(n_1815),
.Y(n_1963)
);

O2A1O1Ixp33_ASAP7_75t_L g1964 ( 
.A1(n_1949),
.A2(n_1768),
.B(n_1775),
.C(n_1782),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_SL g1965 ( 
.A(n_1953),
.B(n_1666),
.Y(n_1965)
);

OAI21xp33_ASAP7_75t_L g1966 ( 
.A1(n_1955),
.A2(n_1814),
.B(n_1642),
.Y(n_1966)
);

AOI21xp5_ASAP7_75t_L g1967 ( 
.A1(n_1960),
.A2(n_1952),
.B(n_1950),
.Y(n_1967)
);

AOI21xp5_ASAP7_75t_L g1968 ( 
.A1(n_1959),
.A2(n_1958),
.B(n_1957),
.Y(n_1968)
);

AOI221xp5_ASAP7_75t_L g1969 ( 
.A1(n_1964),
.A2(n_1784),
.B1(n_1792),
.B2(n_1762),
.C(n_1794),
.Y(n_1969)
);

OAI211xp5_ASAP7_75t_L g1970 ( 
.A1(n_1962),
.A2(n_1624),
.B(n_1745),
.C(n_1750),
.Y(n_1970)
);

AOI221xp5_ASAP7_75t_L g1971 ( 
.A1(n_1963),
.A2(n_1794),
.B1(n_1762),
.B2(n_1788),
.C(n_1792),
.Y(n_1971)
);

XOR2x2_ASAP7_75t_L g1972 ( 
.A(n_1965),
.B(n_1668),
.Y(n_1972)
);

AOI21xp33_ASAP7_75t_L g1973 ( 
.A1(n_1961),
.A2(n_1788),
.B(n_1762),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1967),
.B(n_1966),
.Y(n_1974)
);

NOR2xp67_ASAP7_75t_L g1975 ( 
.A(n_1970),
.B(n_1768),
.Y(n_1975)
);

NOR2x1_ASAP7_75t_L g1976 ( 
.A(n_1968),
.B(n_1972),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1973),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1971),
.Y(n_1978)
);

OR2x2_ASAP7_75t_L g1979 ( 
.A(n_1969),
.B(n_1768),
.Y(n_1979)
);

NOR2x1_ASAP7_75t_L g1980 ( 
.A(n_1976),
.B(n_1775),
.Y(n_1980)
);

NAND2x1p5_ASAP7_75t_L g1981 ( 
.A(n_1974),
.B(n_1633),
.Y(n_1981)
);

AOI222xp33_ASAP7_75t_L g1982 ( 
.A1(n_1978),
.A2(n_1792),
.B1(n_1788),
.B2(n_1762),
.C1(n_1794),
.C2(n_1795),
.Y(n_1982)
);

OAI22xp5_ASAP7_75t_L g1983 ( 
.A1(n_1981),
.A2(n_1975),
.B1(n_1979),
.B2(n_1977),
.Y(n_1983)
);

CKINVDCx20_ASAP7_75t_R g1984 ( 
.A(n_1983),
.Y(n_1984)
);

OAI22xp33_ASAP7_75t_L g1985 ( 
.A1(n_1984),
.A2(n_1980),
.B1(n_1982),
.B2(n_1788),
.Y(n_1985)
);

OAI22xp5_ASAP7_75t_L g1986 ( 
.A1(n_1984),
.A2(n_1769),
.B1(n_1766),
.B2(n_1770),
.Y(n_1986)
);

OAI22xp5_ASAP7_75t_SL g1987 ( 
.A1(n_1985),
.A2(n_1986),
.B1(n_1787),
.B2(n_1801),
.Y(n_1987)
);

OAI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1985),
.A2(n_1817),
.B1(n_1769),
.B2(n_1766),
.Y(n_1988)
);

INVxp67_ASAP7_75t_L g1989 ( 
.A(n_1987),
.Y(n_1989)
);

AOI221xp5_ASAP7_75t_L g1990 ( 
.A1(n_1988),
.A2(n_1792),
.B1(n_1795),
.B2(n_1798),
.C(n_1800),
.Y(n_1990)
);

CKINVDCx20_ASAP7_75t_R g1991 ( 
.A(n_1989),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1990),
.B(n_1795),
.Y(n_1992)
);

AOI22xp33_ASAP7_75t_L g1993 ( 
.A1(n_1991),
.A2(n_1795),
.B1(n_1798),
.B2(n_1800),
.Y(n_1993)
);

XOR2xp5_ASAP7_75t_L g1994 ( 
.A(n_1993),
.B(n_1992),
.Y(n_1994)
);

AOI221xp5_ASAP7_75t_L g1995 ( 
.A1(n_1994),
.A2(n_1798),
.B1(n_1800),
.B2(n_1787),
.C(n_1636),
.Y(n_1995)
);

AOI211xp5_ASAP7_75t_L g1996 ( 
.A1(n_1995),
.A2(n_1640),
.B(n_1645),
.C(n_1637),
.Y(n_1996)
);


endmodule