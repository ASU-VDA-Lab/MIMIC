module real_jpeg_22869_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_2),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_2),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_2),
.B(n_36),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_2),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_2),
.B(n_61),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_2),
.B(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

INVx8_ASAP7_75t_SL g132 ( 
.A(n_4),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_5),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_5),
.B(n_61),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_5),
.B(n_43),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_5),
.B(n_36),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_5),
.B(n_40),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_5),
.B(n_50),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_5),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_5),
.B(n_166),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_6),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_6),
.B(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_6),
.B(n_43),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_6),
.B(n_61),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_6),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_6),
.B(n_50),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_6),
.B(n_131),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_6),
.B(n_166),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_8),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_8),
.B(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_8),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_8),
.B(n_36),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_8),
.B(n_40),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_8),
.B(n_50),
.Y(n_192)
);

INVxp33_ASAP7_75t_L g221 ( 
.A(n_8),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_8),
.B(n_166),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_9),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_9),
.B(n_61),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_9),
.B(n_43),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_9),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_9),
.B(n_50),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_9),
.B(n_131),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_9),
.B(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_10),
.B(n_17),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_10),
.B(n_61),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_10),
.B(n_43),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_10),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_10),
.B(n_40),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_10),
.B(n_50),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_10),
.B(n_346),
.Y(n_345)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_11),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_12),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_12),
.B(n_61),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_12),
.B(n_43),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_12),
.B(n_36),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_12),
.B(n_40),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_12),
.B(n_50),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_12),
.B(n_131),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_12),
.B(n_346),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_13),
.B(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_13),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_13),
.B(n_43),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_13),
.B(n_36),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_13),
.B(n_40),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_13),
.B(n_50),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_13),
.B(n_131),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_13),
.B(n_346),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_15),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_15),
.B(n_43),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_15),
.B(n_40),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_15),
.B(n_50),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_15),
.B(n_346),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_16),
.B(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_16),
.B(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_16),
.B(n_17),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_16),
.B(n_40),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_16),
.B(n_50),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_16),
.B(n_131),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_16),
.B(n_166),
.Y(n_226)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_17),
.Y(n_107)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_17),
.Y(n_207)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

O2A1O1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_381),
.B(n_382),
.C(n_386),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_372),
.C(n_380),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_357),
.C(n_358),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_332),
.C(n_333),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_301),
.C(n_302),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_276),
.C(n_277),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_245),
.C(n_246),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_210),
.C(n_211),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_173),
.C(n_174),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_139),
.C(n_140),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_112),
.C(n_113),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_72),
.C(n_84),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_53),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_45),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_33),
.B(n_45),
.C(n_53),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_38),
.C(n_41),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_34),
.A2(n_35),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_36),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_38),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_75)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_40),
.Y(n_219)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_46),
.B(n_48),
.C(n_49),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_63),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_54),
.B(n_64),
.C(n_65),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_59),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_83)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_58),
.Y(n_160)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_61),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_65)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_67),
.B(n_71),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_70),
.B(n_231),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.C(n_83),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_76),
.A2(n_77),
.B1(n_83),
.B2(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_88)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_108),
.C(n_109),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_93),
.C(n_98),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_91),
.C(n_92),
.Y(n_108)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.C(n_103),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_101),
.B(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_126),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_127),
.C(n_138),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_122),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_121),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_121),
.C(n_122),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_117),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_120),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx24_ASAP7_75t_SL g392 ( 
.A(n_122),
.Y(n_392)
);

FAx1_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_124),
.CI(n_125),
.CON(n_122),
.SN(n_122)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_124),
.C(n_125),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_138),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_136),
.B2(n_137),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_130),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_131),
.Y(n_222)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_135),
.C(n_137),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_155),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_144),
.C(n_155),
.Y(n_173)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_150),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_151),
.C(n_154),
.Y(n_177)
);

BUFx24_ASAP7_75t_SL g388 ( 
.A(n_146),
.Y(n_388)
);

FAx1_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_148),
.CI(n_149),
.CON(n_146),
.SN(n_146)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_147),
.B(n_148),
.C(n_149),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_156),
.B(n_163),
.C(n_171),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_163),
.B1(n_171),
.B2(n_172),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_158),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_161),
.B(n_162),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_161),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_199),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_162),
.B(n_199),
.C(n_200),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_163),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_168),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_169),
.C(n_170),
.Y(n_194)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx8_ASAP7_75t_L g326 ( 
.A(n_167),
.Y(n_326)
);

INVx6_ASAP7_75t_L g348 ( 
.A(n_167),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_195),
.B2(n_209),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_196),
.C(n_197),
.Y(n_210)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_179),
.C(n_188),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_188),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_180),
.B(n_184),
.C(n_187),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_182),
.B(n_231),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_186),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_194),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_190),
.B(n_193),
.C(n_194),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_192),
.Y(n_193)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_195),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_201),
.B(n_241),
.C(n_242),
.Y(n_265)
);

FAx1_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_205),
.CI(n_208),
.CON(n_201),
.SN(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_204),
.B(n_231),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_243),
.B2(n_244),
.Y(n_211)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_212),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_213),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_235),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_235),
.C(n_243),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_223),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_215),
.B(n_224),
.C(n_225),
.Y(n_264)
);

BUFx24_ASAP7_75t_SL g390 ( 
.A(n_215),
.Y(n_390)
);

FAx1_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_218),
.CI(n_220),
.CON(n_215),
.SN(n_215)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_216),
.B(n_218),
.C(n_220),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_217),
.B(n_222),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_222),
.B(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_222),
.B(n_231),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_234),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_226),
.Y(n_234)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_232),
.B2(n_233),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_229),
.A2(n_230),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_233),
.C(n_234),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_229),
.B(n_252),
.C(n_255),
.Y(n_299)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_238),
.C(n_239),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_249),
.C(n_275),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_263),
.B2(n_275),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_257),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_251),
.B(n_258),
.C(n_259),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_255),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_255),
.A2(n_256),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_SL g316 ( 
.A(n_255),
.B(n_281),
.C(n_284),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

BUFx24_ASAP7_75t_SL g389 ( 
.A(n_259),
.Y(n_389)
);

FAx1_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_261),
.CI(n_262),
.CON(n_259),
.SN(n_259)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_261),
.C(n_262),
.Y(n_286)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_263),
.Y(n_275)
);

BUFx24_ASAP7_75t_SL g394 ( 
.A(n_263),
.Y(n_394)
);

FAx1_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_265),
.CI(n_266),
.CON(n_263),
.SN(n_263)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_264),
.B(n_265),
.C(n_266),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_274),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_270),
.C(n_272),
.Y(n_294)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_269),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_270),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_271),
.A2(n_272),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_272),
.B(n_298),
.C(n_299),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_300),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_291),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_291),
.C(n_300),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_285),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_280),
.B(n_286),
.C(n_287),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_283),
.A2(n_284),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_SL g343 ( 
.A(n_284),
.B(n_309),
.C(n_311),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g393 ( 
.A(n_287),
.Y(n_393)
);

FAx1_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_289),
.CI(n_290),
.CON(n_287),
.SN(n_287)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_289),
.C(n_290),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_294),
.C(n_295),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_299),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_297),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_303),
.B(n_305),
.C(n_318),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_317),
.B2(n_318),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_313),
.B2(n_314),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_315),
.C(n_316),
.Y(n_335)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_311),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g349 ( 
.A1(n_311),
.A2(n_312),
.B1(n_350),
.B2(n_351),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_311),
.B(n_351),
.C(n_352),
.Y(n_364)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_319),
.B(n_321),
.C(n_324),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_323),
.B2(n_324),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_324),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_327),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_325),
.B(n_328),
.C(n_331),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_329),
.B1(n_330),
.B2(n_331),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_329),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_330),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_334),
.A2(n_354),
.B1(n_355),
.B2(n_356),
.Y(n_333)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_334),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_335),
.B(n_336),
.C(n_356),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_342),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_337),
.B(n_343),
.C(n_344),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_338),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_338),
.B(n_361),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_338),
.B(n_359),
.C(n_361),
.Y(n_380)
);

FAx1_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_340),
.CI(n_341),
.CON(n_338),
.SN(n_338)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_349),
.B1(n_352),
.B2(n_353),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_345),
.Y(n_352)
);

INVx8_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx8_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_349),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_350),
.A2(n_351),
.B1(n_368),
.B2(n_369),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_351),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_368),
.C(n_371),
.Y(n_374)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_354),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_362),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_362),
.B(n_373),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_362),
.B(n_374),
.C(n_375),
.Y(n_381)
);

FAx1_ASAP7_75t_SL g362 ( 
.A(n_363),
.B(n_364),
.CI(n_365),
.CON(n_362),
.SN(n_362)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_366),
.A2(n_367),
.B1(n_370),
.B2(n_371),
.Y(n_365)
);

CKINVDCx14_ASAP7_75t_R g366 ( 
.A(n_367),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_368),
.A2(n_369),
.B1(n_378),
.B2(n_379),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_369),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_SL g387 ( 
.A(n_369),
.B(n_376),
.C(n_379),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_370),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_378),
.A2(n_379),
.B1(n_385),
.B2(n_386),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_379),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_383),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g383 ( 
.A(n_384),
.B(n_387),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_385),
.Y(n_386)
);


endmodule