module fake_jpeg_24498_n_303 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_303);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_155;
wire n_207;
wire n_31;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx8_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_7),
.B(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_7),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_39),
.Y(n_57)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_28),
.Y(n_47)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g45 ( 
.A(n_36),
.Y(n_45)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_0),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_11),
.B(n_7),
.Y(n_62)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_42),
.B(n_47),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_27),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_55),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_26),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_29),
.B(n_32),
.C(n_18),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_28),
.B1(n_37),
.B2(n_19),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_29),
.C(n_16),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_19),
.B1(n_28),
.B2(n_24),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_52),
.A2(n_29),
.B1(n_18),
.B2(n_16),
.Y(n_76)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_23),
.B1(n_24),
.B2(n_15),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_54),
.A2(n_56),
.B1(n_61),
.B2(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_27),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_23),
.B1(n_15),
.B2(n_25),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_61)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_68),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_44),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_71),
.A2(n_49),
.B(n_51),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_72),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_20),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_82),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_46),
.B(n_29),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_74),
.A2(n_51),
.B(n_60),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_64),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_75),
.A2(n_76),
.B1(n_50),
.B2(n_45),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_77),
.Y(n_105)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

BUFx2_ASAP7_75t_SL g92 ( 
.A(n_79),
.Y(n_92)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_20),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_50),
.B1(n_45),
.B2(n_57),
.Y(n_96)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_103),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_96),
.B(n_78),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_72),
.B(n_59),
.Y(n_97)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_99),
.A2(n_66),
.B(n_86),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_100),
.A2(n_112),
.B1(n_114),
.B2(n_69),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_46),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_83),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

INVxp33_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_110),
.A2(n_71),
.B(n_78),
.Y(n_117)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_83),
.B(n_17),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_83),
.B(n_17),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_117),
.A2(n_90),
.B1(n_48),
.B2(n_95),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_91),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_120),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_110),
.A2(n_89),
.B1(n_84),
.B2(n_74),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_119),
.A2(n_126),
.B1(n_127),
.B2(n_133),
.Y(n_144)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_124),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_74),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_138),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_91),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_125),
.A2(n_109),
.B1(n_101),
.B2(n_48),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_89),
.B1(n_96),
.B2(n_108),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_106),
.A2(n_74),
.B1(n_50),
.B2(n_82),
.Y(n_127)
);

FAx1_ASAP7_75t_SL g160 ( 
.A(n_128),
.B(n_137),
.CI(n_39),
.CON(n_160),
.SN(n_160)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_130),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_108),
.A2(n_53),
.B1(n_83),
.B2(n_90),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_135),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_0),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_36),
.Y(n_140)
);

MAJx2_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_92),
.C(n_36),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_97),
.Y(n_143)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

OAI32xp33_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_111),
.A3(n_114),
.B1(n_105),
.B2(n_107),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_127),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_158),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_148),
.B(n_151),
.Y(n_184)
);

AO22x1_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_92),
.B1(n_105),
.B2(n_68),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_149),
.A2(n_153),
.B(n_165),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_160),
.Y(n_171)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_137),
.B(n_107),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_117),
.A2(n_90),
.B1(n_66),
.B2(n_85),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_157),
.A2(n_113),
.B1(n_95),
.B2(n_48),
.Y(n_178)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_161),
.Y(n_179)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_163),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_164),
.B(n_104),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_128),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_180),
.C(n_143),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_141),
.B(n_131),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_167),
.B(n_145),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_169),
.A2(n_176),
.B1(n_183),
.B2(n_156),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_170),
.A2(n_174),
.B(n_153),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_162),
.A2(n_116),
.B(n_138),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_175),
.B(n_182),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_116),
.B1(n_138),
.B2(n_123),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_178),
.A2(n_185),
.B1(n_189),
.B2(n_45),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_123),
.Y(n_180)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_154),
.A2(n_140),
.B(n_21),
.C(n_22),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_155),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_149),
.A2(n_70),
.B1(n_80),
.B2(n_81),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_187),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_147),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_144),
.A2(n_80),
.B1(n_87),
.B2(n_64),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_192),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_144),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_200),
.Y(n_223)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_172),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_201),
.Y(n_217)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_196),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_188),
.A2(n_153),
.B1(n_160),
.B2(n_148),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_197),
.A2(n_212),
.B1(n_183),
.B2(n_169),
.Y(n_219)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_160),
.B(n_156),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_168),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_171),
.B(n_150),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_173),
.C(n_176),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_203),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_156),
.C(n_163),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_204),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_206),
.A2(n_189),
.B1(n_186),
.B2(n_170),
.Y(n_225)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_168),
.Y(n_207)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_207),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_175),
.B(n_21),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_209),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_184),
.Y(n_211)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_190),
.Y(n_213)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_220),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_219),
.A2(n_218),
.B1(n_214),
.B2(n_216),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_171),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_225),
.A2(n_212),
.B1(n_203),
.B2(n_202),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_206),
.B(n_200),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_231),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_229),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_193),
.B(n_177),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_208),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_213),
.Y(n_237)
);

OAI22x1_ASAP7_75t_L g233 ( 
.A1(n_215),
.A2(n_192),
.B1(n_197),
.B2(n_177),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_233),
.A2(n_248),
.B1(n_249),
.B2(n_18),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_235),
.A2(n_222),
.B1(n_220),
.B2(n_226),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_217),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_242),
.Y(n_261)
);

FAx1_ASAP7_75t_SL g239 ( 
.A(n_225),
.B(n_182),
.CI(n_210),
.CON(n_239),
.SN(n_239)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_244),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_205),
.C(n_194),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_247),
.C(n_31),
.Y(n_254)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_195),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_245),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_201),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_204),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_231),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_9),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_223),
.C(n_221),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_224),
.A2(n_31),
.B1(n_22),
.B2(n_18),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_245),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_259),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_233),
.A2(n_94),
.B1(n_64),
.B2(n_3),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_255),
.A2(n_262),
.B1(n_8),
.B2(n_14),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_256),
.Y(n_273)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_257),
.A2(n_260),
.B(n_263),
.Y(n_270)
);

MAJx2_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_9),
.C(n_14),
.Y(n_258)
);

OAI21x1_ASAP7_75t_SL g271 ( 
.A1(n_258),
.A2(n_8),
.B(n_14),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_94),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_94),
.C(n_2),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_261),
.B(n_253),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_264),
.B(n_265),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_250),
.B(n_239),
.Y(n_266)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_266),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_243),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_269),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_234),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_271),
.A2(n_275),
.B(n_258),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_274),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_254),
.B(n_241),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_263),
.B(n_12),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_270),
.A2(n_255),
.B(n_268),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_276),
.B(n_10),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_9),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_252),
.C(n_2),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_280),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_1),
.C(n_2),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_267),
.A2(n_11),
.B(n_10),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_8),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_273),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_285),
.B(n_287),
.Y(n_293)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_286),
.Y(n_292)
);

NOR3xp33_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_291),
.C(n_3),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_1),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_278),
.C(n_284),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_1),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_286),
.C(n_282),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_295),
.A2(n_296),
.B(n_3),
.Y(n_297)
);

AO21x1_ASAP7_75t_L g296 ( 
.A1(n_290),
.A2(n_282),
.B(n_4),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_297),
.B(n_298),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_292),
.Y(n_300)
);

OA21x2_ASAP7_75t_L g301 ( 
.A1(n_300),
.A2(n_293),
.B(n_5),
.Y(n_301)
);

O2A1O1Ixp33_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_4),
.B(n_6),
.C(n_286),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_302),
.A2(n_6),
.B(n_297),
.Y(n_303)
);


endmodule