module fake_jpeg_1560_n_35 (n_3, n_2, n_1, n_0, n_4, n_5, n_35);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_35;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

INVx6_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

BUFx12_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_6),
.B(n_0),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_12),
.A2(n_8),
.B(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_11),
.B(n_9),
.C(n_10),
.Y(n_14)
);

OAI32xp33_ASAP7_75t_L g21 ( 
.A1(n_14),
.A2(n_8),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_11),
.B(n_3),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_15),
.A2(n_16),
.B1(n_17),
.B2(n_1),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_22),
.C(n_4),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_12),
.A2(n_8),
.B1(n_1),
.B2(n_0),
.Y(n_19)
);

AO22x1_ASAP7_75t_SL g23 ( 
.A1(n_19),
.A2(n_13),
.B1(n_15),
.B2(n_14),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_22),
.Y(n_28)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_26),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_25),
.B(n_19),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_28),
.Y(n_31)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

MAJx2_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_23),
.C(n_17),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_31),
.Y(n_33)
);

AO21x2_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_31),
.B(n_5),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_5),
.Y(n_35)
);


endmodule