module real_aes_8924_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g249 ( .A1(n_0), .A2(n_250), .B(n_251), .C(n_254), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_1), .B(n_238), .Y(n_255) );
INVx1_ASAP7_75t_L g441 ( .A(n_2), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_3), .B(n_166), .Y(n_165) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_4), .A2(n_127), .B(n_130), .C(n_513), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_5), .A2(n_122), .B(n_537), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_6), .A2(n_122), .B(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_7), .B(n_238), .Y(n_543) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_8), .A2(n_157), .B(n_194), .Y(n_193) );
AND2x6_ASAP7_75t_L g127 ( .A(n_9), .B(n_128), .Y(n_127) );
A2O1A1Ixp33_ASAP7_75t_L g210 ( .A1(n_10), .A2(n_127), .B(n_130), .C(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g481 ( .A(n_11), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_12), .B(n_40), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_13), .B(n_214), .Y(n_515) );
INVx1_ASAP7_75t_L g148 ( .A(n_14), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_15), .B(n_166), .Y(n_200) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_16), .A2(n_167), .B(n_499), .C(n_501), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_17), .B(n_238), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_18), .B(n_142), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g129 ( .A1(n_19), .A2(n_130), .B(n_133), .C(n_141), .Y(n_129) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_20), .A2(n_202), .B(n_253), .C(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_21), .B(n_214), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_22), .A2(n_54), .B1(n_745), .B2(n_746), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_22), .Y(n_745) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_23), .B(n_214), .Y(n_454) );
CKINVDCx16_ASAP7_75t_R g528 ( .A(n_24), .Y(n_528) );
INVx1_ASAP7_75t_L g453 ( .A(n_25), .Y(n_453) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_26), .A2(n_130), .B(n_141), .C(n_197), .Y(n_196) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_27), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_28), .Y(n_511) );
INVx1_ASAP7_75t_L g469 ( .A(n_29), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_30), .A2(n_122), .B(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g125 ( .A(n_31), .Y(n_125) );
A2O1A1Ixp33_ASAP7_75t_L g178 ( .A1(n_32), .A2(n_170), .B(n_179), .C(n_181), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_33), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g539 ( .A1(n_34), .A2(n_253), .B(n_540), .C(n_542), .Y(n_539) );
INVxp67_ASAP7_75t_L g470 ( .A(n_35), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_36), .B(n_199), .Y(n_198) );
A2O1A1Ixp33_ASAP7_75t_L g451 ( .A1(n_37), .A2(n_130), .B(n_141), .C(n_452), .Y(n_451) );
CKINVDCx14_ASAP7_75t_R g538 ( .A(n_38), .Y(n_538) );
AOI222xp33_ASAP7_75t_SL g104 ( .A1(n_39), .A2(n_105), .B1(n_111), .B2(n_720), .C1(n_721), .C2(n_725), .Y(n_104) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_41), .A2(n_254), .B(n_479), .C(n_480), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_42), .B(n_121), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_43), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_44), .B(n_166), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_45), .B(n_122), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_46), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_47), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_48), .A2(n_170), .B(n_179), .C(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g252 ( .A(n_49), .Y(n_252) );
OAI22xp5_ASAP7_75t_SL g742 ( .A1(n_50), .A2(n_743), .B1(n_744), .B2(n_747), .Y(n_742) );
CKINVDCx16_ASAP7_75t_R g747 ( .A(n_50), .Y(n_747) );
INVx1_ASAP7_75t_L g224 ( .A(n_51), .Y(n_224) );
INVx1_ASAP7_75t_L g487 ( .A(n_52), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_53), .B(n_122), .Y(n_221) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_54), .A2(n_103), .B1(n_729), .B2(n_738), .C1(n_752), .C2(n_758), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_54), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g150 ( .A(n_55), .Y(n_150) );
CKINVDCx14_ASAP7_75t_R g477 ( .A(n_56), .Y(n_477) );
INVx1_ASAP7_75t_L g128 ( .A(n_57), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_58), .B(n_122), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_59), .B(n_238), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_60), .A2(n_140), .B(n_163), .C(n_235), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_61), .Y(n_751) );
INVx1_ASAP7_75t_L g147 ( .A(n_62), .Y(n_147) );
OAI22xp5_ASAP7_75t_L g106 ( .A1(n_63), .A2(n_101), .B1(n_107), .B2(n_108), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_63), .Y(n_108) );
INVx1_ASAP7_75t_SL g541 ( .A(n_64), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_65), .Y(n_734) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_66), .B(n_166), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_67), .B(n_238), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_68), .B(n_167), .Y(n_212) );
INVx1_ASAP7_75t_L g531 ( .A(n_69), .Y(n_531) );
CKINVDCx16_ASAP7_75t_R g248 ( .A(n_70), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_71), .B(n_135), .Y(n_134) );
A2O1A1Ixp33_ASAP7_75t_L g160 ( .A1(n_72), .A2(n_130), .B(n_161), .C(n_170), .Y(n_160) );
CKINVDCx16_ASAP7_75t_R g233 ( .A(n_73), .Y(n_233) );
INVx1_ASAP7_75t_L g733 ( .A(n_74), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_75), .A2(n_122), .B(n_476), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_76), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_77), .A2(n_122), .B(n_496), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_78), .A2(n_121), .B(n_465), .Y(n_464) );
CKINVDCx16_ASAP7_75t_R g450 ( .A(n_79), .Y(n_450) );
INVx1_ASAP7_75t_L g497 ( .A(n_80), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g137 ( .A(n_81), .B(n_138), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_82), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_83), .A2(n_122), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g500 ( .A(n_84), .Y(n_500) );
INVx2_ASAP7_75t_L g145 ( .A(n_85), .Y(n_145) );
INVx1_ASAP7_75t_L g514 ( .A(n_86), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_87), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_88), .B(n_214), .Y(n_213) );
OR2x2_ASAP7_75t_L g439 ( .A(n_89), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g719 ( .A(n_89), .Y(n_719) );
OR2x2_ASAP7_75t_L g737 ( .A(n_89), .B(n_728), .Y(n_737) );
OAI22xp5_ASAP7_75t_SL g105 ( .A1(n_90), .A2(n_106), .B1(n_109), .B2(n_110), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_90), .Y(n_110) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_91), .A2(n_130), .B(n_170), .C(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_92), .B(n_122), .Y(n_177) );
INVx1_ASAP7_75t_L g182 ( .A(n_93), .Y(n_182) );
INVxp67_ASAP7_75t_L g236 ( .A(n_94), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_95), .B(n_157), .Y(n_482) );
INVx1_ASAP7_75t_L g162 ( .A(n_96), .Y(n_162) );
INVx1_ASAP7_75t_L g208 ( .A(n_97), .Y(n_208) );
INVx2_ASAP7_75t_L g490 ( .A(n_98), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_99), .B(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g226 ( .A(n_100), .B(n_144), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_101), .Y(n_107) );
INVxp67_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g720 ( .A(n_105), .Y(n_720) );
INVx1_ASAP7_75t_L g109 ( .A(n_106), .Y(n_109) );
OAI22xp5_ASAP7_75t_SL g111 ( .A1(n_112), .A2(n_437), .B1(n_443), .B2(n_716), .Y(n_111) );
OAI22xp5_ASAP7_75t_SL g740 ( .A1(n_112), .A2(n_723), .B1(n_741), .B2(n_742), .Y(n_740) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g723 ( .A(n_113), .Y(n_723) );
AND3x1_ASAP7_75t_L g113 ( .A(n_114), .B(n_341), .C(n_398), .Y(n_113) );
NOR3xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_286), .C(n_322), .Y(n_114) );
OAI211xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_188), .B(n_240), .C(n_273), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_152), .Y(n_116) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x4_ASAP7_75t_L g243 ( .A(n_118), .B(n_244), .Y(n_243) );
INVx5_ASAP7_75t_L g272 ( .A(n_118), .Y(n_272) );
AND2x2_ASAP7_75t_L g345 ( .A(n_118), .B(n_261), .Y(n_345) );
AND2x2_ASAP7_75t_L g383 ( .A(n_118), .B(n_289), .Y(n_383) );
AND2x2_ASAP7_75t_L g403 ( .A(n_118), .B(n_245), .Y(n_403) );
OR2x6_ASAP7_75t_L g118 ( .A(n_119), .B(n_149), .Y(n_118) );
AOI21xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_129), .B(n_142), .Y(n_119) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x4_ASAP7_75t_L g122 ( .A(n_123), .B(n_127), .Y(n_122) );
NAND2x1p5_ASAP7_75t_L g209 ( .A(n_123), .B(n_127), .Y(n_209) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_126), .Y(n_123) );
INVx1_ASAP7_75t_L g140 ( .A(n_124), .Y(n_140) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g131 ( .A(n_125), .Y(n_131) );
INVx1_ASAP7_75t_L g203 ( .A(n_125), .Y(n_203) );
INVx1_ASAP7_75t_L g132 ( .A(n_126), .Y(n_132) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_126), .Y(n_136) );
INVx3_ASAP7_75t_L g167 ( .A(n_126), .Y(n_167) );
INVx1_ASAP7_75t_L g199 ( .A(n_126), .Y(n_199) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_126), .Y(n_214) );
BUFx3_ASAP7_75t_L g141 ( .A(n_127), .Y(n_141) );
INVx4_ASAP7_75t_SL g171 ( .A(n_127), .Y(n_171) );
INVx5_ASAP7_75t_L g180 ( .A(n_130), .Y(n_180) );
AND2x6_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_131), .Y(n_169) );
BUFx3_ASAP7_75t_L g185 ( .A(n_131), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_137), .B(n_139), .Y(n_133) );
INVx2_ASAP7_75t_L g138 ( .A(n_135), .Y(n_138) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx4_ASAP7_75t_L g164 ( .A(n_136), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_L g181 ( .A1(n_138), .A2(n_182), .B(n_183), .C(n_184), .Y(n_181) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_138), .A2(n_184), .B(n_224), .C(n_225), .Y(n_223) );
O2A1O1Ixp5_ASAP7_75t_L g513 ( .A1(n_138), .A2(n_514), .B(n_515), .C(n_516), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_138), .A2(n_516), .B(n_531), .C(n_532), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_L g452 ( .A1(n_139), .A2(n_166), .B(n_453), .C(n_454), .Y(n_452) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_140), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_143), .B(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g151 ( .A(n_144), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_144), .A2(n_177), .B(n_178), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_144), .A2(n_221), .B(n_222), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_L g449 ( .A1(n_144), .A2(n_209), .B(n_450), .C(n_451), .Y(n_449) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_144), .A2(n_475), .B(n_482), .Y(n_474) );
AND2x2_ASAP7_75t_SL g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AND2x2_ASAP7_75t_L g158 ( .A(n_145), .B(n_146), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
AO21x2_ASAP7_75t_L g509 ( .A1(n_151), .A2(n_510), .B(n_517), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_152), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g152 ( .A(n_153), .B(n_175), .Y(n_152) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_153), .Y(n_284) );
AND2x2_ASAP7_75t_L g298 ( .A(n_153), .B(n_244), .Y(n_298) );
INVx1_ASAP7_75t_L g321 ( .A(n_153), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_153), .B(n_272), .Y(n_360) );
OR2x2_ASAP7_75t_L g397 ( .A(n_153), .B(n_242), .Y(n_397) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_154), .Y(n_333) );
AND2x2_ASAP7_75t_L g340 ( .A(n_154), .B(n_245), .Y(n_340) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AND2x2_ASAP7_75t_L g261 ( .A(n_155), .B(n_245), .Y(n_261) );
BUFx2_ASAP7_75t_L g289 ( .A(n_155), .Y(n_289) );
AO21x2_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_159), .B(n_173), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_156), .B(n_174), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_156), .B(n_187), .Y(n_186) );
AO21x2_ASAP7_75t_L g206 ( .A1(n_156), .A2(n_207), .B(n_215), .Y(n_206) );
INVx3_ASAP7_75t_L g238 ( .A(n_156), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_156), .B(n_456), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_156), .B(n_518), .Y(n_517) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_156), .A2(n_527), .B(n_533), .Y(n_526) );
INVx4_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_157), .A2(n_195), .B(n_196), .Y(n_194) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_157), .Y(n_230) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g217 ( .A(n_158), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_172), .Y(n_159) );
O2A1O1Ixp33_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_165), .C(n_168), .Y(n_161) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
OAI22xp33_ASAP7_75t_L g468 ( .A1(n_164), .A2(n_166), .B1(n_469), .B2(n_470), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_164), .B(n_490), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_164), .B(n_500), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_166), .B(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g250 ( .A(n_166), .Y(n_250) );
INVx5_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_167), .B(n_481), .Y(n_480) );
HB1xp67_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx3_ASAP7_75t_L g542 ( .A(n_169), .Y(n_542) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_171), .A2(n_180), .B(n_233), .C(n_234), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_SL g247 ( .A1(n_171), .A2(n_180), .B(n_248), .C(n_249), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_SL g465 ( .A1(n_171), .A2(n_180), .B(n_466), .C(n_467), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_SL g476 ( .A1(n_171), .A2(n_180), .B(n_477), .C(n_478), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_SL g486 ( .A1(n_171), .A2(n_180), .B(n_487), .C(n_488), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_SL g496 ( .A1(n_171), .A2(n_180), .B(n_497), .C(n_498), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_L g537 ( .A1(n_171), .A2(n_180), .B(n_538), .C(n_539), .Y(n_537) );
INVx5_ASAP7_75t_L g242 ( .A(n_175), .Y(n_242) );
BUFx2_ASAP7_75t_L g265 ( .A(n_175), .Y(n_265) );
AND2x2_ASAP7_75t_L g422 ( .A(n_175), .B(n_276), .Y(n_422) );
OR2x6_ASAP7_75t_L g175 ( .A(n_176), .B(n_186), .Y(n_175) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g254 ( .A(n_185), .Y(n_254) );
INVx1_ASAP7_75t_L g501 ( .A(n_185), .Y(n_501) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NAND2xp33_ASAP7_75t_L g189 ( .A(n_190), .B(n_227), .Y(n_189) );
OAI221xp5_ASAP7_75t_L g322 ( .A1(n_190), .A2(n_323), .B1(n_330), .B2(n_331), .C(n_334), .Y(n_322) );
OR2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_204), .Y(n_190) );
AND2x2_ASAP7_75t_L g228 ( .A(n_191), .B(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_191), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_SL g191 ( .A(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g257 ( .A(n_192), .B(n_205), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_192), .B(n_206), .Y(n_267) );
OR2x2_ASAP7_75t_L g278 ( .A(n_192), .B(n_229), .Y(n_278) );
AND2x2_ASAP7_75t_L g281 ( .A(n_192), .B(n_269), .Y(n_281) );
AND2x2_ASAP7_75t_L g297 ( .A(n_192), .B(n_218), .Y(n_297) );
OR2x2_ASAP7_75t_L g313 ( .A(n_192), .B(n_206), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_192), .B(n_229), .Y(n_375) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_193), .B(n_218), .Y(n_367) );
AND2x2_ASAP7_75t_L g370 ( .A(n_193), .B(n_206), .Y(n_370) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_200), .B(n_201), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_201), .A2(n_212), .B(n_213), .Y(n_211) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
OR2x2_ASAP7_75t_L g291 ( .A(n_204), .B(n_278), .Y(n_291) );
INVx2_ASAP7_75t_L g317 ( .A(n_204), .Y(n_317) );
OR2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_218), .Y(n_204) );
AND2x2_ASAP7_75t_L g239 ( .A(n_205), .B(n_219), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_205), .B(n_229), .Y(n_296) );
OR2x2_ASAP7_75t_L g307 ( .A(n_205), .B(n_219), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_205), .B(n_269), .Y(n_366) );
OAI221xp5_ASAP7_75t_L g399 ( .A1(n_205), .A2(n_400), .B1(n_402), .B2(n_404), .C(n_407), .Y(n_399) );
INVx5_ASAP7_75t_SL g205 ( .A(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_206), .B(n_229), .Y(n_338) );
OAI21xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_210), .Y(n_207) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_209), .A2(n_511), .B(n_512), .Y(n_510) );
OAI21xp5_ASAP7_75t_L g527 ( .A1(n_209), .A2(n_528), .B(n_529), .Y(n_527) );
INVx4_ASAP7_75t_L g253 ( .A(n_214), .Y(n_253) );
INVx2_ASAP7_75t_L g479 ( .A(n_214), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
INVx2_ASAP7_75t_L g462 ( .A(n_217), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_218), .B(n_269), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_218), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g285 ( .A(n_218), .B(n_257), .Y(n_285) );
OR2x2_ASAP7_75t_L g329 ( .A(n_218), .B(n_229), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_218), .B(n_281), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_218), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g394 ( .A(n_218), .B(n_395), .Y(n_394) );
INVx5_ASAP7_75t_SL g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_SL g258 ( .A(n_219), .B(n_228), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_SL g262 ( .A1(n_219), .A2(n_263), .B(n_266), .C(n_270), .Y(n_262) );
OR2x2_ASAP7_75t_L g300 ( .A(n_219), .B(n_296), .Y(n_300) );
OR2x2_ASAP7_75t_L g336 ( .A(n_219), .B(n_278), .Y(n_336) );
OAI311xp33_ASAP7_75t_L g342 ( .A1(n_219), .A2(n_281), .A3(n_343), .B1(n_346), .C1(n_353), .Y(n_342) );
AND2x2_ASAP7_75t_L g393 ( .A(n_219), .B(n_229), .Y(n_393) );
AND2x2_ASAP7_75t_L g401 ( .A(n_219), .B(n_256), .Y(n_401) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_219), .Y(n_419) );
AND2x2_ASAP7_75t_L g436 ( .A(n_219), .B(n_257), .Y(n_436) );
OR2x6_ASAP7_75t_L g219 ( .A(n_220), .B(n_226), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_228), .B(n_239), .Y(n_227) );
AND2x2_ASAP7_75t_L g264 ( .A(n_228), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g420 ( .A(n_228), .Y(n_420) );
AND2x2_ASAP7_75t_L g256 ( .A(n_229), .B(n_257), .Y(n_256) );
INVx3_ASAP7_75t_L g269 ( .A(n_229), .Y(n_269) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_229), .Y(n_312) );
INVxp67_ASAP7_75t_L g351 ( .A(n_229), .Y(n_351) );
OA21x2_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_237), .Y(n_229) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_230), .A2(n_485), .B(n_491), .Y(n_484) );
OA21x2_ASAP7_75t_L g494 ( .A1(n_230), .A2(n_495), .B(n_502), .Y(n_494) );
OA21x2_ASAP7_75t_L g535 ( .A1(n_230), .A2(n_536), .B(n_543), .Y(n_535) );
OA21x2_ASAP7_75t_L g245 ( .A1(n_238), .A2(n_246), .B(n_255), .Y(n_245) );
AND2x2_ASAP7_75t_L g429 ( .A(n_239), .B(n_277), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_256), .B1(n_258), .B2(n_259), .C(n_262), .Y(n_240) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_242), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g282 ( .A(n_242), .B(n_272), .Y(n_282) );
AND2x2_ASAP7_75t_L g290 ( .A(n_242), .B(n_244), .Y(n_290) );
OR2x2_ASAP7_75t_L g302 ( .A(n_242), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g320 ( .A(n_242), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g344 ( .A(n_242), .B(n_345), .Y(n_344) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_242), .Y(n_364) );
AND2x2_ASAP7_75t_L g416 ( .A(n_242), .B(n_340), .Y(n_416) );
OAI31xp33_ASAP7_75t_L g424 ( .A1(n_242), .A2(n_293), .A3(n_392), .B(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_243), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_SL g388 ( .A(n_243), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_243), .B(n_397), .Y(n_396) );
AND2x4_ASAP7_75t_L g276 ( .A(n_244), .B(n_272), .Y(n_276) );
INVx1_ASAP7_75t_L g363 ( .A(n_244), .Y(n_363) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g413 ( .A(n_245), .B(n_272), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_253), .B(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g516 ( .A(n_254), .Y(n_516) );
INVx1_ASAP7_75t_SL g423 ( .A(n_256), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_257), .B(n_328), .Y(n_327) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_258), .A2(n_370), .B1(n_408), .B2(n_411), .Y(n_407) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g271 ( .A(n_261), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g330 ( .A(n_261), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_261), .B(n_282), .Y(n_435) );
INVx1_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g405 ( .A(n_264), .B(n_406), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_265), .A2(n_324), .B(n_326), .Y(n_323) );
OR2x2_ASAP7_75t_L g331 ( .A(n_265), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g352 ( .A(n_265), .B(n_340), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_265), .B(n_363), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_265), .B(n_403), .Y(n_402) );
OAI221xp5_ASAP7_75t_SL g379 ( .A1(n_266), .A2(n_380), .B1(n_385), .B2(n_388), .C(n_389), .Y(n_379) );
OR2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
OR2x2_ASAP7_75t_L g356 ( .A(n_267), .B(n_329), .Y(n_356) );
INVx1_ASAP7_75t_L g395 ( .A(n_267), .Y(n_395) );
INVx2_ASAP7_75t_L g371 ( .A(n_268), .Y(n_371) );
INVx1_ASAP7_75t_L g305 ( .A(n_269), .Y(n_305) );
INVx1_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g310 ( .A(n_272), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_272), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g339 ( .A(n_272), .B(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g427 ( .A(n_272), .B(n_397), .Y(n_427) );
AOI222xp33_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_277), .B1(n_279), .B2(n_282), .C1(n_283), .C2(n_285), .Y(n_273) );
INVxp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g283 ( .A(n_276), .B(n_284), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_276), .A2(n_326), .B1(n_354), .B2(n_355), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_276), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
OAI21xp33_ASAP7_75t_SL g314 ( .A1(n_285), .A2(n_315), .B(n_318), .Y(n_314) );
OAI211xp5_ASAP7_75t_SL g286 ( .A1(n_287), .A2(n_291), .B(n_292), .C(n_314), .Y(n_286) );
INVxp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
AOI221xp5_ASAP7_75t_L g292 ( .A1(n_290), .A2(n_293), .B1(n_298), .B2(n_299), .C(n_301), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_290), .B(n_378), .Y(n_377) );
INVxp67_ASAP7_75t_L g384 ( .A(n_290), .Y(n_384) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
AND2x2_ASAP7_75t_L g386 ( .A(n_295), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g303 ( .A(n_298), .Y(n_303) );
AND2x2_ASAP7_75t_L g309 ( .A(n_298), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_304), .B1(n_308), .B2(n_311), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_305), .B(n_317), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_306), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g406 ( .A(n_310), .Y(n_406) );
AND2x2_ASAP7_75t_L g425 ( .A(n_310), .B(n_340), .Y(n_425) );
OR2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_317), .B(n_374), .Y(n_433) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_320), .B(n_388), .Y(n_431) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g354 ( .A(n_332), .Y(n_354) );
BUFx2_ASAP7_75t_L g378 ( .A(n_333), .Y(n_378) );
OAI21xp5_ASAP7_75t_SL g334 ( .A1(n_335), .A2(n_337), .B(n_339), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NOR3xp33_ASAP7_75t_L g341 ( .A(n_342), .B(n_357), .C(n_379), .Y(n_341) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OAI21xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_349), .B(n_352), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
A2O1A1Ixp33_ASAP7_75t_SL g357 ( .A1(n_358), .A2(n_361), .B(n_365), .C(n_368), .Y(n_357) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_358), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NOR2xp67_ASAP7_75t_SL g362 ( .A(n_363), .B(n_364), .Y(n_362) );
OR2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx1_ASAP7_75t_SL g387 ( .A(n_367), .Y(n_387) );
OAI21xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_372), .B(n_376), .Y(n_368) );
AND2x4_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
AND2x2_ASAP7_75t_L g392 ( .A(n_370), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_382), .B(n_384), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_392), .B1(n_394), .B2(n_396), .Y(n_389) );
INVx2_ASAP7_75t_SL g410 ( .A(n_397), .Y(n_410) );
NOR3xp33_ASAP7_75t_L g398 ( .A(n_399), .B(n_414), .C(n_426), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVxp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVxp67_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_410), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OAI221xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_417), .B1(n_421), .B2(n_423), .C(n_424), .Y(n_414) );
A2O1A1Ixp33_ASAP7_75t_L g426 ( .A1(n_415), .A2(n_427), .B(n_428), .C(n_430), .Y(n_426) );
INVx1_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_432), .B1(n_434), .B2(n_436), .Y(n_430) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g722 ( .A(n_438), .Y(n_722) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OR2x2_ASAP7_75t_L g718 ( .A(n_440), .B(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g728 ( .A(n_440), .Y(n_728) );
AND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
INVx1_ASAP7_75t_SL g724 ( .A(n_443), .Y(n_724) );
OR5x1_ASAP7_75t_L g443 ( .A(n_444), .B(n_610), .C(n_674), .D(n_690), .E(n_705), .Y(n_443) );
NAND4xp25_ASAP7_75t_L g444 ( .A(n_445), .B(n_544), .C(n_571), .D(n_594), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_492), .B(n_503), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_447), .B(n_457), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx3_ASAP7_75t_SL g523 ( .A(n_448), .Y(n_523) );
AND2x4_ASAP7_75t_L g557 ( .A(n_448), .B(n_546), .Y(n_557) );
OR2x2_ASAP7_75t_L g567 ( .A(n_448), .B(n_525), .Y(n_567) );
OR2x2_ASAP7_75t_L g613 ( .A(n_448), .B(n_460), .Y(n_613) );
AND2x2_ASAP7_75t_L g627 ( .A(n_448), .B(n_524), .Y(n_627) );
AND2x2_ASAP7_75t_L g670 ( .A(n_448), .B(n_560), .Y(n_670) );
AND2x2_ASAP7_75t_L g677 ( .A(n_448), .B(n_535), .Y(n_677) );
AND2x2_ASAP7_75t_L g696 ( .A(n_448), .B(n_586), .Y(n_696) );
AND2x2_ASAP7_75t_L g714 ( .A(n_448), .B(n_556), .Y(n_714) );
OR2x6_ASAP7_75t_L g448 ( .A(n_449), .B(n_455), .Y(n_448) );
INVx1_ASAP7_75t_L g679 ( .A(n_457), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_473), .Y(n_457) );
AND2x2_ASAP7_75t_L g589 ( .A(n_458), .B(n_524), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_458), .B(n_609), .Y(n_608) );
AOI32xp33_ASAP7_75t_L g622 ( .A1(n_458), .A2(n_623), .A3(n_626), .B1(n_628), .B2(n_632), .Y(n_622) );
AND2x2_ASAP7_75t_L g692 ( .A(n_458), .B(n_586), .Y(n_692) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g556 ( .A(n_460), .B(n_525), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_460), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g598 ( .A(n_460), .B(n_545), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_460), .B(n_677), .Y(n_676) );
AO21x2_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_463), .B(n_471), .Y(n_460) );
INVx1_ASAP7_75t_L g561 ( .A(n_461), .Y(n_561) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OA21x2_ASAP7_75t_L g560 ( .A1(n_464), .A2(n_472), .B(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g563 ( .A(n_473), .B(n_507), .Y(n_563) );
AND2x2_ASAP7_75t_L g639 ( .A(n_473), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_SL g711 ( .A(n_473), .Y(n_711) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_483), .Y(n_473) );
OR2x2_ASAP7_75t_L g506 ( .A(n_474), .B(n_484), .Y(n_506) );
AND2x2_ASAP7_75t_L g520 ( .A(n_474), .B(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_474), .B(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g570 ( .A(n_474), .Y(n_570) );
AND2x2_ASAP7_75t_L g597 ( .A(n_474), .B(n_484), .Y(n_597) );
BUFx3_ASAP7_75t_L g600 ( .A(n_474), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_474), .B(n_575), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_474), .B(n_694), .Y(n_693) );
INVx2_ASAP7_75t_L g551 ( .A(n_483), .Y(n_551) );
AND2x2_ASAP7_75t_L g569 ( .A(n_483), .B(n_549), .Y(n_569) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g580 ( .A(n_484), .B(n_494), .Y(n_580) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_484), .Y(n_593) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_493), .B(n_600), .Y(n_650) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_SL g521 ( .A(n_494), .Y(n_521) );
NAND3xp33_ASAP7_75t_L g568 ( .A(n_494), .B(n_569), .C(n_570), .Y(n_568) );
OR2x2_ASAP7_75t_L g576 ( .A(n_494), .B(n_549), .Y(n_576) );
AND2x2_ASAP7_75t_L g596 ( .A(n_494), .B(n_549), .Y(n_596) );
AND2x2_ASAP7_75t_L g640 ( .A(n_494), .B(n_509), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_519), .B(n_522), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_505), .B(n_507), .Y(n_504) );
AND2x2_ASAP7_75t_L g715 ( .A(n_505), .B(n_640), .Y(n_715) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_506), .A2(n_613), .B1(n_655), .B2(n_657), .Y(n_654) );
OR2x2_ASAP7_75t_L g661 ( .A(n_506), .B(n_576), .Y(n_661) );
OR2x2_ASAP7_75t_L g685 ( .A(n_506), .B(n_686), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_506), .B(n_605), .Y(n_698) );
AND2x2_ASAP7_75t_L g591 ( .A(n_507), .B(n_592), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g678 ( .A1(n_507), .A2(n_664), .B(n_679), .Y(n_678) );
AOI32xp33_ASAP7_75t_L g699 ( .A1(n_507), .A2(n_589), .A3(n_700), .B1(n_702), .B2(n_703), .Y(n_699) );
OR2x2_ASAP7_75t_L g710 ( .A(n_507), .B(n_711), .Y(n_710) );
CKINVDCx16_ASAP7_75t_R g507 ( .A(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g578 ( .A(n_508), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_508), .B(n_592), .Y(n_657) );
BUFx3_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx4_ASAP7_75t_L g549 ( .A(n_509), .Y(n_549) );
AND2x2_ASAP7_75t_L g615 ( .A(n_509), .B(n_580), .Y(n_615) );
AND3x2_ASAP7_75t_L g624 ( .A(n_509), .B(n_520), .C(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g550 ( .A(n_521), .B(n_551), .Y(n_550) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_521), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_521), .B(n_549), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
AND2x2_ASAP7_75t_L g545 ( .A(n_523), .B(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g585 ( .A(n_523), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g603 ( .A(n_523), .B(n_535), .Y(n_603) );
AND2x2_ASAP7_75t_L g621 ( .A(n_523), .B(n_525), .Y(n_621) );
OR2x2_ASAP7_75t_L g635 ( .A(n_523), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g681 ( .A(n_523), .B(n_609), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_524), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_535), .Y(n_524) );
AND2x2_ASAP7_75t_L g582 ( .A(n_525), .B(n_560), .Y(n_582) );
OR2x2_ASAP7_75t_L g636 ( .A(n_525), .B(n_560), .Y(n_636) );
AND2x2_ASAP7_75t_L g689 ( .A(n_525), .B(n_546), .Y(n_689) );
INVx2_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
BUFx2_ASAP7_75t_L g587 ( .A(n_526), .Y(n_587) );
AND2x2_ASAP7_75t_L g609 ( .A(n_526), .B(n_535), .Y(n_609) );
INVx2_ASAP7_75t_L g546 ( .A(n_535), .Y(n_546) );
INVx1_ASAP7_75t_L g566 ( .A(n_535), .Y(n_566) );
AOI211xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_547), .B(n_552), .C(n_564), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_545), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g708 ( .A(n_545), .Y(n_708) );
AND2x2_ASAP7_75t_L g586 ( .A(n_546), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_549), .B(n_550), .Y(n_558) );
INVx1_ASAP7_75t_L g643 ( .A(n_549), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_549), .B(n_570), .Y(n_667) );
AND2x2_ASAP7_75t_L g683 ( .A(n_549), .B(n_597), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_550), .B(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g574 ( .A(n_551), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_558), .B1(n_559), .B2(n_562), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_557), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_555), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_556), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g581 ( .A(n_557), .B(n_582), .Y(n_581) );
AOI221xp5_ASAP7_75t_SL g646 ( .A1(n_557), .A2(n_599), .B1(n_647), .B2(n_652), .C(n_654), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_557), .B(n_620), .Y(n_653) );
INVx1_ASAP7_75t_L g713 ( .A(n_559), .Y(n_713) );
BUFx3_ASAP7_75t_L g620 ( .A(n_560), .Y(n_620) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AOI21xp33_ASAP7_75t_SL g564 ( .A1(n_565), .A2(n_567), .B(n_568), .Y(n_564) );
INVx1_ASAP7_75t_L g629 ( .A(n_566), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_566), .B(n_620), .Y(n_673) );
INVx1_ASAP7_75t_L g630 ( .A(n_567), .Y(n_630) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_567), .B(n_620), .Y(n_631) );
INVxp67_ASAP7_75t_L g651 ( .A(n_569), .Y(n_651) );
AND2x2_ASAP7_75t_L g592 ( .A(n_570), .B(n_593), .Y(n_592) );
O2A1O1Ixp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_577), .B(n_581), .C(n_583), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
INVx1_ASAP7_75t_SL g606 ( .A(n_574), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_575), .B(n_606), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_575), .B(n_597), .Y(n_648) );
INVx2_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_578), .A2(n_584), .B1(n_588), .B2(n_590), .Y(n_583) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g599 ( .A(n_580), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g644 ( .A(n_580), .B(n_645), .Y(n_644) );
OAI21xp33_ASAP7_75t_L g647 ( .A1(n_582), .A2(n_648), .B(n_649), .Y(n_647) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
AOI221xp5_ASAP7_75t_L g594 ( .A1(n_586), .A2(n_595), .B1(n_598), .B2(n_599), .C(n_601), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_586), .B(n_620), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_586), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g702 ( .A(n_592), .Y(n_702) );
INVxp67_ASAP7_75t_L g625 ( .A(n_593), .Y(n_625) );
INVx1_ASAP7_75t_L g632 ( .A(n_595), .Y(n_632) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
AND2x2_ASAP7_75t_L g671 ( .A(n_596), .B(n_600), .Y(n_671) );
INVx1_ASAP7_75t_L g645 ( .A(n_600), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_600), .B(n_615), .Y(n_675) );
OAI32xp33_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_604), .A3(n_606), .B1(n_607), .B2(n_608), .Y(n_601) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_SL g614 ( .A(n_609), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_609), .B(n_641), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_609), .B(n_670), .Y(n_701) );
NAND2x1p5_ASAP7_75t_L g709 ( .A(n_609), .B(n_620), .Y(n_709) );
NAND5xp2_ASAP7_75t_L g610 ( .A(n_611), .B(n_633), .C(n_646), .D(n_658), .E(n_659), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_615), .B1(n_616), .B2(n_618), .C(n_622), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp33_ASAP7_75t_SL g637 ( .A(n_617), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_620), .B(n_689), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_621), .A2(n_634), .B1(n_637), .B2(n_641), .Y(n_633) );
INVx2_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
OAI211xp5_ASAP7_75t_SL g628 ( .A1(n_624), .A2(n_629), .B(n_630), .C(n_631), .Y(n_628) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_SL g656 ( .A(n_636), .Y(n_656) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_645), .B(n_694), .Y(n_704) );
OR2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AOI222xp33_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_662), .B1(n_664), .B2(n_668), .C1(n_671), .C2(n_672), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_676), .B1(n_678), .B2(n_680), .C(n_682), .Y(n_674) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
OAI21xp33_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_684), .B(n_687), .Y(n_682) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g694 ( .A(n_686), .Y(n_694) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
OAI221xp5_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_693), .B1(n_695), .B2(n_697), .C(n_699), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
INVxp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
A2O1A1Ixp33_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_709), .B(n_710), .C(n_712), .Y(n_705) );
INVxp67_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OAI21xp33_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_714), .B(n_715), .Y(n_712) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_718), .A2(n_722), .B1(n_723), .B2(n_724), .Y(n_721) );
NOR2x2_ASAP7_75t_L g727 ( .A(n_719), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
NAND2xp33_ASAP7_75t_L g730 ( .A(n_731), .B(n_735), .Y(n_730) );
NOR2xp33_ASAP7_75t_SL g731 ( .A(n_732), .B(n_734), .Y(n_731) );
INVx1_ASAP7_75t_SL g757 ( .A(n_732), .Y(n_757) );
INVx1_ASAP7_75t_L g756 ( .A(n_734), .Y(n_756) );
OA21x2_ASAP7_75t_L g759 ( .A1(n_734), .A2(n_748), .B(n_757), .Y(n_759) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
BUFx2_ASAP7_75t_L g748 ( .A(n_737), .Y(n_748) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_737), .Y(n_750) );
INVxp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_748), .B(n_749), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
NOR2xp33_ASAP7_75t_SL g749 ( .A(n_750), .B(n_751), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_753), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_L g754 ( .A(n_755), .B(n_757), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_759), .Y(n_758) );
endmodule