module fake_jpeg_3739_n_321 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_29),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_20),
.B(n_23),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_33),
.Y(n_54)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_41),
.B(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_42),
.B(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_31),
.A2(n_27),
.B1(n_23),
.B2(n_20),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_55),
.A2(n_27),
.B1(n_18),
.B2(n_15),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_56),
.A2(n_57),
.B1(n_73),
.B2(n_14),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_27),
.B1(n_18),
.B2(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_65),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_39),
.A2(n_27),
.B1(n_34),
.B2(n_32),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_43),
.B1(n_48),
.B2(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_64),
.B(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_67),
.Y(n_83)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_69),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_32),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_41),
.Y(n_80)
);

NOR2x1_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_24),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_SL g95 ( 
.A(n_71),
.B(n_24),
.C(n_16),
.Y(n_95)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_39),
.A2(n_18),
.B1(n_19),
.B2(n_14),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_74),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_19),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_78),
.A2(n_88),
.B1(n_76),
.B2(n_58),
.Y(n_118)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_86),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_89),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_48),
.C(n_50),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_93),
.C(n_59),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_61),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_42),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_71),
.A2(n_43),
.B1(n_50),
.B2(n_24),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_43),
.C(n_40),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_97),
.B(n_75),
.C(n_65),
.Y(n_101)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_71),
.A2(n_16),
.B1(n_19),
.B2(n_17),
.Y(n_97)
);

AO22x2_ASAP7_75t_L g98 ( 
.A1(n_56),
.A2(n_36),
.B1(n_38),
.B2(n_53),
.Y(n_98)
);

OA21x2_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_47),
.B(n_49),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_51),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_101),
.B(n_81),
.Y(n_129)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_107),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_106),
.Y(n_133)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_110),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_98),
.A2(n_57),
.B1(n_62),
.B2(n_67),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_118),
.B1(n_98),
.B2(n_93),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_115),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_60),
.B(n_73),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_113),
.A2(n_88),
.B(n_98),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_94),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_40),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_116),
.A2(n_69),
.B(n_72),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_119),
.Y(n_147)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_122),
.Y(n_130)
);

OAI22x1_ASAP7_75t_SL g135 ( 
.A1(n_121),
.A2(n_98),
.B1(n_90),
.B2(n_36),
.Y(n_135)
);

AND2x6_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_40),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_128),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_92),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_126),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_92),
.B(n_81),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_125),
.A2(n_145),
.B(n_101),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_96),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_127),
.A2(n_129),
.B(n_15),
.Y(n_172)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_131),
.A2(n_135),
.B1(n_137),
.B2(n_144),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_115),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_111),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_91),
.C(n_86),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_138),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_122),
.A2(n_97),
.B1(n_91),
.B2(n_95),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_85),
.C(n_77),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_139),
.A2(n_102),
.B(n_105),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_49),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_140),
.B(n_109),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_85),
.C(n_77),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_102),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_76),
.B1(n_87),
.B2(n_79),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_119),
.A2(n_58),
.B1(n_112),
.B2(n_74),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_58),
.B1(n_17),
.B2(n_15),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_146),
.A2(n_68),
.B1(n_28),
.B2(n_25),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_149),
.A2(n_157),
.B(n_160),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_130),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_135),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_151),
.B(n_153),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_124),
.B(n_107),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_138),
.C(n_143),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_142),
.B(n_108),
.Y(n_156)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

INVx13_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_159),
.Y(n_181)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

AO21x1_ASAP7_75t_L g160 ( 
.A1(n_135),
.A2(n_121),
.B(n_103),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_164),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_141),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_162),
.Y(n_187)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_111),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_167),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_111),
.Y(n_168)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_110),
.Y(n_169)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_17),
.Y(n_170)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_100),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_171),
.B(n_174),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_172),
.A2(n_173),
.B(n_132),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_100),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_82),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_175),
.A2(n_159),
.B1(n_167),
.B2(n_162),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_195),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_174),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_184),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_178),
.A2(n_201),
.B(n_170),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_182),
.C(n_155),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_136),
.C(n_140),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_164),
.A2(n_127),
.B1(n_144),
.B2(n_146),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_154),
.B(n_132),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_188),
.B(n_189),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_154),
.B(n_137),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_158),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_168),
.A2(n_130),
.B1(n_131),
.B2(n_139),
.Y(n_194)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_194),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_150),
.Y(n_195)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_199),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_150),
.B(n_47),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_157),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_172),
.A2(n_26),
.B(n_22),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_208),
.C(n_219),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_149),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_206),
.B(n_25),
.Y(n_244)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_207),
.B(n_214),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_148),
.Y(n_209)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_210),
.A2(n_217),
.B(n_25),
.Y(n_239)
);

INVxp33_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_148),
.Y(n_212)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_192),
.A2(n_152),
.B1(n_151),
.B2(n_173),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_216),
.A2(n_198),
.B1(n_190),
.B2(n_191),
.Y(n_226)
);

AOI21xp33_ASAP7_75t_L g217 ( 
.A1(n_185),
.A2(n_153),
.B(n_166),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_156),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_218),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_152),
.C(n_161),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_169),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_201),
.C(n_197),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_158),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_221),
.B(n_223),
.Y(n_229)
);

FAx1_ASAP7_75t_SL g223 ( 
.A(n_194),
.B(n_165),
.CI(n_151),
.CON(n_223),
.SN(n_223)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_215),
.A2(n_192),
.B1(n_185),
.B2(n_198),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_225),
.A2(n_228),
.B1(n_230),
.B2(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_226),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_215),
.A2(n_182),
.B1(n_191),
.B2(n_196),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_202),
.A2(n_196),
.B1(n_160),
.B2(n_178),
.Y(n_230)
);

XNOR2x1_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_179),
.Y(n_232)
);

NOR2xp67_ASAP7_75t_SL g261 ( 
.A(n_232),
.B(n_244),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_223),
.A2(n_160),
.B1(n_186),
.B2(n_197),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_238),
.C(n_219),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_165),
.C(n_175),
.Y(n_238)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_117),
.Y(n_240)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_203),
.A2(n_117),
.B1(n_68),
.B2(n_22),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_241),
.B(n_216),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_223),
.A2(n_68),
.B1(n_22),
.B2(n_26),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_210),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_220),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_256),
.C(n_259),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_28),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_231),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_252),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_218),
.Y(n_248)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_248),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_249),
.A2(n_258),
.B1(n_243),
.B2(n_239),
.Y(n_267)
);

NAND3xp33_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_208),
.C(n_222),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_250),
.B(n_246),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_212),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_255),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_225),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_235),
.B(n_209),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_204),
.C(n_45),
.Y(n_256)
);

AO221x1_ASAP7_75t_L g258 ( 
.A1(n_237),
.A2(n_45),
.B1(n_44),
.B2(n_22),
.C(n_26),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_204),
.C(n_45),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_228),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_26),
.C(n_22),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_226),
.C(n_236),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_264),
.A2(n_1),
.B(n_2),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_267),
.Y(n_287)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_274),
.C(n_1),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_269),
.A2(n_270),
.B(n_279),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_233),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_273),
.C(n_278),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_230),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_227),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_251),
.A2(n_233),
.B1(n_25),
.B2(n_12),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_260),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_44),
.C(n_26),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_263),
.C(n_259),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_0),
.Y(n_279)
);

NOR2xp67_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_245),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_280),
.A2(n_284),
.B1(n_274),
.B2(n_276),
.Y(n_294)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_281),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_283),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_257),
.Y(n_283)
);

NOR2xp67_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_0),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_289),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_272),
.C(n_277),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_290),
.A2(n_2),
.B(n_3),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_2),
.C(n_3),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_3),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_2),
.C(n_3),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_4),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_SL g310 ( 
.A1(n_294),
.A2(n_297),
.B(n_295),
.C(n_9),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_301),
.C(n_6),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_298),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_287),
.A2(n_38),
.B1(n_36),
.B2(n_6),
.Y(n_299)
);

AOI322xp5_ASAP7_75t_L g306 ( 
.A1(n_299),
.A2(n_300),
.A3(n_303),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_306)
);

NAND4xp25_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_4),
.C(n_5),
.D(n_6),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_4),
.Y(n_301)
);

OAI21x1_ASAP7_75t_L g303 ( 
.A1(n_290),
.A2(n_281),
.B(n_291),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_307),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_306),
.B(n_308),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_7),
.C(n_8),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_296),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_309),
.B(n_297),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_8),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_312),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_314),
.B(n_310),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_305),
.C(n_313),
.Y(n_317)
);

AOI322xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_315),
.C2(n_316),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_318),
.B(n_10),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_10),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_11),
.Y(n_321)
);


endmodule