module fake_jpeg_30562_n_35 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_35);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_35;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_13),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_10),
.B(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_21),
.B1(n_18),
.B2(n_6),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_17),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_15),
.B(n_4),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_4),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_25),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_27),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_22),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_16),
.C(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_18),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_30),
.B2(n_24),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_SL g32 ( 
.A(n_28),
.B(n_25),
.C(n_14),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_5),
.B1(n_6),
.B2(n_11),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_34),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_35)
);


endmodule