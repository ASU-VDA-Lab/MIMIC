module fake_netlist_1_8635_n_1168 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_1168);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1168;
wire n_663;
wire n_791;
wire n_707;
wire n_361;
wire n_513;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_667;
wire n_496;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_1158;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_1122;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_1161;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_1163;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_786;
wire n_724;
wire n_857;
wire n_345;
wire n_360;
wire n_1090;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1024;
wire n_1016;
wire n_1097;
wire n_572;
wire n_1017;
wire n_324;
wire n_1078;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_1060;
wire n_279;
wire n_303;
wire n_975;
wire n_968;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_1025;
wire n_1011;
wire n_1132;
wire n_880;
wire n_1101;
wire n_1155;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_255;
wire n_426;
wire n_624;
wire n_769;
wire n_725;
wire n_818;
wire n_844;
wire n_1160;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_293;
wire n_1138;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_1154;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_935;
wire n_427;
wire n_910;
wire n_950;
wire n_460;
wire n_1046;
wire n_478;
wire n_415;
wire n_482;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_805;
wire n_729;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_1145;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_1167;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_1157;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_990;
wire n_751;
wire n_800;
wire n_626;
wire n_941;
wire n_1147;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_875;
wire n_832;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_649;
wire n_526;
wire n_276;
wire n_527;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_446;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_666;
wire n_621;
wire n_799;
wire n_1089;
wire n_1058;
wire n_370;
wire n_1050;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_899;
wire n_260;
wire n_806;
wire n_881;
wire n_539;
wire n_1066;
wire n_1055;
wire n_974;
wire n_1153;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_315;
wire n_409;
wire n_363;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_1144;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_1152;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_1149;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_419;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_1125;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_955;
wire n_1133;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_1159;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_1110;
wire n_327;
wire n_944;
wire n_325;
wire n_1131;
wire n_1102;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_1156;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_947;
wire n_620;
wire n_841;
wire n_924;
wire n_912;
wire n_1043;
wire n_1141;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1142;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1117;
wire n_1040;
wire n_1165;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_1143;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_901;
wire n_834;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1164;
wire n_1038;
wire n_341;
wire n_1162;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_1073;
wire n_323;
wire n_868;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_1150;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_1104;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_287;
wire n_1146;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_1137;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_1148;
wire n_709;
wire n_739;
wire n_1166;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_257;
wire n_992;
wire n_1127;
wire n_269;
CKINVDCx16_ASAP7_75t_R g255 ( .A(n_144), .Y(n_255) );
INVx1_ASAP7_75t_SL g256 ( .A(n_126), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_199), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_147), .Y(n_258) );
CKINVDCx20_ASAP7_75t_R g259 ( .A(n_217), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_54), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_190), .Y(n_261) );
CKINVDCx20_ASAP7_75t_R g262 ( .A(n_138), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_186), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_60), .Y(n_264) );
OR2x2_ASAP7_75t_L g265 ( .A(n_12), .B(n_120), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_79), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_149), .Y(n_267) );
INVx1_ASAP7_75t_SL g268 ( .A(n_60), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_115), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_119), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_24), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_91), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_162), .Y(n_273) );
CKINVDCx16_ASAP7_75t_R g274 ( .A(n_168), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_209), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_183), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_195), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_57), .Y(n_278) );
INVx3_ASAP7_75t_L g279 ( .A(n_202), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_150), .Y(n_280) );
BUFx3_ASAP7_75t_L g281 ( .A(n_182), .Y(n_281) );
BUFx10_ASAP7_75t_L g282 ( .A(n_49), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_237), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_243), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_77), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_16), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_63), .Y(n_287) );
CKINVDCx16_ASAP7_75t_R g288 ( .A(n_110), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_53), .Y(n_289) );
INVx1_ASAP7_75t_SL g290 ( .A(n_28), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_141), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_214), .Y(n_292) );
INVxp67_ASAP7_75t_L g293 ( .A(n_49), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_127), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_246), .Y(n_295) );
BUFx2_ASAP7_75t_L g296 ( .A(n_94), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_113), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_124), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_234), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_188), .Y(n_300) );
CKINVDCx20_ASAP7_75t_R g301 ( .A(n_122), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_201), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_128), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_142), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_114), .Y(n_305) );
CKINVDCx20_ASAP7_75t_R g306 ( .A(n_3), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_139), .Y(n_307) );
BUFx2_ASAP7_75t_L g308 ( .A(n_143), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_205), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_121), .Y(n_310) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_38), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_35), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_247), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_250), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_31), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_16), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_107), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_223), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_148), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_92), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_11), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_85), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_174), .Y(n_323) );
BUFx3_ASAP7_75t_L g324 ( .A(n_67), .Y(n_324) );
CKINVDCx20_ASAP7_75t_R g325 ( .A(n_75), .Y(n_325) );
CKINVDCx20_ASAP7_75t_R g326 ( .A(n_169), .Y(n_326) );
XOR2xp5_ASAP7_75t_L g327 ( .A(n_135), .B(n_134), .Y(n_327) );
INVx1_ASAP7_75t_SL g328 ( .A(n_11), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_1), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_40), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_43), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_230), .Y(n_332) );
BUFx3_ASAP7_75t_L g333 ( .A(n_133), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_117), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_24), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_7), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_198), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_61), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_69), .B(n_10), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_215), .Y(n_340) );
CKINVDCx16_ASAP7_75t_R g341 ( .A(n_27), .Y(n_341) );
INVx2_ASAP7_75t_SL g342 ( .A(n_104), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_28), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_218), .Y(n_344) );
CKINVDCx20_ASAP7_75t_R g345 ( .A(n_55), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_232), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_69), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_164), .Y(n_348) );
CKINVDCx20_ASAP7_75t_R g349 ( .A(n_225), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_57), .Y(n_350) );
CKINVDCx20_ASAP7_75t_R g351 ( .A(n_90), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_185), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_140), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_1), .Y(n_354) );
CKINVDCx20_ASAP7_75t_R g355 ( .A(n_109), .Y(n_355) );
INVx2_ASAP7_75t_SL g356 ( .A(n_118), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_17), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_248), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_166), .Y(n_359) );
BUFx5_ASAP7_75t_L g360 ( .A(n_13), .Y(n_360) );
BUFx3_ASAP7_75t_L g361 ( .A(n_8), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_44), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_108), .Y(n_363) );
CKINVDCx20_ASAP7_75t_R g364 ( .A(n_123), .Y(n_364) );
BUFx2_ASAP7_75t_SL g365 ( .A(n_229), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_91), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_146), .Y(n_367) );
INVx2_ASAP7_75t_SL g368 ( .A(n_33), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_116), .Y(n_369) );
INVx2_ASAP7_75t_SL g370 ( .A(n_204), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_112), .Y(n_371) );
INVx1_ASAP7_75t_SL g372 ( .A(n_101), .Y(n_372) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_206), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_153), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_111), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_56), .Y(n_376) );
CKINVDCx20_ASAP7_75t_R g377 ( .A(n_242), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_167), .Y(n_378) );
CKINVDCx14_ASAP7_75t_R g379 ( .A(n_207), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_180), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_231), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_178), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_203), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_62), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_20), .Y(n_385) );
CKINVDCx16_ASAP7_75t_R g386 ( .A(n_165), .Y(n_386) );
INVxp33_ASAP7_75t_SL g387 ( .A(n_125), .Y(n_387) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_65), .Y(n_388) );
INVx1_ASAP7_75t_SL g389 ( .A(n_22), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_89), .Y(n_390) );
CKINVDCx16_ASAP7_75t_R g391 ( .A(n_216), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_145), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_59), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_252), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_35), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_81), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_254), .Y(n_397) );
NOR2x1_ASAP7_75t_L g398 ( .A(n_324), .B(n_0), .Y(n_398) );
NOR2x1_ASAP7_75t_L g399 ( .A(n_324), .B(n_0), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_279), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_279), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_341), .A2(n_4), .B1(n_2), .B2(n_3), .Y(n_402) );
BUFx2_ASAP7_75t_L g403 ( .A(n_296), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_303), .Y(n_404) );
BUFx12f_ASAP7_75t_L g405 ( .A(n_308), .Y(n_405) );
INVx5_ASAP7_75t_L g406 ( .A(n_303), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_303), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_306), .A2(n_345), .B1(n_351), .B2(n_325), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_303), .Y(n_409) );
NOR2xp33_ASAP7_75t_SL g410 ( .A(n_255), .B(n_98), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_379), .B(n_2), .Y(n_411) );
INVx3_ASAP7_75t_L g412 ( .A(n_360), .Y(n_412) );
AND2x4_ASAP7_75t_L g413 ( .A(n_361), .B(n_4), .Y(n_413) );
OAI21x1_ASAP7_75t_L g414 ( .A1(n_269), .A2(n_100), .B(n_99), .Y(n_414) );
INVxp33_ASAP7_75t_SL g415 ( .A(n_266), .Y(n_415) );
BUFx2_ASAP7_75t_L g416 ( .A(n_361), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_368), .B(n_5), .Y(n_417) );
OAI21x1_ASAP7_75t_L g418 ( .A1(n_269), .A2(n_103), .B(n_102), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_360), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_379), .B(n_5), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_274), .B(n_6), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_360), .Y(n_422) );
INVx5_ASAP7_75t_L g423 ( .A(n_342), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_360), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_356), .B(n_6), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_360), .Y(n_426) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_281), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_370), .B(n_7), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_360), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_293), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_360), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_283), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_283), .Y(n_433) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_281), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_260), .B(n_8), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_264), .B(n_9), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_288), .B(n_9), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_313), .Y(n_438) );
CKINVDCx16_ASAP7_75t_R g439 ( .A(n_386), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_313), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_412), .Y(n_441) );
CKINVDCx11_ASAP7_75t_R g442 ( .A(n_439), .Y(n_442) );
OAI22xp33_ASAP7_75t_SL g443 ( .A1(n_410), .A2(n_387), .B1(n_391), .B2(n_265), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_412), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_439), .Y(n_445) );
INVx3_ASAP7_75t_L g446 ( .A(n_413), .Y(n_446) );
INVx3_ASAP7_75t_L g447 ( .A(n_413), .Y(n_447) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_414), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_412), .Y(n_449) );
CKINVDCx5p33_ASAP7_75t_R g450 ( .A(n_415), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_412), .Y(n_451) );
INVx4_ASAP7_75t_L g452 ( .A(n_413), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_419), .Y(n_453) );
INVxp33_ASAP7_75t_L g454 ( .A(n_403), .Y(n_454) );
NAND2xp33_ASAP7_75t_L g455 ( .A(n_411), .B(n_397), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_419), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_423), .B(n_387), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_424), .Y(n_458) );
BUFx2_ASAP7_75t_L g459 ( .A(n_411), .Y(n_459) );
AO21x2_ASAP7_75t_L g460 ( .A1(n_414), .A2(n_263), .B(n_258), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_423), .B(n_273), .Y(n_461) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_403), .A2(n_262), .B1(n_267), .B2(n_259), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_416), .B(n_282), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_416), .B(n_271), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_429), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_429), .Y(n_466) );
AND2x4_ASAP7_75t_L g467 ( .A(n_413), .B(n_385), .Y(n_467) );
INVx3_ASAP7_75t_L g468 ( .A(n_400), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_424), .Y(n_469) );
INVx2_ASAP7_75t_SL g470 ( .A(n_420), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_431), .Y(n_471) );
INVx4_ASAP7_75t_L g472 ( .A(n_422), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_422), .B(n_272), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_431), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_426), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_420), .B(n_257), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_423), .B(n_261), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_426), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_426), .Y(n_479) );
OAI22xp33_ASAP7_75t_L g480 ( .A1(n_402), .A2(n_325), .B1(n_345), .B2(n_306), .Y(n_480) );
XNOR2xp5_ASAP7_75t_L g481 ( .A(n_408), .B(n_351), .Y(n_481) );
INVx2_ASAP7_75t_SL g482 ( .A(n_423), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_432), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_423), .B(n_270), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_421), .B(n_287), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_405), .B(n_277), .Y(n_486) );
OR2x6_ASAP7_75t_L g487 ( .A(n_421), .B(n_365), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_472), .B(n_437), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_467), .Y(n_489) );
AO22x1_ASAP7_75t_L g490 ( .A1(n_462), .A2(n_437), .B1(n_430), .B2(n_399), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_454), .B(n_405), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_463), .B(n_408), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_473), .B(n_425), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_472), .B(n_428), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_472), .B(n_417), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_476), .B(n_435), .Y(n_496) );
BUFx3_ASAP7_75t_L g497 ( .A(n_442), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_467), .Y(n_498) );
INVx3_ASAP7_75t_L g499 ( .A(n_452), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_452), .B(n_284), .Y(n_500) );
AND3x2_ASAP7_75t_L g501 ( .A(n_459), .B(n_339), .C(n_327), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_463), .A2(n_402), .B1(n_262), .B2(n_301), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_470), .A2(n_267), .B1(n_326), .B2(n_301), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_446), .A2(n_433), .B1(n_438), .B2(n_432), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_472), .B(n_398), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_464), .B(n_436), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_470), .A2(n_459), .B1(n_485), .B2(n_487), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_443), .B(n_275), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_467), .Y(n_509) );
OAI22xp5_ASAP7_75t_SL g510 ( .A1(n_481), .A2(n_349), .B1(n_355), .B2(n_326), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_443), .B(n_276), .Y(n_511) );
BUFx12f_ASAP7_75t_L g512 ( .A(n_487), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_446), .B(n_399), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_446), .B(n_400), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_447), .B(n_400), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_441), .A2(n_418), .B(n_401), .Y(n_516) );
INVxp67_ASAP7_75t_L g517 ( .A(n_487), .Y(n_517) );
INVxp33_ASAP7_75t_L g518 ( .A(n_481), .Y(n_518) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_487), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_447), .B(n_401), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_486), .B(n_447), .Y(n_521) );
NOR2xp33_ASAP7_75t_SL g522 ( .A(n_487), .B(n_349), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_455), .A2(n_364), .B1(n_377), .B2(n_355), .Y(n_523) );
INVxp67_ASAP7_75t_L g524 ( .A(n_483), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_468), .Y(n_525) );
INVxp67_ASAP7_75t_L g526 ( .A(n_457), .Y(n_526) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_460), .Y(n_527) );
BUFx3_ASAP7_75t_L g528 ( .A(n_445), .Y(n_528) );
INVx3_ASAP7_75t_L g529 ( .A(n_448), .Y(n_529) );
INVx2_ASAP7_75t_SL g530 ( .A(n_460), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_448), .B(n_291), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_441), .B(n_401), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_448), .B(n_292), .Y(n_533) );
INVx3_ASAP7_75t_L g534 ( .A(n_448), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_478), .B(n_282), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_444), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_L g537 ( .A1(n_461), .A2(n_433), .B(n_440), .C(n_438), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_444), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_458), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_477), .B(n_295), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_484), .B(n_297), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_449), .A2(n_418), .B(n_440), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_480), .B(n_268), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_451), .B(n_280), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_444), .Y(n_545) );
AND2x2_ASAP7_75t_SL g546 ( .A(n_448), .B(n_339), .Y(n_546) );
BUFx3_ASAP7_75t_L g547 ( .A(n_478), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_465), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_465), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_466), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_466), .B(n_471), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_460), .A2(n_278), .B1(n_286), .B2(n_285), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_479), .A2(n_289), .B1(n_315), .B2(n_312), .Y(n_553) );
NOR2x1_ASAP7_75t_L g554 ( .A(n_479), .B(n_364), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_471), .B(n_298), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_474), .B(n_294), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_453), .B(n_302), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_453), .B(n_304), .Y(n_558) );
INVx5_ASAP7_75t_L g559 ( .A(n_482), .Y(n_559) );
INVx3_ASAP7_75t_L g560 ( .A(n_456), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_456), .B(n_305), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_469), .B(n_299), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_482), .B(n_300), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_475), .B(n_309), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_475), .B(n_310), .Y(n_565) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_448), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_506), .B(n_493), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_522), .A2(n_377), .B1(n_322), .B2(n_336), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_488), .A2(n_321), .B1(n_329), .B2(n_316), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_510), .B(n_290), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_491), .B(n_320), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_493), .B(n_343), .Y(n_572) );
AO32x1_ASAP7_75t_L g573 ( .A1(n_530), .A2(n_409), .A3(n_407), .B1(n_404), .B2(n_314), .Y(n_573) );
INVx4_ASAP7_75t_L g574 ( .A(n_512), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_489), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_507), .A2(n_362), .B1(n_366), .B2(n_357), .Y(n_576) );
AO21x2_ASAP7_75t_L g577 ( .A1(n_516), .A2(n_323), .B(n_307), .Y(n_577) );
INVx1_ASAP7_75t_SL g578 ( .A(n_535), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_519), .A2(n_330), .B1(n_335), .B2(n_331), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_517), .B(n_376), .Y(n_580) );
A2O1A1Ixp33_ASAP7_75t_L g581 ( .A1(n_548), .A2(n_338), .B(n_350), .C(n_347), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_495), .B(n_393), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_494), .B(n_496), .Y(n_583) );
INVx3_ASAP7_75t_L g584 ( .A(n_547), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_554), .A2(n_389), .B1(n_328), .B2(n_384), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_524), .A2(n_390), .B1(n_395), .B2(n_354), .Y(n_586) );
INVx3_ASAP7_75t_SL g587 ( .A(n_497), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_519), .A2(n_396), .B1(n_385), .B2(n_388), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_498), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_503), .B(n_311), .Y(n_590) );
A2O1A1Ixp33_ASAP7_75t_L g591 ( .A1(n_549), .A2(n_353), .B(n_358), .C(n_352), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_508), .B(n_256), .Y(n_592) );
NOR2x1_ASAP7_75t_L g593 ( .A(n_511), .B(n_367), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_521), .B(n_372), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_551), .A2(n_388), .B1(n_311), .B2(n_374), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_523), .B(n_490), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_502), .B(n_311), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_500), .A2(n_382), .B(n_381), .Y(n_598) );
A2O1A1Ixp33_ASAP7_75t_L g599 ( .A1(n_550), .A2(n_383), .B(n_318), .C(n_346), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_509), .Y(n_600) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_528), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_518), .B(n_317), .Y(n_602) );
O2A1O1Ixp33_ASAP7_75t_L g603 ( .A1(n_543), .A2(n_378), .B(n_363), .C(n_333), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_505), .B(n_319), .Y(n_604) );
AO21x1_ASAP7_75t_L g605 ( .A1(n_563), .A2(n_513), .B(n_562), .Y(n_605) );
O2A1O1Ixp33_ASAP7_75t_L g606 ( .A1(n_537), .A2(n_407), .B(n_409), .C(n_404), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_514), .Y(n_607) );
OAI21xp33_ASAP7_75t_L g608 ( .A1(n_552), .A2(n_434), .B(n_427), .Y(n_608) );
NAND2x1p5_ASAP7_75t_L g609 ( .A(n_499), .B(n_311), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_526), .B(n_332), .Y(n_610) );
CKINVDCx10_ASAP7_75t_R g611 ( .A(n_501), .Y(n_611) );
OAI21xp33_ASAP7_75t_L g612 ( .A1(n_552), .A2(n_434), .B(n_427), .Y(n_612) );
A2O1A1Ixp33_ASAP7_75t_L g613 ( .A1(n_563), .A2(n_388), .B(n_434), .C(n_427), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_499), .B(n_334), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_546), .B(n_337), .Y(n_615) );
AOI33xp33_ASAP7_75t_L g616 ( .A1(n_553), .A2(n_388), .A3(n_12), .B1(n_13), .B2(n_14), .B3(n_15), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_501), .B(n_10), .Y(n_617) );
AND2x4_ASAP7_75t_L g618 ( .A(n_559), .B(n_15), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_546), .B(n_340), .Y(n_619) );
NOR2xp33_ASAP7_75t_SL g620 ( .A(n_559), .B(n_344), .Y(n_620) );
A2O1A1Ixp33_ASAP7_75t_L g621 ( .A1(n_515), .A2(n_359), .B(n_369), .C(n_348), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_504), .A2(n_373), .B1(n_375), .B2(n_371), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_520), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_532), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_504), .A2(n_392), .B1(n_394), .B2(n_380), .Y(n_625) );
AOI221xp5_ASAP7_75t_L g626 ( .A1(n_555), .A2(n_406), .B1(n_19), .B2(n_20), .C(n_21), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_536), .Y(n_627) );
AND2x4_ASAP7_75t_SL g628 ( .A(n_560), .B(n_18), .Y(n_628) );
AOI21xp33_ASAP7_75t_L g629 ( .A1(n_556), .A2(n_18), .B(n_19), .Y(n_629) );
O2A1O1Ixp33_ASAP7_75t_L g630 ( .A1(n_555), .A2(n_26), .B(n_23), .C(n_25), .Y(n_630) );
NAND2x1p5_ASAP7_75t_L g631 ( .A(n_560), .B(n_406), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_538), .Y(n_632) );
NOR2xp33_ASAP7_75t_R g633 ( .A(n_540), .B(n_23), .Y(n_633) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_566), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_545), .Y(n_635) );
OR2x6_ASAP7_75t_L g636 ( .A(n_564), .B(n_26), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_544), .A2(n_106), .B(n_105), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_557), .B(n_29), .Y(n_638) );
O2A1O1Ixp33_ASAP7_75t_L g639 ( .A1(n_558), .A2(n_31), .B(n_29), .C(n_30), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_540), .B(n_30), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_539), .A2(n_34), .B1(n_32), .B2(n_33), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_541), .B(n_32), .Y(n_642) );
A2O1A1Ixp33_ASAP7_75t_L g643 ( .A1(n_541), .A2(n_34), .B(n_36), .C(n_37), .Y(n_643) );
BUFx2_ASAP7_75t_L g644 ( .A(n_561), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_565), .B(n_36), .Y(n_645) );
NAND3xp33_ASAP7_75t_SL g646 ( .A(n_525), .B(n_38), .C(n_39), .Y(n_646) );
OR2x6_ASAP7_75t_L g647 ( .A(n_512), .B(n_39), .Y(n_647) );
CKINVDCx10_ASAP7_75t_R g648 ( .A(n_497), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_491), .B(n_40), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_506), .B(n_41), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_547), .Y(n_651) );
OAI21x1_ASAP7_75t_L g652 ( .A1(n_542), .A2(n_130), .B(n_129), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_489), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_506), .B(n_42), .Y(n_654) );
OAI21xp5_ASAP7_75t_L g655 ( .A1(n_516), .A2(n_132), .B(n_131), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_522), .A2(n_42), .B1(n_43), .B2(n_44), .Y(n_656) );
A2O1A1Ixp33_ASAP7_75t_L g657 ( .A1(n_506), .A2(n_45), .B(n_46), .C(n_47), .Y(n_657) );
BUFx6f_ASAP7_75t_L g658 ( .A(n_547), .Y(n_658) );
NOR3xp33_ASAP7_75t_L g659 ( .A(n_510), .B(n_45), .C(n_46), .Y(n_659) );
O2A1O1Ixp33_ASAP7_75t_L g660 ( .A1(n_543), .A2(n_47), .B(n_48), .C(n_50), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_491), .B(n_50), .Y(n_661) );
OR2x2_ASAP7_75t_L g662 ( .A(n_510), .B(n_51), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_547), .Y(n_663) );
AO21x1_ASAP7_75t_L g664 ( .A1(n_516), .A2(n_51), .B(n_52), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_531), .A2(n_137), .B(n_136), .Y(n_665) );
A2O1A1Ixp33_ASAP7_75t_L g666 ( .A1(n_506), .A2(n_52), .B(n_53), .C(n_54), .Y(n_666) );
CKINVDCx11_ASAP7_75t_R g667 ( .A(n_497), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_547), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_490), .A2(n_55), .B1(n_56), .B2(n_58), .C(n_59), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_506), .B(n_61), .Y(n_670) );
CKINVDCx5p33_ASAP7_75t_R g671 ( .A(n_497), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_489), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_506), .B(n_63), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_519), .A2(n_64), .B1(n_65), .B2(n_66), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_491), .B(n_64), .Y(n_675) );
BUFx2_ASAP7_75t_SL g676 ( .A(n_618), .Y(n_676) );
AND2x4_ASAP7_75t_L g677 ( .A(n_578), .B(n_66), .Y(n_677) );
A2O1A1Ixp33_ASAP7_75t_L g678 ( .A1(n_603), .A2(n_67), .B(n_68), .C(n_70), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_632), .Y(n_679) );
NAND2xp5_ASAP7_75t_SL g680 ( .A(n_658), .B(n_68), .Y(n_680) );
A2O1A1Ixp33_ASAP7_75t_L g681 ( .A1(n_650), .A2(n_70), .B(n_71), .C(n_72), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_624), .A2(n_71), .B1(n_72), .B2(n_73), .Y(n_682) );
OAI221xp5_ASAP7_75t_L g683 ( .A1(n_596), .A2(n_73), .B1(n_74), .B2(n_75), .C(n_76), .Y(n_683) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_634), .Y(n_684) );
BUFx2_ASAP7_75t_L g685 ( .A(n_647), .Y(n_685) );
NAND3x1_ASAP7_75t_L g686 ( .A(n_659), .B(n_76), .C(n_77), .Y(n_686) );
AO31x2_ASAP7_75t_L g687 ( .A1(n_664), .A2(n_78), .A3(n_79), .B(n_80), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_597), .B(n_78), .Y(n_688) );
O2A1O1Ixp33_ASAP7_75t_SL g689 ( .A1(n_613), .A2(n_200), .B(n_253), .C(n_251), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g690 ( .A(n_667), .Y(n_690) );
NAND3xp33_ASAP7_75t_L g691 ( .A(n_639), .B(n_81), .C(n_82), .Y(n_691) );
BUFx3_ASAP7_75t_L g692 ( .A(n_587), .Y(n_692) );
INVxp67_ASAP7_75t_L g693 ( .A(n_647), .Y(n_693) );
OR2x2_ASAP7_75t_L g694 ( .A(n_570), .B(n_82), .Y(n_694) );
NOR2x1_ASAP7_75t_SL g695 ( .A(n_647), .B(n_83), .Y(n_695) );
OAI21xp5_ASAP7_75t_L g696 ( .A1(n_608), .A2(n_83), .B(n_84), .Y(n_696) );
AO31x2_ASAP7_75t_L g697 ( .A1(n_605), .A2(n_84), .A3(n_85), .B(n_86), .Y(n_697) );
A2O1A1Ixp33_ASAP7_75t_L g698 ( .A1(n_654), .A2(n_87), .B(n_88), .C(n_89), .Y(n_698) );
AO31x2_ASAP7_75t_L g699 ( .A1(n_599), .A2(n_87), .A3(n_88), .B(n_90), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_572), .B(n_92), .Y(n_700) );
AOI221x1_ASAP7_75t_L g701 ( .A1(n_612), .A2(n_93), .B1(n_94), .B2(n_95), .C(n_96), .Y(n_701) );
A2O1A1Ixp33_ASAP7_75t_L g702 ( .A1(n_670), .A2(n_93), .B(n_95), .C(n_96), .Y(n_702) );
OAI22x1_ASAP7_75t_L g703 ( .A1(n_568), .A2(n_97), .B1(n_151), .B2(n_152), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_579), .B(n_97), .Y(n_704) );
AOI221x1_ASAP7_75t_L g705 ( .A1(n_612), .A2(n_154), .B1(n_155), .B2(n_156), .C(n_157), .Y(n_705) );
CKINVDCx5p33_ASAP7_75t_R g706 ( .A(n_648), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_673), .Y(n_707) );
INVx2_ASAP7_75t_SL g708 ( .A(n_671), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_649), .A2(n_158), .B1(n_159), .B2(n_160), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_571), .B(n_161), .Y(n_710) );
INVx2_ASAP7_75t_SL g711 ( .A(n_601), .Y(n_711) );
NOR2xp67_ASAP7_75t_L g712 ( .A(n_618), .B(n_163), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_569), .B(n_170), .Y(n_713) );
BUFx10_ASAP7_75t_L g714 ( .A(n_628), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g715 ( .A(n_620), .B(n_171), .Y(n_715) );
A2O1A1Ixp33_ASAP7_75t_L g716 ( .A1(n_660), .A2(n_172), .B(n_173), .C(n_175), .Y(n_716) );
OAI21xp5_ASAP7_75t_L g717 ( .A1(n_607), .A2(n_176), .B(n_177), .Y(n_717) );
BUFx3_ASAP7_75t_L g718 ( .A(n_574), .Y(n_718) );
BUFx8_ASAP7_75t_SL g719 ( .A(n_617), .Y(n_719) );
INVxp67_ASAP7_75t_L g720 ( .A(n_636), .Y(n_720) );
AO31x2_ASAP7_75t_L g721 ( .A1(n_591), .A2(n_179), .A3(n_181), .B(n_184), .Y(n_721) );
NOR2xp67_ASAP7_75t_L g722 ( .A(n_584), .B(n_187), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_662), .B(n_189), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_590), .A2(n_191), .B1(n_192), .B2(n_193), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_582), .B(n_194), .Y(n_725) );
OAI21xp5_ASAP7_75t_L g726 ( .A1(n_623), .A2(n_196), .B(n_197), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_575), .Y(n_727) );
AOI21xp5_ASAP7_75t_SL g728 ( .A1(n_609), .A2(n_249), .B(n_210), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_576), .B(n_644), .Y(n_729) );
AOI221x1_ASAP7_75t_L g730 ( .A1(n_629), .A2(n_208), .B1(n_211), .B2(n_212), .C(n_213), .Y(n_730) );
OAI21xp5_ASAP7_75t_L g731 ( .A1(n_606), .A2(n_219), .B(n_220), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_585), .B(n_589), .Y(n_732) );
AO31x2_ASAP7_75t_L g733 ( .A1(n_657), .A2(n_221), .A3(n_222), .B(n_224), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_627), .A2(n_226), .B1(n_227), .B2(n_228), .Y(n_734) );
AO21x1_ASAP7_75t_L g735 ( .A1(n_637), .A2(n_233), .B(n_235), .Y(n_735) );
CKINVDCx5p33_ASAP7_75t_R g736 ( .A(n_611), .Y(n_736) );
INVx3_ASAP7_75t_L g737 ( .A(n_651), .Y(n_737) );
INVx5_ASAP7_75t_L g738 ( .A(n_636), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g739 ( .A1(n_577), .A2(n_236), .B(n_238), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g740 ( .A1(n_577), .A2(n_239), .B(n_240), .Y(n_740) );
OAI21xp5_ASAP7_75t_L g741 ( .A1(n_635), .A2(n_241), .B(n_244), .Y(n_741) );
NOR2xp33_ASAP7_75t_SL g742 ( .A(n_636), .B(n_245), .Y(n_742) );
AO22x2_ASAP7_75t_L g743 ( .A1(n_646), .A2(n_641), .B1(n_586), .B2(n_645), .Y(n_743) );
AND2x4_ASAP7_75t_L g744 ( .A(n_593), .B(n_663), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g745 ( .A1(n_615), .A2(n_619), .B(n_614), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_640), .A2(n_642), .B(n_598), .Y(n_746) );
NOR3xp33_ASAP7_75t_L g747 ( .A(n_661), .B(n_675), .C(n_669), .Y(n_747) );
NAND2xp5_ASAP7_75t_SL g748 ( .A(n_633), .B(n_625), .Y(n_748) );
NAND2xp33_ASAP7_75t_SL g749 ( .A(n_668), .B(n_616), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_600), .B(n_653), .Y(n_750) );
O2A1O1Ixp33_ASAP7_75t_L g751 ( .A1(n_581), .A2(n_666), .B(n_643), .C(n_638), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_672), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_580), .B(n_592), .Y(n_753) );
XNOR2xp5_ASAP7_75t_L g754 ( .A(n_656), .B(n_588), .Y(n_754) );
NAND3xp33_ASAP7_75t_L g755 ( .A(n_626), .B(n_630), .C(n_674), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_610), .B(n_594), .Y(n_756) );
AO21x1_ASAP7_75t_L g757 ( .A1(n_665), .A2(n_595), .B(n_573), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_602), .B(n_604), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_621), .B(n_622), .Y(n_759) );
BUFx2_ASAP7_75t_L g760 ( .A(n_631), .Y(n_760) );
AOI21xp5_ASAP7_75t_L g761 ( .A1(n_573), .A2(n_567), .B(n_583), .Y(n_761) );
AOI21xp5_ASAP7_75t_L g762 ( .A1(n_631), .A2(n_567), .B(n_583), .Y(n_762) );
OAI21xp5_ASAP7_75t_L g763 ( .A1(n_583), .A2(n_527), .B(n_552), .Y(n_763) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_567), .B(n_492), .Y(n_764) );
O2A1O1Ixp33_ASAP7_75t_SL g765 ( .A1(n_613), .A2(n_537), .B(n_599), .C(n_650), .Y(n_765) );
OAI22xp5_ASAP7_75t_L g766 ( .A1(n_567), .A2(n_624), .B1(n_488), .B2(n_524), .Y(n_766) );
AOI21xp5_ASAP7_75t_L g767 ( .A1(n_567), .A2(n_583), .B(n_533), .Y(n_767) );
AND2x2_ASAP7_75t_L g768 ( .A(n_567), .B(n_578), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_567), .B(n_583), .Y(n_769) );
OAI21x1_ASAP7_75t_L g770 ( .A1(n_652), .A2(n_534), .B(n_529), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_567), .B(n_583), .Y(n_771) );
BUFx2_ASAP7_75t_R g772 ( .A(n_587), .Y(n_772) );
AOI21xp5_ASAP7_75t_L g773 ( .A1(n_567), .A2(n_583), .B(n_533), .Y(n_773) );
OAI22xp5_ASAP7_75t_L g774 ( .A1(n_567), .A2(n_624), .B1(n_488), .B2(n_524), .Y(n_774) );
BUFx4f_ASAP7_75t_L g775 ( .A(n_587), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_567), .Y(n_776) );
AOI21xp5_ASAP7_75t_L g777 ( .A1(n_567), .A2(n_583), .B(n_533), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_567), .Y(n_778) );
CKINVDCx6p67_ASAP7_75t_R g779 ( .A(n_648), .Y(n_779) );
OAI21xp5_ASAP7_75t_L g780 ( .A1(n_583), .A2(n_527), .B(n_552), .Y(n_780) );
INVx2_ASAP7_75t_SL g781 ( .A(n_648), .Y(n_781) );
AND2x2_ASAP7_75t_L g782 ( .A(n_567), .B(n_578), .Y(n_782) );
INVx5_ASAP7_75t_L g783 ( .A(n_647), .Y(n_783) );
AOI21xp5_ASAP7_75t_L g784 ( .A1(n_567), .A2(n_583), .B(n_533), .Y(n_784) );
BUFx6f_ASAP7_75t_L g785 ( .A(n_634), .Y(n_785) );
OAI22xp5_ASAP7_75t_L g786 ( .A1(n_567), .A2(n_624), .B1(n_488), .B2(n_524), .Y(n_786) );
AOI21xp5_ASAP7_75t_L g787 ( .A1(n_567), .A2(n_583), .B(n_533), .Y(n_787) );
AND2x2_ASAP7_75t_L g788 ( .A(n_567), .B(n_578), .Y(n_788) );
AOI221x1_ASAP7_75t_L g789 ( .A1(n_608), .A2(n_612), .B1(n_655), .B2(n_629), .C(n_646), .Y(n_789) );
AND2x2_ASAP7_75t_L g790 ( .A(n_567), .B(n_578), .Y(n_790) );
HB1xp67_ASAP7_75t_L g791 ( .A(n_658), .Y(n_791) );
AND2x2_ASAP7_75t_L g792 ( .A(n_567), .B(n_578), .Y(n_792) );
BUFx3_ASAP7_75t_L g793 ( .A(n_587), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_567), .B(n_583), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_567), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_567), .Y(n_796) );
BUFx6f_ASAP7_75t_L g797 ( .A(n_634), .Y(n_797) );
OAI21xp5_ASAP7_75t_L g798 ( .A1(n_567), .A2(n_527), .B(n_583), .Y(n_798) );
INVx2_ASAP7_75t_SL g799 ( .A(n_648), .Y(n_799) );
OR2x6_ASAP7_75t_L g800 ( .A(n_647), .B(n_512), .Y(n_800) );
INVx4_ASAP7_75t_L g801 ( .A(n_658), .Y(n_801) );
A2O1A1Ixp33_ASAP7_75t_L g802 ( .A1(n_567), .A2(n_603), .B(n_583), .C(n_506), .Y(n_802) );
NAND2xp33_ASAP7_75t_R g803 ( .A(n_671), .B(n_450), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_567), .B(n_583), .Y(n_804) );
AND2x2_ASAP7_75t_SL g805 ( .A(n_618), .B(n_522), .Y(n_805) );
AOI21xp5_ASAP7_75t_L g806 ( .A1(n_567), .A2(n_583), .B(n_533), .Y(n_806) );
INVx2_ASAP7_75t_L g807 ( .A(n_679), .Y(n_807) );
OA21x2_ASAP7_75t_L g808 ( .A1(n_761), .A2(n_789), .B(n_770), .Y(n_808) );
NAND2x1p5_ASAP7_75t_L g809 ( .A(n_738), .B(n_783), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g810 ( .A(n_764), .B(n_769), .Y(n_810) );
INVx1_ASAP7_75t_SL g811 ( .A(n_676), .Y(n_811) );
BUFx3_ASAP7_75t_L g812 ( .A(n_692), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_768), .Y(n_813) );
BUFx4f_ASAP7_75t_SL g814 ( .A(n_779), .Y(n_814) );
HB1xp67_ASAP7_75t_L g815 ( .A(n_677), .Y(n_815) );
A2O1A1Ixp33_ASAP7_75t_L g816 ( .A1(n_751), .A2(n_802), .B(n_762), .C(n_759), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_782), .Y(n_817) );
NAND2xp5_ASAP7_75t_SL g818 ( .A(n_742), .B(n_696), .Y(n_818) );
AO31x2_ASAP7_75t_L g819 ( .A1(n_757), .A2(n_701), .A3(n_705), .B(n_735), .Y(n_819) );
INVx5_ASAP7_75t_SL g820 ( .A(n_800), .Y(n_820) );
AND2x2_ASAP7_75t_L g821 ( .A(n_788), .B(n_790), .Y(n_821) );
HB1xp67_ASAP7_75t_L g822 ( .A(n_760), .Y(n_822) );
AOI21xp5_ASAP7_75t_SL g823 ( .A1(n_696), .A2(n_774), .B(n_766), .Y(n_823) );
OR2x6_ASAP7_75t_L g824 ( .A(n_800), .B(n_793), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_795), .B(n_796), .Y(n_825) );
INVx3_ASAP7_75t_L g826 ( .A(n_801), .Y(n_826) );
AO31x2_ASAP7_75t_L g827 ( .A1(n_730), .A2(n_739), .A3(n_740), .B(n_746), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_771), .B(n_794), .Y(n_828) );
OAI21xp5_ASAP7_75t_L g829 ( .A1(n_767), .A2(n_777), .B(n_773), .Y(n_829) );
NAND2x1p5_ASAP7_75t_L g830 ( .A(n_738), .B(n_783), .Y(n_830) );
AND2x4_ASAP7_75t_L g831 ( .A(n_804), .B(n_738), .Y(n_831) );
INVx3_ASAP7_75t_L g832 ( .A(n_801), .Y(n_832) );
OA21x2_ASAP7_75t_L g833 ( .A1(n_731), .A2(n_717), .B(n_726), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_792), .Y(n_834) );
AND2x4_ASAP7_75t_L g835 ( .A(n_783), .B(n_800), .Y(n_835) );
OAI21xp5_ASAP7_75t_L g836 ( .A1(n_784), .A2(n_806), .B(n_787), .Y(n_836) );
HB1xp67_ASAP7_75t_L g837 ( .A(n_791), .Y(n_837) );
AO21x2_ASAP7_75t_L g838 ( .A1(n_741), .A2(n_763), .B(n_780), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_805), .A2(n_786), .B1(n_754), .B2(n_763), .Y(n_839) );
OR2x2_ASAP7_75t_L g840 ( .A(n_729), .B(n_694), .Y(n_840) );
OAI21x1_ASAP7_75t_SL g841 ( .A1(n_709), .A2(n_780), .B(n_734), .Y(n_841) );
BUFx2_ASAP7_75t_R g842 ( .A(n_706), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_707), .B(n_727), .Y(n_843) );
NAND3xp33_ASAP7_75t_L g844 ( .A(n_691), .B(n_747), .C(n_678), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_752), .B(n_750), .Y(n_845) );
HB1xp67_ASAP7_75t_L g846 ( .A(n_684), .Y(n_846) );
AO31x2_ASAP7_75t_L g847 ( .A1(n_716), .A2(n_703), .A3(n_681), .B(n_698), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_682), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_732), .B(n_756), .Y(n_849) );
AOI21xp5_ASAP7_75t_L g850 ( .A1(n_765), .A2(n_725), .B(n_700), .Y(n_850) );
OAI21x1_ASAP7_75t_SL g851 ( .A1(n_709), .A2(n_745), .B(n_713), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_753), .B(n_758), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_699), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_743), .B(n_723), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_743), .B(n_749), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_755), .B(n_688), .Y(n_856) );
BUFx2_ASAP7_75t_L g857 ( .A(n_775), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_699), .Y(n_858) );
AND2x4_ASAP7_75t_L g859 ( .A(n_720), .B(n_737), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_755), .B(n_704), .Y(n_860) );
OAI21x1_ASAP7_75t_SL g861 ( .A1(n_724), .A2(n_712), .B(n_728), .Y(n_861) );
AOI21xp33_ASAP7_75t_L g862 ( .A1(n_691), .A2(n_748), .B(n_683), .Y(n_862) );
INVxp67_ASAP7_75t_L g863 ( .A(n_685), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_687), .Y(n_864) );
AOI21xp5_ASAP7_75t_L g865 ( .A1(n_689), .A2(n_710), .B(n_797), .Y(n_865) );
BUFx3_ASAP7_75t_L g866 ( .A(n_775), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_697), .Y(n_867) );
BUFx2_ASAP7_75t_R g868 ( .A(n_736), .Y(n_868) );
OAI21x1_ASAP7_75t_L g869 ( .A1(n_722), .A2(n_715), .B(n_680), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_702), .Y(n_870) );
BUFx2_ASAP7_75t_SL g871 ( .A(n_690), .Y(n_871) );
OR2x2_ASAP7_75t_L g872 ( .A(n_708), .B(n_693), .Y(n_872) );
AND2x2_ASAP7_75t_L g873 ( .A(n_714), .B(n_711), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_744), .A2(n_719), .B1(n_714), .B2(n_718), .Y(n_874) );
NOR2x1_ASAP7_75t_SL g875 ( .A(n_785), .B(n_772), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_686), .A2(n_781), .B1(n_799), .B2(n_733), .Y(n_876) );
AND2x2_ASAP7_75t_L g877 ( .A(n_733), .B(n_721), .Y(n_877) );
INVx5_ASAP7_75t_L g878 ( .A(n_803), .Y(n_878) );
AO222x2_ASAP7_75t_L g879 ( .A1(n_721), .A2(n_481), .B1(n_611), .B2(n_617), .C1(n_779), .C2(n_480), .Y(n_879) );
OAI21xp5_ASAP7_75t_L g880 ( .A1(n_721), .A2(n_761), .B(n_802), .Y(n_880) );
OA21x2_ASAP7_75t_L g881 ( .A1(n_761), .A2(n_789), .B(n_770), .Y(n_881) );
O2A1O1Ixp33_ASAP7_75t_L g882 ( .A1(n_802), .A2(n_683), .B(n_666), .C(n_657), .Y(n_882) );
OA21x2_ASAP7_75t_L g883 ( .A1(n_761), .A2(n_789), .B(n_770), .Y(n_883) );
AOI21xp5_ASAP7_75t_L g884 ( .A1(n_746), .A2(n_761), .B(n_767), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_747), .A2(n_805), .B1(n_596), .B2(n_707), .Y(n_885) );
BUFx3_ASAP7_75t_L g886 ( .A(n_692), .Y(n_886) );
NAND2x1p5_ASAP7_75t_L g887 ( .A(n_738), .B(n_783), .Y(n_887) );
OAI21xp5_ASAP7_75t_L g888 ( .A1(n_761), .A2(n_802), .B(n_773), .Y(n_888) );
NAND2x1p5_ASAP7_75t_L g889 ( .A(n_738), .B(n_783), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_768), .B(n_782), .Y(n_890) );
AND2x2_ASAP7_75t_L g891 ( .A(n_768), .B(n_782), .Y(n_891) );
CKINVDCx6p67_ASAP7_75t_R g892 ( .A(n_692), .Y(n_892) );
OA21x2_ASAP7_75t_L g893 ( .A1(n_761), .A2(n_789), .B(n_770), .Y(n_893) );
AND2x4_ASAP7_75t_L g894 ( .A(n_776), .B(n_778), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_768), .Y(n_895) );
OAI21xp5_ASAP7_75t_L g896 ( .A1(n_761), .A2(n_802), .B(n_773), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_768), .Y(n_897) );
OAI21x1_ASAP7_75t_SL g898 ( .A1(n_696), .A2(n_695), .B(n_798), .Y(n_898) );
OAI21xp5_ASAP7_75t_L g899 ( .A1(n_761), .A2(n_802), .B(n_773), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_776), .B(n_778), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_776), .B(n_778), .Y(n_901) );
OAI21xp5_ASAP7_75t_L g902 ( .A1(n_761), .A2(n_802), .B(n_773), .Y(n_902) );
OAI21xp5_ASAP7_75t_L g903 ( .A1(n_761), .A2(n_802), .B(n_773), .Y(n_903) );
BUFx2_ASAP7_75t_L g904 ( .A(n_692), .Y(n_904) );
BUFx3_ASAP7_75t_L g905 ( .A(n_692), .Y(n_905) );
AND2x6_ASAP7_75t_L g906 ( .A(n_684), .B(n_618), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_768), .Y(n_907) );
AND2x2_ASAP7_75t_L g908 ( .A(n_768), .B(n_782), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_768), .B(n_782), .Y(n_909) );
AND2x2_ASAP7_75t_L g910 ( .A(n_821), .B(n_890), .Y(n_910) );
OR2x6_ASAP7_75t_L g911 ( .A(n_823), .B(n_809), .Y(n_911) );
BUFx2_ASAP7_75t_L g912 ( .A(n_906), .Y(n_912) );
HB1xp67_ASAP7_75t_L g913 ( .A(n_891), .Y(n_913) );
AND2x2_ASAP7_75t_L g914 ( .A(n_908), .B(n_909), .Y(n_914) );
AND2x2_ASAP7_75t_L g915 ( .A(n_828), .B(n_894), .Y(n_915) );
AND2x4_ASAP7_75t_L g916 ( .A(n_831), .B(n_835), .Y(n_916) );
AND2x2_ASAP7_75t_L g917 ( .A(n_828), .B(n_810), .Y(n_917) );
AND2x2_ASAP7_75t_L g918 ( .A(n_810), .B(n_807), .Y(n_918) );
INVx3_ASAP7_75t_L g919 ( .A(n_906), .Y(n_919) );
INVx2_ASAP7_75t_SL g920 ( .A(n_904), .Y(n_920) );
BUFx3_ASAP7_75t_L g921 ( .A(n_812), .Y(n_921) );
HB1xp67_ASAP7_75t_L g922 ( .A(n_822), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_864), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_825), .Y(n_924) );
OR2x2_ASAP7_75t_L g925 ( .A(n_840), .B(n_845), .Y(n_925) );
AO21x2_ASAP7_75t_L g926 ( .A1(n_880), .A2(n_884), .B(n_888), .Y(n_926) );
HB1xp67_ASAP7_75t_L g927 ( .A(n_822), .Y(n_927) );
BUFx2_ASAP7_75t_L g928 ( .A(n_906), .Y(n_928) );
BUFx3_ASAP7_75t_L g929 ( .A(n_886), .Y(n_929) );
AO21x2_ASAP7_75t_L g930 ( .A1(n_880), .A2(n_884), .B(n_888), .Y(n_930) );
INVx5_ASAP7_75t_L g931 ( .A(n_906), .Y(n_931) );
NOR2xp33_ASAP7_75t_L g932 ( .A(n_879), .B(n_852), .Y(n_932) );
HB1xp67_ASAP7_75t_L g933 ( .A(n_900), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_853), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_858), .Y(n_935) );
AO21x2_ASAP7_75t_L g936 ( .A1(n_896), .A2(n_902), .B(n_899), .Y(n_936) );
HB1xp67_ASAP7_75t_L g937 ( .A(n_901), .Y(n_937) );
BUFx3_ASAP7_75t_L g938 ( .A(n_905), .Y(n_938) );
AND2x2_ASAP7_75t_L g939 ( .A(n_845), .B(n_813), .Y(n_939) );
AND2x2_ASAP7_75t_L g940 ( .A(n_817), .B(n_834), .Y(n_940) );
INVxp67_ASAP7_75t_L g941 ( .A(n_857), .Y(n_941) );
AO21x2_ASAP7_75t_L g942 ( .A1(n_896), .A2(n_899), .B(n_902), .Y(n_942) );
AO21x1_ASAP7_75t_L g943 ( .A1(n_839), .A2(n_818), .B(n_855), .Y(n_943) );
BUFx3_ASAP7_75t_L g944 ( .A(n_892), .Y(n_944) );
AO31x2_ASAP7_75t_L g945 ( .A1(n_816), .A2(n_867), .A3(n_856), .B(n_855), .Y(n_945) );
BUFx3_ASAP7_75t_L g946 ( .A(n_866), .Y(n_946) );
NOR2xp67_ASAP7_75t_L g947 ( .A(n_878), .B(n_874), .Y(n_947) );
BUFx2_ASAP7_75t_L g948 ( .A(n_846), .Y(n_948) );
AO21x2_ASAP7_75t_L g949 ( .A1(n_903), .A2(n_818), .B(n_829), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_895), .B(n_897), .Y(n_950) );
INVx3_ASAP7_75t_L g951 ( .A(n_809), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_907), .Y(n_952) );
CKINVDCx10_ASAP7_75t_R g953 ( .A(n_824), .Y(n_953) );
AO21x2_ASAP7_75t_L g954 ( .A1(n_829), .A2(n_836), .B(n_841), .Y(n_954) );
HB1xp67_ASAP7_75t_L g955 ( .A(n_837), .Y(n_955) );
INVx3_ASAP7_75t_L g956 ( .A(n_830), .Y(n_956) );
INVx3_ASAP7_75t_L g957 ( .A(n_830), .Y(n_957) );
AO21x2_ASAP7_75t_L g958 ( .A1(n_836), .A2(n_877), .B(n_898), .Y(n_958) );
NAND2x1_ASAP7_75t_L g959 ( .A(n_851), .B(n_861), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_843), .Y(n_960) );
INVx2_ASAP7_75t_SL g961 ( .A(n_824), .Y(n_961) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_849), .B(n_885), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_849), .B(n_885), .Y(n_963) );
OR2x2_ASAP7_75t_L g964 ( .A(n_854), .B(n_815), .Y(n_964) );
OAI21xp5_ASAP7_75t_L g965 ( .A1(n_844), .A2(n_882), .B(n_862), .Y(n_965) );
INVx2_ASAP7_75t_SL g966 ( .A(n_878), .Y(n_966) );
OA21x2_ASAP7_75t_L g967 ( .A1(n_850), .A2(n_865), .B(n_860), .Y(n_967) );
INVx2_ASAP7_75t_SL g968 ( .A(n_931), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_934), .Y(n_969) );
INVx3_ASAP7_75t_SL g970 ( .A(n_931), .Y(n_970) );
INVx4_ASAP7_75t_L g971 ( .A(n_931), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_960), .B(n_848), .Y(n_972) );
AND2x2_ASAP7_75t_L g973 ( .A(n_915), .B(n_838), .Y(n_973) );
AND2x2_ASAP7_75t_L g974 ( .A(n_915), .B(n_808), .Y(n_974) );
OAI22xp5_ASAP7_75t_L g975 ( .A1(n_933), .A2(n_876), .B1(n_820), .B2(n_870), .Y(n_975) );
NAND2x1p5_ASAP7_75t_L g976 ( .A(n_931), .B(n_826), .Y(n_976) );
AND2x2_ASAP7_75t_L g977 ( .A(n_917), .B(n_893), .Y(n_977) );
OR2x2_ASAP7_75t_L g978 ( .A(n_964), .B(n_876), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_935), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_923), .Y(n_980) );
AND2x2_ASAP7_75t_L g981 ( .A(n_917), .B(n_910), .Y(n_981) );
OAI221xp5_ASAP7_75t_L g982 ( .A1(n_932), .A2(n_882), .B1(n_874), .B2(n_811), .C(n_863), .Y(n_982) );
NOR2x1_ASAP7_75t_L g983 ( .A(n_947), .B(n_832), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_910), .B(n_893), .Y(n_984) );
BUFx3_ASAP7_75t_L g985 ( .A(n_931), .Y(n_985) );
AND2x2_ASAP7_75t_L g986 ( .A(n_914), .B(n_881), .Y(n_986) );
AND2x4_ASAP7_75t_L g987 ( .A(n_911), .B(n_875), .Y(n_987) );
NOR2xp33_ASAP7_75t_L g988 ( .A(n_925), .B(n_872), .Y(n_988) );
AND2x4_ASAP7_75t_L g989 ( .A(n_911), .B(n_869), .Y(n_989) );
AND2x2_ASAP7_75t_L g990 ( .A(n_914), .B(n_939), .Y(n_990) );
HB1xp67_ASAP7_75t_L g991 ( .A(n_937), .Y(n_991) );
AND2x2_ASAP7_75t_L g992 ( .A(n_939), .B(n_883), .Y(n_992) );
HB1xp67_ASAP7_75t_L g993 ( .A(n_913), .Y(n_993) );
AND2x2_ASAP7_75t_L g994 ( .A(n_918), .B(n_881), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_936), .B(n_847), .Y(n_995) );
AND2x2_ASAP7_75t_L g996 ( .A(n_936), .B(n_847), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_962), .A2(n_820), .B1(n_878), .B2(n_859), .Y(n_997) );
AND2x2_ASAP7_75t_L g998 ( .A(n_942), .B(n_819), .Y(n_998) );
AND2x2_ASAP7_75t_L g999 ( .A(n_942), .B(n_819), .Y(n_999) );
INVxp67_ASAP7_75t_L g1000 ( .A(n_948), .Y(n_1000) );
AOI222xp33_ASAP7_75t_L g1001 ( .A1(n_963), .A2(n_814), .B1(n_878), .B2(n_859), .C1(n_873), .C2(n_842), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_942), .B(n_819), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_945), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_945), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_954), .B(n_833), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_924), .B(n_827), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_945), .B(n_889), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1008 ( .A(n_945), .B(n_889), .Y(n_1008) );
AND2x2_ASAP7_75t_L g1009 ( .A(n_945), .B(n_887), .Y(n_1009) );
HB1xp67_ASAP7_75t_L g1010 ( .A(n_955), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_990), .B(n_940), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_984), .B(n_958), .Y(n_1012) );
CKINVDCx14_ASAP7_75t_R g1013 ( .A(n_990), .Y(n_1013) );
NOR2xp67_ASAP7_75t_L g1014 ( .A(n_971), .B(n_966), .Y(n_1014) );
BUFx3_ASAP7_75t_L g1015 ( .A(n_970), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_984), .B(n_958), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_986), .B(n_958), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_969), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_986), .B(n_949), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g1020 ( .A(n_981), .B(n_993), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_969), .Y(n_1021) );
AND2x2_ASAP7_75t_L g1022 ( .A(n_973), .B(n_949), .Y(n_1022) );
BUFx2_ASAP7_75t_SL g1023 ( .A(n_971), .Y(n_1023) );
INVx3_ASAP7_75t_L g1024 ( .A(n_989), .Y(n_1024) );
AND2x2_ASAP7_75t_L g1025 ( .A(n_977), .B(n_949), .Y(n_1025) );
AND2x4_ASAP7_75t_L g1026 ( .A(n_989), .B(n_926), .Y(n_1026) );
INVx3_ASAP7_75t_L g1027 ( .A(n_989), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_977), .B(n_926), .Y(n_1028) );
AND2x2_ASAP7_75t_L g1029 ( .A(n_974), .B(n_930), .Y(n_1029) );
NAND2x1p5_ASAP7_75t_L g1030 ( .A(n_971), .B(n_912), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_974), .B(n_930), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_992), .B(n_930), .Y(n_1032) );
NAND2xp5_ASAP7_75t_L g1033 ( .A(n_981), .B(n_940), .Y(n_1033) );
INVxp67_ASAP7_75t_SL g1034 ( .A(n_991), .Y(n_1034) );
OR2x2_ASAP7_75t_L g1035 ( .A(n_978), .B(n_922), .Y(n_1035) );
OR2x2_ASAP7_75t_L g1036 ( .A(n_978), .B(n_994), .Y(n_1036) );
OR2x2_ASAP7_75t_L g1037 ( .A(n_994), .B(n_927), .Y(n_1037) );
INVx3_ASAP7_75t_L g1038 ( .A(n_971), .Y(n_1038) );
BUFx2_ASAP7_75t_SL g1039 ( .A(n_985), .Y(n_1039) );
NOR2x1_ASAP7_75t_L g1040 ( .A(n_985), .B(n_911), .Y(n_1040) );
AND2x4_ASAP7_75t_SL g1041 ( .A(n_987), .B(n_919), .Y(n_1041) );
BUFx2_ASAP7_75t_L g1042 ( .A(n_1000), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_1010), .B(n_950), .Y(n_1043) );
AND2x4_ASAP7_75t_L g1044 ( .A(n_995), .B(n_996), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_979), .B(n_967), .Y(n_1045) );
OR2x2_ASAP7_75t_L g1046 ( .A(n_1036), .B(n_1006), .Y(n_1046) );
INVx1_ASAP7_75t_L g1047 ( .A(n_1018), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1018), .Y(n_1048) );
OR2x2_ASAP7_75t_L g1049 ( .A(n_1036), .B(n_1006), .Y(n_1049) );
OR2x2_ASAP7_75t_L g1050 ( .A(n_1037), .B(n_1003), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1021), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_1044), .B(n_1005), .Y(n_1052) );
AND2x4_ASAP7_75t_L g1053 ( .A(n_1024), .B(n_998), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_1044), .B(n_998), .Y(n_1054) );
NAND2xp5_ASAP7_75t_L g1055 ( .A(n_1013), .B(n_972), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_1044), .B(n_999), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_1029), .B(n_999), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_1029), .B(n_1002), .Y(n_1058) );
OR2x2_ASAP7_75t_L g1059 ( .A(n_1035), .B(n_1004), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_1031), .B(n_1002), .Y(n_1060) );
AND2x2_ASAP7_75t_L g1061 ( .A(n_1031), .B(n_1007), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_1012), .B(n_1008), .Y(n_1062) );
OR2x2_ASAP7_75t_L g1063 ( .A(n_1035), .B(n_1004), .Y(n_1063) );
INVx1_ASAP7_75t_SL g1064 ( .A(n_1020), .Y(n_1064) );
AND2x2_ASAP7_75t_L g1065 ( .A(n_1012), .B(n_1008), .Y(n_1065) );
OR2x6_ASAP7_75t_L g1066 ( .A(n_1023), .B(n_959), .Y(n_1066) );
INVxp67_ASAP7_75t_SL g1067 ( .A(n_1014), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_1016), .B(n_1009), .Y(n_1068) );
AND3x1_ASAP7_75t_L g1069 ( .A(n_1040), .B(n_953), .C(n_814), .Y(n_1069) );
NOR2xp33_ASAP7_75t_L g1070 ( .A(n_1043), .B(n_921), .Y(n_1070) );
NAND2xp5_ASAP7_75t_L g1071 ( .A(n_1034), .B(n_980), .Y(n_1071) );
INVxp33_ASAP7_75t_L g1072 ( .A(n_1070), .Y(n_1072) );
NAND2xp5_ASAP7_75t_L g1073 ( .A(n_1057), .B(n_1022), .Y(n_1073) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_1057), .B(n_1028), .Y(n_1074) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1047), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1058), .B(n_1028), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_1058), .B(n_1032), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_1060), .B(n_1022), .Y(n_1078) );
NAND2xp5_ASAP7_75t_L g1079 ( .A(n_1060), .B(n_1019), .Y(n_1079) );
INVx4_ASAP7_75t_L g1080 ( .A(n_1066), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_1062), .B(n_1032), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1048), .Y(n_1082) );
AND2x4_ASAP7_75t_L g1083 ( .A(n_1053), .B(n_1026), .Y(n_1083) );
HB1xp67_ASAP7_75t_L g1084 ( .A(n_1064), .Y(n_1084) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_1062), .B(n_1016), .Y(n_1085) );
NAND2x1p5_ASAP7_75t_L g1086 ( .A(n_1069), .B(n_1040), .Y(n_1086) );
INVx1_ASAP7_75t_SL g1087 ( .A(n_1055), .Y(n_1087) );
BUFx2_ASAP7_75t_L g1088 ( .A(n_1067), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_1065), .B(n_1017), .Y(n_1089) );
AND2x2_ASAP7_75t_L g1090 ( .A(n_1065), .B(n_1017), .Y(n_1090) );
AND2x4_ASAP7_75t_L g1091 ( .A(n_1053), .B(n_1026), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_1068), .B(n_1025), .Y(n_1092) );
AND2x4_ASAP7_75t_SL g1093 ( .A(n_1066), .B(n_1038), .Y(n_1093) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1051), .Y(n_1094) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_1068), .B(n_1025), .Y(n_1095) );
NAND2xp5_ASAP7_75t_L g1096 ( .A(n_1046), .B(n_1045), .Y(n_1096) );
INVxp67_ASAP7_75t_L g1097 ( .A(n_1084), .Y(n_1097) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1075), .Y(n_1098) );
NOR2xp33_ASAP7_75t_L g1099 ( .A(n_1072), .B(n_1087), .Y(n_1099) );
INVxp67_ASAP7_75t_L g1100 ( .A(n_1088), .Y(n_1100) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1075), .Y(n_1101) );
NAND2xp5_ASAP7_75t_L g1102 ( .A(n_1074), .B(n_1061), .Y(n_1102) );
OR2x2_ASAP7_75t_L g1103 ( .A(n_1096), .B(n_1046), .Y(n_1103) );
NAND2xp5_ASAP7_75t_L g1104 ( .A(n_1074), .B(n_1061), .Y(n_1104) );
NAND2xp5_ASAP7_75t_L g1105 ( .A(n_1076), .B(n_1054), .Y(n_1105) );
INVx2_ASAP7_75t_SL g1106 ( .A(n_1093), .Y(n_1106) );
NAND2xp5_ASAP7_75t_L g1107 ( .A(n_1076), .B(n_1054), .Y(n_1107) );
AOI21xp33_ASAP7_75t_SL g1108 ( .A1(n_1086), .A2(n_1001), .B(n_970), .Y(n_1108) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_1077), .B(n_1056), .Y(n_1109) );
OAI322xp33_ASAP7_75t_L g1110 ( .A1(n_1087), .A2(n_1049), .A3(n_1071), .B1(n_1033), .B2(n_1011), .C1(n_1063), .C2(n_1059), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g1111 ( .A(n_1077), .B(n_1056), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_1081), .B(n_1052), .Y(n_1112) );
INVxp33_ASAP7_75t_L g1113 ( .A(n_1080), .Y(n_1113) );
OAI21xp5_ASAP7_75t_L g1114 ( .A1(n_1088), .A2(n_975), .B(n_982), .Y(n_1114) );
OAI22xp5_ASAP7_75t_L g1115 ( .A1(n_1080), .A2(n_1066), .B1(n_1049), .B2(n_1039), .Y(n_1115) );
OR2x2_ASAP7_75t_L g1116 ( .A(n_1096), .B(n_1050), .Y(n_1116) );
AO32x1_ASAP7_75t_L g1117 ( .A1(n_1115), .A2(n_1080), .A3(n_1093), .B1(n_961), .B2(n_968), .Y(n_1117) );
AOI211xp5_ASAP7_75t_SL g1118 ( .A1(n_1110), .A2(n_987), .B(n_1038), .C(n_1027), .Y(n_1118) );
OAI22x1_ASAP7_75t_L g1119 ( .A1(n_1100), .A2(n_1038), .B1(n_1091), .B2(n_1083), .Y(n_1119) );
OAI322xp33_ASAP7_75t_L g1120 ( .A1(n_1097), .A2(n_1078), .A3(n_1073), .B1(n_1079), .B2(n_1063), .C1(n_1059), .C2(n_1050), .Y(n_1120) );
O2A1O1Ixp33_ASAP7_75t_L g1121 ( .A1(n_1097), .A2(n_1100), .B(n_1099), .C(n_1108), .Y(n_1121) );
INVxp67_ASAP7_75t_L g1122 ( .A(n_1099), .Y(n_1122) );
O2A1O1Ixp33_ASAP7_75t_L g1123 ( .A1(n_1114), .A2(n_944), .B(n_965), .C(n_920), .Y(n_1123) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1098), .Y(n_1124) );
INVx2_ASAP7_75t_SL g1125 ( .A(n_1106), .Y(n_1125) );
OAI21xp5_ASAP7_75t_SL g1126 ( .A1(n_1113), .A2(n_987), .B(n_1041), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_1112), .B(n_1081), .Y(n_1127) );
OAI221xp5_ASAP7_75t_L g1128 ( .A1(n_1113), .A2(n_997), .B1(n_1024), .B2(n_1027), .C(n_1094), .Y(n_1128) );
AOI22xp5_ASAP7_75t_L g1129 ( .A1(n_1103), .A2(n_1083), .B1(n_1091), .B2(n_1053), .Y(n_1129) );
AOI21xp33_ASAP7_75t_L g1130 ( .A1(n_1101), .A2(n_920), .B(n_988), .Y(n_1130) );
OAI22xp5_ASAP7_75t_SL g1131 ( .A1(n_1102), .A2(n_944), .B1(n_871), .B2(n_987), .Y(n_1131) );
AOI21xp33_ASAP7_75t_L g1132 ( .A1(n_1123), .A2(n_941), .B(n_938), .Y(n_1132) );
AOI21xp33_ASAP7_75t_SL g1133 ( .A1(n_1121), .A2(n_970), .B(n_1030), .Y(n_1133) );
OAI21xp5_ASAP7_75t_L g1134 ( .A1(n_1118), .A2(n_1104), .B(n_1116), .Y(n_1134) );
HAxp5_ASAP7_75t_SL g1135 ( .A(n_1129), .B(n_842), .CON(n_1135), .SN(n_1135) );
NOR2xp67_ASAP7_75t_L g1136 ( .A(n_1119), .B(n_1083), .Y(n_1136) );
NAND2xp5_ASAP7_75t_L g1137 ( .A(n_1122), .B(n_1092), .Y(n_1137) );
AOI21xp5_ASAP7_75t_L g1138 ( .A1(n_1117), .A2(n_1066), .B(n_1091), .Y(n_1138) );
AOI322xp5_ASAP7_75t_L g1139 ( .A1(n_1125), .A2(n_1090), .A3(n_1089), .B1(n_1085), .B2(n_1092), .C1(n_1095), .C2(n_1111), .Y(n_1139) );
AOI221xp5_ASAP7_75t_L g1140 ( .A1(n_1120), .A2(n_1109), .B1(n_1107), .B2(n_1105), .C(n_1095), .Y(n_1140) );
OAI221xp5_ASAP7_75t_L g1141 ( .A1(n_1131), .A2(n_1126), .B1(n_1128), .B2(n_1130), .C(n_1124), .Y(n_1141) );
NAND3xp33_ASAP7_75t_L g1142 ( .A(n_1135), .B(n_938), .C(n_929), .Y(n_1142) );
NOR4xp25_ASAP7_75t_SL g1143 ( .A(n_1141), .B(n_1117), .C(n_1042), .D(n_928), .Y(n_1143) );
NOR3xp33_ASAP7_75t_L g1144 ( .A(n_1133), .B(n_946), .C(n_868), .Y(n_1144) );
NOR2x1_ASAP7_75t_L g1145 ( .A(n_1136), .B(n_946), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1134), .B(n_1127), .Y(n_1146) );
NOR3xp33_ASAP7_75t_L g1147 ( .A(n_1132), .B(n_966), .C(n_956), .Y(n_1147) );
AOI211xp5_ASAP7_75t_L g1148 ( .A1(n_1138), .A2(n_943), .B(n_1015), .C(n_1009), .Y(n_1148) );
NOR2xp33_ASAP7_75t_L g1149 ( .A(n_1137), .B(n_1082), .Y(n_1149) );
NAND5xp2_ASAP7_75t_L g1150 ( .A(n_1148), .B(n_1139), .C(n_1140), .D(n_1030), .E(n_976), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1149), .Y(n_1151) );
INVx2_ASAP7_75t_L g1152 ( .A(n_1146), .Y(n_1152) );
INVx3_ASAP7_75t_L g1153 ( .A(n_1145), .Y(n_1153) );
HB1xp67_ASAP7_75t_L g1154 ( .A(n_1142), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1152), .Y(n_1155) );
NAND4xp25_ASAP7_75t_L g1156 ( .A(n_1150), .B(n_1144), .C(n_1147), .D(n_1143), .Y(n_1156) );
AND2x4_ASAP7_75t_L g1157 ( .A(n_1154), .B(n_1052), .Y(n_1157) );
INVx3_ASAP7_75t_L g1158 ( .A(n_1155), .Y(n_1158) );
INVxp67_ASAP7_75t_SL g1159 ( .A(n_1157), .Y(n_1159) );
NOR2xp33_ASAP7_75t_L g1160 ( .A(n_1156), .B(n_1151), .Y(n_1160) );
NOR3xp33_ASAP7_75t_L g1161 ( .A(n_1160), .B(n_1153), .C(n_956), .Y(n_1161) );
INVxp67_ASAP7_75t_L g1162 ( .A(n_1158), .Y(n_1162) );
AOI22x1_ASAP7_75t_L g1163 ( .A1(n_1162), .A2(n_1158), .B1(n_1159), .B2(n_956), .Y(n_1163) );
OAI22xp5_ASAP7_75t_L g1164 ( .A1(n_1163), .A2(n_1161), .B1(n_968), .B2(n_1015), .Y(n_1164) );
AOI22xp5_ASAP7_75t_L g1165 ( .A1(n_1164), .A2(n_957), .B1(n_951), .B2(n_916), .Y(n_1165) );
NAND2x1p5_ASAP7_75t_SL g1166 ( .A(n_1165), .B(n_983), .Y(n_1166) );
OR2x2_ASAP7_75t_L g1167 ( .A(n_1166), .B(n_1042), .Y(n_1167) );
AOI21xp33_ASAP7_75t_SL g1168 ( .A1(n_1167), .A2(n_976), .B(n_952), .Y(n_1168) );
endmodule