module fake_aes_7932_n_31 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_31);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_31;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g9 ( .A(n_7), .Y(n_9) );
CKINVDCx20_ASAP7_75t_R g10 ( .A(n_4), .Y(n_10) );
INVx2_ASAP7_75t_SL g11 ( .A(n_6), .Y(n_11) );
NAND2x1_ASAP7_75t_L g12 ( .A(n_5), .B(n_0), .Y(n_12) );
BUFx6f_ASAP7_75t_L g13 ( .A(n_11), .Y(n_13) );
NOR2xp67_ASAP7_75t_SL g14 ( .A(n_11), .B(n_1), .Y(n_14) );
NOR3xp33_ASAP7_75t_L g15 ( .A(n_12), .B(n_1), .C(n_2), .Y(n_15) );
AOI21xp5_ASAP7_75t_L g16 ( .A1(n_11), .A2(n_2), .B(n_3), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_9), .Y(n_17) );
OR2x6_ASAP7_75t_L g18 ( .A(n_16), .B(n_12), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_13), .Y(n_19) );
AND2x4_ASAP7_75t_L g20 ( .A(n_17), .B(n_9), .Y(n_20) );
INVx1_ASAP7_75t_SL g21 ( .A(n_20), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_20), .B(n_14), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_20), .Y(n_23) );
INVxp67_ASAP7_75t_SL g24 ( .A(n_21), .Y(n_24) );
AOI321xp33_ASAP7_75t_L g25 ( .A1(n_23), .A2(n_15), .A3(n_10), .B1(n_18), .B2(n_14), .C(n_7), .Y(n_25) );
OA22x2_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_18), .B1(n_22), .B2(n_19), .Y(n_26) );
OAI211xp5_ASAP7_75t_SL g27 ( .A1(n_25), .A2(n_19), .B(n_18), .C(n_13), .Y(n_27) );
O2A1O1Ixp33_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_18), .B(n_24), .C(n_13), .Y(n_28) );
INVx1_ASAP7_75t_SL g29 ( .A(n_26), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
AOI22xp5_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_29), .B1(n_28), .B2(n_8), .Y(n_31) );
endmodule