module fake_ariane_2784_n_10217 (n_83, n_8, n_56, n_60, n_64, n_119, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_44, n_30, n_82, n_31, n_42, n_57, n_70, n_10, n_117, n_85, n_6, n_48, n_94, n_101, n_4, n_2, n_32, n_37, n_58, n_65, n_9, n_112, n_45, n_11, n_122, n_52, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_35, n_54, n_25, n_10217);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_70;
input n_10;
input n_117;
input n_85;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_9;
input n_112;
input n_45;
input n_11;
input n_122;
input n_52;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_35;
input n_54;
input n_25;

output n_10217;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_9872;
wire n_9604;
wire n_7329;
wire n_4030;
wire n_7029;
wire n_6790;
wire n_4770;
wire n_8165;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_6603;
wire n_2679;
wire n_6557;
wire n_5402;
wire n_6581;
wire n_2182;
wire n_5553;
wire n_6002;
wire n_7277;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_5717;
wire n_2993;
wire n_4283;
wire n_9297;
wire n_2879;
wire n_4403;
wire n_8139;
wire n_416;
wire n_4962;
wire n_1430;
wire n_7832;
wire n_8438;
wire n_2002;
wire n_1238;
wire n_2729;
wire n_4302;
wire n_5791;
wire n_7127;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_8321;
wire n_864;
wire n_5302;
wire n_1096;
wire n_1379;
wire n_10000;
wire n_2376;
wire n_7922;
wire n_7805;
wire n_9807;
wire n_2790;
wire n_7542;
wire n_2207;
wire n_7053;
wire n_9892;
wire n_5712;
wire n_3954;
wire n_6297;
wire n_4982;
wire n_2042;
wire n_462;
wire n_8699;
wire n_9263;
wire n_9734;
wire n_1131;
wire n_8037;
wire n_5479;
wire n_2646;
wire n_8257;
wire n_737;
wire n_2653;
wire n_4610;
wire n_6058;
wire n_10213;
wire n_232;
wire n_3115;
wire n_9886;
wire n_4028;
wire n_5263;
wire n_5565;
wire n_9096;
wire n_6358;
wire n_8546;
wire n_6293;
wire n_8997;
wire n_2482;
wire n_9985;
wire n_9665;
wire n_1682;
wire n_7001;
wire n_10169;
wire n_958;
wire n_6129;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_5590;
wire n_2621;
wire n_6524;
wire n_146;
wire n_9241;
wire n_9286;
wire n_4853;
wire n_8744;
wire n_338;
wire n_9592;
wire n_1909;
wire n_5229;
wire n_6313;
wire n_7464;
wire n_8449;
wire n_9683;
wire n_4260;
wire n_903;
wire n_7626;
wire n_9939;
wire n_3348;
wire n_239;
wire n_3261;
wire n_9358;
wire n_1761;
wire n_9466;
wire n_8953;
wire n_7965;
wire n_7368;
wire n_9787;
wire n_1690;
wire n_8399;
wire n_2807;
wire n_6664;
wire n_8598;
wire n_7562;
wire n_9997;
wire n_7534;
wire n_1018;
wire n_7428;
wire n_4512;
wire n_6190;
wire n_8460;
wire n_4132;
wire n_1364;
wire n_7373;
wire n_2390;
wire n_8068;
wire n_6891;
wire n_4500;
wire n_9318;
wire n_625;
wire n_2322;
wire n_8734;
wire n_1107;
wire n_8720;
wire n_331;
wire n_559;
wire n_2663;
wire n_8097;
wire n_5481;
wire n_6539;
wire n_495;
wire n_8114;
wire n_4824;
wire n_8422;
wire n_7467;
wire n_350;
wire n_8126;
wire n_381;
wire n_5340;
wire n_3545;
wire n_6797;
wire n_7392;
wire n_9714;
wire n_1428;
wire n_1284;
wire n_7526;
wire n_1241;
wire n_8664;
wire n_4741;
wire n_10131;
wire n_561;
wire n_4143;
wire n_4273;
wire n_507;
wire n_901;
wire n_4136;
wire n_9809;
wire n_3144;
wire n_2359;
wire n_9613;
wire n_9354;
wire n_1519;
wire n_7338;
wire n_5896;
wire n_4567;
wire n_9897;
wire n_786;
wire n_9295;
wire n_5833;
wire n_6249;
wire n_6887;
wire n_6253;
wire n_9119;
wire n_6128;
wire n_3552;
wire n_2950;
wire n_9058;
wire n_6197;
wire n_7200;
wire n_8326;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_5589;
wire n_8504;
wire n_3015;
wire n_5744;
wire n_8920;
wire n_3870;
wire n_6808;
wire n_3749;
wire n_1676;
wire n_1085;
wire n_277;
wire n_5691;
wire n_7937;
wire n_8985;
wire n_3482;
wire n_7490;
wire n_6295;
wire n_5403;
wire n_823;
wire n_1900;
wire n_620;
wire n_6096;
wire n_4268;
wire n_6338;
wire n_587;
wire n_863;
wire n_6992;
wire n_303;
wire n_3960;
wire n_2433;
wire n_352;
wire n_899;
wire n_3975;
wire n_8035;
wire n_5830;
wire n_9516;
wire n_365;
wire n_2004;
wire n_4018;
wire n_1495;
wire n_8660;
wire n_334;
wire n_192;
wire n_3325;
wire n_6681;
wire n_661;
wire n_4227;
wire n_5158;
wire n_9917;
wire n_5152;
wire n_8939;
wire n_533;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_1924;
wire n_6542;
wire n_9202;
wire n_1811;
wire n_6161;
wire n_3612;
wire n_273;
wire n_4505;
wire n_6452;
wire n_1840;
wire n_5247;
wire n_9512;
wire n_9923;
wire n_8469;
wire n_8715;
wire n_5464;
wire n_7306;
wire n_10070;
wire n_4476;
wire n_6740;
wire n_6978;
wire n_579;
wire n_7507;
wire n_844;
wire n_1267;
wire n_8176;
wire n_9677;
wire n_2956;
wire n_7441;
wire n_7215;
wire n_149;
wire n_1213;
wire n_2382;
wire n_7379;
wire n_5210;
wire n_237;
wire n_780;
wire n_5292;
wire n_1918;
wire n_8327;
wire n_8991;
wire n_7438;
wire n_8855;
wire n_4119;
wire n_4443;
wire n_9811;
wire n_4000;
wire n_9508;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_6136;
wire n_1140;
wire n_3458;
wire n_570;
wire n_5843;
wire n_7874;
wire n_8539;
wire n_8630;
wire n_9308;
wire n_8533;
wire n_7108;
wire n_3511;
wire n_2077;
wire n_9638;
wire n_1121;
wire n_490;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_575;
wire n_8435;
wire n_7695;
wire n_6156;
wire n_1216;
wire n_4908;
wire n_8098;
wire n_3754;
wire n_8204;
wire n_5060;
wire n_9199;
wire n_7162;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_9808;
wire n_7331;
wire n_5913;
wire n_8958;
wire n_4530;
wire n_9821;
wire n_1432;
wire n_2245;
wire n_5614;
wire n_5391;
wire n_5452;
wire n_3359;
wire n_7944;
wire n_3841;
wire n_5249;
wire n_249;
wire n_851;
wire n_123;
wire n_444;
wire n_3900;
wire n_3413;
wire n_7850;
wire n_5076;
wire n_3539;
wire n_5757;
wire n_9265;
wire n_6872;
wire n_6644;
wire n_9143;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_930;
wire n_4912;
wire n_9845;
wire n_4226;
wire n_10112;
wire n_4311;
wire n_3284;
wire n_8542;
wire n_8572;
wire n_5046;
wire n_7607;
wire n_7642;
wire n_8373;
wire n_8424;
wire n_8442;
wire n_1386;
wire n_9304;
wire n_6236;
wire n_7104;
wire n_8147;
wire n_3506;
wire n_4827;
wire n_6801;
wire n_1842;
wire n_7397;
wire n_4993;
wire n_3678;
wire n_7205;
wire n_10080;
wire n_366;
wire n_2791;
wire n_1661;
wire n_555;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_6563;
wire n_5968;
wire n_992;
wire n_966;
wire n_3549;
wire n_3914;
wire n_6398;
wire n_5586;
wire n_7461;
wire n_8519;
wire n_1692;
wire n_2611;
wire n_8075;
wire n_5468;
wire n_3029;
wire n_4745;
wire n_7638;
wire n_2398;
wire n_4791;
wire n_4233;
wire n_5971;
wire n_6319;
wire n_8642;
wire n_8648;
wire n_7224;
wire n_6966;
wire n_9791;
wire n_5056;
wire n_9449;
wire n_9934;
wire n_9149;
wire n_9686;
wire n_1178;
wire n_2015;
wire n_7259;
wire n_7838;
wire n_8556;
wire n_5984;
wire n_9844;
wire n_5204;
wire n_6724;
wire n_6705;
wire n_2877;
wire n_7307;
wire n_6776;
wire n_203;
wire n_9458;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_150;
wire n_2930;
wire n_7840;
wire n_8585;
wire n_9717;
wire n_2745;
wire n_8455;
wire n_2087;
wire n_8444;
wire n_619;
wire n_9128;
wire n_2161;
wire n_746;
wire n_6624;
wire n_1357;
wire n_7888;
wire n_8560;
wire n_292;
wire n_6710;
wire n_1787;
wire n_6883;
wire n_9558;
wire n_8108;
wire n_1389;
wire n_8158;
wire n_3172;
wire n_2659;
wire n_4033;
wire n_3747;
wire n_6553;
wire n_9715;
wire n_4905;
wire n_9016;
wire n_4508;
wire n_5897;
wire n_4045;
wire n_6261;
wire n_3651;
wire n_1812;
wire n_6659;
wire n_4894;
wire n_9399;
wire n_428;
wire n_7351;
wire n_3614;
wire n_7256;
wire n_959;
wire n_2257;
wire n_1101;
wire n_1343;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_6893;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_8814;
wire n_5778;
wire n_7021;
wire n_5179;
wire n_2435;
wire n_6337;
wire n_6210;
wire n_1932;
wire n_7583;
wire n_5680;
wire n_1780;
wire n_2825;
wire n_5685;
wire n_5974;
wire n_5723;
wire n_542;
wire n_5922;
wire n_6378;
wire n_5549;
wire n_1087;
wire n_632;
wire n_9094;
wire n_2388;
wire n_2273;
wire n_8130;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_9510;
wire n_7488;
wire n_3700;
wire n_7690;
wire n_4307;
wire n_2795;
wire n_6044;
wire n_1841;
wire n_1680;
wire n_6206;
wire n_7893;
wire n_2954;
wire n_382;
wire n_9429;
wire n_489;
wire n_4438;
wire n_6538;
wire n_7966;
wire n_251;
wire n_974;
wire n_506;
wire n_3814;
wire n_6996;
wire n_5831;
wire n_9653;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_7599;
wire n_9648;
wire n_7231;
wire n_4195;
wire n_7007;
wire n_7717;
wire n_6579;
wire n_5091;
wire n_4866;
wire n_7230;
wire n_1447;
wire n_8675;
wire n_1220;
wire n_9095;
wire n_7900;
wire n_2019;
wire n_5708;
wire n_8123;
wire n_698;
wire n_9048;
wire n_9003;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_124;
wire n_5454;
wire n_307;
wire n_1209;
wire n_4254;
wire n_646;
wire n_8913;
wire n_9932;
wire n_3438;
wire n_8220;
wire n_404;
wire n_2625;
wire n_9309;
wire n_8355;
wire n_9661;
wire n_9799;
wire n_5373;
wire n_7403;
wire n_1578;
wire n_6665;
wire n_8883;
wire n_3147;
wire n_299;
wire n_3661;
wire n_7168;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_133;
wire n_1029;
wire n_2649;
wire n_6461;
wire n_6033;
wire n_10138;
wire n_1247;
wire n_6860;
wire n_9063;
wire n_522;
wire n_1568;
wire n_2919;
wire n_7322;
wire n_6060;
wire n_3108;
wire n_5983;
wire n_5788;
wire n_9895;
wire n_367;
wire n_6709;
wire n_2632;
wire n_5557;
wire n_6914;
wire n_8816;
wire n_4314;
wire n_8418;
wire n_2980;
wire n_5951;
wire n_1728;
wire n_4315;
wire n_5647;
wire n_6117;
wire n_7287;
wire n_7789;
wire n_3239;
wire n_2631;
wire n_9110;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_424;
wire n_4857;
wire n_8739;
wire n_9969;
wire n_8927;
wire n_1651;
wire n_3087;
wire n_6009;
wire n_7221;
wire n_4637;
wire n_5523;
wire n_2697;
wire n_1263;
wire n_1817;
wire n_8243;
wire n_3704;
wire n_8798;
wire n_7963;
wire n_8423;
wire n_6382;
wire n_9028;
wire n_670;
wire n_2677;
wire n_4296;
wire n_379;
wire n_162;
wire n_138;
wire n_9654;
wire n_2483;
wire n_7938;
wire n_5088;
wire n_6615;
wire n_9810;
wire n_441;
wire n_7294;
wire n_6192;
wire n_7414;
wire n_5773;
wire n_1032;
wire n_1592;
wire n_9701;
wire n_5392;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_9270;
wire n_3589;
wire n_6418;
wire n_1743;
wire n_8548;
wire n_9437;
wire n_8996;
wire n_207;
wire n_9483;
wire n_720;
wire n_6263;
wire n_1943;
wire n_6731;
wire n_8156;
wire n_5138;
wire n_8845;
wire n_4588;
wire n_6048;
wire n_7185;
wire n_194;
wire n_5149;
wire n_9256;
wire n_1163;
wire n_3054;
wire n_4970;
wire n_5280;
wire n_6234;
wire n_4153;
wire n_8992;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_7141;
wire n_2373;
wire n_3881;
wire n_6224;
wire n_8510;
wire n_5089;
wire n_5775;
wire n_9854;
wire n_2099;
wire n_3759;
wire n_9737;
wire n_8961;
wire n_9964;
wire n_3323;
wire n_4643;
wire n_9719;
wire n_6142;
wire n_2617;
wire n_6119;
wire n_6619;
wire n_808;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_1439;
wire n_6759;
wire n_6903;
wire n_3466;
wire n_7416;
wire n_2074;
wire n_5031;
wire n_6768;
wire n_1665;
wire n_7092;
wire n_7233;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_9679;
wire n_9669;
wire n_5082;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_4555;
wire n_5230;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_8402;
wire n_8978;
wire n_7191;
wire n_2117;
wire n_6189;
wire n_1053;
wire n_5796;
wire n_9105;
wire n_9699;
wire n_5296;
wire n_5398;
wire n_1906;
wire n_6761;
wire n_9673;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_8685;
wire n_1828;
wire n_9240;
wire n_1304;
wire n_7202;
wire n_3335;
wire n_5960;
wire n_3007;
wire n_2267;
wire n_7445;
wire n_5858;
wire n_9212;
wire n_5985;
wire n_8595;
wire n_604;
wire n_478;
wire n_9040;
wire n_1349;
wire n_9478;
wire n_1061;
wire n_2102;
wire n_4157;
wire n_9742;
wire n_3477;
wire n_7868;
wire n_10124;
wire n_3370;
wire n_874;
wire n_7654;
wire n_3949;
wire n_2286;
wire n_8779;
wire n_5192;
wire n_4247;
wire n_707;
wire n_5051;
wire n_10132;
wire n_5336;
wire n_129;
wire n_126;
wire n_3036;
wire n_2783;
wire n_8520;
wire n_4583;
wire n_8555;
wire n_9456;
wire n_6366;
wire n_1015;
wire n_1162;
wire n_6304;
wire n_4292;
wire n_2118;
wire n_9146;
wire n_688;
wire n_7176;
wire n_636;
wire n_8565;
wire n_8334;
wire n_1490;
wire n_5552;
wire n_6074;
wire n_7547;
wire n_442;
wire n_3764;
wire n_1553;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_1086;
wire n_3025;
wire n_9573;
wire n_3051;
wire n_986;
wire n_1104;
wire n_2802;
wire n_8030;
wire n_8513;
wire n_887;
wire n_9379;
wire n_9219;
wire n_2125;
wire n_1156;
wire n_5123;
wire n_8245;
wire n_6689;
wire n_2861;
wire n_4974;
wire n_7942;
wire n_4344;
wire n_5242;
wire n_3130;
wire n_8753;
wire n_1188;
wire n_1498;
wire n_7527;
wire n_9706;
wire n_7948;
wire n_2618;
wire n_4856;
wire n_7096;
wire n_4216;
wire n_957;
wire n_1242;
wire n_9206;
wire n_2707;
wire n_8485;
wire n_5596;
wire n_6482;
wire n_10118;
wire n_8106;
wire n_2849;
wire n_1489;
wire n_8325;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_6335;
wire n_5742;
wire n_5127;
wire n_4313;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_1119;
wire n_9434;
wire n_3713;
wire n_6229;
wire n_1863;
wire n_5933;
wire n_5536;
wire n_4798;
wire n_1500;
wire n_616;
wire n_7293;
wire n_9874;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_1189;
wire n_5810;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_9082;
wire n_7144;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_4991;
wire n_7316;
wire n_7508;
wire n_9596;
wire n_3070;
wire n_1005;
wire n_8677;
wire n_5818;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_9559;
wire n_9709;
wire n_2452;
wire n_4182;
wire n_8626;
wire n_2827;
wire n_7869;
wire n_3214;
wire n_10069;
wire n_8166;
wire n_9356;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5539;
wire n_5009;
wire n_3710;
wire n_1844;
wire n_6943;
wire n_1957;
wire n_1953;
wire n_1219;
wire n_710;
wire n_6631;
wire n_5889;
wire n_8602;
wire n_9609;
wire n_7151;
wire n_3944;
wire n_7762;
wire n_5632;
wire n_4729;
wire n_8002;
wire n_6728;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_5613;
wire n_7472;
wire n_9342;
wire n_4800;
wire n_1373;
wire n_7075;
wire n_1540;
wire n_5427;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_6770;
wire n_5450;
wire n_7611;
wire n_7796;
wire n_6508;
wire n_832;
wire n_7989;
wire n_8047;
wire n_744;
wire n_2821;
wire n_9233;
wire n_3696;
wire n_7936;
wire n_215;
wire n_1331;
wire n_4781;
wire n_6031;
wire n_1529;
wire n_3531;
wire n_5124;
wire n_655;
wire n_4237;
wire n_8751;
wire n_5297;
wire n_4828;
wire n_3333;
wire n_8800;
wire n_4652;
wire n_4114;
wire n_7105;
wire n_7013;
wire n_7655;
wire n_1007;
wire n_9435;
wire n_1580;
wire n_3135;
wire n_4925;
wire n_5719;
wire n_7254;
wire n_2448;
wire n_9557;
wire n_2211;
wire n_8955;
wire n_9551;
wire n_951;
wire n_8039;
wire n_8193;
wire n_9073;
wire n_7546;
wire n_8432;
wire n_5904;
wire n_6628;
wire n_5318;
wire n_5374;
wire n_8684;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_6456;
wire n_722;
wire n_7407;
wire n_9388;
wire n_3277;
wire n_9721;
wire n_4863;
wire n_1766;
wire n_5463;
wire n_1338;
wire n_2978;
wire n_6328;
wire n_6929;
wire n_4859;
wire n_4568;
wire n_8628;
wire n_3617;
wire n_6012;
wire n_704;
wire n_2958;
wire n_7481;
wire n_1044;
wire n_1714;
wire n_4429;
wire n_5435;
wire n_6484;
wire n_3340;
wire n_5053;
wire n_7182;
wire n_9507;
wire n_5476;
wire n_5483;
wire n_9539;
wire n_8617;
wire n_7605;
wire n_8591;
wire n_8090;
wire n_1243;
wire n_9268;
wire n_5511;
wire n_9718;
wire n_8661;
wire n_10068;
wire n_3486;
wire n_6639;
wire n_358;
wire n_608;
wire n_9672;
wire n_9890;
wire n_9187;
wire n_2457;
wire n_9572;
wire n_2992;
wire n_6124;
wire n_9527;
wire n_317;
wire n_3197;
wire n_9949;
wire n_7423;
wire n_3256;
wire n_1878;
wire n_7375;
wire n_7076;
wire n_7689;
wire n_6344;
wire n_8189;
wire n_8811;
wire n_266;
wire n_9952;
wire n_7736;
wire n_6435;
wire n_3646;
wire n_5829;
wire n_2520;
wire n_7419;
wire n_811;
wire n_6600;
wire n_7010;
wire n_791;
wire n_5881;
wire n_9798;
wire n_3864;
wire n_4694;
wire n_8192;
wire n_9251;
wire n_1025;
wire n_4664;
wire n_6201;
wire n_3450;
wire n_8573;
wire n_687;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_480;
wire n_7918;
wire n_642;
wire n_9546;
wire n_1406;
wire n_5073;
wire n_6555;
wire n_4306;
wire n_6360;
wire n_6735;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_9181;
wire n_9602;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_6803;
wire n_4288;
wire n_3452;
wire n_474;
wire n_4098;
wire n_2691;
wire n_5894;
wire n_9635;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_695;
wire n_2991;
wire n_5419;
wire n_8339;
wire n_386;
wire n_1596;
wire n_4289;
wire n_4972;
wire n_197;
wire n_2723;
wire n_1476;
wire n_6036;
wire n_7346;
wire n_9405;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_8775;
wire n_678;
wire n_10158;
wire n_651;
wire n_2850;
wire n_1874;
wire n_5077;
wire n_6102;
wire n_3780;
wire n_1657;
wire n_9726;
wire n_8804;
wire n_9577;
wire n_6650;
wire n_10024;
wire n_6573;
wire n_6904;
wire n_3753;
wire n_6329;
wire n_7385;
wire n_9802;
wire n_1488;
wire n_6244;
wire n_4846;
wire n_9250;
wire n_1330;
wire n_906;
wire n_6204;
wire n_9540;
wire n_10191;
wire n_2295;
wire n_5225;
wire n_283;
wire n_7295;
wire n_4076;
wire n_7824;
wire n_7148;
wire n_3142;
wire n_9171;
wire n_7169;
wire n_3129;
wire n_9350;
wire n_374;
wire n_3495;
wire n_3843;
wire n_6756;
wire n_4805;
wire n_2606;
wire n_9441;
wire n_7600;
wire n_9124;
wire n_2386;
wire n_8697;
wire n_5826;
wire n_9626;
wire n_4822;
wire n_6946;
wire n_7947;
wire n_8645;
wire n_5931;
wire n_8820;
wire n_8146;
wire n_9408;
wire n_1829;
wire n_4635;
wire n_7847;
wire n_8154;
wire n_1450;
wire n_5532;
wire n_7311;
wire n_3740;
wire n_6804;
wire n_5441;
wire n_6179;
wire n_2417;
wire n_6059;
wire n_1815;
wire n_7039;
wire n_8027;
wire n_7807;
wire n_1493;
wire n_2911;
wire n_515;
wire n_8063;
wire n_3313;
wire n_8406;
wire n_2354;
wire n_6427;
wire n_4281;
wire n_3945;
wire n_5994;
wire n_3726;
wire n_8480;
wire n_9754;
wire n_4419;
wire n_8849;
wire n_5405;
wire n_9750;
wire n_7660;
wire n_1256;
wire n_9529;
wire n_9566;
wire n_3560;
wire n_3345;
wire n_5772;
wire n_5365;
wire n_6442;
wire n_8241;
wire n_140;
wire n_6188;
wire n_3421;
wire n_1448;
wire n_10066;
wire n_1009;
wire n_230;
wire n_3548;
wire n_4906;
wire n_6846;
wire n_10054;
wire n_4630;
wire n_8261;
wire n_6840;
wire n_142;
wire n_6645;
wire n_8535;
wire n_8348;
wire n_4829;
wire n_6749;
wire n_6915;
wire n_7831;
wire n_8138;
wire n_2612;
wire n_5259;
wire n_3236;
wire n_8702;
wire n_1995;
wire n_7455;
wire n_8273;
wire n_1397;
wire n_6247;
wire n_5921;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_4966;
wire n_2250;
wire n_8235;
wire n_1117;
wire n_6104;
wire n_3321;
wire n_9940;
wire n_8294;
wire n_1303;
wire n_4188;
wire n_10016;
wire n_2001;
wire n_9036;
wire n_9165;
wire n_7509;
wire n_9283;
wire n_6205;
wire n_2506;
wire n_8349;
wire n_2413;
wire n_4825;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_9822;
wire n_10036;
wire n_2626;
wire n_9443;
wire n_9607;
wire n_7497;
wire n_7315;
wire n_10166;
wire n_8429;
wire n_2892;
wire n_6939;
wire n_2605;
wire n_7887;
wire n_2804;
wire n_9298;
wire n_5884;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_10006;
wire n_5728;
wire n_1035;
wire n_3475;
wire n_4878;
wire n_8486;
wire n_9052;
wire n_2070;
wire n_426;
wire n_6706;
wire n_7431;
wire n_8140;
wire n_398;
wire n_3842;
wire n_1367;
wire n_4202;
wire n_6909;
wire n_2044;
wire n_6487;
wire n_5679;
wire n_166;
wire n_8117;
wire n_3886;
wire n_825;
wire n_732;
wire n_2619;
wire n_7521;
wire n_10058;
wire n_1192;
wire n_5141;
wire n_3098;
wire n_6627;
wire n_4503;
wire n_8129;
wire n_1291;
wire n_7253;
wire n_9535;
wire n_5208;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_9943;
wire n_7569;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_7452;
wire n_6551;
wire n_3386;
wire n_400;
wire n_7972;
wire n_8672;
wire n_7505;
wire n_3921;
wire n_282;
wire n_467;
wire n_2177;
wire n_6516;
wire n_2766;
wire n_10060;
wire n_7524;
wire n_4196;
wire n_1197;
wire n_8934;
wire n_7318;
wire n_2613;
wire n_9977;
wire n_7411;
wire n_7326;
wire n_5667;
wire n_168;
wire n_9555;
wire n_1517;
wire n_2647;
wire n_8847;
wire n_8005;
wire n_5508;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_5879;
wire n_1671;
wire n_6500;
wire n_5027;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_3380;
wire n_5688;
wire n_2826;
wire n_9030;
wire n_5825;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_8221;
wire n_7573;
wire n_6630;
wire n_5629;
wire n_5759;
wire n_2411;
wire n_4631;
wire n_8191;
wire n_6798;
wire n_5999;
wire n_1504;
wire n_9590;
wire n_2110;
wire n_7498;
wire n_7895;
wire n_6421;
wire n_5377;
wire n_6180;
wire n_8225;
wire n_3822;
wire n_889;
wire n_4355;
wire n_7453;
wire n_3818;
wire n_7932;
wire n_9651;
wire n_7890;
wire n_5599;
wire n_3587;
wire n_2608;
wire n_6004;
wire n_9583;
wire n_9763;
wire n_9944;
wire n_1948;
wire n_6652;
wire n_9888;
wire n_7183;
wire n_4155;
wire n_810;
wire n_4278;
wire n_10040;
wire n_4710;
wire n_1959;
wire n_6275;
wire n_6403;
wire n_3497;
wire n_6395;
wire n_9862;
wire n_4542;
wire n_5451;
wire n_6578;
wire n_3243;
wire n_4326;
wire n_9966;
wire n_2121;
wire n_3865;
wire n_6350;
wire n_5460;
wire n_4685;
wire n_9936;
wire n_565;
wire n_3927;
wire n_6141;
wire n_8559;
wire n_2068;
wire n_3595;
wire n_6875;
wire n_7189;
wire n_1194;
wire n_9617;
wire n_4060;
wire n_1647;
wire n_9341;
wire n_6194;
wire n_1454;
wire n_2459;
wire n_941;
wire n_8689;
wire n_3396;
wire n_9749;
wire n_5517;
wire n_9629;
wire n_5807;
wire n_5426;
wire n_6475;
wire n_4093;
wire n_452;
wire n_5693;
wire n_5695;
wire n_4123;
wire n_4294;
wire n_8330;
wire n_10011;
wire n_1521;
wire n_1940;
wire n_3683;
wire n_6502;
wire n_10030;
wire n_6944;
wire n_4452;
wire n_284;
wire n_3887;
wire n_3195;
wire n_8304;
wire n_9349;
wire n_5587;
wire n_4722;
wire n_6318;
wire n_10119;
wire n_8163;
wire n_6805;
wire n_3048;
wire n_3339;
wire n_4164;
wire n_4126;
wire n_7240;
wire n_5030;
wire n_8907;
wire n_409;
wire n_2963;
wire n_5674;
wire n_2561;
wire n_7499;
wire n_9423;
wire n_1056;
wire n_526;
wire n_5584;
wire n_674;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_6075;
wire n_10063;
wire n_6559;
wire n_4088;
wire n_9038;
wire n_8777;
wire n_2669;
wire n_8698;
wire n_3911;
wire n_6068;
wire n_3802;
wire n_4366;
wire n_1584;
wire n_6248;
wire n_6541;
wire n_9034;
wire n_848;
wire n_5125;
wire n_4922;
wire n_6066;
wire n_6080;
wire n_629;
wire n_4733;
wire n_7927;
wire n_161;
wire n_8928;
wire n_1814;
wire n_7219;
wire n_2441;
wire n_8081;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_216;
wire n_6150;
wire n_6638;
wire n_7063;
wire n_7402;
wire n_9676;
wire n_6351;
wire n_4509;
wire n_4935;
wire n_2073;
wire n_7382;
wire n_8384;
wire n_4004;
wire n_5238;
wire n_750;
wire n_834;
wire n_8650;
wire n_3630;
wire n_1612;
wire n_800;
wire n_1910;
wire n_5906;
wire n_7767;
wire n_2189;
wire n_5732;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_2602;
wire n_5780;
wire n_724;
wire n_2931;
wire n_3433;
wire n_8284;
wire n_8374;
wire n_5556;
wire n_6006;
wire n_3597;
wire n_6474;
wire n_5743;
wire n_6481;
wire n_10078;
wire n_1956;
wire n_1589;
wire n_5633;
wire n_4111;
wire n_7510;
wire n_9041;
wire n_3786;
wire n_875;
wire n_9995;
wire n_6022;
wire n_6991;
wire n_2828;
wire n_7434;
wire n_1626;
wire n_5950;
wire n_1335;
wire n_9035;
wire n_9011;
wire n_1715;
wire n_4204;
wire n_7691;
wire n_296;
wire n_3553;
wire n_5323;
wire n_7745;
wire n_9135;
wire n_6744;
wire n_3645;
wire n_9776;
wire n_793;
wire n_5705;
wire n_6927;
wire n_7335;
wire n_132;
wire n_9413;
wire n_9107;
wire n_4996;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_7735;
wire n_8531;
wire n_6116;
wire n_9548;
wire n_8074;
wire n_494;
wire n_3550;
wire n_8780;
wire n_7956;
wire n_5510;
wire n_7495;
wire n_7651;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_9775;
wire n_1805;
wire n_8580;
wire n_4068;
wire n_5440;
wire n_9288;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_2443;
wire n_3610;
wire n_185;
wire n_5011;
wire n_6757;
wire n_7536;
wire n_1554;
wire n_3279;
wire n_5513;
wire n_5875;
wire n_8358;
wire n_972;
wire n_7734;
wire n_4262;
wire n_2923;
wire n_164;
wire n_2843;
wire n_3714;
wire n_9305;
wire n_9093;
wire n_184;
wire n_7671;
wire n_10043;
wire n_4832;
wire n_8033;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_6485;
wire n_5848;
wire n_1679;
wire n_5834;
wire n_7926;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_5784;
wire n_3125;
wire n_5128;
wire n_8643;
wire n_2356;
wire n_5618;
wire n_10134;
wire n_6495;
wire n_7528;
wire n_6209;
wire n_4672;
wire n_8094;
wire n_2564;
wire n_3558;
wire n_9425;
wire n_3034;
wire n_3502;
wire n_783;
wire n_4053;
wire n_1127;
wire n_7413;
wire n_7993;
wire n_7821;
wire n_160;
wire n_7620;
wire n_1008;
wire n_3963;
wire n_581;
wire n_3091;
wire n_6274;
wire n_1024;
wire n_176;
wire n_5157;
wire n_4496;
wire n_9347;
wire n_2518;
wire n_936;
wire n_4596;
wire n_5178;
wire n_9420;
wire n_3105;
wire n_6237;
wire n_1525;
wire n_4628;
wire n_6802;
wire n_7343;
wire n_5982;
wire n_8477;
wire n_1775;
wire n_908;
wire n_1036;
wire n_9344;
wire n_7109;
wire n_8028;
wire n_341;
wire n_4083;
wire n_1270;
wire n_1272;
wire n_549;
wire n_2794;
wire n_6155;
wire n_2901;
wire n_7506;
wire n_3940;
wire n_9530;
wire n_6809;
wire n_10160;
wire n_6099;
wire n_3225;
wire n_8530;
wire n_9446;
wire n_3621;
wire n_5529;
wire n_244;
wire n_7561;
wire n_3473;
wire n_6349;
wire n_3680;
wire n_8500;
wire n_6716;
wire n_8713;
wire n_3565;
wire n_7885;
wire n_8297;
wire n_6905;
wire n_8926;
wire n_9865;
wire n_8456;
wire n_7722;
wire n_5388;
wire n_7470;
wire n_5824;
wire n_8025;
wire n_5354;
wire n_2453;
wire n_7898;
wire n_3331;
wire n_1788;
wire n_6203;
wire n_2138;
wire n_6407;
wire n_3040;
wire n_4230;
wire n_6899;
wire n_7980;
wire n_7817;
wire n_6413;
wire n_445;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_7070;
wire n_9025;
wire n_2000;
wire n_5276;
wire n_4037;
wire n_9713;
wire n_3804;
wire n_4659;
wire n_8293;
wire n_3211;
wire n_7299;
wire n_917;
wire n_5196;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_8029;
wire n_2215;
wire n_9314;
wire n_3847;
wire n_6960;
wire n_4073;
wire n_8880;
wire n_1261;
wire n_7249;
wire n_9660;
wire n_5763;
wire n_3633;
wire n_857;
wire n_363;
wire n_6061;
wire n_1235;
wire n_9769;
wire n_2584;
wire n_4001;
wire n_8471;
wire n_1462;
wire n_5701;
wire n_7002;
wire n_1064;
wire n_633;
wire n_1446;
wire n_9902;
wire n_1701;
wire n_6273;
wire n_7094;
wire n_7396;
wire n_3111;
wire n_8726;
wire n_731;
wire n_8977;
wire n_1813;
wire n_315;
wire n_2997;
wire n_7018;
wire n_1573;
wire n_6746;
wire n_3258;
wire n_758;
wire n_3691;
wire n_2252;
wire n_8316;
wire n_6174;
wire n_6545;
wire n_7773;
wire n_6763;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_7297;
wire n_784;
wire n_4339;
wire n_5907;
wire n_7730;
wire n_8134;
wire n_6013;
wire n_6182;
wire n_6754;
wire n_4690;
wire n_2987;
wire n_6279;
wire n_1473;
wire n_1076;
wire n_1348;
wire n_5895;
wire n_9410;
wire n_2651;
wire n_753;
wire n_9588;
wire n_2445;
wire n_2733;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_8610;
wire n_4023;
wire n_10071;
wire n_4253;
wire n_7637;
wire n_2522;
wire n_3632;
wire n_309;
wire n_1344;
wire n_485;
wire n_4064;
wire n_6131;
wire n_3351;
wire n_5478;
wire n_10176;
wire n_435;
wire n_6113;
wire n_1141;
wire n_3457;
wire n_9740;
wire n_5384;
wire n_6477;
wire n_7486;
wire n_840;
wire n_2324;
wire n_6575;
wire n_5283;
wire n_9910;
wire n_3454;
wire n_7544;
wire n_5961;
wire n_2139;
wire n_7613;
wire n_9061;
wire n_7995;
wire n_9941;
wire n_8113;
wire n_9579;
wire n_2521;
wire n_5686;
wire n_6391;
wire n_2740;
wire n_1991;
wire n_8724;
wire n_7140;
wire n_614;
wire n_4066;
wire n_9668;
wire n_6252;
wire n_6426;
wire n_4681;
wire n_8253;
wire n_9258;
wire n_9228;
wire n_3303;
wire n_7910;
wire n_6592;
wire n_4414;
wire n_10214;
wire n_2541;
wire n_5094;
wire n_10195;
wire n_3232;
wire n_1113;
wire n_9598;
wire n_248;
wire n_7741;
wire n_3768;
wire n_4295;
wire n_1615;
wire n_4100;
wire n_228;
wire n_6668;
wire n_9311;
wire n_1265;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_4087;
wire n_8232;
wire n_1409;
wire n_1684;
wire n_1588;
wire n_1148;
wire n_8803;
wire n_1673;
wire n_4473;
wire n_4619;
wire n_6670;
wire n_5371;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_7679;
wire n_3018;
wire n_8818;
wire n_7698;
wire n_1875;
wire n_10073;
wire n_6962;
wire n_2429;
wire n_6779;
wire n_9608;
wire n_5286;
wire n_10164;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_10205;
wire n_1039;
wire n_5676;
wire n_5949;
wire n_5040;
wire n_6901;
wire n_1150;
wire n_7800;
wire n_4266;
wire n_6336;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_6503;
wire n_7835;
wire n_1136;
wire n_458;
wire n_1190;
wire n_6049;
wire n_5885;
wire n_3628;
wire n_9818;
wire n_7100;
wire n_4777;
wire n_7243;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_7415;
wire n_8823;
wire n_5399;
wire n_8536;
wire n_9433;
wire n_658;
wire n_362;
wire n_8795;
wire n_2846;
wire n_3371;
wire n_9599;
wire n_8674;
wire n_9186;
wire n_4918;
wire n_5856;
wire n_8016;
wire n_3872;
wire n_5760;
wire n_7747;
wire n_9935;
wire n_4415;
wire n_5110;
wire n_8966;
wire n_1964;
wire n_3659;
wire n_7552;
wire n_3928;
wire n_10018;
wire n_9537;
wire n_1777;
wire n_9552;
wire n_9421;
wire n_3366;
wire n_6998;
wire n_7395;
wire n_5844;
wire n_6298;
wire n_8132;
wire n_7650;
wire n_3441;
wire n_199;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_7535;
wire n_708;
wire n_6609;
wire n_2545;
wire n_2513;
wire n_7635;
wire n_4408;
wire n_2115;
wire n_8567;
wire n_8259;
wire n_2017;
wire n_1810;
wire n_1347;
wire n_4976;
wire n_9473;
wire n_860;
wire n_6525;
wire n_10208;
wire n_3555;
wire n_9469;
wire n_5938;
wire n_7274;
wire n_3534;
wire n_450;
wire n_8578;
wire n_4548;
wire n_7819;
wire n_8495;
wire n_2670;
wire n_6494;
wire n_3556;
wire n_896;
wire n_4574;
wire n_8160;
wire n_8980;
wire n_2644;
wire n_6132;
wire n_4557;
wire n_3071;
wire n_8336;
wire n_1698;
wire n_1337;
wire n_774;
wire n_2148;
wire n_5548;
wire n_7788;
wire n_6974;
wire n_1168;
wire n_4663;
wire n_219;
wire n_5840;
wire n_6882;
wire n_3296;
wire n_9909;
wire n_3794;
wire n_3762;
wire n_4624;
wire n_656;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_6498;
wire n_6562;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_8600;
wire n_8229;
wire n_415;
wire n_4686;
wire n_9236;
wire n_9751;
wire n_2384;
wire n_7794;
wire n_1705;
wire n_768;
wire n_3707;
wire n_1091;
wire n_3895;
wire n_9369;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_5917;
wire n_9757;
wire n_6965;
wire n_2058;
wire n_3231;
wire n_8761;
wire n_1846;
wire n_7630;
wire n_4161;
wire n_304;
wire n_9076;
wire n_6168;
wire n_5304;
wire n_5437;
wire n_6963;
wire n_6951;
wire n_1581;
wire n_946;
wire n_757;
wire n_2047;
wire n_3058;
wire n_375;
wire n_1655;
wire n_3398;
wire n_5355;
wire n_1146;
wire n_9729;
wire n_3709;
wire n_6284;
wire n_998;
wire n_3592;
wire n_5321;
wire n_7454;
wire n_2536;
wire n_1604;
wire n_3399;
wire n_8473;
wire n_9366;
wire n_4772;
wire n_6931;
wire n_6521;
wire n_8351;
wire n_5915;
wire n_7276;
wire n_174;
wire n_6379;
wire n_9647;
wire n_1368;
wire n_963;
wire n_7085;
wire n_6306;
wire n_4120;
wire n_925;
wire n_7753;
wire n_6834;
wire n_2880;
wire n_1313;
wire n_1001;
wire n_3722;
wire n_4716;
wire n_1115;
wire n_4654;
wire n_8948;
wire n_1339;
wire n_1051;
wire n_5116;
wire n_3771;
wire n_7225;
wire n_719;
wire n_7541;
wire n_3158;
wire n_3221;
wire n_10062;
wire n_2316;
wire n_7913;
wire n_10128;
wire n_8020;
wire n_7946;
wire n_8944;
wire n_1010;
wire n_2830;
wire n_5500;
wire n_9275;
wire n_4622;
wire n_4757;
wire n_803;
wire n_1871;
wire n_9520;
wire n_6949;
wire n_6471;
wire n_5669;
wire n_5672;
wire n_4016;
wire n_3334;
wire n_5621;
wire n_9493;
wire n_6760;
wire n_2940;
wire n_548;
wire n_3427;
wire n_8875;
wire n_3162;
wire n_5569;
wire n_4591;
wire n_9102;
wire n_5966;
wire n_5515;
wire n_6589;
wire n_3083;
wire n_4570;
wire n_7014;
wire n_9801;
wire n_2491;
wire n_7920;
wire n_1931;
wire n_5559;
wire n_8649;
wire n_2259;
wire n_5337;
wire n_849;
wire n_5059;
wire n_4655;
wire n_7459;
wire n_1820;
wire n_7841;
wire n_9424;
wire n_10013;
wire n_7160;
wire n_7324;
wire n_9333;
wire n_8205;
wire n_6046;
wire n_7054;
wire n_1233;
wire n_4493;
wire n_8975;
wire n_6055;
wire n_7161;
wire n_9004;
wire n_1808;
wire n_6364;
wire n_8919;
wire n_6091;
wire n_6348;
wire n_9987;
wire n_1635;
wire n_8440;
wire n_1704;
wire n_4896;
wire n_8041;
wire n_4851;
wire n_6848;
wire n_2479;
wire n_9860;
wire n_886;
wire n_7837;
wire n_359;
wire n_9670;
wire n_6788;
wire n_1308;
wire n_6144;
wire n_1451;
wire n_1487;
wire n_675;
wire n_9200;
wire n_5528;
wire n_7806;
wire n_5605;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_9417;
wire n_6896;
wire n_2484;
wire n_5753;
wire n_8076;
wire n_5358;
wire n_1469;
wire n_4901;
wire n_3480;
wire n_8757;
wire n_1355;
wire n_10020;
wire n_7201;
wire n_4213;
wire n_4127;
wire n_6221;
wire n_2500;
wire n_9386;
wire n_8897;
wire n_7676;
wire n_8177;
wire n_2334;
wire n_5467;
wire n_7241;
wire n_1169;
wire n_789;
wire n_3181;
wire n_5493;
wire n_9207;
wire n_1916;
wire n_6285;
wire n_610;
wire n_7644;
wire n_9276;
wire n_4602;
wire n_1713;
wire n_7816;
wire n_8829;
wire n_1436;
wire n_2818;
wire n_4900;
wire n_10110;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_3745;
wire n_6748;
wire n_7430;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_8638;
wire n_1515;
wire n_817;
wire n_5901;
wire n_9980;
wire n_1566;
wire n_2837;
wire n_717;
wire n_952;
wire n_2446;
wire n_6582;
wire n_4116;
wire n_7724;
wire n_5360;
wire n_7269;
wire n_7047;
wire n_2671;
wire n_2702;
wire n_9176;
wire n_6937;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_1138;
wire n_214;
wire n_9728;
wire n_4103;
wire n_2529;
wire n_8101;
wire n_2374;
wire n_5439;
wire n_8687;
wire n_6115;
wire n_1225;
wire n_3154;
wire n_9866;
wire n_137;
wire n_8721;
wire n_1366;
wire n_8749;
wire n_9465;
wire n_3938;
wire n_8937;
wire n_2278;
wire n_6272;
wire n_7067;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_4416;
wire n_7879;
wire n_8730;
wire n_9702;
wire n_6607;
wire n_4439;
wire n_520;
wire n_870;
wire n_4985;
wire n_9000;
wire n_3382;
wire n_7117;
wire n_3930;
wire n_3808;
wire n_9610;
wire n_5471;
wire n_2248;
wire n_813;
wire n_4660;
wire n_8503;
wire n_10082;
wire n_3081;
wire n_6446;
wire n_5497;
wire n_9139;
wire n_5519;
wire n_6071;
wire n_995;
wire n_2579;
wire n_8315;
wire n_1961;
wire n_1535;
wire n_6849;
wire n_2960;
wire n_3270;
wire n_871;
wire n_6807;
wire n_2844;
wire n_8197;
wire n_402;
wire n_1979;
wire n_9407;
wire n_6616;
wire n_6719;
wire n_829;
wire n_4814;
wire n_8019;
wire n_8801;
wire n_339;
wire n_6178;
wire n_8707;
wire n_6677;
wire n_2221;
wire n_7875;
wire n_5502;
wire n_8962;
wire n_8931;
wire n_8248;
wire n_1283;
wire n_7550;
wire n_8554;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_7302;
wire n_2781;
wire n_6191;
wire n_9357;
wire n_2442;
wire n_9477;
wire n_7238;
wire n_6862;
wire n_8501;
wire n_3657;
wire n_5706;
wire n_2634;
wire n_2746;
wire n_7292;
wire n_242;
wire n_645;
wire n_7804;
wire n_5098;
wire n_721;
wire n_1084;
wire n_6000;
wire n_6774;
wire n_9289;
wire n_6443;
wire n_9828;
wire n_1276;
wire n_8263;
wire n_5145;
wire n_6072;
wire n_2878;
wire n_7248;
wire n_3830;
wire n_3252;
wire n_6647;
wire n_8040;
wire n_5466;
wire n_1528;
wire n_6941;
wire n_7239;
wire n_9797;
wire n_6552;
wire n_7826;
wire n_9981;
wire n_3315;
wire n_6094;
wire n_3523;
wire n_8102;
wire n_3999;
wire n_9793;
wire n_518;
wire n_8196;
wire n_7112;
wire n_3420;
wire n_3859;
wire n_868;
wire n_8822;
wire n_5213;
wire n_3474;
wire n_5738;
wire n_9514;
wire n_2458;
wire n_7971;
wire n_8885;
wire n_5592;
wire n_5620;
wire n_3150;
wire n_5491;
wire n_1542;
wire n_4831;
wire n_4782;
wire n_9825;
wire n_1539;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_5953;
wire n_1415;
wire n_8474;
wire n_1034;
wire n_1652;
wire n_5703;
wire n_6886;
wire n_7078;
wire n_1636;
wire n_4597;
wire n_9501;
wire n_9043;
wire n_8152;
wire n_8269;
wire n_4546;
wire n_5187;
wire n_7006;
wire n_4031;
wire n_5119;
wire n_1254;
wire n_4147;
wire n_1703;
wire n_10042;
wire n_3073;
wire n_6531;
wire n_9481;
wire n_3571;
wire n_238;
wire n_4576;
wire n_7577;
wire n_7354;
wire n_6098;
wire n_5995;
wire n_3297;
wire n_8144;
wire n_5148;
wire n_3003;
wire n_6726;
wire n_6983;
wire n_7513;
wire n_10098;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_7812;
wire n_5330;
wire n_9351;
wire n_9766;
wire n_6935;
wire n_1560;
wire n_2899;
wire n_6984;
wire n_6778;
wire n_10106;
wire n_8058;
wire n_8909;
wire n_6897;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5526;
wire n_5202;
wire n_3817;
wire n_6345;
wire n_9242;
wire n_6386;
wire n_2722;
wire n_3728;
wire n_6596;
wire n_612;
wire n_333;
wire n_5107;
wire n_7165;
wire n_512;
wire n_9777;
wire n_4680;
wire n_5067;
wire n_9522;
wire n_6830;
wire n_1012;
wire n_2061;
wire n_2685;
wire n_9748;
wire n_5987;
wire n_2512;
wire n_1790;
wire n_9005;
wire n_2788;
wire n_6642;
wire n_6291;
wire n_9666;
wire n_6510;
wire n_1443;
wire n_5264;
wire n_2595;
wire n_1465;
wire n_3084;
wire n_10028;
wire n_705;
wire n_6781;
wire n_7667;
wire n_4593;
wire n_8024;
wire n_7123;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_461;
wire n_3554;
wire n_6509;
wire n_2717;
wire n_6376;
wire n_1391;
wire n_8107;
wire n_9605;
wire n_2981;
wire n_225;
wire n_9947;
wire n_1006;
wire n_546;
wire n_9930;
wire n_4995;
wire n_1159;
wire n_6514;
wire n_5873;
wire n_4498;
wire n_772;
wire n_6741;
wire n_10083;
wire n_1245;
wire n_6434;
wire n_9662;
wire n_5741;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_9768;
wire n_1675;
wire n_2466;
wire n_6593;
wire n_676;
wire n_7827;
wire n_3758;
wire n_7631;
wire n_8748;
wire n_8452;
wire n_6690;
wire n_5423;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_8742;
wire n_3777;
wire n_8393;
wire n_9835;
wire n_1872;
wire n_9656;
wire n_1585;
wire n_3767;
wire n_6056;
wire n_9475;
wire n_5866;
wire n_5926;
wire n_212;
wire n_3692;
wire n_1351;
wire n_3234;
wire n_2216;
wire n_8122;
wire n_9724;
wire n_2426;
wire n_652;
wire n_6947;
wire n_8403;
wire n_8912;
wire n_4850;
wire n_10007;
wire n_9154;
wire n_1260;
wire n_3716;
wire n_7157;
wire n_2926;
wire n_4937;
wire n_798;
wire n_8740;
wire n_5574;
wire n_8310;
wire n_3391;
wire n_5877;
wire n_912;
wire n_10104;
wire n_6375;
wire n_460;
wire n_7781;
wire n_4786;
wire n_6042;
wire n_8238;
wire n_5203;
wire n_7908;
wire n_8296;
wire n_7091;
wire n_9788;
wire n_9833;
wire n_4354;
wire n_6429;
wire n_4235;
wire n_9589;
wire n_3159;
wire n_6315;
wire n_7855;
wire n_8850;
wire n_9861;
wire n_2855;
wire n_794;
wire n_2848;
wire n_7886;
wire n_7675;
wire n_6775;
wire n_8943;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_8993;
wire n_9205;
wire n_9418;
wire n_9946;
wire n_288;
wire n_1292;
wire n_7774;
wire n_8634;
wire n_8831;
wire n_6970;
wire n_1026;
wire n_9979;
wire n_6948;
wire n_3460;
wire n_1610;
wire n_5155;
wire n_8676;
wire n_2202;
wire n_306;
wire n_2952;
wire n_3530;
wire n_6133;
wire n_6920;
wire n_2693;
wire n_7409;
wire n_10087;
wire n_5408;
wire n_8758;
wire n_5812;
wire n_9973;
wire n_5540;
wire n_7381;
wire n_5804;
wire n_9007;
wire n_8544;
wire n_3240;
wire n_7999;
wire n_5066;
wire n_931;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_7087;
wire n_967;
wire n_9020;
wire n_10027;
wire n_9260;
wire n_5130;
wire n_4175;
wire n_10154;
wire n_6241;
wire n_9619;
wire n_1079;
wire n_5200;
wire n_9235;
wire n_3393;
wire n_10161;
wire n_8652;
wire n_9112;
wire n_2836;
wire n_7873;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_9691;
wire n_5992;
wire n_8646;
wire n_2172;
wire n_2601;
wire n_1880;
wire n_2365;
wire n_9133;
wire n_5684;
wire n_1399;
wire n_7228;
wire n_5981;
wire n_7784;
wire n_9752;
wire n_1855;
wire n_6632;
wire n_2333;
wire n_8999;
wire n_3629;
wire n_4948;
wire n_5413;
wire n_1903;
wire n_2147;
wire n_7713;
wire n_6623;
wire n_9395;
wire n_4020;
wire n_5111;
wire n_5150;
wire n_1226;
wire n_2224;
wire n_6933;
wire n_1970;
wire n_3724;
wire n_9353;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_3046;
wire n_2921;
wire n_1240;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_5444;
wire n_8031;
wire n_3257;
wire n_9804;
wire n_5737;
wire n_9125;
wire n_8015;
wire n_8412;
wire n_425;
wire n_3730;
wire n_8439;
wire n_8575;
wire n_6908;
wire n_3979;
wire n_5615;
wire n_5097;
wire n_2695;
wire n_7084;
wire n_2598;
wire n_3727;
wire n_6083;
wire n_6537;
wire n_976;
wire n_4003;
wire n_1832;
wire n_767;
wire n_8499;
wire n_9397;
wire n_6390;
wire n_7640;
wire n_2302;
wire n_6799;
wire n_8772;
wire n_9767;
wire n_3014;
wire n_7912;
wire n_2294;
wire n_6278;
wire n_2274;
wire n_7195;
wire n_5640;
wire n_3342;
wire n_2895;
wire n_6101;
wire n_7298;
wire n_8557;
wire n_3796;
wire n_9384;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_5550;
wire n_397;
wire n_3375;
wire n_2768;
wire n_351;
wire n_155;
wire n_5661;
wire n_3760;
wire n_7641;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_5306;
wire n_5905;
wire n_8815;
wire n_7949;
wire n_6112;
wire n_2728;
wire n_9906;
wire n_2025;
wire n_8679;
wire n_3744;
wire n_5457;
wire n_5159;
wire n_4022;
wire n_7115;
wire n_1020;
wire n_9310;
wire n_7764;
wire n_8446;
wire n_9163;
wire n_172;
wire n_2495;
wire n_1058;
wire n_4336;
wire n_8789;
wire n_8128;
wire n_7520;
wire n_9322;
wire n_5314;
wire n_7616;
wire n_8359;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_6412;
wire n_1279;
wire n_6271;
wire n_9377;
wire n_7235;
wire n_2511;
wire n_564;
wire n_6572;
wire n_9224;
wire n_10211;
wire n_3981;
wire n_7271;
wire n_9055;
wire n_2681;
wire n_7222;
wire n_8678;
wire n_9971;
wire n_1689;
wire n_8605;
wire n_2535;
wire n_1255;
wire n_3031;
wire n_345;
wire n_9624;
wire n_6930;
wire n_10045;
wire n_2335;
wire n_5482;
wire n_9145;
wire n_3215;
wire n_8443;
wire n_8525;
wire n_1401;
wire n_3138;
wire n_8312;
wire n_776;
wire n_2860;
wire n_8901;
wire n_2041;
wire n_1933;
wire n_6584;
wire n_4494;
wire n_9887;
wire n_130;
wire n_6387;
wire n_466;
wire n_9373;
wire n_4201;
wire n_346;
wire n_6470;
wire n_7206;
wire n_8869;
wire n_552;
wire n_9770;
wire n_5287;
wire n_8272;
wire n_4719;
wire n_5651;
wire n_264;
wire n_3577;
wire n_6625;
wire n_4074;
wire n_7383;
wire n_3994;
wire n_4636;
wire n_6826;
wire n_3185;
wire n_4983;
wire n_1217;
wire n_10103;
wire n_327;
wire n_2662;
wire n_4386;
wire n_6341;
wire n_6374;
wire n_3917;
wire n_10183;
wire n_1231;
wire n_5623;
wire n_8870;
wire n_9753;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_9468;
wire n_8178;
wire n_7854;
wire n_5524;
wire n_9517;
wire n_926;
wire n_9544;
wire n_2296;
wire n_5735;
wire n_7959;
wire n_8234;
wire n_6363;
wire n_6588;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_7897;
wire n_186;
wire n_4225;
wire n_6811;
wire n_6687;
wire n_4658;
wire n_7135;
wire n_6037;
wire n_4186;
wire n_1501;
wire n_8488;
wire n_2241;
wire n_6865;
wire n_7211;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_9774;
wire n_2531;
wire n_7132;
wire n_1570;
wire n_7533;
wire n_9586;
wire n_10150;
wire n_3377;
wire n_6722;
wire n_9780;
wire n_1518;
wire n_6420;
wire n_10004;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_7766;
wire n_855;
wire n_8862;
wire n_2059;
wire n_8184;
wire n_4713;
wire n_5787;
wire n_6911;
wire n_10151;
wire n_1287;
wire n_10187;
wire n_1611;
wire n_10171;
wire n_7129;
wire n_7080;
wire n_3374;
wire n_4870;
wire n_6981;
wire n_7776;
wire n_4818;
wire n_8001;
wire n_8695;
wire n_7436;
wire n_8767;
wire n_8571;
wire n_7020;
wire n_8064;
wire n_5935;
wire n_6696;
wire n_4916;
wire n_8472;
wire n_5967;
wire n_6095;
wire n_4323;
wire n_5934;
wire n_529;
wire n_1899;
wire n_6045;
wire n_5376;
wire n_3508;
wire n_6300;
wire n_6653;
wire n_6372;
wire n_4129;
wire n_7120;
wire n_7978;
wire n_10033;
wire n_5488;
wire n_9099;
wire n_1105;
wire n_6900;
wire n_10034;
wire n_5727;
wire n_3599;
wire n_6660;
wire n_8787;
wire n_9543;
wire n_8131;
wire n_5988;
wire n_6424;
wire n_5646;
wire n_7448;
wire n_4480;
wire n_5711;
wire n_3734;
wire n_6787;
wire n_7694;
wire n_8771;
wire n_9245;
wire n_5832;
wire n_6254;
wire n_7460;
wire n_3401;
wire n_983;
wire n_7142;
wire n_6423;
wire n_6526;
wire n_699;
wire n_3542;
wire n_301;
wire n_3263;
wire n_5891;
wire n_8150;
wire n_2523;
wire n_1945;
wire n_9168;
wire n_2418;
wire n_1614;
wire n_1377;
wire n_5328;
wire n_3819;
wire n_9074;
wire n_3222;
wire n_325;
wire n_1740;
wire n_5016;
wire n_6011;
wire n_4616;
wire n_9367;
wire n_9330;
wire n_7465;
wire n_5470;
wire n_8917;
wire n_1092;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_6176;
wire n_1963;
wire n_9300;
wire n_3868;
wire n_729;
wire n_8230;
wire n_6222;
wire n_2218;
wire n_8352;
wire n_1122;
wire n_7760;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_9918;
wire n_6969;
wire n_390;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_9496;
wire n_8914;
wire n_8821;
wire n_8465;
wire n_6587;
wire n_6688;
wire n_8360;
wire n_6505;
wire n_9837;
wire n_5362;
wire n_8209;
wire n_388;
wire n_8986;
wire n_2754;
wire n_4580;
wire n_6762;
wire n_1218;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_7629;
wire n_6987;
wire n_877;
wire n_3995;
wire n_7567;
wire n_8743;
wire n_8963;
wire n_9191;
wire n_3908;
wire n_6453;
wire n_9114;
wire n_6308;
wire n_1055;
wire n_8396;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_8514;
wire n_8550;
wire n_1089;
wire n_7449;
wire n_8151;
wire n_1502;
wire n_3501;
wire n_1478;
wire n_2555;
wire n_3216;
wire n_3568;
wire n_9913;
wire n_2708;
wire n_6187;
wire n_735;
wire n_6597;
wire n_4844;
wire n_9329;
wire n_6220;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_845;
wire n_7479;
wire n_7882;
wire n_1649;
wire n_2470;
wire n_7517;
wire n_1297;
wire n_9627;
wire n_3551;
wire n_417;
wire n_1708;
wire n_5037;
wire n_7305;
wire n_5650;
wire n_5729;
wire n_5581;
wire n_5189;
wire n_4677;
wire n_8070;
wire n_4525;
wire n_8866;
wire n_6149;
wire n_10064;
wire n_3364;
wire n_10137;
wire n_2643;
wire n_755;
wire n_9585;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_7878;
wire n_9376;
wire n_4369;
wire n_3826;
wire n_5648;
wire n_278;
wire n_2266;
wire n_6439;
wire n_4324;
wire n_842;
wire n_148;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_8797;
wire n_6547;
wire n_9524;
wire n_7177;
wire n_7902;
wire n_742;
wire n_5160;
wire n_1719;
wire n_2742;
wire n_769;
wire n_3671;
wire n_2366;
wire n_5762;
wire n_9606;
wire n_1753;
wire n_5484;
wire n_1372;
wire n_476;
wire n_10019;
wire n_1895;
wire n_7353;
wire n_4104;
wire n_8054;
wire n_982;
wire n_3791;
wire n_915;
wire n_10047;
wire n_6478;
wire n_2008;
wire n_454;
wire n_298;
wire n_4989;
wire n_5874;
wire n_3064;
wire n_3199;
wire n_8841;
wire n_9084;
wire n_2127;
wire n_7050;
wire n_3151;
wire n_7590;
wire n_6906;
wire n_403;
wire n_3016;
wire n_2460;
wire n_6739;
wire n_1319;
wire n_3669;
wire n_3367;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_606;
wire n_4528;
wire n_2772;
wire n_1700;
wire n_659;
wire n_1332;
wire n_7818;
wire n_509;
wire n_7645;
wire n_5385;
wire n_7482;
wire n_1747;
wire n_3990;
wire n_5622;
wire n_8618;
wire n_1171;
wire n_5635;
wire n_4069;
wire n_8538;
wire n_3582;
wire n_8590;
wire n_7907;
wire n_9204;
wire n_8970;
wire n_4280;
wire n_1867;
wire n_6034;
wire n_5609;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_8791;
wire n_4811;
wire n_2696;
wire n_5595;
wire n_5256;
wire n_4779;
wire n_521;
wire n_5910;
wire n_2140;
wire n_10165;
wire n_2157;
wire n_1966;
wire n_5380;
wire n_9616;
wire n_9708;
wire n_1400;
wire n_7862;
wire n_10153;
wire n_9130;
wire n_9988;
wire n_3735;
wire n_8703;
wire n_7565;
wire n_7410;
wire n_6422;
wire n_1513;
wire n_1527;
wire n_3656;
wire n_7721;
wire n_4524;
wire n_9209;
wire n_8061;
wire n_2831;
wire n_10173;
wire n_3069;
wire n_4657;
wire n_5568;
wire n_8754;
wire n_8864;
wire n_5941;
wire n_4891;
wire n_8837;
wire n_2629;
wire n_3369;
wire n_8915;
wire n_1257;
wire n_1954;
wire n_8784;
wire n_6604;
wire n_3964;
wire n_6611;
wire n_5364;
wire n_3302;
wire n_5597;
wire n_2486;
wire n_9086;
wire n_1897;
wire n_8768;
wire n_6999;
wire n_8072;
wire n_8086;
wire n_9014;
wire n_5469;
wire n_2137;
wire n_3685;
wire n_6019;
wire n_7539;
wire n_9010;
wire n_6440;
wire n_4977;
wire n_8774;
wire n_2492;
wire n_6976;
wire n_7608;
wire n_7234;
wire n_2939;
wire n_3425;
wire n_4876;
wire n_241;
wire n_5021;
wire n_1449;
wire n_2900;
wire n_797;
wire n_9044;
wire n_2912;
wire n_5936;
wire n_8307;
wire n_595;
wire n_1405;
wire n_3813;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_6784;
wire n_9694;
wire n_1757;
wire n_8470;
wire n_2264;
wire n_1950;
wire n_805;
wire n_5928;
wire n_2032;
wire n_2090;
wire n_7830;
wire n_8050;
wire n_3124;
wire n_3811;
wire n_295;
wire n_4200;
wire n_190;
wire n_2249;
wire n_5785;
wire n_3411;
wire n_5222;
wire n_9633;
wire n_6165;
wire n_10133;
wire n_3463;
wire n_2785;
wire n_730;
wire n_4938;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_6114;
wire n_1856;
wire n_463;
wire n_1524;
wire n_2928;
wire n_5505;
wire n_1118;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_1293;
wire n_961;
wire n_469;
wire n_9261;
wire n_726;
wire n_5504;
wire n_878;
wire n_7348;
wire n_9345;
wire n_4118;
wire n_6829;
wire n_3857;
wire n_3110;
wire n_9375;
wire n_4239;
wire n_9472;
wire n_9764;
wire n_8010;
wire n_3157;
wire n_1180;
wire n_1697;
wire n_2730;
wire n_9448;
wire n_6464;
wire n_8802;
wire n_8950;
wire n_5129;
wire n_806;
wire n_1350;
wire n_7320;
wire n_4704;
wire n_2720;
wire n_649;
wire n_1561;
wire n_8603;
wire n_9487;
wire n_5494;
wire n_5970;
wire n_2405;
wire n_6838;
wire n_2700;
wire n_6368;
wire n_1616;
wire n_7935;
wire n_2416;
wire n_8143;
wire n_2064;
wire n_3640;
wire n_9271;
wire n_5663;
wire n_5161;
wire n_7933;
wire n_1557;
wire n_6640;
wire n_7155;
wire n_9851;
wire n_6166;
wire n_4744;
wire n_5378;
wire n_5626;
wire n_349;
wire n_4706;
wire n_2022;
wire n_3879;
wire n_4343;
wire n_6850;
wire n_1505;
wire n_2408;
wire n_4764;
wire n_5389;
wire n_7743;
wire n_4990;
wire n_2986;
wire n_8584;
wire n_949;
wire n_2454;
wire n_9101;
wire n_6550;
wire n_6656;
wire n_8153;
wire n_6972;
wire n_3591;
wire n_8574;
wire n_198;
wire n_2760;
wire n_4919;
wire n_1208;
wire n_7043;
wire n_7986;
wire n_3317;
wire n_8049;
wire n_9927;
wire n_7266;
wire n_5653;
wire n_4835;
wire n_1151;
wire n_554;
wire n_4420;
wire n_7996;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_354;
wire n_5266;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_5800;
wire n_8509;
wire n_1133;
wire n_883;
wire n_4372;
wire n_5396;
wire n_4097;
wire n_9850;
wire n_4162;
wire n_5766;
wire n_5293;
wire n_779;
wire n_4790;
wire n_594;
wire n_7035;
wire n_4173;
wire n_8354;
wire n_5309;
wire n_6047;
wire n_9432;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_9824;
wire n_422;
wire n_1269;
wire n_8277;
wire n_7442;
wire n_4727;
wire n_1547;
wire n_1438;
wire n_6568;
wire n_3654;
wire n_5627;
wire n_1047;
wire n_3783;
wire n_10055;
wire n_4008;
wire n_2158;
wire n_8583;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_7153;
wire n_8681;
wire n_6258;
wire n_1288;
wire n_8644;
wire n_10148;
wire n_7939;
wire n_9884;
wire n_7715;
wire n_2173;
wire n_3982;
wire n_7350;
wire n_3647;
wire n_7314;
wire n_6026;
wire n_8609;
wire n_1143;
wire n_9144;
wire n_3973;
wire n_8052;
wire n_4799;
wire n_8733;
wire n_9758;
wire n_8082;
wire n_5882;
wire n_6700;
wire n_7136;
wire n_4534;
wire n_5636;
wire n_4960;
wire n_9931;
wire n_7699;
wire n_9693;
wire n_1153;
wire n_9273;
wire n_271;
wire n_465;
wire n_9196;
wire n_1103;
wire n_5707;
wire n_5594;
wire n_9029;
wire n_10086;
wire n_3738;
wire n_894;
wire n_5697;
wire n_1380;
wire n_562;
wire n_2020;
wire n_7580;
wire n_5606;
wire n_6727;
wire n_2310;
wire n_510;
wire n_5911;
wire n_7340;
wire n_8080;
wire n_256;
wire n_3600;
wire n_7303;
wire n_1023;
wire n_9967;
wire n_8819;
wire n_914;
wire n_7870;
wire n_689;
wire n_7568;
wire n_6139;
wire n_7399;
wire n_5382;
wire n_4327;
wire n_7387;
wire n_3190;
wire n_8487;
wire n_3027;
wire n_6454;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_9881;
wire n_2820;
wire n_497;
wire n_3733;
wire n_1165;
wire n_3967;
wire n_6333;
wire n_7004;
wire n_455;
wire n_588;
wire n_638;
wire n_4370;
wire n_5638;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_8382;
wire n_1417;
wire n_9733;
wire n_3096;
wire n_8517;
wire n_7207;
wire n_8827;
wire n_9075;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_7167;
wire n_2234;
wire n_1341;
wire n_5849;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_8906;
wire n_1603;
wire n_5841;
wire n_10109;
wire n_7146;
wire n_7030;
wire n_4478;
wire n_8203;
wire n_413;
wire n_2935;
wire n_9442;
wire n_4246;
wire n_715;
wire n_7618;
wire n_1066;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_685;
wire n_9630;
wire n_4061;
wire n_9898;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_8340;
wire n_4754;
wire n_9582;
wire n_1534;
wire n_8268;
wire n_8171;
wire n_1290;
wire n_4375;
wire n_617;
wire n_9877;
wire n_10179;
wire n_2396;
wire n_3368;
wire n_9986;
wire n_1559;
wire n_8008;
wire n_7633;
wire n_9636;
wire n_3117;
wire n_4684;
wire n_743;
wire n_1546;
wire n_3384;
wire n_5279;
wire n_7159;
wire n_8553;
wire n_2592;
wire n_8824;
wire n_3490;
wire n_7280;
wire n_8369;
wire n_962;
wire n_5043;
wire n_7339;
wire n_7597;
wire n_8884;
wire n_4241;
wire n_1622;
wire n_2751;
wire n_3113;
wire n_9225;
wire n_4183;
wire n_7768;
wire n_918;
wire n_1968;
wire n_5645;
wire n_639;
wire n_6455;
wire n_673;
wire n_5020;
wire n_2842;
wire n_7615;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_10182;
wire n_8271;
wire n_9091;
wire n_3720;
wire n_6183;
wire n_8392;
wire n_8309;
wire n_6107;
wire n_6476;
wire n_5232;
wire n_10046;
wire n_2560;
wire n_9412;
wire n_1164;
wire n_4256;
wire n_8874;
wire n_8228;
wire n_1193;
wire n_1345;
wire n_5035;
wire n_3037;
wire n_1336;
wire n_1033;
wire n_5453;
wire n_4333;
wire n_5339;
wire n_8483;
wire n_6003;
wire n_5443;
wire n_8133;
wire n_7612;
wire n_1166;
wire n_2007;
wire n_3363;
wire n_6636;
wire n_9525;
wire n_1158;
wire n_1803;
wire n_872;
wire n_3522;
wire n_8172;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_6554;
wire n_9575;
wire n_5631;
wire n_3481;
wire n_280;
wire n_6994;
wire n_7401;
wire n_5101;
wire n_9738;
wire n_6020;
wire n_2236;
wire n_9252;
wire n_6185;
wire n_8344;
wire n_692;
wire n_7594;
wire n_7711;
wire n_7321;
wire n_4457;
wire n_223;
wire n_2150;
wire n_8738;
wire n_8936;
wire n_9739;
wire n_6785;
wire n_1816;
wire n_2803;
wire n_9727;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_6870;
wire n_3305;
wire n_6643;
wire n_7574;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_8226;
wire n_6695;
wire n_7529;
wire n_3354;
wire n_5608;
wire n_6501;
wire n_2204;
wire n_9148;
wire n_1481;
wire n_2040;
wire n_6466;
wire n_9958;
wire n_2151;
wire n_2455;
wire n_827;
wire n_3437;
wire n_6467;
wire n_9323;
wire n_2231;
wire n_4212;
wire n_622;
wire n_4584;
wire n_7522;
wire n_7188;
wire n_9779;
wire n_8088;
wire n_5702;
wire n_9545;
wire n_8930;
wire n_9155;
wire n_8662;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_9046;
wire n_9430;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_4477;
wire n_5806;
wire n_4110;
wire n_9625;
wire n_8783;
wire n_8663;
wire n_1221;
wire n_4217;
wire n_5182;
wire n_5277;
wire n_792;
wire n_1262;
wire n_6507;
wire n_1942;
wire n_6618;
wire n_9447;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_6213;
wire n_1579;
wire n_8364;
wire n_9485;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_8490;
wire n_8981;
wire n_229;
wire n_9129;
wire n_923;
wire n_1124;
wire n_7872;
wire n_1326;
wire n_3969;
wire n_6873;
wire n_7958;
wire n_2282;
wire n_4605;
wire n_8118;
wire n_981;
wire n_3873;
wire n_4649;
wire n_5747;
wire n_8671;
wire n_7101;
wire n_8785;
wire n_10210;
wire n_1204;
wire n_7843;
wire n_994;
wire n_2428;
wire n_9047;
wire n_10057;
wire n_1360;
wire n_6063;
wire n_2858;
wire n_3076;
wire n_7578;
wire n_3410;
wire n_5415;
wire n_856;
wire n_7261;
wire n_8982;
wire n_4999;
wire n_4592;
wire n_1564;
wire n_6993;
wire n_9745;
wire n_508;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_8100;
wire n_1858;
wire n_353;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_8522;
wire n_1361;
wire n_8381;
wire n_9320;
wire n_8835;
wire n_6767;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_5687;
wire n_1411;
wire n_1359;
wire n_6558;
wire n_6755;
wire n_9108;
wire n_9457;
wire n_9907;
wire n_6153;
wire n_3536;
wire n_1721;
wire n_7263;
wire n_3782;
wire n_1317;
wire n_6608;
wire n_6202;
wire n_6780;
wire n_7688;
wire n_3594;
wire n_5383;
wire n_2385;
wire n_6635;
wire n_7245;
wire n_7925;
wire n_7310;
wire n_9567;
wire n_294;
wire n_6359;
wire n_5690;
wire n_1980;
wire n_5740;
wire n_7093;
wire n_4177;
wire n_2501;
wire n_7585;
wire n_8356;
wire n_1385;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_9852;
wire n_3855;
wire n_7418;
wire n_6353;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_6577;
wire n_7772;
wire n_8736;
wire n_2028;
wire n_919;
wire n_3114;
wire n_2092;
wire n_6082;
wire n_3622;
wire n_2817;
wire n_2773;
wire n_8918;
wire n_2402;
wire n_1458;
wire n_679;
wire n_220;
wire n_3047;
wire n_3163;
wire n_5361;
wire n_7312;
wire n_9022;
wire n_7514;
wire n_1550;
wire n_1358;
wire n_8616;
wire n_1200;
wire n_6105;
wire n_387;
wire n_826;
wire n_5512;
wire n_7738;
wire n_2808;
wire n_2344;
wire n_8838;
wire n_8908;
wire n_3520;
wire n_2392;
wire n_7609;
wire n_9161;
wire n_3272;
wire n_3122;
wire n_5898;
wire n_7113;
wire n_6548;
wire n_8607;
wire n_607;
wire n_8213;
wire n_5923;
wire n_3687;
wire n_2787;
wire n_6657;
wire n_5617;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_5946;
wire n_1268;
wire n_2676;
wire n_9903;
wire n_9831;
wire n_10032;
wire n_8436;
wire n_7282;
wire n_372;
wire n_8551;
wire n_2770;
wire n_4550;
wire n_9238;
wire n_4347;
wire n_7921;
wire n_702;
wire n_5193;
wire n_4933;
wire n_968;
wire n_4144;
wire n_9248;
wire n_5514;
wire n_5611;
wire n_2375;
wire n_3278;
wire n_5579;
wire n_4167;
wire n_6380;
wire n_3608;
wire n_4895;
wire n_9867;
wire n_1282;
wire n_6163;
wire n_7170;
wire n_4726;
wire n_10005;
wire n_5573;
wire n_5143;
wire n_5836;
wire n_1755;
wire n_5188;
wire n_6674;
wire n_5049;
wire n_2212;
wire n_7489;
wire n_9056;
wire n_6331;
wire n_5308;
wire n_9106;
wire n_311;
wire n_4434;
wire n_5068;
wire n_7863;
wire n_6493;
wire n_7363;
wire n_7281;
wire n_5739;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_7968;
wire n_10061;
wire n_6023;
wire n_7820;
wire n_8437;
wire n_269;
wire n_816;
wire n_7833;
wire n_1322;
wire n_3829;
wire n_4510;
wire n_7750;
wire n_5057;
wire n_446;
wire n_9071;
wire n_6196;
wire n_5425;
wire n_5273;
wire n_10136;
wire n_5839;
wire n_2469;
wire n_7588;
wire n_1125;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_7697;
wire n_10025;
wire n_5887;
wire n_7808;
wire n_3068;
wire n_9519;
wire n_1629;
wire n_9027;
wire n_7603;
wire n_1094;
wire n_6321;
wire n_5683;
wire n_1510;
wire n_8704;
wire n_3002;
wire n_8984;
wire n_9786;
wire n_10194;
wire n_7192;
wire n_1099;
wire n_5248;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_759;
wire n_567;
wire n_4156;
wire n_8613;
wire n_1727;
wire n_3693;
wire n_5880;
wire n_8012;
wire n_3132;
wire n_5002;
wire n_5487;
wire n_5649;
wire n_8881;
wire n_5531;
wire n_9404;
wire n_831;
wire n_3681;
wire n_5666;
wire n_3970;
wire n_778;
wire n_2351;
wire n_1619;
wire n_7988;
wire n_550;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_6824;
wire n_6954;
wire n_8763;
wire n_6450;
wire n_9370;
wire n_1152;
wire n_6995;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_1236;
wire n_4579;
wire n_6347;
wire n_6496;
wire n_4776;
wire n_671;
wire n_8387;
wire n_9352;
wire n_8105;
wire n_10144;
wire n_2704;
wire n_1334;
wire n_6745;
wire n_7943;
wire n_3729;
wire n_6698;
wire n_4471;
wire n_6968;
wire n_7377;
wire n_8900;
wire n_4392;
wire n_3103;
wire n_488;
wire n_6064;
wire n_9681;
wire n_8353;
wire n_505;
wire n_9051;
wire n_2048;
wire n_7723;
wire n_498;
wire n_3028;
wire n_4691;
wire n_7904;
wire n_3148;
wire n_3775;
wire n_5682;
wire n_684;
wire n_5461;
wire n_9098;
wire n_7296;
wire n_3966;
wire n_4397;
wire n_8323;
wire n_6164;
wire n_8711;
wire n_3616;
wire n_4753;
wire n_9484;
wire n_4803;
wire n_8731;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_5730;
wire n_10155;
wire n_6292;
wire n_7759;
wire n_6743;
wire n_4165;
wire n_2056;
wire n_5754;
wire n_2852;
wire n_8597;
wire n_2515;
wire n_6330;
wire n_1600;
wire n_1144;
wire n_7178;
wire n_838;
wire n_1941;
wire n_7045;
wire n_175;
wire n_3637;
wire n_9853;
wire n_8534;
wire n_1017;
wire n_8655;
wire n_9210;
wire n_734;
wire n_4893;
wire n_2240;
wire n_7777;
wire n_8302;
wire n_4258;
wire n_5756;
wire n_310;
wire n_8496;
wire n_7693;
wire n_709;
wire n_2917;
wire n_3194;
wire n_2085;
wire n_2432;
wire n_10156;
wire n_5033;
wire n_6015;
wire n_1686;
wire n_6408;
wire n_4232;
wire n_5075;
wire n_8078;
wire n_2097;
wire n_662;
wire n_3461;
wire n_10215;
wire n_7682;
wire n_7300;
wire n_939;
wire n_1410;
wire n_2297;
wire n_6861;
wire n_10152;
wire n_4203;
wire n_9756;
wire n_5789;
wire n_5400;
wire n_1325;
wire n_7558;
wire n_1223;
wire n_5347;
wire n_2957;
wire n_572;
wire n_9166;
wire n_8103;
wire n_8719;
wire n_1983;
wire n_7798;
wire n_9778;
wire n_8879;
wire n_4767;
wire n_8969;
wire n_9141;
wire n_4569;
wire n_948;
wire n_448;
wire n_6528;
wire n_9700;
wire n_8896;
wire n_3820;
wire n_5144;
wire n_6895;
wire n_3072;
wire n_8335;
wire n_2961;
wire n_4468;
wire n_5509;
wire n_1923;
wire n_3848;
wire n_7400;
wire n_3631;
wire n_7393;
wire n_6590;
wire n_8116;
wire n_6523;
wire n_5169;
wire n_4885;
wire n_7475;
wire n_1479;
wire n_9363;
wire n_4698;
wire n_1031;
wire n_3674;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_5349;
wire n_6472;
wire n_9532;
wire n_3763;
wire n_933;
wire n_6389;
wire n_3499;
wire n_5534;
wire n_1821;
wire n_9307;
wire n_9876;
wire n_3947;
wire n_3910;
wire n_492;
wire n_252;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_2995;
wire n_6073;
wire n_4533;
wire n_4287;
wire n_8462;
wire n_9959;
wire n_3228;
wire n_8834;
wire n_9989;
wire n_8417;
wire n_8286;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_8964;
wire n_1186;
wire n_6869;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_7672;
wire n_4556;
wire n_6137;
wire n_9467;
wire n_2205;
wire n_2183;
wire n_389;
wire n_1724;
wire n_3088;
wire n_1707;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_1126;
wire n_5079;
wire n_8247;
wire n_2761;
wire n_2357;
wire n_9406;
wire n_10089;
wire n_4520;
wire n_895;
wire n_8639;
wire n_1639;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_9160;
wire n_5751;
wire n_626;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_7712;
wire n_6885;
wire n_7681;
wire n_8566;
wire n_1818;
wire n_6580;
wire n_6613;
wire n_8727;
wire n_5039;
wire n_4265;
wire n_8482;
wire n_6404;
wire n_6120;
wire n_3557;
wire n_1598;
wire n_2269;
wire n_7491;
wire n_265;
wire n_1583;
wire n_10094;
wire n_8599;
wire n_4612;
wire n_5997;
wire n_8781;
wire n_5375;
wire n_5438;
wire n_9167;
wire n_7150;
wire n_7954;
wire n_7974;
wire n_1264;
wire n_6530;
wire n_6602;
wire n_7915;
wire n_4958;
wire n_1827;
wire n_4149;
wire n_6135;
wire n_246;
wire n_8839;
wire n_1752;
wire n_2361;
wire n_4538;
wire n_3030;
wire n_3505;
wire n_5563;
wire n_3075;
wire n_8365;
wire n_1102;
wire n_2239;
wire n_6942;
wire n_7860;
wire n_6892;
wire n_1296;
wire n_4730;
wire n_7357;
wire n_8112;
wire n_8489;
wire n_8859;
wire n_8060;
wire n_9290;
wire n_6782;
wire n_4421;
wire n_6230;
wire n_2464;
wire n_3697;
wire n_882;
wire n_8244;
wire n_2304;
wire n_2514;
wire n_6977;
wire n_7229;
wire n_8096;
wire n_7336;
wire n_5932;
wire n_289;
wire n_6598;
wire n_10105;
wire n_6795;
wire n_6121;
wire n_457;
wire n_1299;
wire n_3430;
wire n_5919;
wire n_2063;
wire n_8346;
wire n_3489;
wire n_5012;
wire n_6614;
wire n_6506;
wire n_2079;
wire n_9705;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_8367;
wire n_9113;
wire n_3484;
wire n_6001;
wire n_411;
wire n_4971;
wire n_9521;
wire n_9682;
wire n_2095;
wire n_7493;
wire n_9278;
wire n_5664;
wire n_2738;
wire n_6406;
wire n_5890;
wire n_2590;
wire n_4661;
wire n_2797;
wire n_357;
wire n_3041;
wire n_412;
wire n_8898;
wire n_8658;
wire n_5823;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_5944;
wire n_8905;
wire n_5422;
wire n_9222;
wire n_6989;
wire n_8145;
wire n_8237;
wire n_6299;
wire n_9813;
wire n_7424;
wire n_10216;
wire n_5246;
wire n_8562;
wire n_4376;
wire n_9863;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_9394;
wire n_10170;
wire n_1069;
wire n_4305;
wire n_2037;
wire n_2953;
wire n_573;
wire n_2823;
wire n_7273;
wire n_9663;
wire n_7901;
wire n_3684;
wire n_5725;
wire n_10146;
wire n_5404;
wire n_913;
wire n_10175;
wire n_1681;
wire n_4834;
wire n_9994;
wire n_1507;
wire n_5332;
wire n_7149;
wire n_9723;
wire n_589;
wire n_2866;
wire n_7116;
wire n_3153;
wire n_1174;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_8211;
wire n_3268;
wire n_2559;
wire n_8537;
wire n_8946;
wire n_5616;
wire n_1383;
wire n_603;
wire n_8055;
wire n_373;
wire n_4259;
wire n_7909;
wire n_5870;
wire n_2030;
wire n_6053;
wire n_850;
wire n_6233;
wire n_4299;
wire n_5625;
wire n_245;
wire n_319;
wire n_6758;
wire n_2407;
wire n_690;
wire n_9069;
wire n_5367;
wire n_525;
wire n_2243;
wire n_6629;
wire n_5288;
wire n_2694;
wire n_6356;
wire n_8332;
wire n_5601;
wire n_3742;
wire n_7601;
wire n_8998;
wire n_4965;
wire n_1837;
wire n_7033;
wire n_6010;
wire n_4178;
wire n_189;
wire n_8157;
wire n_2006;
wire n_9284;
wire n_4953;
wire n_8484;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_7147;
wire n_7596;
wire n_9556;
wire n_5294;
wire n_8161;
wire n_5570;
wire n_6411;
wire n_9337;
wire n_2731;
wire n_3703;
wire n_5411;
wire n_5670;
wire n_1246;
wire n_9211;
wire n_5265;
wire n_7549;
wire n_5955;
wire n_2123;
wire n_2238;
wire n_4802;
wire n_4793;
wire n_6032;
wire n_1196;
wire n_5733;
wire n_8692;
wire n_3435;
wire n_410;
wire n_2380;
wire n_1187;
wire n_4897;
wire n_9243;
wire n_6918;
wire n_1298;
wire n_1745;
wire n_9773;
wire n_4674;
wire n_8812;
wire n_568;
wire n_8682;
wire n_4796;
wire n_8290;
wire n_1088;
wire n_7138;
wire n_766;
wire n_6401;
wire n_7279;
wire n_7976;
wire n_5184;
wire n_377;
wire n_9928;
wire n_2750;
wire n_8890;
wire n_2547;
wire n_8747;
wire n_7617;
wire n_279;
wire n_945;
wire n_4575;
wire n_9784;
wire n_3665;
wire n_3063;
wire n_8062;
wire n_3281;
wire n_7137;
wire n_3535;
wire n_5061;
wire n_2288;
wire n_3858;
wire n_7700;
wire n_4653;
wire n_8275;
wire n_7474;
wire n_4589;
wire n_7124;
wire n_5978;
wire n_6853;
wire n_8667;
wire n_3220;
wire n_4581;
wire n_9192;
wire n_6008;
wire n_500;
wire n_665;
wire n_4625;
wire n_7098;
wire n_6181;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_9134;
wire n_3679;
wire n_738;
wire n_5575;
wire n_6654;
wire n_7661;
wire n_672;
wire n_4968;
wire n_7801;
wire n_8807;
wire n_9975;
wire n_9765;
wire n_6907;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_3856;
wire n_4038;
wire n_7876;
wire n_5316;
wire n_2735;
wire n_953;
wire n_4214;
wire n_143;
wire n_1888;
wire n_5290;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_557;
wire n_3419;
wire n_7323;
wire n_989;
wire n_5048;
wire n_2233;
wire n_5363;
wire n_5665;
wire n_6517;
wire n_795;
wire n_4892;
wire n_6339;
wire n_1936;
wire n_9564;
wire n_9127;
wire n_3890;
wire n_6170;
wire n_7247;
wire n_6394;
wire n_8048;
wire n_821;
wire n_770;
wire n_5607;
wire n_1514;
wire n_7929;
wire n_486;
wire n_2782;
wire n_569;
wire n_3929;
wire n_9306;
wire n_971;
wire n_4353;
wire n_2201;
wire n_8212;
wire n_4950;
wire n_1650;
wire n_7755;
wire n_6504;
wire n_9891;
wire n_10022;
wire n_4176;
wire n_9078;
wire n_7556;
wire n_222;
wire n_4124;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_5462;
wire n_6814;
wire n_7216;
wire n_4488;
wire n_10127;
wire n_5278;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_9332;
wire n_3756;
wire n_8043;
wire n_8223;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_8159;
wire n_8868;
wire n_5845;
wire n_9889;
wire n_4608;
wire n_9294;
wire n_6691;
wire n_432;
wire n_293;
wire n_3948;
wire n_4839;
wire n_9174;
wire n_1074;
wire n_5969;
wire n_1765;
wire n_9132;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_206;
wire n_2332;
wire n_9547;
wire n_2391;
wire n_6343;
wire n_6005;
wire n_611;
wire n_1295;
wire n_2060;
wire n_3883;
wire n_1013;
wire n_6686;
wire n_4032;
wire n_2571;
wire n_136;
wire n_6437;
wire n_5736;
wire n_4929;
wire n_2874;
wire n_6029;
wire n_6536;
wire n_6684;
wire n_4117;
wire n_300;
wire n_6025;
wire n_3049;
wire n_8434;
wire n_3634;
wire n_5436;
wire n_7962;
wire n_2341;
wire n_1654;
wire n_6697;
wire n_3066;
wire n_2045;
wire n_10122;
wire n_6085;
wire n_3913;
wire n_9762;
wire n_5341;
wire n_8608;
wire n_2575;
wire n_3739;
wire n_1230;
wire n_5140;
wire n_376;
wire n_1597;
wire n_2942;
wire n_6062;
wire n_1771;
wire n_4541;
wire n_6715;
wire n_3271;
wire n_3164;
wire n_8656;
wire n_3861;
wire n_5096;
wire n_9183;
wire n_2043;
wire n_6771;
wire n_7905;
wire n_4171;
wire n_5847;
wire n_7204;
wire n_9461;
wire n_9117;
wire n_7022;
wire n_6383;
wire n_4815;
wire n_5639;
wire n_4665;
wire n_6877;
wire n_7308;
wire n_7476;
wire n_10116;
wire n_4884;
wire n_3580;
wire n_1437;
wire n_8249;
wire n_4276;
wire n_1378;
wire n_5268;
wire n_5050;
wire n_9062;
wire n_209;
wire n_5503;
wire n_5240;
wire n_1461;
wire n_5718;
wire n_7208;
wire n_9915;
wire n_7718;
wire n_1876;
wire n_1830;
wire n_5001;
wire n_6567;
wire n_503;
wire n_5658;
wire n_1112;
wire n_700;
wire n_4174;
wire n_9001;
wire n_6868;
wire n_7290;
wire n_5131;
wire n_9081;
wire n_6813;
wire n_7756;
wire n_5546;
wire n_9156;
wire n_6294;
wire n_7795;
wire n_7822;
wire n_8717;
wire n_10159;
wire n_5174;
wire n_9024;
wire n_9198;
wire n_10178;
wire n_2145;
wire n_4801;
wire n_6079;
wire n_6260;
wire n_680;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_6520;
wire n_7623;
wire n_380;
wire n_3119;
wire n_6671;
wire n_9335;
wire n_4740;
wire n_1108;
wire n_9488;
wire n_1274;
wire n_7632;
wire n_4394;
wire n_257;
wire n_5544;
wire n_6444;
wire n_6637;
wire n_9725;
wire n_8842;
wire n_475;
wire n_6729;
wire n_5660;
wire n_6958;
wire n_8073;
wire n_10185;
wire n_9526;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_5541;
wire n_6314;
wire n_577;
wire n_5610;
wire n_407;
wire n_9962;
wire n_8576;
wire n_916;
wire n_2810;
wire n_6703;
wire n_1884;
wire n_1555;
wire n_8799;
wire n_762;
wire n_1468;
wire n_1253;
wire n_4378;
wire n_9667;
wire n_5166;
wire n_2683;
wire n_6065;
wire n_7265;
wire n_4180;
wire n_4459;
wire n_6878;
wire n_3624;
wire n_6725;
wire n_8181;
wire n_5808;
wire n_1182;
wire n_6527;
wire n_4594;
wire n_8447;
wire n_8045;
wire n_7289;
wire n_7538;
wire n_2748;
wire n_4642;
wire n_9716;
wire n_6913;
wire n_1376;
wire n_7473;
wire n_7242;
wire n_9253;
wire n_6533;
wire n_513;
wire n_179;
wire n_7164;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_8022;
wire n_3544;
wire n_6845;
wire n_8227;
wire n_5300;
wire n_7853;
wire n_2072;
wire n_3852;
wire n_5233;
wire n_5381;
wire n_436;
wire n_9796;
wire n_5770;
wire n_7483;
wire n_8756;
wire n_5710;
wire n_10021;
wire n_324;
wire n_9953;
wire n_1491;
wire n_2628;
wire n_7389;
wire n_3219;
wire n_10053;
wire n_274;
wire n_1083;
wire n_5333;
wire n_5799;
wire n_6265;
wire n_4914;
wire n_8604;
wire n_8809;
wire n_8976;
wire n_3510;
wire n_7046;
wire n_7834;
wire n_4587;
wire n_1139;
wire n_3688;
wire n_8940;
wire n_5008;
wire n_1312;
wire n_9077;
wire n_3871;
wire n_892;
wire n_3757;
wire n_1567;
wire n_563;
wire n_2219;
wire n_8844;
wire n_6148;
wire n_8995;
wire n_2100;
wire n_8255;
wire n_3666;
wire n_5538;
wire n_990;
wire n_6357;
wire n_867;
wire n_8216;
wire n_8693;
wire n_3479;
wire n_944;
wire n_5499;
wire n_749;
wire n_9123;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_7811;
wire n_6522;
wire n_8669;
wire n_7097;
wire n_4285;
wire n_7000;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_650;
wire n_3741;
wire n_9922;
wire n_5582;
wire n_2567;
wire n_9177;
wire n_2557;
wire n_1908;
wire n_5675;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_7880;
wire n_5109;
wire n_712;
wire n_8769;
wire n_9463;
wire n_909;
wire n_6713;
wire n_8149;
wire n_1392;
wire n_10067;
wire n_2066;
wire n_5281;
wire n_2762;
wire n_6087;
wire n_964;
wire n_7851;
wire n_2220;
wire n_7342;
wire n_7044;
wire n_7810;
wire n_10135;
wire n_6108;
wire n_7664;
wire n_6100;
wire n_6800;
wire n_7364;
wire n_6866;
wire n_7114;
wire n_6373;
wire n_4433;
wire n_2829;
wire n_7332;
wire n_8990;
wire n_5862;
wire n_471;
wire n_7477;
wire n_1914;
wire n_8208;
wire n_2253;
wire n_7468;
wire n_5886;
wire n_9451;
wire n_7714;
wire n_7899;
wire n_8710;
wire n_6415;
wire n_8479;
wire n_6783;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_8512;
wire n_9843;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_9710;
wire n_2507;
wire n_1633;
wire n_9087;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_2328;
wire n_7845;
wire n_347;
wire n_2434;
wire n_183;
wire n_1234;
wire n_3936;
wire n_479;
wire n_5564;
wire n_2261;
wire n_9956;
wire n_3082;
wire n_9079;
wire n_5162;
wire n_5442;
wire n_2473;
wire n_5802;
wire n_9782;
wire n_10049;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_6340;
wire n_9950;
wire n_7858;
wire n_3867;
wire n_3397;
wire n_6103;
wire n_1646;
wire n_6392;
wire n_6513;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_9197;
wire n_1237;
wire n_6720;
wire n_5883;
wire n_9140;
wire n_8401;
wire n_1095;
wire n_3078;
wire n_6078;
wire n_3971;
wire n_370;
wire n_7680;
wire n_5630;
wire n_6666;
wire n_286;
wire n_9364;
wire n_9452;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_9362;
wire n_9398;
wire n_1531;
wire n_2113;
wire n_6815;
wire n_9203;
wire n_1387;
wire n_6207;
wire n_6381;
wire n_3711;
wire n_9712;
wire n_9536;
wire n_8450;
wire n_9848;
wire n_5054;
wire n_6571;
wire n_3171;
wire n_5929;
wire n_9460;
wire n_7710;
wire n_8788;
wire n_5394;
wire n_8324;
wire n_5975;
wire n_4751;
wire n_4242;
wire n_9841;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_9772;
wire n_1496;
wire n_10147;
wire n_2812;
wire n_9057;
wire n_3300;
wire n_7061;
wire n_8104;
wire n_7066;
wire n_9068;
wire n_5496;
wire n_7485;
wire n_3104;
wire n_7174;
wire n_8014;
wire n_4122;
wire n_6661;
wire n_2132;
wire n_4522;
wire n_5991;
wire n_8623;
wire n_4952;
wire n_9634;
wire n_6967;
wire n_4426;
wire n_5956;
wire n_5699;
wire n_4362;
wire n_3267;
wire n_6017;
wire n_9348;
wire n_3946;
wire n_5920;
wire n_2112;
wire n_2640;
wire n_6125;
wire n_8651;
wire n_5000;
wire n_9632;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_9257;
wire n_4089;
wire n_9500;
wire n_3513;
wire n_1173;
wire n_3498;
wire n_5132;
wire n_9747;
wire n_2350;
wire n_9470;
wire n_6414;
wire n_5535;
wire n_1068;
wire n_1198;
wire n_4506;
wire n_6097;
wire n_7783;
wire n_7662;
wire n_6057;
wire n_6936;
wire n_10188;
wire n_9591;
wire n_9049;
wire n_487;
wire n_4728;
wire n_7171;
wire n_7990;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_7003;
wire n_8137;
wire n_2187;
wire n_1413;
wire n_8413;
wire n_2481;
wire n_3863;
wire n_6302;
wire n_2327;
wire n_158;
wire n_3882;
wire n_9471;
wire n_3916;
wire n_6922;
wire n_1365;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_405;
wire n_3332;
wire n_8300;
wire n_8069;
wire n_7501;
wire n_320;
wire n_9409;
wire n_6432;
wire n_7984;
wire n_2055;
wire n_2998;
wire n_7366;
wire n_1423;
wire n_8173;
wire n_4359;
wire n_481;
wire n_1609;
wire n_2822;
wire n_2308;
wire n_1939;
wire n_2242;
wire n_7589;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_218;
wire n_6880;
wire n_6223;
wire n_5176;
wire n_9832;
wire n_4039;
wire n_5793;
wire n_6926;
wire n_1798;
wire n_8091;
wire n_3057;
wire n_1608;
wire n_5761;
wire n_6699;
wire n_547;
wire n_439;
wire n_677;
wire n_3983;
wire n_9067;
wire n_8254;
wire n_703;
wire n_8400;
wire n_10141;
wire n_3318;
wire n_7232;
wire n_3385;
wire n_9858;
wire n_7511;
wire n_326;
wire n_227;
wire n_3773;
wire n_3494;
wire n_9482;
wire n_1278;
wire n_9033;
wire n_6957;
wire n_5074;
wire n_7917;
wire n_3939;
wire n_3788;
wire n_590;
wire n_727;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_8368;
wire n_6694;
wire n_545;
wire n_9247;
wire n_2496;
wire n_3260;
wire n_8463;
wire n_536;
wire n_9965;
wire n_3349;
wire n_6449;
wire n_4348;
wire n_1602;
wire n_7422;
wire n_9299;
wire n_3139;
wire n_8889;
wire n_427;
wire n_3801;
wire n_5681;
wire n_9244;
wire n_9785;
wire n_2338;
wire n_5261;
wire n_1080;
wire n_9195;
wire n_8322;
wire n_3636;
wire n_6591;
wire n_7466;
wire n_8987;
wire n_3653;
wire n_3823;
wire n_9280;
wire n_3403;
wire n_7621;
wire n_9911;
wire n_8274;
wire n_2057;
wire n_6594;
wire n_6342;
wire n_1205;
wire n_6195;
wire n_163;
wire n_2716;
wire n_6441;
wire n_7572;
wire n_7158;
wire n_314;
wire n_2944;
wire n_2780;
wire n_3439;
wire n_1120;
wire n_7500;
wire n_1202;
wire n_4084;
wire n_627;
wire n_7985;
wire n_9687;
wire n_1371;
wire n_4240;
wire n_8657;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_233;
wire n_8954;
wire n_2774;
wire n_6354;
wire n_2799;
wire n_8311;
wire n_5748;
wire n_4393;
wire n_321;
wire n_6662;
wire n_7494;
wire n_9088;
wire n_3984;
wire n_1586;
wire n_8728;
wire n_9580;
wire n_9569;
wire n_1431;
wire n_8994;
wire n_4389;
wire n_6433;
wire n_9680;
wire n_1763;
wire n_8398;
wire n_6200;
wire n_5641;
wire n_8407;
wire n_8071;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_6902;
wire n_4615;
wire n_3044;
wire n_3492;
wire n_7197;
wire n_3737;
wire n_6369;
wire n_8528;
wire n_9227;
wire n_5657;
wire n_8475;
wire n_297;
wire n_9951;
wire n_9855;
wire n_2379;
wire n_3579;
wire n_9072;
wire n_10102;
wire n_1667;
wire n_888;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_1677;
wire n_5244;
wire n_5765;
wire n_5114;
wire n_9054;
wire n_4551;
wire n_178;
wire n_10117;
wire n_551;
wire n_4521;
wire n_6956;
wire n_10126;
wire n_7587;
wire n_2284;
wire n_6451;
wire n_3005;
wire n_7704;
wire n_5420;
wire n_6497;
wire n_8511;
wire n_7865;
wire n_2283;
wire n_5206;
wire n_582;
wire n_2526;
wire n_1097;
wire n_1711;
wire n_4387;
wire n_9584;
wire n_9287;
wire n_534;
wire n_2508;
wire n_3186;
wire n_9459;
wire n_6701;
wire n_2594;
wire n_1239;
wire n_9490;
wire n_5298;
wire n_10209;
wire n_8867;
wire n_3417;
wire n_8246;
wire n_560;
wire n_8558;
wire n_890;
wire n_9655;
wire n_9846;
wire n_3626;
wire n_451;
wire n_9593;
wire n_4598;
wire n_4464;
wire n_8925;
wire n_5106;
wire n_7881;
wire n_9147;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_1081;
wire n_9678;
wire n_2119;
wire n_8641;
wire n_9658;
wire n_2493;
wire n_9560;
wire n_9578;
wire n_5080;
wire n_535;
wire n_9396;
wire n_4565;
wire n_7032;
wire n_9303;
wire n_3392;
wire n_1800;
wire n_7198;
wire n_6884;
wire n_7752;
wire n_5081;
wire n_8201;
wire n_6921;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_7953;
wire n_6106;
wire n_6876;
wire n_3512;
wire n_9553;
wire n_1734;
wire n_1860;
wire n_8046;
wire n_4552;
wire n_7193;
wire n_6287;
wire n_2840;
wire n_6172;
wire n_9942;
wire n_9805;
wire n_4482;
wire n_837;
wire n_812;
wire n_4172;
wire n_5957;
wire n_4040;
wire n_8414;
wire n_3024;
wire n_5567;
wire n_8292;
wire n_9138;
wire n_9879;
wire n_5406;
wire n_8647;
wire n_6362;
wire n_9213;
wire n_4328;
wire n_8543;
wire n_1854;
wire n_666;
wire n_5191;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_6067;
wire n_2893;
wire n_6833;
wire n_4940;
wire n_9374;
wire n_785;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_8331;
wire n_999;
wire n_2280;
wire n_8317;
wire n_7126;
wire n_5867;
wire n_456;
wire n_1394;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_7496;
wire n_6430;
wire n_9179;
wire n_873;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_6296;
wire n_10014;
wire n_4112;
wire n_342;
wire n_5602;
wire n_2035;
wire n_7196;
wire n_4928;
wire n_2614;
wire n_7360;
wire n_5428;
wire n_6325;
wire n_2494;
wire n_1538;
wire n_4865;
wire n_6678;
wire n_7982;
wire n_2128;
wire n_4071;
wire n_6564;
wire n_7268;
wire n_8187;
wire n_8174;
wire n_8929;
wire n_10108;
wire n_4436;
wire n_5786;
wire n_5822;
wire n_3586;
wire n_8846;
wire n_5817;
wire n_9277;
wire n_4160;
wire n_6109;
wire n_9611;
wire n_6385;
wire n_1668;
wire n_9744;
wire n_5798;
wire n_10123;
wire n_4137;
wire n_1078;
wire n_8032;
wire n_9504;
wire n_5417;
wire n_10048;
wire n_4545;
wire n_8200;
wire n_4758;
wire n_1161;
wire n_8036;
wire n_9285;
wire n_4840;
wire n_5713;
wire n_9905;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_9190;
wire n_8586;
wire n_8524;
wire n_618;
wire n_1191;
wire n_4535;
wire n_7518;
wire n_8828;
wire n_9639;
wire n_4385;
wire n_7779;
wire n_9664;
wire n_1215;
wire n_3748;
wire n_4731;
wire n_7575;
wire n_2337;
wire n_7073;
wire n_8092;
wire n_1786;
wire n_6309;
wire n_8370;
wire n_3732;
wire n_9109;
wire n_211;
wire n_1804;
wire n_10189;
wire n_408;
wire n_8135;
wire n_6519;
wire n_4671;
wire n_9741;
wire n_2272;
wire n_5571;
wire n_4766;
wire n_5989;
wire n_592;
wire n_4558;
wire n_1318;
wire n_8764;
wire n_1632;
wire n_1769;
wire n_7349;
wire n_1929;
wire n_9875;
wire n_8502;
wire n_4319;
wire n_9360;
wire n_6585;
wire n_7786;
wire n_9021;
wire n_8454;
wire n_2929;
wire n_4358;
wire n_9122;
wire n_1526;
wire n_7579;
wire n_10099;
wire n_7122;
wire n_10193;
wire n_4874;
wire n_180;
wire n_2656;
wire n_4904;
wire n_516;
wire n_1997;
wire n_10203;
wire n_10140;
wire n_1137;
wire n_1258;
wire n_640;
wire n_1733;
wire n_6490;
wire n_7867;
wire n_4651;
wire n_10149;
wire n_943;
wire n_3167;
wire n_4748;
wire n_7624;
wire n_9803;
wire n_1807;
wire n_1123;
wire n_8776;
wire n_2857;
wire n_8564;
wire n_8343;
wire n_7828;
wire n_1784;
wire n_4618;
wire n_6721;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_8718;
wire n_752;
wire n_985;
wire n_5506;
wire n_7543;
wire n_9659;
wire n_8042;
wire n_5475;
wire n_7727;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_9013;
wire n_1352;
wire n_5908;
wire n_5431;
wire n_9427;
wire n_8379;
wire n_643;
wire n_8034;
wire n_226;
wire n_7778;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_7019;
wire n_682;
wire n_9126;
wire n_5315;
wire n_2633;
wire n_3708;
wire n_5752;
wire n_2907;
wire n_8441;
wire n_9474;
wire n_1429;
wire n_2353;
wire n_7702;
wire n_2528;
wire n_1778;
wire n_5746;
wire n_686;
wire n_1154;
wire n_584;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_1130;
wire n_9538;
wire n_3718;
wire n_6685;
wire n_756;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_8569;
wire n_9574;
wire n_4666;
wire n_4082;
wire n_2320;
wire n_3140;
wire n_979;
wire n_8592;
wire n_8865;
wire n_3976;
wire n_2813;
wire n_897;
wire n_2546;
wire n_3381;
wire n_7952;
wire n_7347;
wire n_9450;
wire n_3736;
wire n_10031;
wire n_4466;
wire n_6016;
wire n_9998;
wire n_891;
wire n_885;
wire n_1659;
wire n_3955;
wire n_5366;
wire n_5322;
wire n_1864;
wire n_5414;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_7791;
wire n_6971;
wire n_8362;
wire n_3336;
wire n_8632;
wire n_10035;
wire n_7739;
wire n_396;
wire n_7945;
wire n_9372;
wire n_9045;
wire n_8361;
wire n_9657;
wire n_7656;
wire n_5903;
wire n_7199;
wire n_10107;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_714;
wire n_3605;
wire n_5307;
wire n_2170;
wire n_4721;
wire n_9904;
wire n_9924;
wire n_9159;
wire n_8561;
wire n_6549;
wire n_725;
wire n_8611;
wire n_9326;
wire n_8410;
wire n_1577;
wire n_5003;
wire n_3840;
wire n_6540;
wire n_7166;
wire n_2198;
wire n_6658;
wire n_5369;
wire n_9476;
wire n_6683;
wire n_3067;
wire n_154;
wire n_3809;
wire n_4921;
wire n_473;
wire n_1852;
wire n_801;
wire n_5912;
wire n_5745;
wire n_7923;
wire n_6086;
wire n_4377;
wire n_818;
wire n_10050;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_5803;
wire n_6327;
wire n_8878;
wire n_5593;
wire n_5270;
wire n_5853;
wire n_6171;
wire n_3468;
wire n_5779;
wire n_1877;
wire n_272;
wire n_8492;
wire n_9301;
wire n_7213;
wire n_5313;
wire n_4301;
wire n_2133;
wire n_8888;
wire n_6820;
wire n_2497;
wire n_879;
wire n_5446;
wire n_7610;
wire n_7107;
wire n_4561;
wire n_1541;
wire n_597;
wire n_3291;
wire n_7456;
wire n_9382;
wire n_8095;
wire n_9921;
wire n_7369;
wire n_1472;
wire n_9325;
wire n_1050;
wire n_9945;
wire n_9643;
wire n_7548;
wire n_2578;
wire n_152;
wire n_1201;
wire n_8735;
wire n_7598;
wire n_1185;
wire n_2475;
wire n_7250;
wire n_8808;
wire n_9201;
wire n_8902;
wire n_7823;
wire n_9771;
wire n_8833;
wire n_4715;
wire n_6157;
wire n_8796;
wire n_2715;
wire n_335;
wire n_2665;
wire n_4879;
wire n_344;
wire n_8794;
wire n_5044;
wire n_210;
wire n_1090;
wire n_4536;
wire n_3755;
wire n_9274;
wire n_9894;
wire n_8549;
wire n_6676;
wire n_4304;
wire n_10095;
wire n_4927;
wire n_4078;
wire n_5459;
wire n_224;
wire n_10088;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_7525;
wire n_4418;
wire n_7924;
wire n_3341;
wire n_9232;
wire n_8690;
wire n_4125;
wire n_5390;
wire n_5351;
wire n_5267;
wire n_1116;
wire n_5024;
wire n_7012;
wire n_3043;
wire n_2747;
wire n_1511;
wire n_8593;
wire n_276;
wire n_9649;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_538;
wire n_2845;
wire n_4151;
wire n_4412;
wire n_2036;
wire n_6923;
wire n_7649;
wire n_843;
wire n_8009;
wire n_8588;
wire n_8195;
wire n_9839;
wire n_3358;
wire n_6704;
wire n_7634;
wire n_9090;
wire n_2003;
wire n_2533;
wire n_1307;
wire n_7406;
wire n_4682;
wire n_1128;
wire n_9346;
wire n_6673;
wire n_9696;
wire n_2419;
wire n_2330;
wire n_9996;
wire n_6534;
wire n_9968;
wire n_8805;
wire n_5078;
wire n_4810;
wire n_7659;
wire n_6162;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_6127;
wire n_1955;
wire n_3289;
wire n_4855;
wire n_9383;
wire n_9498;
wire n_1440;
wire n_6246;
wire n_1370;
wire n_305;
wire n_9836;
wire n_5005;
wire n_6126;
wire n_7372;
wire n_8596;
wire n_9938;
wire n_1549;
wire n_7427;
wire n_6151;
wire n_6828;
wire n_6841;
wire n_10206;
wire n_7844;
wire n_5207;
wire n_7934;
wire n_361;
wire n_2658;
wire n_5624;
wire n_10092;
wire n_3620;
wire n_4601;
wire n_1065;
wire n_4518;
wire n_2767;
wire n_5474;
wire n_7009;
wire n_3376;
wire n_181;
wire n_9743;
wire n_9121;
wire n_7371;
wire n_1362;
wire n_9509;
wire n_3123;
wire n_5447;
wire n_2692;
wire n_683;
wire n_7463;
wire n_9621;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_5755;
wire n_5700;
wire n_9158;
wire n_2862;
wire n_4325;
wire n_1420;
wire n_2645;
wire n_2553;
wire n_4711;
wire n_6889;
wire n_2749;
wire n_5962;
wire n_660;
wire n_464;
wire n_4413;
wire n_8627;
wire n_1210;
wire n_3307;
wire n_8945;
wire n_9142;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_9216;
wire n_9189;
wire n_6723;
wire n_7398;
wire n_1038;
wire n_3723;
wire n_7941;
wire n_4135;
wire n_9563;
wire n_6154;
wire n_5223;
wire n_5662;
wire n_8858;
wire n_414;
wire n_571;
wire n_3880;
wire n_5801;
wire n_3904;
wire n_6054;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_7011;
wire n_3405;
wire n_2313;
wire n_6393;
wire n_7074;
wire n_8916;
wire n_613;
wire n_1022;
wire n_5465;
wire n_171;
wire n_8745;
wire n_3532;
wire n_5154;
wire n_5721;
wire n_2609;
wire n_8169;
wire n_6184;
wire n_8018;
wire n_1767;
wire n_9984;
wire n_4138;
wire n_1040;
wire n_3131;
wire n_7083;
wire n_316;
wire n_125;
wire n_1973;
wire n_1444;
wire n_820;
wire n_8260;
wire n_254;
wire n_2882;
wire n_7143;
wire n_2303;
wire n_7701;
wire n_8688;
wire n_9794;
wire n_7969;
wire n_8279;
wire n_4384;
wire n_8793;
wire n_4639;
wire n_1664;
wire n_4577;
wire n_6312;
wire n_7683;
wire n_9550;
wire n_532;
wire n_2154;
wire n_7669;
wire n_1986;
wire n_8298;
wire n_6711;
wire n_2624;
wire n_6818;
wire n_6438;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_984;
wire n_5087;
wire n_1552;
wire n_2938;
wire n_7209;
wire n_2498;
wire n_6193;
wire n_3992;
wire n_8023;
wire n_9319;
wire n_7330;
wire n_6007;
wire n_621;
wire n_6734;
wire n_6535;
wire n_8053;
wire n_8059;
wire n_1772;
wire n_9871;
wire n_6879;
wire n_9562;
wire n_9896;
wire n_9612;
wire n_493;
wire n_1311;
wire n_3106;
wire n_6208;
wire n_7190;
wire n_9698;
wire n_2881;
wire n_6303;
wire n_3092;
wire n_6014;
wire n_4270;
wire n_7692;
wire n_697;
wire n_9528;
wire n_4620;
wire n_5397;
wire n_6457;
wire n_6255;
wire n_9272;
wire n_9955;
wire n_9645;
wire n_4924;
wire n_4044;
wire n_8372;
wire n_6270;
wire n_2305;
wire n_8737;
wire n_9731;
wire n_10026;
wire n_5996;
wire n_880;
wire n_5566;
wire n_9697;
wire n_3304;
wire n_7288;
wire n_4388;
wire n_7362;
wire n_7082;
wire n_7237;
wire n_8988;
wire n_3247;
wire n_7131;
wire n_6276;
wire n_739;
wire n_1028;
wire n_9642;
wire n_530;
wire n_8723;
wire n_9929;
wire n_9050;
wire n_4406;
wire n_2180;
wire n_4271;
wire n_7042;
wire n_9859;
wire n_8419;
wire n_2809;
wire n_5652;
wire n_8893;
wire n_975;
wire n_1645;
wire n_5805;
wire n_7304;
wire n_932;
wire n_6266;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_9531;
wire n_3785;
wire n_5492;
wire n_8077;
wire n_2465;
wire n_5501;
wire n_6934;
wire n_7386;
wire n_2972;
wire n_7391;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_7754;
wire n_8826;
wire n_3178;
wire n_268;
wire n_7023;
wire n_2251;
wire n_9732;
wire n_5842;
wire n_5758;
wire n_9685;
wire n_3100;
wire n_3721;
wire n_7404;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_8959;
wire n_6147;
wire n_5692;
wire n_6765;
wire n_4973;
wire n_7981;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_191;
wire n_2487;
wire n_5473;
wire n_1834;
wire n_8712;
wire n_1011;
wire n_2534;
wire n_6352;
wire n_2941;
wire n_4286;
wire n_9378;
wire n_3638;
wire n_6211;
wire n_8109;
wire n_3576;
wire n_10074;
wire n_9389;
wire n_5562;
wire n_4858;
wire n_1445;
wire n_6093;
wire n_5370;
wire n_10001;
wire n_7378;
wire n_9623;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_5458;
wire n_7877;
wire n_7787;
wire n_7836;
wire n_8515;
wire n_8725;
wire n_8007;
wire n_2387;
wire n_4318;
wire n_332;
wire n_8910;
wire n_5227;
wire n_830;
wire n_10100;
wire n_5902;
wire n_987;
wire n_2510;
wire n_9164;
wire n_6402;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_2793;
wire n_5282;
wire n_9387;
wire n_8301;
wire n_6764;
wire n_7871;
wire n_541;
wire n_499;
wire n_10162;
wire n_2639;
wire n_9840;
wire n_7016;
wire n_4738;
wire n_2603;
wire n_8892;
wire n_9637;
wire n_5386;
wire n_1167;
wire n_6215;
wire n_4554;
wire n_7571;
wire n_8252;
wire n_4526;
wire n_4105;
wire n_969;
wire n_3663;
wire n_9491;
wire n_1663;
wire n_6955;
wire n_7563;
wire n_5952;
wire n_7180;
wire n_2086;
wire n_1926;
wire n_8972;
wire n_8494;
wire n_6569;
wire n_1630;
wire n_7919;
wire n_9992;
wire n_663;
wire n_1720;
wire n_2966;
wire n_2409;
wire n_8278;
wire n_443;
wire n_3431;
wire n_8180;
wire n_3355;
wire n_7031;
wire n_1738;
wire n_5716;
wire n_8941;
wire n_8891;
wire n_406;
wire n_3897;
wire n_7103;
wire n_139;
wire n_6605;
wire n_1735;
wire n_391;
wire n_9266;
wire n_5888;
wire n_4005;
wire n_8270;
wire n_8231;
wire n_4181;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_6832;
wire n_5980;
wire n_8683;
wire n_956;
wire n_9391;
wire n_765;
wire n_4092;
wire n_4875;
wire n_7771;
wire n_8903;
wire n_4255;
wire n_2758;
wire n_385;
wire n_6544;
wire n_8810;
wire n_6469;
wire n_5036;
wire n_1271;
wire n_6332;
wire n_2186;
wire n_5790;
wire n_399;
wire n_7130;
wire n_10174;
wire n_6680;
wire n_4647;
wire n_3575;
wire n_6310;
wire n_8932;
wire n_8264;
wire n_2471;
wire n_9695;
wire n_7134;
wire n_3042;
wire n_8288;
wire n_1067;
wire n_1323;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_9834;
wire n_900;
wire n_5485;
wire n_9901;
wire n_5525;
wire n_7102;
wire n_10015;
wire n_10076;
wire n_6259;
wire n_3004;
wire n_1551;
wire n_5271;
wire n_4849;
wire n_2039;
wire n_7133;
wire n_9800;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_3838;
wire n_6651;
wire n_6289;
wire n_9255;
wire n_8882;
wire n_4059;
wire n_6565;
wire n_5194;
wire n_8388;
wire n_5445;
wire n_2734;
wire n_8067;
wire n_8385;
wire n_7227;
wire n_5948;
wire n_4499;
wire n_8670;
wire n_4504;
wire n_3598;
wire n_7813;
wire n_7706;
wire n_4917;
wire n_8142;
wire n_2420;
wire n_7992;
wire n_9085;
wire n_7643;
wire n_153;
wire n_648;
wire n_6836;
wire n_3273;
wire n_9120;
wire n_2918;
wire n_6595;
wire n_835;
wire n_9899;
wire n_9136;
wire n_6186;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_401;
wire n_7628;
wire n_1792;
wire n_5628;
wire n_504;
wire n_5245;
wire n_2062;
wire n_483;
wire n_9436;
wire n_4489;
wire n_822;
wire n_1459;
wire n_2153;
wire n_5329;
wire n_8224;
wire n_5472;
wire n_6035;
wire n_9042;
wire n_839;
wire n_1754;
wire n_7236;
wire n_9239;
wire n_9570;
wire n_3394;
wire n_4833;
wire n_6405;
wire n_8345;
wire n_9644;
wire n_2235;
wire n_5850;
wire n_1575;
wire n_9343;
wire n_8614;
wire n_8242;
wire n_6786;
wire n_4564;
wire n_8299;
wire n_1848;
wire n_9131;
wire n_1172;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_9060;
wire n_9792;
wire n_3581;
wire n_8110;
wire n_5072;
wire n_8529;
wire n_3778;
wire n_6769;
wire n_6844;
wire n_4322;
wire n_6361;
wire n_8951;
wire n_2260;
wire n_323;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_2206;
wire n_997;
wire n_635;
wire n_8700;
wire n_6766;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_5940;
wire n_3001;
wire n_5260;
wire n_6751;
wire n_4981;
wire n_6232;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_7519;
wire n_7802;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_7457;
wire n_5372;
wire n_6736;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_5860;
wire n_9982;
wire n_2422;
wire n_6416;
wire n_654;
wire n_2933;
wire n_8468;
wire n_9031;
wire n_7515;
wire n_3387;
wire n_7639;
wire n_8933;
wire n_6214;
wire n_3952;
wire n_8636;
wire n_9006;
wire n_9221;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_1059;
wire n_7049;
wire n_7884;
wire n_6945;
wire n_8378;
wire n_6143;
wire n_2736;
wire n_6491;
wire n_7749;
wire n_7592;
wire n_10091;
wire n_3825;
wire n_4198;
wire n_7172;
wire n_539;
wire n_8283;
wire n_977;
wire n_449;
wire n_2339;
wire n_392;
wire n_6225;
wire n_2532;
wire n_4373;
wire n_7914;
wire n_1866;
wire n_8860;
wire n_2664;
wire n_4154;
wire n_7344;
wire n_5859;
wire n_6447;
wire n_4390;
wire n_459;
wire n_1782;
wire n_7892;
wire n_1558;
wire n_4107;
wire n_2519;
wire n_9523;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_7325;
wire n_2360;
wire n_4453;
wire n_6219;
wire n_723;
wire n_1393;
wire n_7674;
wire n_8686;
wire n_6175;
wire n_6445;
wire n_9829;
wire n_8563;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_809;
wire n_10197;
wire n_3032;
wire n_5612;
wire n_4886;
wire n_8493;
wire n_6198;
wire n_5172;
wire n_881;
wire n_1019;
wire n_1477;
wire n_6499;
wire n_9411;
wire n_1982;
wire n_7983;
wire n_641;
wire n_5311;
wire n_8765;
wire n_910;
wire n_290;
wire n_5164;
wire n_4964;
wire n_10180;
wire n_9153;
wire n_4700;
wire n_6842;
wire n_4002;
wire n_217;
wire n_10079;
wire n_7361;
wire n_1114;
wire n_1742;
wire n_4679;
wire n_6397;
wire n_3815;
wire n_6827;
wire n_201;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_1273;
wire n_2982;
wire n_8653;
wire n_5495;
wire n_6281;
wire n_4483;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_5547;
wire n_4693;
wire n_8601;
wire n_1043;
wire n_9675;
wire n_6822;
wire n_5121;
wire n_4956;
wire n_255;
wire n_2869;
wire n_8333;
wire n_9097;
wire n_9571;
wire n_5379;
wire n_7079;
wire n_4487;
wire n_5878;
wire n_10075;
wire n_9789;
wire n_2674;
wire n_5820;
wire n_9925;
wire n_1737;
wire n_7309;
wire n_7119;
wire n_1613;
wire n_3026;
wire n_7184;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_7696;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_10012;
wire n_3902;
wire n_196;
wire n_3244;
wire n_1779;
wire n_2562;
wire n_954;
wire n_3112;
wire n_2051;
wire n_10008;
wire n_9511;
wire n_9795;
wire n_3196;
wire n_231;
wire n_8708;
wire n_5964;
wire n_2673;
wire n_6076;
wire n_10111;
wire n_4678;
wire n_664;
wire n_1591;
wire n_5301;
wire n_5126;
wire n_8659;
wire n_6732;
wire n_8759;
wire n_2548;
wire n_3488;
wire n_9622;
wire n_2381;
wire n_9761;
wire n_2744;
wire n_6817;
wire n_1967;
wire n_5776;
wire n_2179;
wire n_1280;
wire n_544;
wire n_7646;
wire n_9954;
wire n_3779;
wire n_599;
wire n_6982;
wire n_537;
wire n_1063;
wire n_7291;
wire n_8790;
wire n_991;
wire n_2275;
wire n_7668;
wire n_7435;
wire n_8832;
wire n_4606;
wire n_8305;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_5603;
wire n_938;
wire n_1891;
wire n_8453;
wire n_6560;
wire n_6634;
wire n_5348;
wire n_583;
wire n_9847;
wire n_1000;
wire n_313;
wire n_4868;
wire n_7017;
wire n_378;
wire n_4072;
wire n_7848;
wire n_2792;
wire n_4465;
wire n_9640;
wire n_8127;
wire n_2596;
wire n_5217;
wire n_8337;
wire n_9115;
wire n_3986;
wire n_5558;
wire n_3725;
wire n_7861;
wire n_10190;
wire n_9534;
wire n_472;
wire n_4026;
wire n_4245;
wire n_5520;
wire n_2524;
wire n_7889;
wire n_208;
wire n_3894;
wire n_1702;
wire n_5909;
wire n_4852;
wire n_275;
wire n_7554;
wire n_3202;
wire n_8508;
wire n_4290;
wire n_4945;
wire n_5750;
wire n_7648;
wire n_8968;
wire n_147;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1082;
wire n_1725;
wire n_5654;
wire n_2318;
wire n_866;
wire n_2819;
wire n_1722;
wire n_9594;
wire n_2229;
wire n_7653;
wire n_6400;
wire n_1644;
wire n_7846;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_8347;
wire n_131;
wire n_2255;
wire n_5554;
wire n_9503;
wire n_1252;
wire n_3045;
wire n_9919;
wire n_250;
wire n_773;
wire n_5135;
wire n_7551;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_6655;
wire n_10017;
wire n_718;
wire n_1434;
wire n_8093;
wire n_8899;
wire n_9385;
wire n_1905;
wire n_1569;
wire n_5448;
wire n_2573;
wire n_6480;
wire n_7737;
wire n_5837;
wire n_2336;
wire n_5412;
wire n_523;
wire n_1662;
wire n_8481;
wire n_3249;
wire n_3483;
wire n_6851;
wire n_6621;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_782;
wire n_2915;
wire n_7606;
wire n_9963;
wire n_7420;
wire n_9885;
wire n_8115;
wire n_4869;
wire n_3213;
wire n_5533;
wire n_4047;
wire n_1244;
wire n_1796;
wire n_484;
wire n_2719;
wire n_10115;
wire n_2876;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_6226;
wire n_9827;
wire n_1574;
wire n_3033;
wire n_893;
wire n_9182;
wire n_1582;
wire n_8182;
wire n_9426;
wire n_9293;
wire n_1981;
wire n_2824;
wire n_10065;
wire n_7973;
wire n_7545;
wire n_5327;
wire n_4417;
wire n_796;
wire n_127;
wire n_531;
wire n_1374;
wire n_2089;
wire n_7896;
wire n_6283;
wire n_4688;
wire n_7156;
wire n_4939;
wire n_9581;
wire n_8629;
wire n_5900;
wire n_8186;
wire n_7319;
wire n_1486;
wire n_3619;
wire n_6158;
wire n_9400;
wire n_4013;
wire n_3434;
wire n_9246;
wire n_4342;
wire n_691;
wire n_6819;
wire n_4903;
wire n_6122;
wire n_2131;
wire n_3853;
wire n_8233;
wire n_4382;
wire n_2509;
wire n_423;
wire n_4085;
wire n_6898;
wire n_6570;
wire n_5486;
wire n_2135;
wire n_9445;
wire n_8282;
wire n_7260;
wire n_6894;
wire n_4475;
wire n_6843;
wire n_5432;
wire n_7516;
wire n_5851;
wire n_6317;
wire n_6928;
wire n_6707;
wire n_10009;
wire n_7244;
wire n_187;
wire n_1463;
wire n_4626;
wire n_10072;
wire n_7625;
wire n_8750;
wire n_10130;
wire n_4997;
wire n_8183;
wire n_5065;
wire n_9104;
wire n_6806;
wire n_924;
wire n_7991;
wire n_781;
wire n_8637;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_9542;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_8792;
wire n_6835;
wire n_7286;
wire n_2436;
wire n_3517;
wire n_6269;
wire n_7857;
wire n_7970;
wire n_9302;
wire n_1706;
wire n_2461;
wire n_8258;
wire n_3719;
wire n_7154;
wire n_524;
wire n_634;
wire n_1214;
wire n_3526;
wire n_3888;
wire n_9960;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_5295;
wire n_8390;
wire n_8416;
wire n_6088;
wire n_1181;
wire n_1999;
wire n_7194;
wire n_4841;
wire n_4683;
wire n_5173;
wire n_2873;
wire n_10002;
wire n_8696;
wire n_9185;
wire n_9601;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_5655;
wire n_3383;
wire n_1835;
wire n_7175;
wire n_5855;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_7163;
wire n_3797;
wire n_1836;
wire n_7027;
wire n_3416;
wire n_8552;
wire n_4600;
wire n_5861;
wire n_1453;
wire n_6964;
wire n_3943;
wire n_3145;
wire n_7964;
wire n_5749;
wire n_6320;
wire n_9403;
wire n_6316;
wire n_8619;
wire n_419;
wire n_7068;
wire n_9972;
wire n_2908;
wire n_8594;
wire n_9878;
wire n_10139;
wire n_270;
wire n_4106;
wire n_9541;
wire n_285;
wire n_2156;
wire n_1184;
wire n_202;
wire n_8162;
wire n_9735;
wire n_754;
wire n_9576;
wire n_2323;
wire n_1073;
wire n_4549;
wire n_7327;
wire n_1277;
wire n_1746;
wire n_6610;
wire n_1062;
wire n_5998;
wire n_8318;
wire n_4702;
wire n_5102;
wire n_9974;
wire n_4954;
wire n_740;
wire n_167;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_8425;
wire n_6752;
wire n_6959;
wire n_9704;
wire n_6250;
wire n_3283;
wire n_259;
wire n_4331;
wire n_7317;
wire n_4159;
wire n_7864;
wire n_3451;
wire n_8051;
wire n_4734;
wire n_6675;
wire n_7955;
wire n_2832;
wire n_1688;
wire n_5827;
wire n_2370;
wire n_1944;
wire n_9039;
wire n_7384;
wire n_267;
wire n_2914;
wire n_5656;
wire n_7218;
wire n_1988;
wire n_5678;
wire n_6561;
wire n_6858;
wire n_5865;
wire n_6050;
wire n_7512;
wire n_1718;
wire n_7814;
wire n_8389;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_200;
wire n_10029;
wire n_2539;
wire n_8620;
wire n_10125;
wire n_5555;
wire n_2078;
wire n_8886;
wire n_1145;
wire n_7152;
wire n_4809;
wire n_787;
wire n_4012;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_5212;
wire n_4760;
wire n_1207;
wire n_6823;
wire n_3606;
wire n_7062;
wire n_7090;
wire n_8202;
wire n_2232;
wire n_1847;
wire n_5815;
wire n_4320;
wire n_5084;
wire n_7223;
wire n_5251;
wire n_1314;
wire n_8755;
wire n_1512;
wire n_8668;
wire n_5965;
wire n_884;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_6796;
wire n_8979;
wire n_5407;
wire n_2988;
wire n_4560;
wire n_7761;
wire n_8141;
wire n_3230;
wire n_5042;
wire n_859;
wire n_8199;
wire n_3793;
wire n_7055;
wire n_6024;
wire n_4768;
wire n_1889;
wire n_6090;
wire n_693;
wire n_5368;
wire n_929;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_9908;
wire n_8004;
wire n_8383;
wire n_3607;
wire n_1637;
wire n_9688;
wire n_9864;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_7388;
wire n_1751;
wire n_7056;
wire n_10212;
wire n_7437;
wire n_6489;
wire n_9023;
wire n_5310;
wire n_2769;
wire n_8895;
wire n_438;
wire n_8680;
wire n_1548;
wire n_4987;
wire n_6714;
wire n_8394;
wire n_440;
wire n_7849;
wire n_7726;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_7417;
wire n_2739;
wire n_3962;
wire n_7446;
wire n_4988;
wire n_6038;
wire n_2902;
wire n_6030;
wire n_6620;
wire n_4360;
wire n_1544;
wire n_6791;
wire n_6245;
wire n_4540;
wire n_9220;
wire n_6821;
wire n_9317;
wire n_2094;
wire n_8198;
wire n_3854;
wire n_5588;
wire n_9993;
wire n_1354;
wire n_8665;
wire n_6583;
wire n_2349;
wire n_3652;
wire n_7859;
wire n_3449;
wire n_1021;
wire n_3089;
wire n_4854;
wire n_9561;
wire n_491;
wire n_9444;
wire n_1595;
wire n_8017;
wire n_1142;
wire n_5477;
wire n_260;
wire n_2727;
wire n_942;
wire n_7523;
wire n_5234;
wire n_1416;
wire n_6890;
wire n_9184;
wire n_7559;
wire n_9037;
wire n_7576;
wire n_6988;
wire n_8303;
wire n_1599;
wire n_5871;
wire n_4747;
wire n_8000;
wire n_3472;
wire n_2527;
wire n_6052;
wire n_7769;
wire n_9505;
wire n_9193;
wire n_7257;
wire n_3126;
wire n_2759;
wire n_6973;
wire n_8852;
wire n_5007;
wire n_8709;
wire n_4881;
wire n_2038;
wire n_6488;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_9218;
wire n_9755;
wire n_4357;
wire n_7729;
wire n_2806;
wire n_4502;
wire n_287;
wire n_3191;
wire n_1716;
wire n_302;
wire n_7005;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_8782;
wire n_7081;
wire n_7742;
wire n_5253;
wire n_3588;
wire n_355;
wire n_6280;
wire n_1590;
wire n_3280;
wire n_4115;
wire n_5274;
wire n_6399;
wire n_5418;
wire n_5019;
wire n_5939;
wire n_1819;
wire n_9162;
wire n_9506;
wire n_135;
wire n_3095;
wire n_947;
wire n_7341;
wire n_5792;
wire n_3698;
wire n_4513;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_4775;
wire n_6256;
wire n_482;
wire n_2620;
wire n_1833;
wire n_8716;
wire n_1691;
wire n_8250;
wire n_7264;
wire n_7842;
wire n_2549;
wire n_2499;
wire n_6648;
wire n_9415;
wire n_7492;
wire n_804;
wire n_6649;
wire n_8714;
wire n_1656;
wire n_8357;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_6910;
wire n_9990;
wire n_3885;
wire n_955;
wire n_8466;
wire n_4264;
wire n_9015;
wire n_5954;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_514;
wire n_6431;
wire n_418;
wire n_8589;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_8266;
wire n_3839;
wire n_8587;
wire n_7285;
wire n_5490;
wire n_5694;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_6324;
wire n_5489;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_8876;
wire n_9214;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_8922;
wire n_10090;
wire n_3120;
wire n_6512;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_9070;
wire n_8498;
wire n_4794;
wire n_9933;
wire n_4843;
wire n_669;
wire n_5580;
wire n_5215;
wire n_337;
wire n_437;
wire n_3937;
wire n_4763;
wire n_9339;
wire n_1418;
wire n_9991;
wire n_9486;
wire n_8457;
wire n_6243;
wire n_5795;
wire n_5715;
wire n_4170;
wire n_5561;
wire n_8267;
wire n_2462;
wire n_7051;
wire n_6773;
wire n_2155;
wire n_6231;
wire n_615;
wire n_7503;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_517;
wire n_8124;
wire n_3604;
wire n_8545;
wire n_5430;
wire n_6041;
wire n_8526;
wire n_824;
wire n_159;
wire n_8319;
wire n_7997;
wire n_5659;
wire n_9279;
wire n_6859;
wire n_7716;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_9790;
wire n_144;
wire n_3792;
wire n_7950;
wire n_6323;
wire n_5720;
wire n_4267;
wire n_8581;
wire n_8214;
wire n_7793;
wire n_9053;
wire n_8516;
wire n_2083;
wire n_815;
wire n_5598;
wire n_2753;
wire n_1340;
wire n_470;
wire n_3021;
wire n_8989;
wire n_7746;
wire n_477;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_7570;
wire n_9650;
wire n_9880;
wire n_2898;
wire n_1825;
wire n_6912;
wire n_3567;
wire n_7425;
wire n_2682;
wire n_5854;
wire n_5958;
wire n_5585;
wire n_5112;
wire n_5326;
wire n_1627;
wire n_9217;
wire n_9499;
wire n_5783;
wire n_7829;
wire n_6837;
wire n_6747;
wire n_2903;
wire n_5303;
wire n_10081;
wire n_3812;
wire n_3127;
wire n_6916;
wire n_1731;
wire n_799;
wire n_7894;
wire n_9282;
wire n_1147;
wire n_10145;
wire n_7957;
wire n_8262;
wire n_2378;
wire n_10167;
wire n_5530;
wire n_6718;
wire n_8289;
wire n_965;
wire n_5809;
wire n_934;
wire n_2213;
wire n_7121;
wire n_7531;
wire n_6410;
wire n_356;
wire n_6473;
wire n_8087;
wire n_4056;
wire n_4806;
wire n_7961;
wire n_1674;
wire n_9920;
wire n_5993;
wire n_4015;
wire n_6574;
wire n_2924;
wire n_6492;
wire n_4445;
wire n_7687;
wire n_9948;
wire n_4462;
wire n_5299;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_8863;
wire n_9371;
wire n_4517;
wire n_2896;
wire n_8701;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_1042;
wire n_3170;
wire n_9237;
wire n_2311;
wire n_6857;
wire n_8705;
wire n_1455;
wire n_2287;
wire n_9815;
wire n_836;
wire n_3415;
wire n_6975;
wire n_7763;
wire n_3464;
wire n_6290;
wire n_3414;
wire n_6646;
wire n_205;
wire n_7703;
wire n_7928;
wire n_4234;
wire n_760;
wire n_1483;
wire n_10168;
wire n_1363;
wire n_8722;
wire n_1111;
wire n_970;
wire n_3467;
wire n_5821;
wire n_713;
wire n_3179;
wire n_598;
wire n_6622;
wire n_5522;
wire n_7665;
wire n_3889;
wire n_7677;
wire n_4836;
wire n_5262;
wire n_3262;
wire n_5319;
wire n_927;
wire n_7469;
wire n_261;
wire n_3699;
wire n_10163;
wire n_6118;
wire n_706;
wire n_2120;
wire n_7125;
wire n_7856;
wire n_6028;
wire n_6663;
wire n_6532;
wire n_1419;
wire n_8622;
wire n_3816;
wire n_8099;
wire n_8729;
wire n_9479;
wire n_3528;
wire n_6267;
wire n_6682;
wire n_9480;
wire n_4207;
wire n_8085;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_4725;
wire n_9597;
wire n_348;
wire n_9173;
wire n_2312;
wire n_7203;
wire n_8947;
wire n_9641;
wire n_7797;
wire n_1826;
wire n_9983;
wire n_9267;
wire n_5943;
wire n_6556;
wire n_10039;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_6216;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_637;
wire n_7128;
wire n_9849;
wire n_5335;
wire n_1259;
wire n_6365;
wire n_8459;
wire n_7111;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_8478;
wire n_5284;
wire n_8786;
wire n_9414;
wire n_4978;
wire n_5771;
wire n_3246;
wire n_9419;
wire n_3299;
wire n_8887;
wire n_980;
wire n_1618;
wire n_1869;
wire n_3623;
wire n_905;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_8851;
wire n_6950;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_8540;
wire n_5516;
wire n_7284;
wire n_3615;
wire n_8276;
wire n_7057;
wire n_1802;
wire n_9823;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_9152;
wire n_8706;
wire n_3200;
wire n_6167;
wire n_3642;
wire n_145;
wire n_2146;
wire n_4274;
wire n_5583;
wire n_3276;
wire n_7064;
wire n_8532;
wire n_9533;
wire n_5433;
wire n_3682;
wire n_5429;
wire n_7278;
wire n_9281;
wire n_9103;
wire n_9111;
wire n_6772;
wire n_7088;
wire n_7799;
wire n_9618;
wire n_5698;
wire n_5731;
wire n_8871;
wire n_4007;
wire n_1456;
wire n_8433;
wire n_9065;
wire n_1879;
wire n_6159;
wire n_2129;
wire n_7048;
wire n_5857;
wire n_7979;
wire n_9674;
wire n_6617;
wire n_553;
wire n_7725;
wire n_814;
wire n_578;
wire n_5120;
wire n_3572;
wire n_8371;
wire n_2975;
wire n_2399;
wire n_8547;
wire n_1134;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_8467;
wire n_647;
wire n_2027;
wire n_2932;
wire n_8409;
wire n_6217;
wire n_600;
wire n_3118;
wire n_9157;
wire n_5560;
wire n_9170;
wire n_4441;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_5455;
wire n_502;
wire n_6777;
wire n_8640;
wire n_10196;
wire n_6742;
wire n_1467;
wire n_7447;
wire n_5209;
wire n_247;
wire n_6307;
wire n_5704;
wire n_4889;
wire n_2159;
wire n_8431;
wire n_4458;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_8415;
wire n_5916;
wire n_10184;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_6479;
wire n_5099;
wire n_681;
wire n_3286;
wire n_5781;
wire n_5619;
wire n_2023;
wire n_9416;
wire n_3974;
wire n_9368;
wire n_7365;
wire n_3443;
wire n_8329;
wire n_2599;
wire n_3988;
wire n_7792;
wire n_8089;
wire n_5022;
wire n_9208;
wire n_6370;
wire n_9223;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3996;
wire n_3761;
wire n_7275;
wire n_5353;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_6856;
wire n_1098;
wire n_9781;
wire n_3009;
wire n_8633;
wire n_777;
wire n_7095;
wire n_7390;
wire n_9392;
wire n_6140;
wire n_6111;
wire n_5219;
wire n_9422;
wire n_920;
wire n_8541;
wire n_10084;
wire n_8762;
wire n_3951;
wire n_5518;
wire n_9970;
wire n_3035;
wire n_4261;
wire n_7037;
wire n_1132;
wire n_9338;
wire n_8125;
wire n_501;
wire n_1823;
wire n_6240;
wire n_5236;
wire n_4236;
wire n_10077;
wire n_3942;
wire n_3023;
wire n_9492;
wire n_2254;
wire n_3290;
wire n_6693;
wire n_9226;
wire n_6712;
wire n_7530;
wire n_10129;
wire n_10101;
wire n_1402;
wire n_3957;
wire n_3418;
wire n_1607;
wire n_7471;
wire n_9328;
wire n_6465;
wire n_221;
wire n_8188;
wire n_10192;
wire n_5673;
wire n_861;
wire n_8615;
wire n_5814;
wire n_1666;
wire n_6586;
wire n_7058;
wire n_5103;
wire n_4648;
wire n_8011;
wire n_10207;
wire n_2214;
wire n_6730;
wire n_6367;
wire n_2256;
wire n_8923;
wire n_281;
wire n_3326;
wire n_8624;
wire n_262;
wire n_8222;
wire n_6069;
wire n_2732;
wire n_1883;
wire n_6515;
wire n_8206;
wire n_4094;
wire n_2776;
wire n_6077;
wire n_9513;
wire n_3224;
wire n_9393;
wire n_1969;
wire n_5671;
wire n_7429;
wire n_6940;
wire n_8065;
wire n_9914;
wire n_527;
wire n_2949;
wire n_7008;
wire n_7709;
wire n_6468;
wire n_4269;
wire n_1927;
wire n_7540;
wire n_7581;
wire n_343;
wire n_1222;
wire n_7139;
wire n_8935;
wire n_3803;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_7782;
wire n_7432;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_8155;
wire n_9334;
wire n_2449;
wire n_10093;
wire n_4428;
wire n_745;
wire n_6483;
wire n_1572;
wire n_7770;
wire n_9684;
wire n_8397;
wire n_8568;
wire n_4463;
wire n_8175;
wire n_5357;
wire n_7173;
wire n_3648;
wire n_9254;
wire n_6576;
wire n_6810;
wire n_10003;
wire n_1975;
wire n_5421;
wire n_9083;
wire n_1388;
wire n_1266;
wire n_4396;
wire n_1990;
wire n_6708;
wire n_8026;
wire n_6667;
wire n_9175;
wire n_9838;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1075;
wire n_6040;
wire n_1890;
wire n_6847;
wire n_8974;
wire n_6305;
wire n_8836;
wire n_4034;
wire n_4228;
wire n_1227;
wire n_7251;
wire n_3166;
wire n_7356;
wire n_3649;
wire n_7412;
wire n_3065;
wire n_8168;
wire n_7212;
wire n_5045;
wire n_5237;
wire n_7751;
wire n_7951;
wire n_657;
wire n_7060;
wire n_3924;
wire n_9336;
wire n_3997;
wire n_8873;
wire n_7591;
wire n_3564;
wire n_862;
wire n_6750;
wire n_2637;
wire n_7444;
wire n_5769;
wire n_7911;
wire n_3795;
wire n_7595;
wire n_4931;
wire n_2306;
wire n_7790;
wire n_2071;
wire n_7426;
wire n_430;
wire n_3953;
wire n_4400;
wire n_7502;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_5434;
wire n_1532;
wire n_6855;
wire n_8170;
wire n_1030;
wire n_5181;
wire n_6239;
wire n_10181;
wire n_3208;
wire n_9554;
wire n_5768;
wire n_1342;
wire n_6199;
wire n_2737;
wire n_3282;
wire n_8120;
wire n_9116;
wire n_9315;
wire n_9830;
wire n_8825;
wire n_852;
wire n_9169;
wire n_2916;
wire n_7252;
wire n_1060;
wire n_5963;
wire n_9999;
wire n_4424;
wire n_4351;
wire n_6543;
wire n_7532;
wire n_4192;
wire n_8003;
wire n_9215;
wire n_1748;
wire n_1301;
wire n_6789;
wire n_8395;
wire n_3400;
wire n_5972;
wire n_7065;
wire n_1466;
wire n_8083;
wire n_6177;
wire n_8057;
wire n_2581;
wire n_5937;
wire n_1783;
wire n_9259;
wire n_5146;
wire n_7367;
wire n_8164;
wire n_7405;
wire n_7267;
wire n_4646;
wire n_4221;
wire n_1037;
wire n_3650;
wire n_8877;
wire n_1329;
wire n_6825;
wire n_7614;
wire n_1993;
wire n_1545;
wire n_6460;
wire n_134;
wire n_4035;
wire n_9150;
wire n_6952;
wire n_9595;
wire n_1480;
wire n_3670;
wire n_8366;
wire n_6173;
wire n_2540;
wire n_4190;
wire n_8476;
wire n_1605;
wire n_3060;
wire n_6218;
wire n_7685;
wire n_6486;
wire n_2984;
wire n_4009;
wire n_157;
wire n_7619;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_6852;
wire n_624;
wire n_5577;
wire n_876;
wire n_9100;
wire n_7883;
wire n_5872;
wire n_6692;
wire n_9707;
wire n_5017;
wire n_8854;
wire n_736;
wire n_10202;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_7220;
wire n_7560;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_9262;
wire n_5976;
wire n_4717;
wire n_9249;
wire n_6888;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_602;
wire n_854;
wire n_8256;
wire n_2091;
wire n_393;
wire n_4312;
wire n_5424;
wire n_3789;
wire n_7270;
wire n_1658;
wire n_1072;
wire n_8621;
wire n_1305;
wire n_4750;
wire n_2348;
wire n_9806;
wire n_1873;
wire n_8577;
wire n_9019;
wire n_10097;
wire n_2725;
wire n_2667;
wire n_9361;
wire n_3746;
wire n_7731;
wire n_6626;
wire n_4537;
wire n_1046;
wire n_5838;
wire n_7034;
wire n_8654;
wire n_3694;
wire n_6854;
wire n_7940;
wire n_771;
wire n_6793;
wire n_5456;
wire n_3893;
wire n_4847;
wire n_5846;
wire n_9814;
wire n_2307;
wire n_421;
wire n_3702;
wire n_5930;
wire n_8952;
wire n_1984;
wire n_3453;
wire n_9438;
wire n_1556;
wire n_7537;
wire n_6980;
wire n_7040;
wire n_5345;
wire n_2815;
wire n_7458;
wire n_4427;
wire n_1824;
wire n_7740;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_6794;
wire n_819;
wire n_1971;
wire n_2945;
wire n_586;
wire n_1324;
wire n_3543;
wire n_8421;
wire n_9856;
wire n_7179;
wire n_1776;
wire n_3448;
wire n_7433;
wire n_4279;
wire n_9327;
wire n_9313;
wire n_605;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_6334;
wire n_6257;
wire n_10142;
wire n_4152;
wire n_6874;
wire n_8911;
wire n_5537;
wire n_9518;
wire n_2698;
wire n_5572;
wire n_4783;
wire n_7658;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_5409;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_807;
wire n_5142;
wire n_10177;
wire n_8971;
wire n_7015;
wire n_6355;
wire n_6039;
wire n_6286;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_7226;
wire n_7987;
wire n_9291;
wire n_1987;
wire n_7217;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_9009;
wire n_2368;
wire n_9882;
wire n_6377;
wire n_802;
wire n_5401;
wire n_4595;
wire n_960;
wire n_7272;
wire n_8215;
wire n_2352;
wire n_5201;
wire n_5816;
wire n_790;
wire n_5551;
wire n_9722;
wire n_5416;
wire n_4404;
wire n_2377;
wire n_151;
wire n_7906;
wire n_2652;
wire n_5498;
wire n_5543;
wire n_4054;
wire n_9760;
wire n_6018;
wire n_7765;
wire n_1286;
wire n_6021;
wire n_4617;
wire n_1685;
wire n_2477;
wire n_4611;
wire n_10037;
wire n_8949;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_5797;
wire n_9454;
wire n_6511;
wire n_7815;
wire n_1052;
wire n_4732;
wire n_2076;
wire n_2203;
wire n_5942;
wire n_5764;
wire n_1426;
wire n_8983;
wire n_4969;
wire n_8121;
wire n_5252;
wire n_5777;
wire n_8942;
wire n_7785;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_6867;
wire n_4140;
wire n_5171;
wire n_566;
wire n_7728;
wire n_8280;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_7255;
wire n_3309;
wire n_169;
wire n_7181;
wire n_173;
wire n_2796;
wire n_858;
wire n_5393;
wire n_8328;
wire n_4817;
wire n_8861;
wire n_6863;
wire n_7352;
wire n_7355;
wire n_8427;
wire n_2136;
wire n_433;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_7328;
wire n_2771;
wire n_7359;
wire n_6322;
wire n_2403;
wire n_2947;
wire n_5643;
wire n_9826;
wire n_253;
wire n_928;
wire n_9937;
wire n_3769;
wire n_7825;
wire n_1565;
wire n_4437;
wire n_6419;
wire n_128;
wire n_7916;
wire n_3055;
wire n_8194;
wire n_420;
wire n_4070;
wire n_7283;
wire n_5346;
wire n_9453;
wire n_748;
wire n_7903;
wire n_9900;
wire n_7089;
wire n_1045;
wire n_8217;
wire n_9331;
wire n_1881;
wire n_2635;
wire n_7604;
wire n_7647;
wire n_2999;
wire n_988;
wire n_4139;
wire n_4769;
wire n_6130;
wire n_330;
wire n_5868;
wire n_6417;
wire n_328;
wire n_368;
wire n_8285;
wire n_7145;
wire n_8521;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_9178;
wire n_7803;
wire n_9689;
wire n_2713;
wire n_1422;
wire n_8448;
wire n_1965;
wire n_644;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_6979;
wire n_5986;
wire n_9355;
wire n_9489;
wire n_6932;
wire n_2934;
wire n_7258;
wire n_5104;
wire n_6961;
wire n_576;
wire n_8732;
wire n_511;
wire n_7622;
wire n_9359;
wire n_429;
wire n_7839;
wire n_6792;
wire n_7720;
wire n_2210;
wire n_4368;
wire n_5794;
wire n_8136;
wire n_3141;
wire n_2053;
wire n_5272;
wire n_3476;
wire n_6919;
wire n_1049;
wire n_8420;
wire n_141;
wire n_4430;
wire n_8386;
wire n_6123;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_7440;
wire n_1356;
wire n_9568;
wire n_6831;
wire n_1773;
wire n_3175;
wire n_4544;
wire n_2666;
wire n_5578;
wire n_312;
wire n_728;
wire n_4409;
wire n_4191;
wire n_2401;
wire n_7809;
wire n_3255;
wire n_2588;
wire n_5722;
wire n_5811;
wire n_935;
wire n_7072;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_911;
wire n_623;
wire n_3509;
wire n_8746;
wire n_10051;
wire n_1403;
wire n_5395;
wire n_453;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_6458;
wire n_9401;
wire n_8857;
wire n_543;
wire n_6986;
wire n_9495;
wire n_3456;
wire n_4532;
wire n_236;
wire n_601;
wire n_7564;
wire n_628;
wire n_5863;
wire n_8185;
wire n_8313;
wire n_6633;
wire n_3790;
wire n_7775;
wire n_907;
wire n_7118;
wire n_9234;
wire n_7960;
wire n_6152;
wire n_9431;
wire n_5734;
wire n_10023;
wire n_8281;
wire n_847;
wire n_747;
wire n_1135;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_6169;
wire n_5774;
wire n_7069;
wire n_5199;
wire n_6546;
wire n_4257;
wire n_4282;
wire n_7636;
wire n_4341;
wire n_10199;
wire n_1694;
wire n_6925;
wire n_7186;
wire n_593;
wire n_8766;
wire n_1695;
wire n_4027;
wire n_4650;
wire n_4309;
wire n_5480;
wire n_6428;
wire n_609;
wire n_6924;
wire n_3077;
wire n_4944;
wire n_8066;
wire n_9340;
wire n_9380;
wire n_7666;
wire n_6425;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_9976;
wire n_4994;
wire n_7967;
wire n_5977;
wire n_519;
wire n_8314;
wire n_384;
wire n_3533;
wire n_5175;
wire n_7246;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_9064;
wire n_3409;
wire n_4381;
wire n_8239;
wire n_9092;
wire n_3583;
wire n_4316;
wire n_7301;
wire n_4860;
wire n_4469;
wire n_9746;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_8497;
wire n_1157;
wire n_7262;
wire n_234;
wire n_5959;
wire n_8056;
wire n_8210;
wire n_3563;
wire n_5945;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_3689;
wire n_7584;
wire n_7748;
wire n_1789;
wire n_9066;
wire n_763;
wire n_6301;
wire n_2174;
wire n_540;
wire n_5668;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_1687;
wire n_7686;
wire n_6282;
wire n_4934;
wire n_4703;
wire n_9870;
wire n_9817;
wire n_2638;
wire n_2046;
wire n_7059;
wire n_6985;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_5600;
wire n_395;
wire n_6737;
wire n_1587;
wire n_213;
wire n_2340;
wire n_9857;
wire n_4804;
wire n_8404;
wire n_2444;
wire n_4888;
wire n_1014;
wire n_5767;
wire n_9455;
wire n_10056;
wire n_6459;
wire n_1427;
wire n_7670;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_8505;
wire n_2199;
wire n_6384;
wire n_4669;
wire n_5228;
wire n_1100;
wire n_585;
wire n_9916;
wire n_1617;
wire n_10157;
wire n_2600;
wire n_8606;
wire n_7443;
wire n_3436;
wire n_5973;
wire n_7484;
wire n_1962;
wire n_3806;
wire n_9440;
wire n_4759;
wire n_10038;
wire n_9059;
wire n_9812;
wire n_5869;
wire n_6753;
wire n_2114;
wire n_5914;
wire n_9690;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_9912;
wire n_1175;
wire n_4887;
wire n_3751;
wire n_9002;
wire n_3402;
wire n_9620;
wire n_1621;
wire n_6448;
wire n_9229;
wire n_5186;
wire n_7930;
wire n_7487;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_580;
wire n_3664;
wire n_4218;
wire n_9464;
wire n_434;
wire n_4687;
wire n_7077;
wire n_394;
wire n_1381;
wire n_3686;
wire n_1183;
wire n_8518;
wire n_4720;
wire n_2889;
wire n_6043;
wire n_6268;
wire n_9497;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_5604;
wire n_3470;
wire n_243;
wire n_7663;
wire n_8350;
wire n_8741;
wire n_7024;
wire n_8148;
wire n_1407;
wire n_5221;
wire n_8408;
wire n_6145;
wire n_2865;
wire n_5925;
wire n_6529;
wire n_973;
wire n_5591;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_8236;
wire n_7214;
wire n_8806;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_8295;
wire n_1176;
wire n_9587;
wire n_3677;
wire n_1054;
wire n_7977;
wire n_5387;
wire n_3292;
wire n_6311;
wire n_8167;
wire n_8377;
wire n_3989;
wire n_7652;
wire n_9783;
wire n_4644;
wire n_8956;
wire n_4752;
wire n_8673;
wire n_4746;
wire n_7566;
wire n_1057;
wire n_4131;
wire n_5449;
wire n_8760;
wire n_4215;
wire n_978;
wire n_2488;
wire n_1509;
wire n_828;
wire n_6134;
wire n_322;
wire n_4158;
wire n_6812;
wire n_3079;
wire n_10044;
wire n_5190;
wire n_6733;
wire n_3269;
wire n_558;
wire n_5325;
wire n_4231;
wire n_8960;
wire n_8957;
wire n_9008;
wire n_10143;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_653;
wire n_6262;
wire n_4926;
wire n_2050;
wire n_8207;
wire n_6938;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_5876;
wire n_5344;
wire n_2550;
wire n_556;
wire n_170;
wire n_1536;
wire n_3177;
wire n_6160;
wire n_10186;
wire n_4667;
wire n_5813;
wire n_10113;
wire n_6235;
wire n_1471;
wire n_6212;
wire n_3440;
wire n_9381;
wire n_9194;
wire n_6816;
wire n_8904;
wire n_3658;
wire n_7374;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1620;
wire n_2542;
wire n_10120;
wire n_5892;
wire n_9549;
wire n_7678;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_788;
wire n_7110;
wire n_5714;
wire n_2169;
wire n_6953;
wire n_9652;
wire n_7975;
wire n_9957;
wire n_8451;
wire n_6089;
wire n_591;
wire n_5634;
wire n_5133;
wire n_7553;
wire n_8527;
wire n_5990;
wire n_7086;
wire n_2175;
wire n_1625;
wire n_7732;
wire n_5689;
wire n_5305;
wire n_7891;
wire n_9089;
wire n_4578;
wire n_318;
wire n_8840;
wire n_5644;
wire n_9137;
wire n_9390;
wire n_3644;
wire n_8038;
wire n_8190;
wire n_9439;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_6138;
wire n_528;
wire n_9080;
wire n_1922;
wire n_9296;
wire n_940;
wire n_1537;
wire n_4877;
wire n_9312;
wire n_2065;
wire n_9151;
wire n_8179;
wire n_7038;
wire n_7994;
wire n_4470;
wire n_4187;
wire n_9883;
wire n_8287;
wire n_1904;
wire n_8111;
wire n_8341;
wire n_8830;
wire n_4998;
wire n_10200;
wire n_5576;
wire n_2395;
wire n_2868;
wire n_7345;
wire n_9324;
wire n_9631;
wire n_8308;
wire n_1530;
wire n_4057;
wire n_6070;
wire n_5852;
wire n_5918;
wire n_631;
wire n_8021;
wire n_1170;
wire n_2724;
wire n_8965;
wire n_9736;
wire n_2258;
wire n_7041;
wire n_9365;
wire n_6717;
wire n_7593;
wire n_8265;
wire n_898;
wire n_6881;
wire n_10085;
wire n_3328;
wire n_2012;
wire n_9600;
wire n_3182;
wire n_6871;
wire n_2967;
wire n_9816;
wire n_6672;
wire n_5343;
wire n_9869;
wire n_7757;
wire n_1093;
wire n_8251;
wire n_9402;
wire n_7866;
wire n_7334;
wire n_6518;
wire n_4021;
wire n_7028;
wire n_6396;
wire n_3379;
wire n_4379;
wire n_8773;
wire n_6242;
wire n_5947;
wire n_336;
wire n_6601;
wire n_8570;
wire n_2268;
wire n_3469;
wire n_10041;
wire n_1452;
wire n_2835;
wire n_5835;
wire n_10096;
wire n_668;
wire n_8579;
wire n_2111;
wire n_3743;
wire n_8079;
wire n_5542;
wire n_9615;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_5527;
wire n_2897;
wire n_9711;
wire n_9759;
wire n_4812;
wire n_8506;
wire n_8973;
wire n_4497;
wire n_6606;
wire n_2583;
wire n_8291;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_9820;
wire n_1770;
wire n_701;
wire n_1003;
wire n_7758;
wire n_8320;
wire n_8635;
wire n_9703;
wire n_4472;
wire n_9819;
wire n_9118;
wire n_2699;
wire n_9321;
wire n_5819;
wire n_3901;
wire n_291;
wire n_5180;
wire n_1640;
wire n_8375;
wire n_2973;
wire n_9428;
wire n_8612;
wire n_10198;
wire n_8778;
wire n_5893;
wire n_9292;
wire n_2710;
wire n_7705;
wire n_6092;
wire n_6462;
wire n_2505;
wire n_4519;
wire n_9018;
wire n_5025;
wire n_2397;
wire n_8872;
wire n_240;
wire n_369;
wire n_7333;
wire n_3878;
wire n_4197;
wire n_6669;
wire n_8006;
wire n_9565;
wire n_2721;
wire n_1892;
wire n_6251;
wire n_2615;
wire n_4787;
wire n_8491;
wire n_8218;
wire n_1212;
wire n_7337;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_7439;
wire n_5726;
wire n_4371;
wire n_188;
wire n_1902;
wire n_7744;
wire n_2784;
wire n_7210;
wire n_5828;
wire n_3898;
wire n_694;
wire n_6228;
wire n_6702;
wire n_7358;
wire n_8240;
wire n_10059;
wire n_9961;
wire n_4749;
wire n_7707;
wire n_5924;
wire n_1845;
wire n_7733;
wire n_921;
wire n_5545;
wire n_8458;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_8853;
wire n_9603;
wire n_5083;
wire n_7684;
wire n_3253;
wire n_8306;
wire n_2088;
wire n_1275;
wire n_6997;
wire n_9692;
wire n_4238;
wire n_6371;
wire n_904;
wire n_7673;
wire n_2005;
wire n_1696;
wire n_7187;
wire n_8013;
wire n_2108;
wire n_3824;
wire n_8342;
wire n_2246;
wire n_7313;
wire n_5899;
wire n_9012;
wire n_3846;
wire n_5122;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_6641;
wire n_3845;
wire n_6463;
wire n_10172;
wire n_3203;
wire n_383;
wire n_4986;
wire n_1316;
wire n_4668;
wire n_950;
wire n_9868;
wire n_711;
wire n_6264;
wire n_5782;
wire n_8119;
wire n_9264;
wire n_630;
wire n_4168;
wire n_1369;
wire n_8582;
wire n_7036;
wire n_4298;
wire n_7370;
wire n_7931;
wire n_4743;
wire n_8445;
wire n_1781;
wire n_9720;
wire n_4250;
wire n_3143;
wire n_8044;
wire n_3690;
wire n_3229;
wire n_5864;
wire n_8363;
wire n_8464;
wire n_8921;
wire n_235;
wire n_2188;
wire n_10010;
wire n_2430;
wire n_2504;
wire n_5637;
wire n_4211;
wire n_6084;
wire n_3094;
wire n_741;
wire n_9646;
wire n_7480;
wire n_8843;
wire n_371;
wire n_5185;
wire n_8405;
wire n_2964;
wire n_8376;
wire n_308;
wire n_5032;
wire n_6990;
wire n_865;
wire n_5034;
wire n_3312;
wire n_7071;
wire n_1041;
wire n_2451;
wire n_8694;
wire n_2913;
wire n_8848;
wire n_6288;
wire n_993;
wire n_1862;
wire n_3752;
wire n_8752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_8625;
wire n_8894;
wire n_7380;
wire n_2839;
wire n_8813;
wire n_3237;
wire n_7708;
wire n_9842;
wire n_4128;
wire n_4036;
wire n_9671;
wire n_5269;
wire n_8430;
wire n_3655;
wire n_2955;
wire n_5709;
wire n_1764;
wire n_4807;
wire n_8770;
wire n_6277;
wire n_8426;
wire n_5115;
wire n_7376;
wire n_8411;
wire n_902;
wire n_8817;
wire n_8461;
wire n_1723;
wire n_3918;
wire n_9230;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_596;
wire n_9893;
wire n_6409;
wire n_4095;
wire n_8391;
wire n_8507;
wire n_1310;
wire n_5927;
wire n_8691;
wire n_9188;
wire n_4485;
wire n_9032;
wire n_7657;
wire n_6388;
wire n_574;
wire n_3593;
wire n_6839;
wire n_5163;
wire n_9614;
wire n_8967;
wire n_1229;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_9628;
wire n_1896;
wire n_9231;
wire n_6864;
wire n_1516;
wire n_4890;
wire n_10204;
wire n_8084;
wire n_8856;
wire n_2485;
wire n_6679;
wire n_10201;
wire n_8631;
wire n_6051;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_8219;
wire n_9730;
wire n_5507;
wire n_195;
wire n_4573;
wire n_1328;
wire n_4943;
wire n_2875;
wire n_6599;
wire n_3519;
wire n_2209;
wire n_7504;
wire n_4042;
wire n_7099;
wire n_7586;
wire n_4244;
wire n_1928;
wire n_5642;
wire n_4708;
wire n_4883;
wire n_6227;
wire n_4553;
wire n_7052;
wire n_8428;
wire n_9172;
wire n_1634;
wire n_1203;
wire n_9926;
wire n_1699;
wire n_6738;
wire n_5226;
wire n_2081;
wire n_937;
wire n_1474;
wire n_8338;
wire n_1631;
wire n_7602;
wire n_9180;
wire n_9017;
wire n_156;
wire n_9269;
wire n_6566;
wire n_9026;
wire n_1794;
wire n_9462;
wire n_5696;
wire n_7998;
wire n_8666;
wire n_1375;
wire n_3053;
wire n_5014;
wire n_7106;
wire n_6346;
wire n_204;
wire n_7557;
wire n_3772;
wire n_7408;
wire n_2891;
wire n_496;
wire n_4335;
wire n_7026;
wire n_3128;
wire n_10052;
wire n_6146;
wire n_5677;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_1002;
wire n_7394;
wire n_9515;
wire n_9502;
wire n_263;
wire n_4516;
wire n_5235;
wire n_360;
wire n_1129;
wire n_7627;
wire n_6436;
wire n_1464;
wire n_7719;
wire n_2798;
wire n_7450;
wire n_165;
wire n_9316;
wire n_3217;
wire n_8938;
wire n_6081;
wire n_1249;
wire n_329;
wire n_7852;
wire n_5724;
wire n_3821;
wire n_340;
wire n_3201;
wire n_7462;
wire n_7780;
wire n_3503;
wire n_8523;
wire n_5979;
wire n_6027;
wire n_1870;
wire n_10121;
wire n_4467;
wire n_177;
wire n_364;
wire n_258;
wire n_7582;
wire n_5521;
wire n_431;
wire n_2654;
wire n_3935;
wire n_7421;
wire n_1861;
wire n_9873;
wire n_1228;
wire n_2319;
wire n_8924;
wire n_2965;
wire n_4955;
wire n_7555;
wire n_10114;
wire n_5410;
wire n_1251;
wire n_1989;
wire n_447;
wire n_2689;
wire n_6110;
wire n_1762;
wire n_6238;
wire n_7025;
wire n_3798;
wire n_3080;
wire n_8380;
wire n_9978;
wire n_5241;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_5331;
wire n_7478;
wire n_3308;
wire n_6326;
wire n_841;
wire n_3204;
wire n_7451;
wire n_9494;
wire n_4134;
wire n_5018;
wire n_6917;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;
wire n_6612;
wire n_5258;

INVx1_ASAP7_75t_L g123 ( 
.A(n_20),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_65),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_63),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_84),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_34),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_93),
.Y(n_129)
);

BUFx10_ASAP7_75t_L g130 ( 
.A(n_22),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_20),
.Y(n_131)
);

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_119),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_102),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_37),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_111),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_120),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_80),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_42),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_114),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_52),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_61),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_5),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_104),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_118),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_8),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_2),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_9),
.Y(n_151)
);

BUFx10_ASAP7_75t_L g152 ( 
.A(n_110),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_78),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_98),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_70),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_6),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_22),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_29),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_23),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_55),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_91),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_108),
.Y(n_162)
);

BUFx8_ASAP7_75t_SL g163 ( 
.A(n_82),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_116),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_11),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_31),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_16),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_50),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_57),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_87),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_51),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_86),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_38),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_97),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_58),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_45),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_117),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_18),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_33),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_69),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_113),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_95),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_23),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_60),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_100),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_27),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_6),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_48),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_89),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_44),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_122),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_17),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g193 ( 
.A(n_88),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_11),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_40),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_43),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_41),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_64),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_101),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_109),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_0),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_24),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_81),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_3),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_54),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_107),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_19),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_56),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_15),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_92),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_1),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_83),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_16),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g214 ( 
.A(n_46),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_99),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_24),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_4),
.Y(n_217)
);

BUFx10_ASAP7_75t_L g218 ( 
.A(n_21),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_94),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_90),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_5),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_27),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_12),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_49),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_72),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_13),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_121),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_14),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_53),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_112),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_71),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_30),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_8),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_13),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_115),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_77),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_3),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_67),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_85),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_26),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_14),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_39),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_9),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_225),
.Y(n_246)
);

INVxp33_ASAP7_75t_L g247 ( 
.A(n_123),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_163),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_159),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_186),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_129),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_163),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

BUFx2_ASAP7_75t_SL g255 ( 
.A(n_129),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_141),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_141),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_142),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_173),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_142),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_162),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_152),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_162),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_138),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_172),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_165),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_172),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_220),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_220),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_178),
.Y(n_270)
);

INVxp67_ASAP7_75t_SL g271 ( 
.A(n_156),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_233),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_131),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_232),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_231),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_146),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_231),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_149),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_256),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_251),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_256),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_257),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

NOR2xp67_ASAP7_75t_L g284 ( 
.A(n_248),
.B(n_128),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_258),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_252),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_264),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_258),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_260),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_255),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_255),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_R g292 ( 
.A(n_259),
.B(n_138),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_273),
.Y(n_293)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_266),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_276),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_278),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_249),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_262),
.B(n_195),
.Y(n_299)
);

BUFx6f_ASAP7_75t_SL g300 ( 
.A(n_244),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_270),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_259),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_262),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_260),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_261),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_262),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_261),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_263),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_263),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_262),
.B(n_271),
.Y(n_310)
);

NOR2xp67_ASAP7_75t_L g311 ( 
.A(n_278),
.B(n_128),
.Y(n_311)
);

INVxp33_ASAP7_75t_L g312 ( 
.A(n_247),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_244),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_244),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_265),
.Y(n_315)
);

NOR2xp67_ASAP7_75t_L g316 ( 
.A(n_246),
.B(n_124),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_246),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_279),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_303),
.A2(n_196),
.B1(n_203),
.B2(n_182),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_299),
.B(n_274),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_274),
.Y(n_322)
);

AND2x4_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_156),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_292),
.Y(n_324)
);

CKINVDCx11_ASAP7_75t_R g325 ( 
.A(n_280),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_297),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_279),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_312),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_281),
.Y(n_329)
);

AND2x4_ASAP7_75t_L g330 ( 
.A(n_311),
.B(n_150),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_293),
.A2(n_233),
.B1(n_211),
.B2(n_209),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_281),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_282),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_282),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_294),
.B(n_265),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_298),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_283),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_283),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_296),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_285),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_301),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_285),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_288),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_287),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_290),
.B(n_267),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_288),
.Y(n_346)
);

NOR2x1_ASAP7_75t_L g347 ( 
.A(n_284),
.B(n_166),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_289),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_289),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_304),
.Y(n_350)
);

AND2x4_ASAP7_75t_L g351 ( 
.A(n_316),
.B(n_150),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_313),
.B(n_244),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_304),
.Y(n_353)
);

AND2x4_ASAP7_75t_L g354 ( 
.A(n_315),
.B(n_217),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_305),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_305),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_307),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_291),
.B(n_267),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_302),
.Y(n_359)
);

INVxp33_ASAP7_75t_SL g360 ( 
.A(n_295),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_307),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_308),
.B(n_245),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_308),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_309),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_314),
.B(n_244),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_309),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_315),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_300),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_286),
.B(n_245),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_300),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_300),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_279),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_298),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_299),
.B(n_244),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_310),
.B(n_217),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_310),
.B(n_250),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_293),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_297),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_279),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_279),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_279),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_303),
.A2(n_166),
.B1(n_180),
.B2(n_182),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_297),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_299),
.B(n_268),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_297),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_297),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_280),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_292),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_297),
.Y(n_389)
);

AND2x2_ASAP7_75t_SL g390 ( 
.A(n_299),
.B(n_167),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_297),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_312),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_293),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_279),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_310),
.B(n_250),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_303),
.A2(n_180),
.B1(n_196),
.B2(n_203),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_297),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_317),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_279),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_293),
.Y(n_400)
);

BUFx12f_ASAP7_75t_L g401 ( 
.A(n_293),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_297),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_279),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_312),
.B(n_253),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_299),
.B(n_268),
.Y(n_405)
);

BUFx8_ASAP7_75t_L g406 ( 
.A(n_300),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_279),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_279),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_297),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_317),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_279),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_292),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_312),
.B(n_253),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_297),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_297),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_280),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_280),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_279),
.Y(n_418)
);

BUFx8_ASAP7_75t_L g419 ( 
.A(n_300),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_292),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_312),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_312),
.B(n_254),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_279),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_312),
.B(n_254),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_310),
.B(n_277),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_297),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_279),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_279),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_310),
.B(n_277),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_297),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_279),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_279),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_297),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_279),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_293),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_279),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_279),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_408),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_318),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_318),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_318),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_361),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_361),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_373),
.B(n_328),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_354),
.B(n_187),
.Y(n_445)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_392),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_361),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_418),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_421),
.B(n_159),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_418),
.Y(n_450)
);

AOI21x1_ASAP7_75t_L g451 ( 
.A1(n_374),
.A2(n_275),
.B(n_269),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_337),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_418),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_390),
.B(n_269),
.Y(n_454)
);

AO22x2_ASAP7_75t_L g455 ( 
.A1(n_375),
.A2(n_275),
.B1(n_243),
.B2(n_241),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_434),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_434),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_344),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_390),
.B(n_125),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g460 ( 
.A(n_336),
.Y(n_460)
);

INVxp33_ASAP7_75t_SL g461 ( 
.A(n_339),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_434),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_436),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_436),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_436),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_327),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_327),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_332),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_332),
.Y(n_469)
);

AND3x2_ASAP7_75t_L g470 ( 
.A(n_324),
.B(n_194),
.C(n_213),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_342),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_342),
.Y(n_472)
);

BUFx10_ASAP7_75t_L g473 ( 
.A(n_339),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_346),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_346),
.Y(n_475)
);

INVx8_ASAP7_75t_L g476 ( 
.A(n_425),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_337),
.Y(n_477)
);

NAND2xp33_ASAP7_75t_L g478 ( 
.A(n_377),
.B(n_193),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_404),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_408),
.B(n_134),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_348),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_348),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_350),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_425),
.B(n_169),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_350),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_353),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_353),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_408),
.B(n_135),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_366),
.Y(n_489)
);

BUFx16f_ASAP7_75t_R g490 ( 
.A(n_325),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_425),
.B(n_198),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_366),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_377),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_408),
.B(n_136),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_367),
.Y(n_495)
);

NAND2xp33_ASAP7_75t_L g496 ( 
.A(n_393),
.B(n_400),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_367),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_360),
.B(n_151),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_406),
.Y(n_499)
);

NAND2xp33_ASAP7_75t_L g500 ( 
.A(n_393),
.B(n_400),
.Y(n_500)
);

AND3x2_ASAP7_75t_L g501 ( 
.A(n_324),
.B(n_234),
.C(n_222),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_372),
.Y(n_502)
);

NOR2x1p5_ASAP7_75t_L g503 ( 
.A(n_401),
.B(n_157),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_429),
.B(n_183),
.Y(n_504)
);

BUFx10_ASAP7_75t_L g505 ( 
.A(n_435),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_372),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_379),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_379),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_380),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_380),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_381),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_381),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_337),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_408),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_394),
.Y(n_515)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_337),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_394),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_399),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_399),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_403),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_403),
.Y(n_521)
);

AND2x2_ASAP7_75t_SL g522 ( 
.A(n_375),
.B(n_139),
.Y(n_522)
);

AOI21x1_ASAP7_75t_L g523 ( 
.A1(n_352),
.A2(n_170),
.B(n_238),
.Y(n_523)
);

NOR2x1p5_ASAP7_75t_L g524 ( 
.A(n_401),
.B(n_192),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_360),
.B(n_201),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_407),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_336),
.B(n_202),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_407),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_411),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_411),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_356),
.B(n_140),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_356),
.B(n_145),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_406),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_423),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_423),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_356),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_404),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_356),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_413),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_427),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_427),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_429),
.B(n_153),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_413),
.B(n_130),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_428),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_429),
.B(n_155),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_428),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_322),
.B(n_204),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_321),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_431),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_345),
.B(n_207),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_431),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_321),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_432),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_432),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_376),
.B(n_160),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_437),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_437),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_358),
.B(n_216),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_376),
.B(n_221),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_329),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_362),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_369),
.B(n_388),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_333),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_362),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_334),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_422),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_338),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_340),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_321),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_376),
.B(n_223),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_343),
.Y(n_571)
);

BUFx6f_ASAP7_75t_SL g572 ( 
.A(n_359),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_321),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_349),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_355),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_435),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_357),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_363),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_369),
.B(n_226),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_422),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_398),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_395),
.B(n_168),
.Y(n_582)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_398),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_364),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_406),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_395),
.B(n_228),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_326),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_398),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_398),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_395),
.B(n_171),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_388),
.B(n_237),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_410),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_378),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_412),
.B(n_130),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_375),
.B(n_177),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_383),
.Y(n_596)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_319),
.B(n_382),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_410),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_410),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_410),
.Y(n_600)
);

NAND3xp33_ASAP7_75t_L g601 ( 
.A(n_331),
.B(n_242),
.C(n_179),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_354),
.B(n_184),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_320),
.B(n_126),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_424),
.B(n_130),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_384),
.B(n_127),
.Y(n_605)
);

INVx1_ASAP7_75t_SL g606 ( 
.A(n_344),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_385),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_405),
.B(n_132),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_386),
.Y(n_609)
);

AOI21x1_ASAP7_75t_L g610 ( 
.A1(n_365),
.A2(n_235),
.B(n_189),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_323),
.B(n_133),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_389),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_424),
.B(n_218),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_391),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_397),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_412),
.B(n_218),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_402),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_409),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_414),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_415),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_426),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_430),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_323),
.B(n_137),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_433),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_368),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_368),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_371),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_371),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_370),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_354),
.A2(n_230),
.B1(n_219),
.B2(n_215),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_323),
.B(n_148),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_335),
.B(n_218),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_419),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_351),
.B(n_208),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_351),
.B(n_193),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_330),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_330),
.Y(n_637)
);

INVxp67_ASAP7_75t_L g638 ( 
.A(n_341),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_351),
.B(n_193),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_330),
.Y(n_640)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_420),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_347),
.B(n_193),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_419),
.Y(n_643)
);

AO21x2_ASAP7_75t_L g644 ( 
.A1(n_396),
.A2(n_214),
.B(n_152),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_419),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_420),
.Y(n_646)
);

NAND3xp33_ASAP7_75t_L g647 ( 
.A(n_359),
.B(n_147),
.C(n_236),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_387),
.B(n_193),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_325),
.B(n_152),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_387),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_416),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_416),
.B(n_143),
.Y(n_652)
);

INVx5_ASAP7_75t_L g653 ( 
.A(n_417),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_417),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_318),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_390),
.B(n_193),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_318),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_318),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_390),
.B(n_144),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_390),
.B(n_239),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_408),
.Y(n_661)
);

BUFx2_ASAP7_75t_L g662 ( 
.A(n_328),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_390),
.B(n_214),
.Y(n_663)
);

CKINVDCx6p67_ASAP7_75t_R g664 ( 
.A(n_401),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_318),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_390),
.B(n_154),
.Y(n_666)
);

NAND2xp33_ASAP7_75t_SL g667 ( 
.A(n_339),
.B(n_212),
.Y(n_667)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_328),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_408),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_354),
.B(n_232),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_318),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_318),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_373),
.B(n_214),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_318),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_390),
.B(n_229),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_390),
.B(n_0),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_318),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_318),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_337),
.Y(n_679)
);

OAI22xp33_ASAP7_75t_L g680 ( 
.A1(n_339),
.A2(n_227),
.B1(n_224),
.B2(n_210),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_404),
.Y(n_681)
);

AND2x6_ASAP7_75t_L g682 ( 
.A(n_368),
.B(n_193),
.Y(n_682)
);

INVx5_ASAP7_75t_L g683 ( 
.A(n_408),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_390),
.B(n_206),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_318),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_318),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_318),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_337),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_408),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_390),
.B(n_205),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_318),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_390),
.B(n_1),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_318),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_408),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_336),
.B(n_2),
.Y(n_695)
);

INVxp33_ASAP7_75t_SL g696 ( 
.A(n_339),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_390),
.B(n_200),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_318),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_354),
.B(n_4),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_390),
.B(n_7),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_318),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_390),
.B(n_199),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_318),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_318),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_318),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_318),
.Y(n_706)
);

NAND3xp33_ASAP7_75t_L g707 ( 
.A(n_322),
.B(n_176),
.C(n_191),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_390),
.B(n_197),
.Y(n_708)
);

OR2x6_ASAP7_75t_L g709 ( 
.A(n_401),
.B(n_7),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_318),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_318),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_318),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_390),
.B(n_190),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_404),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_318),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_373),
.B(n_188),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_318),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_318),
.Y(n_718)
);

OR2x6_ASAP7_75t_L g719 ( 
.A(n_401),
.B(n_10),
.Y(n_719)
);

NAND3xp33_ASAP7_75t_L g720 ( 
.A(n_322),
.B(n_181),
.C(n_175),
.Y(n_720)
);

INVxp67_ASAP7_75t_L g721 ( 
.A(n_328),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_318),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_390),
.B(n_185),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_318),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_318),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_318),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_452),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_499),
.B(n_10),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_466),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_607),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_516),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_607),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_516),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_461),
.B(n_174),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_476),
.B(n_164),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_476),
.B(n_562),
.Y(n_736)
);

INVx4_ASAP7_75t_L g737 ( 
.A(n_476),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_476),
.B(n_158),
.Y(n_738)
);

BUFx4f_ASAP7_75t_L g739 ( 
.A(n_664),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_653),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_466),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_516),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_468),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_468),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_469),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_461),
.B(n_161),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_560),
.B(n_12),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_469),
.Y(n_748)
);

INVx1_ASAP7_75t_SL g749 ( 
.A(n_446),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_696),
.B(n_15),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_471),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_452),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_493),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_452),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_696),
.B(n_17),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_460),
.B(n_18),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_498),
.B(n_19),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_615),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_560),
.B(n_21),
.Y(n_759)
);

AND2x6_ASAP7_75t_L g760 ( 
.A(n_699),
.B(n_62),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_662),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_676),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_653),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_471),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_474),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_452),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_615),
.Y(n_767)
);

INVx4_ASAP7_75t_L g768 ( 
.A(n_653),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_477),
.Y(n_769)
);

INVx5_ASAP7_75t_L g770 ( 
.A(n_477),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_543),
.B(n_25),
.Y(n_771)
);

INVx4_ASAP7_75t_L g772 ( 
.A(n_653),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_617),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_522),
.B(n_28),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_617),
.Y(n_775)
);

BUFx8_ASAP7_75t_SL g776 ( 
.A(n_493),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_522),
.B(n_32),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_525),
.B(n_35),
.Y(n_778)
);

CKINVDCx20_ASAP7_75t_R g779 ( 
.A(n_576),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_543),
.B(n_36),
.Y(n_780)
);

INVxp67_ASAP7_75t_L g781 ( 
.A(n_668),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_444),
.B(n_47),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_606),
.B(n_68),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_620),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_576),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_621),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_653),
.Y(n_787)
);

AND2x6_ASAP7_75t_L g788 ( 
.A(n_699),
.B(n_75),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_621),
.Y(n_789)
);

AND2x6_ASAP7_75t_L g790 ( 
.A(n_699),
.B(n_676),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_604),
.B(n_76),
.Y(n_791)
);

NAND3xp33_ASAP7_75t_L g792 ( 
.A(n_550),
.B(n_79),
.C(n_96),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_477),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_692),
.A2(n_103),
.B1(n_106),
.B2(n_700),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_477),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_474),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_664),
.Y(n_797)
);

BUFx2_ASAP7_75t_L g798 ( 
.A(n_458),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_473),
.Y(n_799)
);

INVx4_ASAP7_75t_SL g800 ( 
.A(n_682),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_613),
.B(n_632),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_563),
.B(n_567),
.Y(n_802)
);

INVxp67_ASAP7_75t_L g803 ( 
.A(n_632),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_622),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_475),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_622),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_624),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_563),
.B(n_567),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_475),
.Y(n_809)
);

INVx5_ASAP7_75t_L g810 ( 
.A(n_513),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_481),
.Y(n_811)
);

AND2x4_ASAP7_75t_L g812 ( 
.A(n_499),
.B(n_533),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_624),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_568),
.B(n_574),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_568),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_574),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_575),
.B(n_577),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_575),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_577),
.B(n_578),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_513),
.Y(n_820)
);

INVx4_ASAP7_75t_L g821 ( 
.A(n_683),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_473),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_663),
.B(n_479),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_578),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_449),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_663),
.B(n_638),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_479),
.B(n_537),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_692),
.A2(n_700),
.B1(n_459),
.B2(n_708),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_584),
.Y(n_829)
);

INVx5_ASAP7_75t_L g830 ( 
.A(n_513),
.Y(n_830)
);

CKINVDCx16_ASAP7_75t_R g831 ( 
.A(n_473),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_533),
.B(n_585),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_537),
.B(n_539),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_481),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_482),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_584),
.Y(n_836)
);

CKINVDCx16_ASAP7_75t_R g837 ( 
.A(n_505),
.Y(n_837)
);

INVx8_ASAP7_75t_L g838 ( 
.A(n_572),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_587),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_539),
.B(n_566),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_558),
.B(n_721),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_439),
.B(n_440),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_513),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_482),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_593),
.Y(n_845)
);

AND2x6_ASAP7_75t_L g846 ( 
.A(n_585),
.B(n_439),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_505),
.Y(n_847)
);

AND2x6_ASAP7_75t_L g848 ( 
.A(n_440),
.B(n_442),
.Y(n_848)
);

BUFx10_ASAP7_75t_L g849 ( 
.A(n_572),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_596),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_459),
.A2(n_597),
.B1(n_713),
.B2(n_708),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_566),
.B(n_580),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_505),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_713),
.B(n_652),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_679),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_609),
.Y(n_856)
);

INVx4_ASAP7_75t_L g857 ( 
.A(n_683),
.Y(n_857)
);

OR2x2_ASAP7_75t_L g858 ( 
.A(n_650),
.B(n_651),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_SL g859 ( 
.A1(n_455),
.A2(n_579),
.B1(n_660),
.B2(n_659),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_612),
.Y(n_860)
);

INVx6_ASAP7_75t_L g861 ( 
.A(n_503),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_580),
.B(n_681),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_679),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_681),
.B(n_714),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_679),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_442),
.B(n_443),
.Y(n_866)
);

NAND3xp33_ASAP7_75t_SL g867 ( 
.A(n_527),
.B(n_547),
.C(n_591),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_656),
.A2(n_714),
.B1(n_545),
.B2(n_555),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_641),
.B(n_679),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_650),
.Y(n_870)
);

INVx6_ASAP7_75t_L g871 ( 
.A(n_524),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_614),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_618),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_688),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_656),
.A2(n_590),
.B1(n_545),
.B2(n_555),
.Y(n_875)
);

INVx4_ASAP7_75t_L g876 ( 
.A(n_683),
.Y(n_876)
);

CKINVDCx16_ASAP7_75t_R g877 ( 
.A(n_572),
.Y(n_877)
);

INVx3_ASAP7_75t_L g878 ( 
.A(n_688),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_485),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_619),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_651),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_688),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_688),
.B(n_695),
.Y(n_883)
);

INVx1_ASAP7_75t_SL g884 ( 
.A(n_654),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_443),
.B(n_448),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_666),
.B(n_675),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_633),
.B(n_643),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_448),
.B(n_453),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_667),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_565),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_625),
.Y(n_891)
);

NAND2xp33_ASAP7_75t_SL g892 ( 
.A(n_684),
.B(n_690),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_453),
.B(n_456),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_571),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_487),
.Y(n_895)
);

NAND2x1_ASAP7_75t_L g896 ( 
.A(n_583),
.B(n_438),
.Y(n_896)
);

AO21x2_ASAP7_75t_L g897 ( 
.A1(n_642),
.A2(n_610),
.B(n_523),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_467),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_487),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_456),
.B(n_457),
.Y(n_900)
);

AND2x6_ASAP7_75t_L g901 ( 
.A(n_457),
.B(n_462),
.Y(n_901)
);

INVx5_ASAP7_75t_L g902 ( 
.A(n_682),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_697),
.B(n_702),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_581),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_489),
.Y(n_905)
);

AND2x6_ASAP7_75t_L g906 ( 
.A(n_462),
.B(n_463),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_463),
.B(n_464),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_625),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_594),
.B(n_616),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_625),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_472),
.Y(n_911)
);

AND2x2_ASAP7_75t_SL g912 ( 
.A(n_496),
.B(n_500),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_625),
.Y(n_913)
);

INVx5_ASAP7_75t_L g914 ( 
.A(n_682),
.Y(n_914)
);

INVxp67_ASAP7_75t_SL g915 ( 
.A(n_581),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_483),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_489),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_581),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_486),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_723),
.B(n_648),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_496),
.B(n_500),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_648),
.B(n_673),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_492),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_502),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_646),
.B(n_629),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_495),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_628),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_506),
.Y(n_928)
);

CKINVDCx16_ASAP7_75t_R g929 ( 
.A(n_649),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_629),
.B(n_484),
.Y(n_930)
);

INVx4_ASAP7_75t_SL g931 ( 
.A(n_682),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_508),
.Y(n_932)
);

INVx1_ASAP7_75t_SL g933 ( 
.A(n_454),
.Y(n_933)
);

INVx4_ASAP7_75t_L g934 ( 
.A(n_683),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_509),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_512),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_515),
.Y(n_937)
);

INVx6_ASAP7_75t_L g938 ( 
.A(n_709),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_491),
.B(n_716),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_683),
.B(n_581),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_633),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_634),
.B(n_542),
.Y(n_942)
);

INVxp67_ASAP7_75t_L g943 ( 
.A(n_542),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_582),
.A2(n_590),
.B1(n_478),
.B2(n_595),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_445),
.B(n_561),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_517),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_643),
.B(n_645),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_464),
.B(n_465),
.Y(n_948)
);

BUFx4f_ASAP7_75t_L g949 ( 
.A(n_709),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_645),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_628),
.Y(n_951)
);

INVx2_ASAP7_75t_SL g952 ( 
.A(n_670),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_465),
.B(n_655),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_634),
.B(n_582),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_640),
.B(n_636),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_640),
.B(n_595),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_564),
.B(n_637),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_455),
.A2(n_534),
.B1(n_530),
.B2(n_529),
.Y(n_958)
);

OR2x2_ASAP7_75t_L g959 ( 
.A(n_504),
.B(n_559),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_667),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_628),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_445),
.B(n_570),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_655),
.B(n_657),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_495),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_586),
.B(n_602),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_628),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_520),
.Y(n_967)
);

NAND3xp33_ASAP7_75t_SL g968 ( 
.A(n_601),
.B(n_630),
.C(n_605),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_521),
.Y(n_969)
);

INVx1_ASAP7_75t_SL g970 ( 
.A(n_670),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_526),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_535),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_445),
.B(n_455),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_657),
.B(n_658),
.Y(n_974)
);

OR2x2_ASAP7_75t_L g975 ( 
.A(n_670),
.B(n_602),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_583),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_541),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_546),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_649),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_551),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_583),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_658),
.B(n_672),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_611),
.B(n_623),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_631),
.B(n_680),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_470),
.B(n_501),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_709),
.B(n_719),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_672),
.B(n_677),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_536),
.B(n_538),
.Y(n_988)
);

INVxp67_ASAP7_75t_SL g989 ( 
.A(n_536),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_497),
.Y(n_990)
);

OR2x6_ASAP7_75t_L g991 ( 
.A(n_709),
.B(n_719),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_719),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_536),
.B(n_538),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_719),
.B(n_644),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_497),
.Y(n_995)
);

NOR2x1p5_ASAP7_75t_L g996 ( 
.A(n_490),
.B(n_647),
.Y(n_996)
);

BUFx2_ASAP7_75t_L g997 ( 
.A(n_644),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_677),
.B(n_678),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_626),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_678),
.B(n_686),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_626),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_556),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_507),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_627),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_686),
.B(n_698),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_507),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_538),
.B(n_438),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_608),
.B(n_603),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_510),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_510),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_698),
.B(n_701),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_438),
.B(n_514),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_514),
.B(n_661),
.Y(n_1013)
);

OR2x2_ASAP7_75t_L g1014 ( 
.A(n_635),
.B(n_639),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_701),
.B(n_703),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_557),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_511),
.Y(n_1017)
);

NAND3x1_ASAP7_75t_L g1018 ( 
.A(n_548),
.B(n_600),
.C(n_552),
.Y(n_1018)
);

BUFx3_ASAP7_75t_L g1019 ( 
.A(n_627),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_511),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_514),
.B(n_669),
.Y(n_1021)
);

INVx4_ASAP7_75t_SL g1022 ( 
.A(n_682),
.Y(n_1022)
);

NAND3xp33_ASAP7_75t_L g1023 ( 
.A(n_478),
.B(n_441),
.C(n_447),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_703),
.B(n_725),
.Y(n_1024)
);

BUFx3_ASAP7_75t_L g1025 ( 
.A(n_548),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_518),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_588),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_635),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_661),
.Y(n_1029)
);

OR2x2_ASAP7_75t_L g1030 ( 
.A(n_639),
.B(n_544),
.Y(n_1030)
);

INVx5_ASAP7_75t_L g1031 ( 
.A(n_682),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_642),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_450),
.B(n_726),
.Y(n_1033)
);

INVx1_ASAP7_75t_SL g1034 ( 
.A(n_588),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_518),
.B(n_534),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_519),
.Y(n_1036)
);

AND2x6_ASAP7_75t_L g1037 ( 
.A(n_705),
.B(n_725),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_519),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_661),
.B(n_669),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_528),
.Y(n_1040)
);

AND2x6_ASAP7_75t_L g1041 ( 
.A(n_705),
.B(n_724),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_669),
.B(n_694),
.Y(n_1042)
);

BUFx10_ASAP7_75t_L g1043 ( 
.A(n_665),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_689),
.Y(n_1044)
);

CKINVDCx20_ASAP7_75t_R g1045 ( 
.A(n_531),
.Y(n_1045)
);

INVx2_ASAP7_75t_SL g1046 ( 
.A(n_548),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_528),
.Y(n_1047)
);

BUFx10_ASAP7_75t_L g1048 ( 
.A(n_671),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_706),
.B(n_724),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_674),
.B(n_722),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_529),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_706),
.B(n_715),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_710),
.B(n_715),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_530),
.B(n_540),
.Y(n_1054)
);

NOR2x1p5_ASAP7_75t_L g1055 ( 
.A(n_707),
.B(n_720),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_685),
.B(n_693),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_540),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_544),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_710),
.B(n_718),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_549),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_549),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_717),
.B(n_718),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_717),
.B(n_712),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_553),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_553),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_554),
.Y(n_1066)
);

INVx1_ASAP7_75t_SL g1067 ( 
.A(n_589),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_589),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_552),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_687),
.B(n_711),
.Y(n_1070)
);

OR2x2_ASAP7_75t_L g1071 ( 
.A(n_554),
.B(n_531),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_592),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_691),
.A2(n_704),
.B1(n_694),
.B2(n_689),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_552),
.B(n_573),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_569),
.Y(n_1075)
);

AO22x2_ASAP7_75t_L g1076 ( 
.A1(n_592),
.A2(n_599),
.B1(n_598),
.B2(n_532),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_569),
.B(n_573),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_598),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_569),
.B(n_573),
.Y(n_1079)
);

INVx4_ASAP7_75t_L g1080 ( 
.A(n_689),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_694),
.B(n_599),
.Y(n_1081)
);

INVx4_ASAP7_75t_SL g1082 ( 
.A(n_480),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_532),
.B(n_480),
.Y(n_1083)
);

AOI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_488),
.A2(n_676),
.B1(n_700),
.B2(n_692),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_494),
.B(n_488),
.Y(n_1085)
);

BUFx2_ASAP7_75t_L g1086 ( 
.A(n_494),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_451),
.B(n_360),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_607),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_461),
.B(n_360),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_607),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_607),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_821),
.Y(n_1092)
);

OR2x6_ASAP7_75t_L g1093 ( 
.A(n_737),
.B(n_838),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_841),
.B(n_933),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1089),
.B(n_826),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_729),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_909),
.B(n_939),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_794),
.B(n_912),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_839),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_825),
.B(n_867),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_794),
.B(n_851),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_845),
.Y(n_1102)
);

INVxp33_ASAP7_75t_L g1103 ( 
.A(n_798),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_933),
.B(n_801),
.Y(n_1104)
);

AND2x6_ASAP7_75t_SL g1105 ( 
.A(n_991),
.B(n_750),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_851),
.B(n_944),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_757),
.A2(n_778),
.B(n_984),
.C(n_922),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_886),
.B(n_903),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_850),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_856),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_944),
.B(n_828),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_828),
.B(n_902),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_867),
.A2(n_825),
.B(n_803),
.C(n_774),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_761),
.B(n_803),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_1084),
.A2(n_1008),
.B1(n_854),
.B2(n_989),
.Y(n_1115)
);

BUFx8_ASAP7_75t_L g1116 ( 
.A(n_790),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_860),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_790),
.B(n_945),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_902),
.B(n_914),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_790),
.B(n_930),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_761),
.B(n_970),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_989),
.A2(n_875),
.B1(n_959),
.B2(n_868),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_790),
.B(n_823),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_872),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_973),
.B(n_749),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_965),
.B(n_962),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_920),
.A2(n_762),
.B(n_983),
.C(n_875),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_776),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_942),
.B(n_954),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_902),
.B(n_914),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_762),
.A2(n_968),
.B(n_755),
.C(n_868),
.Y(n_1131)
);

NOR3xp33_ASAP7_75t_L g1132 ( 
.A(n_968),
.B(n_746),
.C(n_734),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_859),
.A2(n_1045),
.B1(n_870),
.B2(n_955),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_821),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_741),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_873),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_943),
.B(n_833),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_770),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_739),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_736),
.A2(n_890),
.B1(n_894),
.B2(n_859),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_902),
.B(n_914),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_743),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_744),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_914),
.B(n_1031),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_943),
.B(n_840),
.Y(n_1145)
);

BUFx8_ASAP7_75t_L g1146 ( 
.A(n_921),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_880),
.Y(n_1147)
);

AOI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_889),
.A2(n_960),
.B1(n_1087),
.B2(n_753),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_730),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_1031),
.B(n_770),
.Y(n_1150)
);

NOR3xp33_ASAP7_75t_L g1151 ( 
.A(n_756),
.B(n_777),
.C(n_929),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_862),
.B(n_925),
.Y(n_1152)
);

NOR2x1p5_ASAP7_75t_L g1153 ( 
.A(n_797),
.B(n_785),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_779),
.A2(n_749),
.B1(n_884),
.B2(n_781),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_732),
.Y(n_1155)
);

AOI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_955),
.A2(n_970),
.B1(n_884),
.B2(n_958),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_957),
.B(n_771),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_781),
.B(n_728),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1031),
.B(n_770),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_745),
.Y(n_1160)
);

NAND2xp33_ASAP7_75t_SL g1161 ( 
.A(n_737),
.B(n_1055),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_975),
.B(n_952),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_956),
.B(n_802),
.Y(n_1163)
);

INVxp67_ASAP7_75t_L g1164 ( 
.A(n_858),
.Y(n_1164)
);

INVx2_ASAP7_75t_SL g1165 ( 
.A(n_739),
.Y(n_1165)
);

INVx2_ASAP7_75t_SL g1166 ( 
.A(n_838),
.Y(n_1166)
);

AND2x2_ASAP7_75t_SL g1167 ( 
.A(n_949),
.B(n_994),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_979),
.B(n_847),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_802),
.B(n_808),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_758),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_748),
.Y(n_1171)
);

OAI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_991),
.A2(n_949),
.B1(n_837),
.B2(n_831),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_751),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_767),
.Y(n_1174)
);

INVxp67_ASAP7_75t_L g1175 ( 
.A(n_881),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_764),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_958),
.A2(n_950),
.B1(n_947),
.B2(n_775),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_1031),
.B(n_770),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_810),
.B(n_830),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_810),
.B(n_830),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_808),
.B(n_814),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_765),
.Y(n_1182)
);

A2O1A1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_780),
.A2(n_792),
.B(n_892),
.C(n_791),
.Y(n_1183)
);

INVxp67_ASAP7_75t_L g1184 ( 
.A(n_783),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_796),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_814),
.B(n_817),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_812),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_773),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_810),
.B(n_830),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_817),
.B(n_819),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_792),
.A2(n_747),
.B(n_759),
.C(n_1033),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_784),
.B(n_786),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_728),
.B(n_991),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1023),
.A2(n_1069),
.B1(n_1056),
.B2(n_1050),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_789),
.B(n_804),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_810),
.B(n_830),
.Y(n_1196)
);

OAI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1023),
.A2(n_1081),
.B(n_866),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_806),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_904),
.B(n_918),
.Y(n_1199)
);

INVx8_ASAP7_75t_L g1200 ( 
.A(n_838),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_853),
.B(n_877),
.Y(n_1201)
);

NOR2xp67_ASAP7_75t_L g1202 ( 
.A(n_822),
.B(n_763),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_807),
.B(n_813),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1088),
.Y(n_1204)
);

NAND3xp33_ASAP7_75t_L g1205 ( 
.A(n_747),
.B(n_759),
.C(n_782),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_842),
.A2(n_885),
.B(n_866),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_805),
.Y(n_1207)
);

INVx8_ASAP7_75t_L g1208 ( 
.A(n_760),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1090),
.B(n_1091),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_986),
.B(n_812),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_904),
.B(n_918),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_809),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_904),
.B(n_918),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_827),
.B(n_852),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_999),
.B(n_1001),
.Y(n_1215)
);

INVx8_ASAP7_75t_L g1216 ( 
.A(n_760),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_815),
.B(n_816),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_811),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_818),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_834),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_727),
.B(n_754),
.Y(n_1221)
);

OAI221xp5_ASAP7_75t_L g1222 ( 
.A1(n_864),
.A2(n_992),
.B1(n_938),
.B2(n_799),
.C(n_941),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_887),
.B(n_938),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_824),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_835),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_887),
.B(n_947),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_832),
.B(n_988),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_832),
.B(n_985),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_844),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_735),
.B(n_738),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_727),
.B(n_754),
.Y(n_1231)
);

NAND2xp33_ASAP7_75t_L g1232 ( 
.A(n_760),
.B(n_788),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_SL g1233 ( 
.A(n_727),
.B(n_754),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_SL g1234 ( 
.A(n_763),
.B(n_768),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1086),
.B(n_996),
.Y(n_1235)
);

XNOR2xp5_ASAP7_75t_L g1236 ( 
.A(n_997),
.B(n_1032),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_829),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_836),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1034),
.B(n_1067),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1034),
.B(n_1067),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1081),
.A2(n_885),
.B(n_842),
.Y(n_1241)
);

NOR3xp33_ASAP7_75t_L g1242 ( 
.A(n_883),
.B(n_869),
.C(n_738),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1004),
.A2(n_1019),
.B1(n_788),
.B2(n_760),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_788),
.A2(n_980),
.B1(n_971),
.B2(n_969),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_861),
.B(n_871),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_898),
.Y(n_1246)
);

NOR2x1p5_ASAP7_75t_L g1247 ( 
.A(n_768),
.B(n_772),
.Y(n_1247)
);

INVxp67_ASAP7_75t_L g1248 ( 
.A(n_1027),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_911),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_735),
.B(n_988),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_766),
.B(n_769),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_888),
.A2(n_900),
.B(n_893),
.Y(n_1252)
);

NOR2xp67_ASAP7_75t_L g1253 ( 
.A(n_772),
.B(n_740),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_916),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_766),
.B(n_769),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_766),
.B(n_769),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_788),
.A2(n_977),
.B1(n_972),
.B2(n_967),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_879),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_919),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_793),
.B(n_795),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_793),
.B(n_795),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_923),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_846),
.B(n_924),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_895),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_976),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_899),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_928),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_857),
.Y(n_1268)
);

OR2x2_ASAP7_75t_L g1269 ( 
.A(n_932),
.B(n_935),
.Y(n_1269)
);

INVx2_ASAP7_75t_SL g1270 ( 
.A(n_849),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_993),
.B(n_1007),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_793),
.B(n_795),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_846),
.B(n_936),
.Y(n_1273)
);

INVxp67_ASAP7_75t_SL g1274 ( 
.A(n_915),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_905),
.Y(n_1275)
);

NOR2xp67_ASAP7_75t_L g1276 ( 
.A(n_787),
.B(n_752),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_917),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_937),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_820),
.B(n_843),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_846),
.B(n_946),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_978),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_846),
.B(n_1002),
.Y(n_1282)
);

INVxp33_ASAP7_75t_L g1283 ( 
.A(n_993),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1016),
.B(n_1035),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1068),
.B(n_1007),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_926),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_976),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1012),
.B(n_1013),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1012),
.B(n_1013),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_820),
.B(n_843),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1020),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_SL g1292 ( 
.A(n_849),
.Y(n_1292)
);

INVxp67_ASAP7_75t_L g1293 ( 
.A(n_1021),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_861),
.B(n_871),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1036),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1038),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1021),
.B(n_1039),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1039),
.B(n_1042),
.Y(n_1298)
);

OAI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1014),
.A2(n_1085),
.B1(n_1028),
.B2(n_1070),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1083),
.B(n_1042),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1040),
.Y(n_1301)
);

INVx2_ASAP7_75t_SL g1302 ( 
.A(n_1025),
.Y(n_1302)
);

NAND2xp33_ASAP7_75t_L g1303 ( 
.A(n_848),
.B(n_901),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_900),
.B(n_907),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_964),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1047),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_990),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1051),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1029),
.B(n_1075),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1057),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_820),
.B(n_843),
.Y(n_1311)
);

INVxp33_ASAP7_75t_L g1312 ( 
.A(n_1074),
.Y(n_1312)
);

OAI221xp5_ASAP7_75t_L g1313 ( 
.A1(n_1073),
.A2(n_1085),
.B1(n_1070),
.B2(n_1063),
.C(n_1079),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_855),
.B(n_865),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_907),
.B(n_948),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_948),
.B(n_953),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_953),
.B(n_963),
.Y(n_1317)
);

NOR2xp67_ASAP7_75t_L g1318 ( 
.A(n_752),
.B(n_863),
.Y(n_1318)
);

AND2x4_ASAP7_75t_SL g1319 ( 
.A(n_976),
.B(n_857),
.Y(n_1319)
);

BUFx2_ASAP7_75t_L g1320 ( 
.A(n_915),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_963),
.B(n_974),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_974),
.B(n_982),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_982),
.B(n_987),
.Y(n_1323)
);

AOI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_848),
.A2(n_1041),
.B1(n_906),
.B2(n_901),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1054),
.B(n_1060),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1065),
.B(n_1066),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_987),
.B(n_998),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_998),
.B(n_1000),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_995),
.Y(n_1329)
);

INVx4_ASAP7_75t_L g1330 ( 
.A(n_876),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1003),
.B(n_1006),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1009),
.Y(n_1332)
);

AO22x2_ASAP7_75t_L g1333 ( 
.A1(n_1082),
.A2(n_1073),
.B1(n_1017),
.B2(n_1026),
.Y(n_1333)
);

INVxp67_ASAP7_75t_L g1334 ( 
.A(n_1072),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1000),
.B(n_1011),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_855),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1010),
.Y(n_1337)
);

A2O1A1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1005),
.A2(n_1015),
.B(n_1011),
.C(n_1052),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1005),
.B(n_1015),
.Y(n_1339)
);

OAI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1063),
.A2(n_1030),
.B1(n_1052),
.B2(n_1053),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1053),
.B(n_1059),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1058),
.Y(n_1342)
);

INVxp33_ASAP7_75t_L g1343 ( 
.A(n_1077),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_855),
.B(n_865),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1059),
.B(n_731),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1061),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_731),
.B(n_733),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_865),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1064),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_733),
.B(n_742),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1071),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_SL g1352 ( 
.A(n_874),
.B(n_882),
.Y(n_1352)
);

OAI22x1_ASAP7_75t_R g1353 ( 
.A1(n_1043),
.A2(n_1048),
.B1(n_1018),
.B2(n_1044),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_742),
.B(n_981),
.Y(n_1354)
);

AOI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_848),
.A2(n_906),
.B1(n_901),
.B2(n_1037),
.Y(n_1355)
);

AOI221xp5_ASAP7_75t_L g1356 ( 
.A1(n_1024),
.A2(n_1062),
.B1(n_1049),
.B2(n_1046),
.C(n_1076),
.Y(n_1356)
);

NAND2xp33_ASAP7_75t_L g1357 ( 
.A(n_848),
.B(n_906),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_981),
.B(n_1029),
.Y(n_1358)
);

BUFx5_ASAP7_75t_L g1359 ( 
.A(n_901),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_906),
.B(n_1037),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1078),
.A2(n_1076),
.B1(n_1041),
.B2(n_1037),
.Y(n_1361)
);

INVx8_ASAP7_75t_L g1362 ( 
.A(n_1037),
.Y(n_1362)
);

NAND2x1p5_ASAP7_75t_L g1363 ( 
.A(n_876),
.B(n_934),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1041),
.B(n_1080),
.Y(n_1364)
);

INVx8_ASAP7_75t_L g1365 ( 
.A(n_1041),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1044),
.B(n_1080),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_SL g1367 ( 
.A(n_874),
.B(n_882),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1043),
.Y(n_1368)
);

AOI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_863),
.A2(n_878),
.B1(n_891),
.B2(n_927),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_SL g1370 ( 
.A(n_874),
.B(n_882),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1044),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_878),
.Y(n_1372)
);

O2A1O1Ixp5_ASAP7_75t_L g1373 ( 
.A1(n_940),
.A2(n_896),
.B(n_934),
.C(n_891),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_951),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_951),
.Y(n_1375)
);

NAND2x1p5_ASAP7_75t_L g1376 ( 
.A(n_951),
.B(n_961),
.Y(n_1376)
);

INVx1_ASAP7_75t_SL g1377 ( 
.A(n_1082),
.Y(n_1377)
);

NOR2xp67_ASAP7_75t_SL g1378 ( 
.A(n_961),
.B(n_927),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1082),
.B(n_966),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_908),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_908),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1048),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_910),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_SL g1384 ( 
.A(n_800),
.B(n_931),
.Y(n_1384)
);

INVxp67_ASAP7_75t_L g1385 ( 
.A(n_961),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_910),
.B(n_913),
.Y(n_1386)
);

NOR2xp67_ASAP7_75t_L g1387 ( 
.A(n_913),
.B(n_966),
.Y(n_1387)
);

AOI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_800),
.A2(n_931),
.B1(n_1022),
.B2(n_897),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_897),
.Y(n_1389)
);

AND2x6_ASAP7_75t_L g1390 ( 
.A(n_800),
.B(n_931),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1022),
.B(n_841),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1022),
.A2(n_939),
.B1(n_841),
.B2(n_390),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_841),
.B(n_933),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_737),
.B(n_921),
.Y(n_1394)
);

INVxp67_ASAP7_75t_L g1395 ( 
.A(n_749),
.Y(n_1395)
);

BUFx6f_ASAP7_75t_SL g1396 ( 
.A(n_812),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_841),
.B(n_933),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_794),
.B(n_912),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_757),
.A2(n_377),
.B1(n_393),
.B2(n_339),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_841),
.B(n_933),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_841),
.B(n_933),
.Y(n_1401)
);

BUFx2_ASAP7_75t_L g1402 ( 
.A(n_761),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_SL g1403 ( 
.A(n_794),
.B(n_912),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_821),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_839),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_841),
.B(n_933),
.Y(n_1406)
);

NOR3xp33_ASAP7_75t_L g1407 ( 
.A(n_867),
.B(n_757),
.C(n_841),
.Y(n_1407)
);

INVx2_ASAP7_75t_SL g1408 ( 
.A(n_739),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_839),
.Y(n_1409)
);

INVx3_ASAP7_75t_L g1410 ( 
.A(n_821),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_841),
.B(n_461),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_839),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1089),
.B(n_312),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_859),
.A2(n_597),
.B1(n_663),
.B2(n_676),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_841),
.B(n_933),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_841),
.B(n_461),
.Y(n_1416)
);

AO22x2_ASAP7_75t_L g1417 ( 
.A1(n_994),
.A2(n_663),
.B1(n_692),
.B2(n_676),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_841),
.B(n_933),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_SL g1419 ( 
.A(n_794),
.B(n_912),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_839),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_841),
.B(n_461),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_729),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_839),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_841),
.B(n_461),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_SL g1425 ( 
.A(n_794),
.B(n_912),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_770),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_739),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_794),
.B(n_912),
.Y(n_1428)
);

INVx2_ASAP7_75t_SL g1429 ( 
.A(n_739),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_839),
.Y(n_1430)
);

BUFx6f_ASAP7_75t_SL g1431 ( 
.A(n_812),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_841),
.B(n_933),
.Y(n_1432)
);

NAND2xp33_ASAP7_75t_L g1433 ( 
.A(n_760),
.B(n_788),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_841),
.B(n_933),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_SL g1435 ( 
.A(n_794),
.B(n_912),
.Y(n_1435)
);

INVx4_ASAP7_75t_L g1436 ( 
.A(n_737),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_939),
.A2(n_841),
.B1(n_390),
.B2(n_778),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_SL g1438 ( 
.A(n_794),
.B(n_912),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_939),
.A2(n_841),
.B1(n_390),
.B2(n_778),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_SL g1440 ( 
.A(n_794),
.B(n_912),
.Y(n_1440)
);

INVxp67_ASAP7_75t_L g1441 ( 
.A(n_749),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_729),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_729),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_SL g1444 ( 
.A(n_794),
.B(n_912),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_839),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_841),
.B(n_933),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_859),
.A2(n_597),
.B1(n_663),
.B2(n_676),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_SL g1448 ( 
.A(n_794),
.B(n_912),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_SL g1449 ( 
.A(n_794),
.B(n_912),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_839),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1089),
.B(n_312),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_761),
.Y(n_1452)
);

NAND3xp33_ASAP7_75t_L g1453 ( 
.A(n_757),
.B(n_841),
.C(n_558),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_841),
.B(n_933),
.Y(n_1454)
);

INVx2_ASAP7_75t_SL g1455 ( 
.A(n_739),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_729),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_SL g1457 ( 
.A(n_812),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_841),
.B(n_461),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_839),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_SL g1460 ( 
.A(n_794),
.B(n_912),
.Y(n_1460)
);

NOR3xp33_ASAP7_75t_L g1461 ( 
.A(n_867),
.B(n_757),
.C(n_841),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_841),
.B(n_933),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_839),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_SL g1464 ( 
.A(n_794),
.B(n_912),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_729),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_729),
.Y(n_1466)
);

INVxp67_ASAP7_75t_L g1467 ( 
.A(n_749),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_841),
.B(n_933),
.Y(n_1468)
);

INVxp33_ASAP7_75t_L g1469 ( 
.A(n_826),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_SL g1470 ( 
.A(n_794),
.B(n_912),
.Y(n_1470)
);

AOI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_757),
.A2(n_377),
.B1(n_393),
.B2(n_339),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1089),
.B(n_312),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_SL g1473 ( 
.A(n_794),
.B(n_912),
.Y(n_1473)
);

INVxp67_ASAP7_75t_L g1474 ( 
.A(n_749),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_794),
.B(n_912),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_841),
.B(n_933),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1089),
.B(n_312),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_841),
.B(n_933),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_729),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_841),
.B(n_933),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_729),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_794),
.B(n_912),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_839),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_841),
.B(n_933),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_841),
.B(n_933),
.Y(n_1485)
);

INVxp67_ASAP7_75t_L g1486 ( 
.A(n_749),
.Y(n_1486)
);

INVxp67_ASAP7_75t_L g1487 ( 
.A(n_749),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_729),
.Y(n_1488)
);

INVx2_ASAP7_75t_SL g1489 ( 
.A(n_739),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_841),
.B(n_933),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_729),
.Y(n_1491)
);

O2A1O1Ixp33_ASAP7_75t_L g1492 ( 
.A1(n_757),
.A2(n_867),
.B(n_841),
.C(n_558),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_841),
.B(n_933),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_729),
.Y(n_1494)
);

NAND3xp33_ASAP7_75t_SL g1495 ( 
.A(n_757),
.B(n_377),
.C(n_339),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_839),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_739),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_839),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_839),
.Y(n_1499)
);

NOR2xp67_ASAP7_75t_L g1500 ( 
.A(n_797),
.B(n_401),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_841),
.B(n_933),
.Y(n_1501)
);

AND2x4_ASAP7_75t_SL g1502 ( 
.A(n_737),
.B(n_812),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1089),
.B(n_312),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_841),
.B(n_461),
.Y(n_1504)
);

INVx3_ASAP7_75t_L g1505 ( 
.A(n_821),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_SL g1506 ( 
.A(n_797),
.B(n_401),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_841),
.B(n_933),
.Y(n_1507)
);

NOR2x1p5_ASAP7_75t_L g1508 ( 
.A(n_797),
.B(n_664),
.Y(n_1508)
);

NAND2xp33_ASAP7_75t_L g1509 ( 
.A(n_760),
.B(n_788),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_841),
.B(n_933),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_SL g1511 ( 
.A(n_794),
.B(n_912),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_839),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_841),
.B(n_933),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_SL g1514 ( 
.A(n_794),
.B(n_912),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_841),
.B(n_933),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_729),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_841),
.B(n_933),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_761),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_757),
.A2(n_377),
.B1(n_393),
.B2(n_339),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_841),
.B(n_933),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_729),
.Y(n_1521)
);

CKINVDCx8_ASAP7_75t_R g1522 ( 
.A(n_797),
.Y(n_1522)
);

NOR2xp67_ASAP7_75t_L g1523 ( 
.A(n_797),
.B(n_401),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_839),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1089),
.B(n_312),
.Y(n_1525)
);

INVx3_ASAP7_75t_L g1526 ( 
.A(n_821),
.Y(n_1526)
);

AOI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1008),
.A2(n_1023),
.B(n_476),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_839),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_839),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_841),
.B(n_933),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_729),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_841),
.B(n_933),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_841),
.B(n_933),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_859),
.A2(n_597),
.B1(n_663),
.B2(n_676),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_841),
.B(n_933),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_SL g1536 ( 
.A(n_794),
.B(n_912),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_729),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1089),
.B(n_312),
.Y(n_1538)
);

NAND3xp33_ASAP7_75t_L g1539 ( 
.A(n_757),
.B(n_841),
.C(n_558),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_841),
.B(n_933),
.Y(n_1540)
);

AOI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_757),
.A2(n_377),
.B1(n_393),
.B2(n_339),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_729),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_737),
.B(n_921),
.Y(n_1543)
);

NOR3xp33_ASAP7_75t_L g1544 ( 
.A(n_867),
.B(n_757),
.C(n_841),
.Y(n_1544)
);

AOI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_757),
.A2(n_377),
.B1(n_393),
.B2(n_339),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_SL g1546 ( 
.A(n_794),
.B(n_912),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_729),
.Y(n_1547)
);

INVx3_ASAP7_75t_L g1548 ( 
.A(n_821),
.Y(n_1548)
);

INVxp67_ASAP7_75t_L g1549 ( 
.A(n_749),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1089),
.B(n_312),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_841),
.B(n_933),
.Y(n_1551)
);

O2A1O1Ixp33_ASAP7_75t_L g1552 ( 
.A1(n_757),
.A2(n_867),
.B(n_841),
.C(n_558),
.Y(n_1552)
);

NOR2xp33_ASAP7_75t_L g1553 ( 
.A(n_841),
.B(n_461),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_776),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_839),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_761),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_729),
.Y(n_1557)
);

INVxp33_ASAP7_75t_L g1558 ( 
.A(n_826),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_841),
.B(n_933),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_729),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_839),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_SL g1562 ( 
.A(n_794),
.B(n_912),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_729),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_841),
.B(n_933),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_839),
.Y(n_1565)
);

O2A1O1Ixp5_ASAP7_75t_L g1566 ( 
.A1(n_778),
.A2(n_757),
.B(n_892),
.C(n_939),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_841),
.B(n_933),
.Y(n_1567)
);

AND2x6_ASAP7_75t_L g1568 ( 
.A(n_794),
.B(n_699),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_841),
.B(n_933),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_841),
.B(n_933),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_841),
.B(n_933),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_841),
.B(n_461),
.Y(n_1572)
);

NAND2xp33_ASAP7_75t_L g1573 ( 
.A(n_760),
.B(n_788),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_729),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_SL g1575 ( 
.A(n_794),
.B(n_912),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_839),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_839),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_761),
.B(n_606),
.Y(n_1578)
);

INVx6_ASAP7_75t_L g1579 ( 
.A(n_849),
.Y(n_1579)
);

INVx2_ASAP7_75t_SL g1580 ( 
.A(n_739),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_SL g1581 ( 
.A(n_794),
.B(n_912),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_839),
.Y(n_1582)
);

INVxp67_ASAP7_75t_L g1583 ( 
.A(n_749),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_776),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_841),
.B(n_461),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_794),
.B(n_912),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_841),
.B(n_933),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_841),
.B(n_461),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_841),
.B(n_933),
.Y(n_1589)
);

INVxp67_ASAP7_75t_SL g1590 ( 
.A(n_989),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_841),
.B(n_933),
.Y(n_1591)
);

NOR3xp33_ASAP7_75t_L g1592 ( 
.A(n_867),
.B(n_757),
.C(n_841),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_841),
.B(n_933),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_841),
.B(n_933),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_839),
.Y(n_1595)
);

BUFx5_ASAP7_75t_L g1596 ( 
.A(n_848),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_729),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_737),
.B(n_921),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_729),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_841),
.B(n_933),
.Y(n_1600)
);

NAND2x1p5_ASAP7_75t_L g1601 ( 
.A(n_737),
.B(n_770),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_839),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_729),
.Y(n_1603)
);

AO21x2_ASAP7_75t_L g1604 ( 
.A1(n_897),
.A2(n_610),
.B(n_523),
.Y(n_1604)
);

OAI221xp5_ASAP7_75t_L g1605 ( 
.A1(n_841),
.A2(n_498),
.B1(n_525),
.B2(n_757),
.C(n_825),
.Y(n_1605)
);

OAI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1008),
.A2(n_939),
.B(n_903),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_841),
.B(n_933),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_841),
.B(n_933),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_729),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_841),
.B(n_933),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_SL g1611 ( 
.A(n_794),
.B(n_912),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_729),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_839),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_841),
.B(n_933),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1568),
.A2(n_1437),
.B1(n_1439),
.B2(n_1101),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1402),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1129),
.B(n_1606),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1108),
.B(n_1107),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1107),
.A2(n_1453),
.B1(n_1539),
.B2(n_1097),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_SL g1620 ( 
.A(n_1094),
.B(n_1393),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1291),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1295),
.Y(n_1622)
);

BUFx6f_ASAP7_75t_L g1623 ( 
.A(n_1390),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1296),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1394),
.B(n_1543),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_SL g1626 ( 
.A(n_1397),
.B(n_1400),
.Y(n_1626)
);

BUFx4f_ASAP7_75t_L g1627 ( 
.A(n_1568),
.Y(n_1627)
);

OAI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1131),
.A2(n_1127),
.B1(n_1605),
.B2(n_1398),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1568),
.B(n_1163),
.Y(n_1629)
);

AOI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1568),
.A2(n_1101),
.B1(n_1132),
.B2(n_1115),
.Y(n_1630)
);

BUFx6f_ASAP7_75t_L g1631 ( 
.A(n_1390),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1200),
.Y(n_1632)
);

INVx3_ASAP7_75t_L g1633 ( 
.A(n_1390),
.Y(n_1633)
);

INVx1_ASAP7_75t_SL g1634 ( 
.A(n_1578),
.Y(n_1634)
);

INVx5_ASAP7_75t_L g1635 ( 
.A(n_1390),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_L g1636 ( 
.A(n_1411),
.B(n_1416),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1301),
.Y(n_1637)
);

NAND2x1p5_ASAP7_75t_L g1638 ( 
.A(n_1384),
.B(n_1112),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_L g1639 ( 
.A(n_1421),
.B(n_1424),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1568),
.B(n_1127),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_R g1641 ( 
.A(n_1522),
.B(n_1506),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1200),
.Y(n_1642)
);

INVxp67_ASAP7_75t_L g1643 ( 
.A(n_1452),
.Y(n_1643)
);

AND2x6_ASAP7_75t_SL g1644 ( 
.A(n_1458),
.B(n_1504),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1389),
.Y(n_1645)
);

AOI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1568),
.A2(n_1398),
.B1(n_1403),
.B2(n_1098),
.Y(n_1646)
);

INVx3_ASAP7_75t_L g1647 ( 
.A(n_1390),
.Y(n_1647)
);

NAND3xp33_ASAP7_75t_SL g1648 ( 
.A(n_1492),
.B(n_1552),
.C(n_1461),
.Y(n_1648)
);

AOI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1098),
.A2(n_1419),
.B1(n_1425),
.B2(n_1403),
.Y(n_1649)
);

O2A1O1Ixp5_ASAP7_75t_SL g1650 ( 
.A1(n_1106),
.A2(n_1419),
.B(n_1428),
.C(n_1425),
.Y(n_1650)
);

BUFx2_ASAP7_75t_L g1651 ( 
.A(n_1590),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1306),
.Y(n_1652)
);

INVx1_ASAP7_75t_SL g1653 ( 
.A(n_1518),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_SL g1654 ( 
.A(n_1401),
.B(n_1406),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1126),
.B(n_1169),
.Y(n_1655)
);

BUFx2_ASAP7_75t_L g1656 ( 
.A(n_1320),
.Y(n_1656)
);

AOI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1428),
.A2(n_1435),
.B1(n_1440),
.B2(n_1438),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1415),
.B(n_1418),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1308),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1432),
.B(n_1434),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1310),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1446),
.B(n_1454),
.Y(n_1662)
);

NAND2xp33_ASAP7_75t_SL g1663 ( 
.A(n_1095),
.B(n_1436),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1300),
.B(n_1417),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_SL g1665 ( 
.A(n_1462),
.B(n_1468),
.Y(n_1665)
);

INVx3_ASAP7_75t_L g1666 ( 
.A(n_1390),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1192),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1195),
.Y(n_1668)
);

OR2x6_ASAP7_75t_L g1669 ( 
.A(n_1208),
.B(n_1216),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1181),
.B(n_1186),
.Y(n_1670)
);

INVx3_ASAP7_75t_L g1671 ( 
.A(n_1362),
.Y(n_1671)
);

NAND2x1p5_ASAP7_75t_L g1672 ( 
.A(n_1384),
.B(n_1112),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1183),
.A2(n_1191),
.B(n_1566),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1203),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1209),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1417),
.B(n_1414),
.Y(n_1676)
);

NAND2x1p5_ASAP7_75t_L g1677 ( 
.A(n_1324),
.B(n_1355),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1217),
.Y(n_1678)
);

AND3x2_ASAP7_75t_SL g1679 ( 
.A(n_1435),
.B(n_1440),
.C(n_1438),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1553),
.B(n_1572),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1585),
.B(n_1588),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1111),
.B(n_1106),
.Y(n_1682)
);

INVx3_ASAP7_75t_L g1683 ( 
.A(n_1362),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1096),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1190),
.B(n_1122),
.Y(n_1685)
);

BUFx6f_ASAP7_75t_L g1686 ( 
.A(n_1362),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1476),
.B(n_1478),
.Y(n_1687)
);

AND2x4_ASAP7_75t_L g1688 ( 
.A(n_1394),
.B(n_1543),
.Y(n_1688)
);

OAI22xp5_ASAP7_75t_SL g1689 ( 
.A1(n_1100),
.A2(n_1447),
.B1(n_1534),
.B2(n_1471),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1096),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1135),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1135),
.Y(n_1692)
);

BUFx6f_ASAP7_75t_L g1693 ( 
.A(n_1362),
.Y(n_1693)
);

AND2x2_ASAP7_75t_SL g1694 ( 
.A(n_1232),
.B(n_1433),
.Y(n_1694)
);

XNOR2xp5_ASAP7_75t_L g1695 ( 
.A(n_1413),
.B(n_1451),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_SL g1696 ( 
.A1(n_1417),
.A2(n_1140),
.B1(n_1392),
.B2(n_1157),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1288),
.B(n_1111),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1472),
.B(n_1477),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1230),
.B(n_1131),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1120),
.B(n_1407),
.Y(n_1700)
);

AOI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1183),
.A2(n_1191),
.B(n_1444),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_SL g1702 ( 
.A(n_1480),
.B(n_1484),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1142),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1544),
.B(n_1592),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1444),
.A2(n_1449),
.B1(n_1460),
.B2(n_1448),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1142),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1503),
.B(n_1525),
.Y(n_1707)
);

INVx3_ASAP7_75t_L g1708 ( 
.A(n_1365),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_1556),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1394),
.B(n_1543),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1143),
.Y(n_1711)
);

BUFx4f_ASAP7_75t_L g1712 ( 
.A(n_1208),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1304),
.B(n_1315),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1316),
.B(n_1317),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1321),
.B(n_1322),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1323),
.B(n_1327),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1143),
.Y(n_1717)
);

BUFx4f_ASAP7_75t_L g1718 ( 
.A(n_1208),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1160),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1160),
.Y(n_1720)
);

INVx3_ASAP7_75t_L g1721 ( 
.A(n_1365),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1171),
.Y(n_1722)
);

OR2x6_ASAP7_75t_L g1723 ( 
.A(n_1208),
.B(n_1216),
.Y(n_1723)
);

INVxp67_ASAP7_75t_SL g1724 ( 
.A(n_1239),
.Y(n_1724)
);

AOI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1448),
.A2(n_1449),
.B1(n_1464),
.B2(n_1460),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1171),
.Y(n_1726)
);

NOR2x2_ASAP7_75t_L g1727 ( 
.A(n_1093),
.B(n_1153),
.Y(n_1727)
);

BUFx3_ASAP7_75t_L g1728 ( 
.A(n_1200),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1173),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1328),
.B(n_1335),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1176),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1339),
.B(n_1341),
.Y(n_1732)
);

INVx3_ASAP7_75t_L g1733 ( 
.A(n_1365),
.Y(n_1733)
);

AND2x2_ASAP7_75t_SL g1734 ( 
.A(n_1232),
.B(n_1433),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1598),
.B(n_1299),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_SL g1736 ( 
.A(n_1485),
.B(n_1490),
.Y(n_1736)
);

OR2x2_ASAP7_75t_SL g1737 ( 
.A(n_1495),
.B(n_1391),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1598),
.B(n_1288),
.Y(n_1738)
);

NOR3xp33_ASAP7_75t_SL g1739 ( 
.A(n_1128),
.B(n_1584),
.C(n_1554),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1598),
.B(n_1493),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_SL g1741 ( 
.A(n_1501),
.B(n_1507),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1614),
.B(n_1510),
.Y(n_1742)
);

OR2x6_ASAP7_75t_SL g1743 ( 
.A(n_1194),
.B(n_1513),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1288),
.B(n_1271),
.Y(n_1744)
);

BUFx8_ASAP7_75t_L g1745 ( 
.A(n_1292),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1515),
.B(n_1517),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1182),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1158),
.Y(n_1748)
);

INVx2_ASAP7_75t_SL g1749 ( 
.A(n_1200),
.Y(n_1749)
);

BUFx2_ASAP7_75t_L g1750 ( 
.A(n_1146),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1520),
.B(n_1530),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_SL g1752 ( 
.A(n_1532),
.B(n_1533),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1185),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1538),
.B(n_1550),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1535),
.B(n_1540),
.Y(n_1755)
);

INVxp67_ASAP7_75t_L g1756 ( 
.A(n_1114),
.Y(n_1756)
);

OAI22xp5_ASAP7_75t_SL g1757 ( 
.A1(n_1399),
.A2(n_1519),
.B1(n_1545),
.B2(n_1541),
.Y(n_1757)
);

CKINVDCx11_ASAP7_75t_R g1758 ( 
.A(n_1105),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1271),
.B(n_1125),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_SL g1760 ( 
.A(n_1551),
.B(n_1559),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1133),
.A2(n_1464),
.B1(n_1473),
.B2(n_1470),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_SL g1762 ( 
.A(n_1564),
.B(n_1567),
.Y(n_1762)
);

O2A1O1Ixp33_ASAP7_75t_L g1763 ( 
.A1(n_1470),
.A2(n_1473),
.B(n_1482),
.C(n_1475),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1569),
.B(n_1570),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1207),
.Y(n_1765)
);

NAND2xp33_ASAP7_75t_SL g1766 ( 
.A(n_1436),
.B(n_1469),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1571),
.B(n_1587),
.Y(n_1767)
);

AND2x4_ASAP7_75t_L g1768 ( 
.A(n_1271),
.B(n_1093),
.Y(n_1768)
);

INVx2_ASAP7_75t_SL g1769 ( 
.A(n_1502),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1207),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1212),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1212),
.Y(n_1772)
);

INVx4_ASAP7_75t_L g1773 ( 
.A(n_1216),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1218),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1589),
.B(n_1591),
.Y(n_1775)
);

AOI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1475),
.A2(n_1511),
.B(n_1482),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_SL g1777 ( 
.A(n_1593),
.B(n_1594),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1220),
.Y(n_1778)
);

INVx2_ASAP7_75t_SL g1779 ( 
.A(n_1502),
.Y(n_1779)
);

BUFx3_ASAP7_75t_L g1780 ( 
.A(n_1227),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1225),
.Y(n_1781)
);

NOR3xp33_ASAP7_75t_L g1782 ( 
.A(n_1113),
.B(n_1514),
.C(n_1511),
.Y(n_1782)
);

BUFx6f_ASAP7_75t_L g1783 ( 
.A(n_1365),
.Y(n_1783)
);

NOR2xp33_ASAP7_75t_L g1784 ( 
.A(n_1469),
.B(n_1558),
.Y(n_1784)
);

BUFx2_ASAP7_75t_L g1785 ( 
.A(n_1146),
.Y(n_1785)
);

CKINVDCx20_ASAP7_75t_R g1786 ( 
.A(n_1128),
.Y(n_1786)
);

OR2x6_ASAP7_75t_L g1787 ( 
.A(n_1333),
.B(n_1514),
.Y(n_1787)
);

NOR2x1_ASAP7_75t_L g1788 ( 
.A(n_1509),
.B(n_1573),
.Y(n_1788)
);

INVx2_ASAP7_75t_SL g1789 ( 
.A(n_1579),
.Y(n_1789)
);

BUFx3_ASAP7_75t_L g1790 ( 
.A(n_1227),
.Y(n_1790)
);

OR2x2_ASAP7_75t_SL g1791 ( 
.A(n_1600),
.B(n_1607),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1229),
.Y(n_1792)
);

BUFx2_ASAP7_75t_L g1793 ( 
.A(n_1146),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_1292),
.Y(n_1794)
);

AND2x6_ASAP7_75t_SL g1795 ( 
.A(n_1201),
.B(n_1168),
.Y(n_1795)
);

OR2x6_ASAP7_75t_L g1796 ( 
.A(n_1333),
.B(n_1536),
.Y(n_1796)
);

AOI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1536),
.A2(n_1562),
.B1(n_1575),
.B2(n_1546),
.Y(n_1797)
);

AND2x4_ASAP7_75t_L g1798 ( 
.A(n_1093),
.B(n_1227),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1229),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1608),
.B(n_1610),
.Y(n_1800)
);

INVx3_ASAP7_75t_L g1801 ( 
.A(n_1138),
.Y(n_1801)
);

NOR2x1_ASAP7_75t_L g1802 ( 
.A(n_1509),
.B(n_1573),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1148),
.B(n_1154),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1152),
.B(n_1546),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1258),
.Y(n_1805)
);

NOR2xp33_ASAP7_75t_SL g1806 ( 
.A(n_1116),
.B(n_1500),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_SL g1807 ( 
.A(n_1558),
.B(n_1104),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1258),
.Y(n_1808)
);

AOI22xp33_ASAP7_75t_L g1809 ( 
.A1(n_1562),
.A2(n_1575),
.B1(n_1586),
.B2(n_1581),
.Y(n_1809)
);

INVx2_ASAP7_75t_SL g1810 ( 
.A(n_1579),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1264),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1264),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1266),
.Y(n_1813)
);

CKINVDCx6p67_ASAP7_75t_R g1814 ( 
.A(n_1139),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1266),
.Y(n_1815)
);

HB1xp67_ASAP7_75t_L g1816 ( 
.A(n_1248),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1275),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1326),
.B(n_1193),
.Y(n_1818)
);

AOI22xp33_ASAP7_75t_L g1819 ( 
.A1(n_1581),
.A2(n_1586),
.B1(n_1611),
.B2(n_1156),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1275),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1277),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1611),
.B(n_1351),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1277),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1286),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1286),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1305),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1305),
.Y(n_1827)
);

INVx3_ASAP7_75t_L g1828 ( 
.A(n_1138),
.Y(n_1828)
);

BUFx6f_ASAP7_75t_L g1829 ( 
.A(n_1138),
.Y(n_1829)
);

INVx3_ASAP7_75t_L g1830 ( 
.A(n_1426),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1307),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_SL g1832 ( 
.A(n_1527),
.B(n_1250),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1340),
.B(n_1284),
.Y(n_1833)
);

O2A1O1Ixp33_ASAP7_75t_L g1834 ( 
.A1(n_1151),
.A2(n_1214),
.B(n_1343),
.C(n_1312),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1307),
.Y(n_1835)
);

OR2x6_ASAP7_75t_SL g1836 ( 
.A(n_1123),
.B(n_1118),
.Y(n_1836)
);

INVx2_ASAP7_75t_SL g1837 ( 
.A(n_1579),
.Y(n_1837)
);

INVxp33_ASAP7_75t_SL g1838 ( 
.A(n_1245),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_1312),
.B(n_1343),
.Y(n_1839)
);

AOI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1235),
.A2(n_1161),
.B1(n_1172),
.B2(n_1121),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1240),
.B(n_1241),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1184),
.A2(n_1177),
.B1(n_1226),
.B2(n_1329),
.Y(n_1842)
);

INVx1_ASAP7_75t_SL g1843 ( 
.A(n_1285),
.Y(n_1843)
);

AOI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1161),
.A2(n_1145),
.B1(n_1137),
.B2(n_1116),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1331),
.B(n_1149),
.Y(n_1845)
);

BUFx4f_ASAP7_75t_L g1846 ( 
.A(n_1426),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1244),
.B(n_1257),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1103),
.B(n_1283),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_L g1849 ( 
.A(n_1103),
.B(n_1283),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1395),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_1396),
.Y(n_1851)
);

OAI22xp33_ASAP7_75t_L g1852 ( 
.A1(n_1523),
.A2(n_1222),
.B1(n_1269),
.B2(n_1441),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1155),
.B(n_1170),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1293),
.B(n_1289),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1332),
.Y(n_1855)
);

AND2x4_ASAP7_75t_L g1856 ( 
.A(n_1093),
.B(n_1247),
.Y(n_1856)
);

AOI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1342),
.A2(n_1346),
.B1(n_1167),
.B2(n_1236),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_R g1858 ( 
.A(n_1139),
.B(n_1427),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1174),
.B(n_1188),
.Y(n_1859)
);

BUFx6f_ASAP7_75t_L g1860 ( 
.A(n_1426),
.Y(n_1860)
);

CKINVDCx5p33_ASAP7_75t_R g1861 ( 
.A(n_1396),
.Y(n_1861)
);

BUFx6f_ASAP7_75t_L g1862 ( 
.A(n_1426),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1332),
.Y(n_1863)
);

OR2x6_ASAP7_75t_L g1864 ( 
.A(n_1333),
.B(n_1379),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1337),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1337),
.Y(n_1866)
);

INVx4_ASAP7_75t_L g1867 ( 
.A(n_1436),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1198),
.B(n_1204),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1349),
.Y(n_1869)
);

AOI22xp33_ASAP7_75t_L g1870 ( 
.A1(n_1167),
.A2(n_1228),
.B1(n_1422),
.B2(n_1349),
.Y(n_1870)
);

BUFx3_ASAP7_75t_L g1871 ( 
.A(n_1116),
.Y(n_1871)
);

INVxp67_ASAP7_75t_L g1872 ( 
.A(n_1467),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1297),
.B(n_1298),
.Y(n_1873)
);

AND2x4_ASAP7_75t_L g1874 ( 
.A(n_1330),
.B(n_1319),
.Y(n_1874)
);

INVx3_ASAP7_75t_L g1875 ( 
.A(n_1330),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1219),
.B(n_1224),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1422),
.Y(n_1877)
);

BUFx6f_ASAP7_75t_L g1878 ( 
.A(n_1374),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1237),
.B(n_1238),
.Y(n_1879)
);

BUFx12f_ASAP7_75t_L g1880 ( 
.A(n_1508),
.Y(n_1880)
);

INVx4_ASAP7_75t_L g1881 ( 
.A(n_1330),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1325),
.B(n_1099),
.Y(n_1882)
);

BUFx2_ASAP7_75t_L g1883 ( 
.A(n_1274),
.Y(n_1883)
);

AOI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1313),
.A2(n_1243),
.B1(n_1242),
.B2(n_1303),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_L g1885 ( 
.A(n_1474),
.B(n_1486),
.Y(n_1885)
);

INVx2_ASAP7_75t_SL g1886 ( 
.A(n_1427),
.Y(n_1886)
);

AND2x4_ASAP7_75t_L g1887 ( 
.A(n_1319),
.B(n_1092),
.Y(n_1887)
);

NOR3xp33_ASAP7_75t_SL g1888 ( 
.A(n_1309),
.B(n_1382),
.C(n_1368),
.Y(n_1888)
);

NOR2xp33_ASAP7_75t_R g1889 ( 
.A(n_1497),
.B(n_1165),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1442),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1102),
.B(n_1613),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1265),
.B(n_1287),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_SL g1893 ( 
.A(n_1265),
.B(n_1287),
.Y(n_1893)
);

BUFx12f_ASAP7_75t_L g1894 ( 
.A(n_1408),
.Y(n_1894)
);

AOI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1303),
.A2(n_1357),
.B(n_1205),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1109),
.B(n_1110),
.Y(n_1896)
);

AND2x6_ASAP7_75t_SL g1897 ( 
.A(n_1294),
.B(n_1223),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_SL g1898 ( 
.A(n_1265),
.B(n_1287),
.Y(n_1898)
);

AOI21xp33_ASAP7_75t_L g1899 ( 
.A1(n_1357),
.A2(n_1361),
.B(n_1377),
.Y(n_1899)
);

INVx5_ASAP7_75t_L g1900 ( 
.A(n_1374),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1117),
.B(n_1124),
.Y(n_1901)
);

OR2x2_ASAP7_75t_SL g1902 ( 
.A(n_1263),
.B(n_1273),
.Y(n_1902)
);

BUFx2_ASAP7_75t_L g1903 ( 
.A(n_1197),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1136),
.B(n_1147),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1443),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1443),
.Y(n_1906)
);

HB1xp67_ASAP7_75t_L g1907 ( 
.A(n_1487),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1210),
.B(n_1405),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_1431),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1456),
.Y(n_1910)
);

AOI22xp33_ASAP7_75t_L g1911 ( 
.A1(n_1465),
.A2(n_1612),
.B1(n_1488),
.B2(n_1547),
.Y(n_1911)
);

AOI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1162),
.A2(n_1431),
.B1(n_1457),
.B2(n_1498),
.Y(n_1912)
);

INVx2_ASAP7_75t_SL g1913 ( 
.A(n_1497),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_SL g1914 ( 
.A(n_1265),
.B(n_1287),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1164),
.B(n_1549),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1465),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1466),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1466),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1479),
.Y(n_1919)
);

BUFx3_ASAP7_75t_L g1920 ( 
.A(n_1601),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_SL g1921 ( 
.A(n_1366),
.B(n_1336),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1479),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1481),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1481),
.Y(n_1924)
);

NOR2xp33_ASAP7_75t_L g1925 ( 
.A(n_1583),
.B(n_1187),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1488),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1409),
.B(n_1412),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1420),
.B(n_1423),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1491),
.Y(n_1929)
);

INVx2_ASAP7_75t_SL g1930 ( 
.A(n_1353),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1092),
.B(n_1134),
.Y(n_1931)
);

AOI21xp5_ASAP7_75t_L g1932 ( 
.A1(n_1338),
.A2(n_1252),
.B(n_1206),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_SL g1933 ( 
.A(n_1336),
.B(n_1348),
.Y(n_1933)
);

AOI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1491),
.A2(n_1612),
.B1(n_1609),
.B2(n_1494),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1494),
.Y(n_1935)
);

INVx4_ASAP7_75t_L g1936 ( 
.A(n_1601),
.Y(n_1936)
);

OR2x2_ASAP7_75t_SL g1937 ( 
.A(n_1280),
.B(n_1282),
.Y(n_1937)
);

AND2x2_ASAP7_75t_SL g1938 ( 
.A(n_1388),
.B(n_1234),
.Y(n_1938)
);

OAI22xp5_ASAP7_75t_L g1939 ( 
.A1(n_1430),
.A2(n_1450),
.B1(n_1602),
.B2(n_1595),
.Y(n_1939)
);

AOI22xp33_ASAP7_75t_L g1940 ( 
.A1(n_1516),
.A2(n_1609),
.B1(n_1603),
.B2(n_1599),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1516),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1521),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1521),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1445),
.B(n_1459),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1463),
.B(n_1483),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_1457),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1531),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_1270),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1496),
.B(n_1499),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1531),
.Y(n_1950)
);

BUFx6f_ASAP7_75t_L g1951 ( 
.A(n_1374),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1512),
.B(n_1524),
.Y(n_1952)
);

NOR2x2_ASAP7_75t_L g1953 ( 
.A(n_1371),
.B(n_1372),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1528),
.B(n_1529),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1555),
.B(n_1561),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1537),
.Y(n_1956)
);

AND2x4_ASAP7_75t_SL g1957 ( 
.A(n_1092),
.B(n_1134),
.Y(n_1957)
);

INVx2_ASAP7_75t_SL g1958 ( 
.A(n_1336),
.Y(n_1958)
);

A2O1A1Ixp33_ASAP7_75t_L g1959 ( 
.A1(n_1338),
.A2(n_1356),
.B(n_1249),
.C(n_1267),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1537),
.Y(n_1960)
);

AND2x4_ASAP7_75t_L g1961 ( 
.A(n_1134),
.B(n_1268),
.Y(n_1961)
);

INVx3_ASAP7_75t_L g1962 ( 
.A(n_1359),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1565),
.B(n_1576),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1542),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1542),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1547),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1557),
.Y(n_1967)
);

BUFx3_ASAP7_75t_L g1968 ( 
.A(n_1376),
.Y(n_1968)
);

BUFx3_ASAP7_75t_L g1969 ( 
.A(n_1376),
.Y(n_1969)
);

BUFx6f_ASAP7_75t_L g1970 ( 
.A(n_1374),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1557),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1577),
.B(n_1582),
.Y(n_1972)
);

BUFx6f_ASAP7_75t_L g1973 ( 
.A(n_1336),
.Y(n_1973)
);

NOR2xp33_ASAP7_75t_L g1974 ( 
.A(n_1429),
.B(n_1455),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1560),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1560),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1246),
.B(n_1254),
.Y(n_1977)
);

BUFx2_ASAP7_75t_L g1978 ( 
.A(n_1380),
.Y(n_1978)
);

INVxp67_ASAP7_75t_SL g1979 ( 
.A(n_1215),
.Y(n_1979)
);

INVx3_ASAP7_75t_L g1980 ( 
.A(n_1359),
.Y(n_1980)
);

CKINVDCx5p33_ASAP7_75t_R g1981 ( 
.A(n_1489),
.Y(n_1981)
);

CKINVDCx20_ASAP7_75t_R g1982 ( 
.A(n_1580),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1259),
.B(n_1262),
.Y(n_1983)
);

BUFx6f_ASAP7_75t_L g1984 ( 
.A(n_1348),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1563),
.Y(n_1985)
);

OR2x6_ASAP7_75t_SL g1986 ( 
.A(n_1360),
.B(n_1364),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_SL g1987 ( 
.A(n_1348),
.B(n_1202),
.Y(n_1987)
);

BUFx2_ASAP7_75t_L g1988 ( 
.A(n_1380),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1563),
.Y(n_1989)
);

AOI21xp5_ASAP7_75t_L g1990 ( 
.A1(n_1119),
.A2(n_1130),
.B(n_1141),
.Y(n_1990)
);

HB1xp67_ASAP7_75t_L g1991 ( 
.A(n_1175),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1278),
.B(n_1281),
.Y(n_1992)
);

NAND2xp33_ASAP7_75t_SL g1993 ( 
.A(n_1166),
.B(n_1378),
.Y(n_1993)
);

AND2x4_ASAP7_75t_L g1994 ( 
.A(n_1268),
.B(n_1404),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1574),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1371),
.B(n_1386),
.Y(n_1996)
);

A2O1A1Ixp33_ASAP7_75t_L g1997 ( 
.A1(n_1345),
.A2(n_1387),
.B(n_1276),
.C(n_1253),
.Y(n_1997)
);

OAI22xp33_ASAP7_75t_L g1998 ( 
.A1(n_1302),
.A2(n_1369),
.B1(n_1347),
.B2(n_1354),
.Y(n_1998)
);

NOR2xp33_ASAP7_75t_L g1999 ( 
.A(n_1385),
.B(n_1372),
.Y(n_1999)
);

AOI22xp33_ASAP7_75t_SL g2000 ( 
.A1(n_1359),
.A2(n_1596),
.B1(n_1334),
.B2(n_1599),
.Y(n_2000)
);

AOI22xp33_ASAP7_75t_L g2001 ( 
.A1(n_1574),
.A2(n_1603),
.B1(n_1597),
.B2(n_1383),
.Y(n_2001)
);

BUFx6f_ASAP7_75t_L g2002 ( 
.A(n_1348),
.Y(n_2002)
);

INVx3_ASAP7_75t_L g2003 ( 
.A(n_1359),
.Y(n_2003)
);

BUFx3_ASAP7_75t_L g2004 ( 
.A(n_1375),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_1375),
.Y(n_2005)
);

AND2x4_ASAP7_75t_L g2006 ( 
.A(n_1268),
.B(n_1526),
.Y(n_2006)
);

INVx1_ASAP7_75t_SL g2007 ( 
.A(n_1381),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_SL g2008 ( 
.A(n_1318),
.B(n_1410),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1597),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1381),
.B(n_1383),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1604),
.Y(n_2011)
);

BUFx3_ASAP7_75t_L g2012 ( 
.A(n_1375),
.Y(n_2012)
);

AND3x1_ASAP7_75t_L g2013 ( 
.A(n_1404),
.B(n_1410),
.C(n_1548),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1604),
.Y(n_2014)
);

NOR2xp33_ASAP7_75t_L g2015 ( 
.A(n_1358),
.B(n_1260),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1404),
.B(n_1548),
.Y(n_2016)
);

BUFx4f_ASAP7_75t_L g2017 ( 
.A(n_1363),
.Y(n_2017)
);

NOR2xp33_ASAP7_75t_L g2018 ( 
.A(n_1199),
.B(n_1260),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1410),
.B(n_1505),
.Y(n_2019)
);

OAI21xp5_ASAP7_75t_L g2020 ( 
.A1(n_1373),
.A2(n_1350),
.B(n_1130),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1596),
.Y(n_2021)
);

AOI22xp5_ASAP7_75t_L g2022 ( 
.A1(n_1359),
.A2(n_1596),
.B1(n_1159),
.B2(n_1150),
.Y(n_2022)
);

CKINVDCx8_ASAP7_75t_R g2023 ( 
.A(n_1179),
.Y(n_2023)
);

OAI22xp5_ASAP7_75t_L g2024 ( 
.A1(n_1505),
.A2(n_1526),
.B1(n_1548),
.B2(n_1363),
.Y(n_2024)
);

HB1xp67_ASAP7_75t_L g2025 ( 
.A(n_1199),
.Y(n_2025)
);

INVx3_ASAP7_75t_L g2026 ( 
.A(n_1359),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1596),
.Y(n_2027)
);

BUFx6f_ASAP7_75t_L g2028 ( 
.A(n_1119),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1596),
.B(n_1150),
.Y(n_2029)
);

AOI22xp33_ASAP7_75t_L g2030 ( 
.A1(n_1596),
.A2(n_1141),
.B1(n_1144),
.B2(n_1251),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1596),
.B(n_1159),
.Y(n_2031)
);

BUFx2_ASAP7_75t_L g2032 ( 
.A(n_1211),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_SL g2033 ( 
.A(n_1179),
.B(n_1196),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1178),
.B(n_1196),
.Y(n_2034)
);

HB1xp67_ASAP7_75t_L g2035 ( 
.A(n_1211),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1370),
.Y(n_2036)
);

OAI22xp5_ASAP7_75t_SL g2037 ( 
.A1(n_1213),
.A2(n_1261),
.B1(n_1367),
.B2(n_1352),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1370),
.Y(n_2038)
);

HB1xp67_ASAP7_75t_L g2039 ( 
.A(n_1213),
.Y(n_2039)
);

AND2x4_ASAP7_75t_L g2040 ( 
.A(n_1178),
.B(n_1180),
.Y(n_2040)
);

AND2x4_ASAP7_75t_L g2041 ( 
.A(n_1180),
.B(n_1189),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1367),
.Y(n_2042)
);

INVx3_ASAP7_75t_L g2043 ( 
.A(n_1144),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_SL g2044 ( 
.A(n_1189),
.B(n_1221),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1221),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1352),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_SL g2047 ( 
.A(n_1231),
.B(n_1233),
.Y(n_2047)
);

BUFx3_ASAP7_75t_L g2048 ( 
.A(n_1231),
.Y(n_2048)
);

AOI22xp33_ASAP7_75t_L g2049 ( 
.A1(n_1233),
.A2(n_1251),
.B1(n_1255),
.B2(n_1256),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1344),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1255),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1256),
.Y(n_2052)
);

BUFx6f_ASAP7_75t_L g2053 ( 
.A(n_1261),
.Y(n_2053)
);

OAI22xp5_ASAP7_75t_L g2054 ( 
.A1(n_1272),
.A2(n_1279),
.B1(n_1290),
.B2(n_1311),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1272),
.Y(n_2055)
);

OAI22xp5_ASAP7_75t_SL g2056 ( 
.A1(n_1279),
.A2(n_1290),
.B1(n_1311),
.B2(n_1314),
.Y(n_2056)
);

NOR2xp33_ASAP7_75t_L g2057 ( 
.A(n_1314),
.B(n_1344),
.Y(n_2057)
);

NAND2xp33_ASAP7_75t_L g2058 ( 
.A(n_1568),
.B(n_1107),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1291),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1291),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1291),
.Y(n_2061)
);

INVx5_ASAP7_75t_L g2062 ( 
.A(n_1390),
.Y(n_2062)
);

HB1xp67_ASAP7_75t_L g2063 ( 
.A(n_1402),
.Y(n_2063)
);

A2O1A1Ixp33_ASAP7_75t_L g2064 ( 
.A1(n_1107),
.A2(n_1552),
.B(n_1492),
.C(n_1437),
.Y(n_2064)
);

AOI22xp33_ASAP7_75t_L g2065 ( 
.A1(n_1568),
.A2(n_1447),
.B1(n_1534),
.B2(n_1414),
.Y(n_2065)
);

INVx1_ASAP7_75t_SL g2066 ( 
.A(n_1402),
.Y(n_2066)
);

HB1xp67_ASAP7_75t_L g2067 ( 
.A(n_1402),
.Y(n_2067)
);

BUFx2_ASAP7_75t_L g2068 ( 
.A(n_1568),
.Y(n_2068)
);

NAND2x1p5_ASAP7_75t_L g2069 ( 
.A(n_1384),
.B(n_1112),
.Y(n_2069)
);

BUFx4f_ASAP7_75t_L g2070 ( 
.A(n_1568),
.Y(n_2070)
);

NOR2xp33_ASAP7_75t_R g2071 ( 
.A(n_1522),
.B(n_344),
.Y(n_2071)
);

A2O1A1Ixp33_ASAP7_75t_L g2072 ( 
.A1(n_1107),
.A2(n_1552),
.B(n_1492),
.C(n_1437),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2073)
);

CKINVDCx5p33_ASAP7_75t_R g2074 ( 
.A(n_1128),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1291),
.Y(n_2075)
);

AOI22xp33_ASAP7_75t_SL g2076 ( 
.A1(n_1568),
.A2(n_264),
.B1(n_251),
.B2(n_1437),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2077)
);

AOI22xp33_ASAP7_75t_L g2078 ( 
.A1(n_1568),
.A2(n_1447),
.B1(n_1534),
.B2(n_1414),
.Y(n_2078)
);

XOR2x2_ASAP7_75t_L g2079 ( 
.A(n_1437),
.B(n_1439),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1389),
.Y(n_2081)
);

INVx8_ASAP7_75t_L g2082 ( 
.A(n_1568),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1291),
.Y(n_2083)
);

NOR2xp33_ASAP7_75t_L g2084 ( 
.A(n_1453),
.B(n_1539),
.Y(n_2084)
);

CKINVDCx20_ASAP7_75t_R g2085 ( 
.A(n_1128),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1291),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1291),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1291),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1291),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2090)
);

AOI21xp5_ASAP7_75t_L g2091 ( 
.A1(n_1107),
.A2(n_1183),
.B(n_1437),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_SL g2092 ( 
.A(n_1107),
.B(n_1437),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1291),
.Y(n_2093)
);

AOI22xp5_ASAP7_75t_L g2094 ( 
.A1(n_1568),
.A2(n_1437),
.B1(n_1439),
.B2(n_1101),
.Y(n_2094)
);

AND2x4_ASAP7_75t_L g2095 ( 
.A(n_1394),
.B(n_1543),
.Y(n_2095)
);

NOR2xp33_ASAP7_75t_L g2096 ( 
.A(n_1453),
.B(n_1539),
.Y(n_2096)
);

BUFx3_ASAP7_75t_L g2097 ( 
.A(n_1200),
.Y(n_2097)
);

INVx2_ASAP7_75t_SL g2098 ( 
.A(n_1200),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1291),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_SL g2100 ( 
.A(n_1107),
.B(n_1437),
.Y(n_2100)
);

AOI21xp5_ASAP7_75t_L g2101 ( 
.A1(n_1107),
.A2(n_1183),
.B(n_1437),
.Y(n_2101)
);

AOI22xp5_ASAP7_75t_L g2102 ( 
.A1(n_1568),
.A2(n_1437),
.B1(n_1439),
.B2(n_1101),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_1129),
.B(n_1300),
.Y(n_2105)
);

NOR2xp67_ASAP7_75t_L g2106 ( 
.A(n_1375),
.B(n_770),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2107)
);

HB1xp67_ASAP7_75t_L g2108 ( 
.A(n_1402),
.Y(n_2108)
);

AOI22xp33_ASAP7_75t_L g2109 ( 
.A1(n_1568),
.A2(n_1447),
.B1(n_1534),
.B2(n_1414),
.Y(n_2109)
);

AND2x4_ASAP7_75t_L g2110 ( 
.A(n_1394),
.B(n_1543),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1291),
.Y(n_2111)
);

NAND3xp33_ASAP7_75t_SL g2112 ( 
.A(n_1605),
.B(n_1552),
.C(n_1492),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1291),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1389),
.Y(n_2116)
);

NAND2xp33_ASAP7_75t_L g2117 ( 
.A(n_1568),
.B(n_1107),
.Y(n_2117)
);

BUFx12f_ASAP7_75t_L g2118 ( 
.A(n_1128),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_1129),
.B(n_1300),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2122)
);

AND2x4_ASAP7_75t_L g2123 ( 
.A(n_1394),
.B(n_1543),
.Y(n_2123)
);

AOI22xp5_ASAP7_75t_L g2124 ( 
.A1(n_1568),
.A2(n_1437),
.B1(n_1439),
.B2(n_1101),
.Y(n_2124)
);

AOI22xp5_ASAP7_75t_L g2125 ( 
.A1(n_1568),
.A2(n_1437),
.B1(n_1439),
.B2(n_1101),
.Y(n_2125)
);

BUFx12f_ASAP7_75t_L g2126 ( 
.A(n_1128),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_1129),
.B(n_1300),
.Y(n_2127)
);

CKINVDCx5p33_ASAP7_75t_R g2128 ( 
.A(n_1128),
.Y(n_2128)
);

BUFx6f_ASAP7_75t_SL g2129 ( 
.A(n_1568),
.Y(n_2129)
);

AOI22xp5_ASAP7_75t_L g2130 ( 
.A1(n_1568),
.A2(n_1437),
.B1(n_1439),
.B2(n_1101),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1389),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2132)
);

AOI22xp5_ASAP7_75t_L g2133 ( 
.A1(n_1568),
.A2(n_1437),
.B1(n_1439),
.B2(n_1101),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2134)
);

NAND2xp33_ASAP7_75t_SL g2135 ( 
.A(n_1437),
.B(n_1439),
.Y(n_2135)
);

BUFx6f_ASAP7_75t_L g2136 ( 
.A(n_1390),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_1389),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1291),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1291),
.Y(n_2139)
);

BUFx6f_ASAP7_75t_L g2140 ( 
.A(n_1390),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1291),
.Y(n_2141)
);

AOI22xp33_ASAP7_75t_L g2142 ( 
.A1(n_1568),
.A2(n_1447),
.B1(n_1534),
.B2(n_1414),
.Y(n_2142)
);

OAI21xp5_ASAP7_75t_L g2143 ( 
.A1(n_1107),
.A2(n_1439),
.B(n_1437),
.Y(n_2143)
);

INVx2_ASAP7_75t_SL g2144 ( 
.A(n_1200),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_1389),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1389),
.Y(n_2146)
);

OAI22xp5_ASAP7_75t_L g2147 ( 
.A1(n_1437),
.A2(n_1439),
.B1(n_1107),
.B2(n_1453),
.Y(n_2147)
);

NOR2xp67_ASAP7_75t_L g2148 ( 
.A(n_1375),
.B(n_770),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1291),
.Y(n_2151)
);

HB1xp67_ASAP7_75t_L g2152 ( 
.A(n_1402),
.Y(n_2152)
);

OAI21xp33_ASAP7_75t_L g2153 ( 
.A1(n_1107),
.A2(n_1539),
.B(n_1453),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1291),
.Y(n_2154)
);

AOI22xp5_ASAP7_75t_L g2155 ( 
.A1(n_1568),
.A2(n_1437),
.B1(n_1439),
.B2(n_1101),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1291),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1291),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_SL g2159 ( 
.A(n_1107),
.B(n_1437),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2161)
);

NOR2xp33_ASAP7_75t_L g2162 ( 
.A(n_1453),
.B(n_1539),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1291),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_1389),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_SL g2165 ( 
.A(n_1107),
.B(n_1437),
.Y(n_2165)
);

AND2x6_ASAP7_75t_L g2166 ( 
.A(n_1568),
.B(n_1324),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1291),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1291),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_1389),
.Y(n_2169)
);

INVx2_ASAP7_75t_SL g2170 ( 
.A(n_1200),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_1389),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1291),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_SL g2173 ( 
.A(n_1107),
.B(n_1437),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_1389),
.Y(n_2174)
);

BUFx6f_ASAP7_75t_SL g2175 ( 
.A(n_1568),
.Y(n_2175)
);

AOI22xp33_ASAP7_75t_L g2176 ( 
.A1(n_1568),
.A2(n_1447),
.B1(n_1534),
.B2(n_1414),
.Y(n_2176)
);

BUFx6f_ASAP7_75t_L g2177 ( 
.A(n_1390),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_SL g2178 ( 
.A(n_1107),
.B(n_1437),
.Y(n_2178)
);

BUFx3_ASAP7_75t_L g2179 ( 
.A(n_1200),
.Y(n_2179)
);

CKINVDCx11_ASAP7_75t_R g2180 ( 
.A(n_1522),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_SL g2181 ( 
.A(n_1107),
.B(n_1437),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_1129),
.B(n_1300),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2183)
);

AND2x4_ASAP7_75t_L g2184 ( 
.A(n_1394),
.B(n_1543),
.Y(n_2184)
);

OR2x6_ASAP7_75t_L g2185 ( 
.A(n_1208),
.B(n_1216),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2186)
);

BUFx6f_ASAP7_75t_L g2187 ( 
.A(n_1390),
.Y(n_2187)
);

INVx2_ASAP7_75t_SL g2188 ( 
.A(n_1200),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2189)
);

O2A1O1Ixp5_ASAP7_75t_L g2190 ( 
.A1(n_1107),
.A2(n_1439),
.B(n_1437),
.C(n_1566),
.Y(n_2190)
);

NOR2xp33_ASAP7_75t_L g2191 ( 
.A(n_1453),
.B(n_1539),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_SL g2192 ( 
.A(n_1107),
.B(n_1437),
.Y(n_2192)
);

NAND2xp33_ASAP7_75t_L g2193 ( 
.A(n_1568),
.B(n_1107),
.Y(n_2193)
);

INVx2_ASAP7_75t_SL g2194 ( 
.A(n_1200),
.Y(n_2194)
);

AOI22xp5_ASAP7_75t_L g2195 ( 
.A1(n_1568),
.A2(n_1437),
.B1(n_1439),
.B2(n_1101),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1291),
.Y(n_2196)
);

OR2x2_ASAP7_75t_SL g2197 ( 
.A(n_1453),
.B(n_1539),
.Y(n_2197)
);

NOR2xp33_ASAP7_75t_L g2198 ( 
.A(n_1453),
.B(n_1539),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_1389),
.Y(n_2199)
);

OR2x2_ASAP7_75t_L g2200 ( 
.A(n_1111),
.B(n_1129),
.Y(n_2200)
);

NAND2x1p5_ASAP7_75t_L g2201 ( 
.A(n_1384),
.B(n_1112),
.Y(n_2201)
);

NOR2x1p5_ASAP7_75t_L g2202 ( 
.A(n_1139),
.B(n_664),
.Y(n_2202)
);

AND2x6_ASAP7_75t_SL g2203 ( 
.A(n_1411),
.B(n_991),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1291),
.Y(n_2204)
);

AOI21xp5_ASAP7_75t_L g2205 ( 
.A1(n_1107),
.A2(n_1183),
.B(n_1437),
.Y(n_2205)
);

NOR2xp33_ASAP7_75t_L g2206 ( 
.A(n_1453),
.B(n_1539),
.Y(n_2206)
);

INVx2_ASAP7_75t_SL g2207 ( 
.A(n_1200),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_SL g2208 ( 
.A(n_1107),
.B(n_1437),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1291),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1291),
.Y(n_2210)
);

O2A1O1Ixp33_ASAP7_75t_L g2211 ( 
.A1(n_1107),
.A2(n_1437),
.B(n_1439),
.C(n_1605),
.Y(n_2211)
);

OAI22xp33_ASAP7_75t_L g2212 ( 
.A1(n_1437),
.A2(n_1439),
.B1(n_1605),
.B2(n_1539),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_1389),
.Y(n_2213)
);

AND2x4_ASAP7_75t_L g2214 ( 
.A(n_1394),
.B(n_1543),
.Y(n_2214)
);

AND2x4_ASAP7_75t_L g2215 ( 
.A(n_1394),
.B(n_1543),
.Y(n_2215)
);

AOI22xp33_ASAP7_75t_L g2216 ( 
.A1(n_1568),
.A2(n_1447),
.B1(n_1534),
.B2(n_1414),
.Y(n_2216)
);

BUFx3_ASAP7_75t_L g2217 ( 
.A(n_1200),
.Y(n_2217)
);

NAND3xp33_ASAP7_75t_L g2218 ( 
.A(n_1107),
.B(n_1539),
.C(n_1453),
.Y(n_2218)
);

AND2x4_ASAP7_75t_L g2219 ( 
.A(n_1394),
.B(n_1543),
.Y(n_2219)
);

BUFx3_ASAP7_75t_L g2220 ( 
.A(n_1200),
.Y(n_2220)
);

AOI22xp33_ASAP7_75t_L g2221 ( 
.A1(n_1568),
.A2(n_1447),
.B1(n_1534),
.B2(n_1414),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2223)
);

NOR2xp33_ASAP7_75t_L g2224 ( 
.A(n_1453),
.B(n_1539),
.Y(n_2224)
);

AOI22xp33_ASAP7_75t_L g2225 ( 
.A1(n_1568),
.A2(n_1447),
.B1(n_1534),
.B2(n_1414),
.Y(n_2225)
);

HB1xp67_ASAP7_75t_L g2226 ( 
.A(n_1402),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2227)
);

NAND2x1p5_ASAP7_75t_L g2228 ( 
.A(n_1384),
.B(n_1112),
.Y(n_2228)
);

OR2x6_ASAP7_75t_L g2229 ( 
.A(n_1208),
.B(n_1216),
.Y(n_2229)
);

HB1xp67_ASAP7_75t_L g2230 ( 
.A(n_1402),
.Y(n_2230)
);

OAI22xp5_ASAP7_75t_L g2231 ( 
.A1(n_1437),
.A2(n_1439),
.B1(n_1107),
.B2(n_1453),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1291),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1291),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1291),
.Y(n_2234)
);

NAND3xp33_ASAP7_75t_SL g2235 ( 
.A(n_1605),
.B(n_1552),
.C(n_1492),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1291),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1291),
.Y(n_2237)
);

OR2x2_ASAP7_75t_SL g2238 ( 
.A(n_1453),
.B(n_1539),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_1389),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2240)
);

AND2x2_ASAP7_75t_L g2241 ( 
.A(n_1129),
.B(n_1300),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_1291),
.Y(n_2242)
);

INVx2_ASAP7_75t_SL g2243 ( 
.A(n_1200),
.Y(n_2243)
);

BUFx8_ASAP7_75t_L g2244 ( 
.A(n_1292),
.Y(n_2244)
);

NOR2xp33_ASAP7_75t_L g2245 ( 
.A(n_1453),
.B(n_1539),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2246)
);

AND2x4_ASAP7_75t_L g2247 ( 
.A(n_1394),
.B(n_1543),
.Y(n_2247)
);

HB1xp67_ASAP7_75t_L g2248 ( 
.A(n_1402),
.Y(n_2248)
);

OR2x2_ASAP7_75t_L g2249 ( 
.A(n_1111),
.B(n_1129),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_1389),
.Y(n_2250)
);

AND2x4_ASAP7_75t_L g2251 ( 
.A(n_1394),
.B(n_1543),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1291),
.Y(n_2252)
);

OAI22xp5_ASAP7_75t_L g2253 ( 
.A1(n_1437),
.A2(n_1439),
.B1(n_1107),
.B2(n_1453),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_1389),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1291),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1291),
.Y(n_2256)
);

OAI22xp33_ASAP7_75t_L g2257 ( 
.A1(n_1437),
.A2(n_1439),
.B1(n_1605),
.B2(n_1539),
.Y(n_2257)
);

AO22x1_ASAP7_75t_L g2258 ( 
.A1(n_1568),
.A2(n_1437),
.B1(n_1439),
.B2(n_1132),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2259)
);

INVx5_ASAP7_75t_L g2260 ( 
.A(n_1390),
.Y(n_2260)
);

NAND2x1_ASAP7_75t_L g2261 ( 
.A(n_1568),
.B(n_1390),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_1389),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_SL g2263 ( 
.A(n_1107),
.B(n_1437),
.Y(n_2263)
);

HB1xp67_ASAP7_75t_L g2264 ( 
.A(n_1402),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_SL g2265 ( 
.A(n_1107),
.B(n_1437),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1291),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1389),
.Y(n_2267)
);

CKINVDCx20_ASAP7_75t_R g2268 ( 
.A(n_1128),
.Y(n_2268)
);

INVx2_ASAP7_75t_SL g2269 ( 
.A(n_1200),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1291),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_1389),
.Y(n_2271)
);

CKINVDCx8_ASAP7_75t_R g2272 ( 
.A(n_1105),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_1389),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_SL g2274 ( 
.A(n_1107),
.B(n_1437),
.Y(n_2274)
);

OR2x2_ASAP7_75t_SL g2275 ( 
.A(n_1453),
.B(n_1539),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_1291),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1291),
.Y(n_2278)
);

AND2x2_ASAP7_75t_L g2279 ( 
.A(n_1129),
.B(n_1300),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_1129),
.B(n_1300),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_SL g2281 ( 
.A(n_1107),
.B(n_1437),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_1291),
.Y(n_2282)
);

AOI22xp33_ASAP7_75t_L g2283 ( 
.A1(n_1568),
.A2(n_1447),
.B1(n_1534),
.B2(n_1414),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2284)
);

BUFx3_ASAP7_75t_L g2285 ( 
.A(n_1200),
.Y(n_2285)
);

INVxp67_ASAP7_75t_SL g2286 ( 
.A(n_1590),
.Y(n_2286)
);

AND2x4_ASAP7_75t_L g2287 ( 
.A(n_1394),
.B(n_1543),
.Y(n_2287)
);

HB1xp67_ASAP7_75t_L g2288 ( 
.A(n_1402),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_1291),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_1389),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_SL g2292 ( 
.A(n_1107),
.B(n_1437),
.Y(n_2292)
);

AOI21xp5_ASAP7_75t_L g2293 ( 
.A1(n_1107),
.A2(n_1183),
.B(n_1437),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_1129),
.B(n_1300),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2295)
);

BUFx8_ASAP7_75t_L g2296 ( 
.A(n_1292),
.Y(n_2296)
);

AOI22xp5_ASAP7_75t_L g2297 ( 
.A1(n_1568),
.A2(n_1437),
.B1(n_1439),
.B2(n_1101),
.Y(n_2297)
);

OR2x2_ASAP7_75t_L g2298 ( 
.A(n_1111),
.B(n_1129),
.Y(n_2298)
);

INVx1_ASAP7_75t_SL g2299 ( 
.A(n_1402),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_SL g2300 ( 
.A(n_1107),
.B(n_1437),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_1389),
.Y(n_2301)
);

NOR2x1p5_ASAP7_75t_L g2302 ( 
.A(n_1139),
.B(n_664),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_1389),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_1291),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_SL g2307 ( 
.A(n_1107),
.B(n_1437),
.Y(n_2307)
);

AOI22xp5_ASAP7_75t_L g2308 ( 
.A1(n_1568),
.A2(n_1437),
.B1(n_1439),
.B2(n_1101),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_1291),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_1129),
.B(n_1300),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_1129),
.B(n_1606),
.Y(n_2311)
);

AND2x2_ASAP7_75t_L g2312 ( 
.A(n_1129),
.B(n_1300),
.Y(n_2312)
);

AND2x4_ASAP7_75t_L g2313 ( 
.A(n_1394),
.B(n_1543),
.Y(n_2313)
);

BUFx6f_ASAP7_75t_L g2314 ( 
.A(n_1390),
.Y(n_2314)
);

HB1xp67_ASAP7_75t_L g2315 ( 
.A(n_1402),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_1291),
.Y(n_2316)
);

HB1xp67_ASAP7_75t_L g2317 ( 
.A(n_1402),
.Y(n_2317)
);

CKINVDCx5p33_ASAP7_75t_R g2318 ( 
.A(n_1128),
.Y(n_2318)
);

INVx2_ASAP7_75t_SL g2319 ( 
.A(n_1200),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_1389),
.Y(n_2320)
);

OAI21xp33_ASAP7_75t_L g2321 ( 
.A1(n_2079),
.A2(n_2143),
.B(n_2147),
.Y(n_2321)
);

CKINVDCx10_ASAP7_75t_R g2322 ( 
.A(n_2180),
.Y(n_2322)
);

AND2x4_ASAP7_75t_L g2323 ( 
.A(n_2068),
.B(n_1625),
.Y(n_2323)
);

HB1xp67_ASAP7_75t_L g2324 ( 
.A(n_2315),
.Y(n_2324)
);

OAI21x1_ASAP7_75t_L g2325 ( 
.A1(n_1932),
.A2(n_1673),
.B(n_1895),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_2143),
.B(n_2068),
.Y(n_2326)
);

BUFx6f_ASAP7_75t_L g2327 ( 
.A(n_1623),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_1658),
.B(n_1660),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_1645),
.Y(n_2329)
);

NOR2xp33_ASAP7_75t_L g2330 ( 
.A(n_1636),
.B(n_1639),
.Y(n_2330)
);

NOR2xp67_ASAP7_75t_L g2331 ( 
.A(n_1635),
.B(n_2062),
.Y(n_2331)
);

A2O1A1Ixp33_ASAP7_75t_L g2332 ( 
.A1(n_2211),
.A2(n_2135),
.B(n_2094),
.C(n_2124),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_1742),
.B(n_1746),
.Y(n_2333)
);

AOI21xp5_ASAP7_75t_L g2334 ( 
.A1(n_2058),
.A2(n_2193),
.B(n_2117),
.Y(n_2334)
);

AO21x2_ASAP7_75t_L g2335 ( 
.A1(n_2011),
.A2(n_2014),
.B(n_2091),
.Y(n_2335)
);

INVx3_ASAP7_75t_L g2336 ( 
.A(n_1878),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_1645),
.Y(n_2337)
);

OAI21xp5_ASAP7_75t_L g2338 ( 
.A1(n_2190),
.A2(n_2205),
.B(n_2101),
.Y(n_2338)
);

AOI21xp5_ASAP7_75t_L g2339 ( 
.A1(n_2293),
.A2(n_2100),
.B(n_2092),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_SL g2340 ( 
.A(n_2076),
.B(n_2212),
.Y(n_2340)
);

AOI21xp5_ASAP7_75t_L g2341 ( 
.A1(n_2159),
.A2(n_2173),
.B(n_2165),
.Y(n_2341)
);

OAI22xp5_ASAP7_75t_L g2342 ( 
.A1(n_1615),
.A2(n_2102),
.B1(n_2124),
.B2(n_2094),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_1742),
.B(n_1746),
.Y(n_2343)
);

NOR2xp33_ASAP7_75t_L g2344 ( 
.A(n_1680),
.B(n_1681),
.Y(n_2344)
);

AND2x2_ASAP7_75t_L g2345 ( 
.A(n_1615),
.B(n_2102),
.Y(n_2345)
);

OAI21xp5_ASAP7_75t_L g2346 ( 
.A1(n_2064),
.A2(n_2072),
.B(n_2147),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_1751),
.B(n_1755),
.Y(n_2347)
);

AOI21xp5_ASAP7_75t_L g2348 ( 
.A1(n_2178),
.A2(n_2192),
.B(n_2181),
.Y(n_2348)
);

A2O1A1Ixp33_ASAP7_75t_L g2349 ( 
.A1(n_2125),
.A2(n_2195),
.B(n_2297),
.C(n_2133),
.Y(n_2349)
);

OAI21xp5_ASAP7_75t_L g2350 ( 
.A1(n_2231),
.A2(n_2253),
.B(n_2257),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_1618),
.B(n_1685),
.Y(n_2351)
);

OAI22xp5_ASAP7_75t_L g2352 ( 
.A1(n_2125),
.A2(n_2133),
.B1(n_2155),
.B2(n_2130),
.Y(n_2352)
);

BUFx3_ASAP7_75t_L g2353 ( 
.A(n_1798),
.Y(n_2353)
);

AOI21x1_ASAP7_75t_L g2354 ( 
.A1(n_2258),
.A2(n_2263),
.B(n_2208),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2081),
.Y(n_2355)
);

BUFx6f_ASAP7_75t_L g2356 ( 
.A(n_1623),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_1618),
.B(n_1685),
.Y(n_2357)
);

AOI21xp5_ASAP7_75t_L g2358 ( 
.A1(n_2265),
.A2(n_2292),
.B(n_2281),
.Y(n_2358)
);

AOI21xp5_ASAP7_75t_L g2359 ( 
.A1(n_2300),
.A2(n_2307),
.B(n_2274),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2200),
.B(n_2249),
.Y(n_2360)
);

BUFx8_ASAP7_75t_L g2361 ( 
.A(n_2129),
.Y(n_2361)
);

AOI21xp5_ASAP7_75t_L g2362 ( 
.A1(n_1627),
.A2(n_2070),
.B(n_2258),
.Y(n_2362)
);

BUFx6f_ASAP7_75t_L g2363 ( 
.A(n_1623),
.Y(n_2363)
);

NOR2xp33_ASAP7_75t_L g2364 ( 
.A(n_1644),
.B(n_1838),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_SL g2365 ( 
.A(n_1840),
.B(n_1844),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_SL g2366 ( 
.A(n_1840),
.B(n_1844),
.Y(n_2366)
);

INVxp67_ASAP7_75t_L g2367 ( 
.A(n_1698),
.Y(n_2367)
);

NAND2x1_ASAP7_75t_L g2368 ( 
.A(n_1788),
.B(n_1802),
.Y(n_2368)
);

O2A1O1Ixp33_ASAP7_75t_L g2369 ( 
.A1(n_1619),
.A2(n_2235),
.B(n_2112),
.C(n_2231),
.Y(n_2369)
);

NAND3xp33_ASAP7_75t_L g2370 ( 
.A(n_2253),
.B(n_2218),
.C(n_1628),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_2130),
.B(n_2155),
.Y(n_2371)
);

NOR2xp33_ASAP7_75t_L g2372 ( 
.A(n_1644),
.B(n_1756),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_2081),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_1751),
.B(n_1755),
.Y(n_2374)
);

NAND3xp33_ASAP7_75t_L g2375 ( 
.A(n_2218),
.B(n_1628),
.C(n_2153),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_1764),
.B(n_1767),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2081),
.Y(n_2377)
);

NOR2xp33_ASAP7_75t_L g2378 ( 
.A(n_1707),
.B(n_1754),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_SL g2379 ( 
.A(n_1699),
.B(n_1617),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_SL g2380 ( 
.A(n_1699),
.B(n_1617),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_1764),
.B(n_1767),
.Y(n_2381)
);

CKINVDCx8_ASAP7_75t_R g2382 ( 
.A(n_2203),
.Y(n_2382)
);

AND2x4_ASAP7_75t_L g2383 ( 
.A(n_1625),
.B(n_1688),
.Y(n_2383)
);

BUFx6f_ASAP7_75t_L g2384 ( 
.A(n_1623),
.Y(n_2384)
);

OR2x2_ASAP7_75t_L g2385 ( 
.A(n_1682),
.B(n_1640),
.Y(n_2385)
);

O2A1O1Ixp33_ASAP7_75t_L g2386 ( 
.A1(n_1619),
.A2(n_2153),
.B(n_1704),
.C(n_1648),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_1775),
.B(n_1800),
.Y(n_2387)
);

AOI22xp5_ASAP7_75t_L g2388 ( 
.A1(n_2079),
.A2(n_1689),
.B1(n_2297),
.B2(n_2195),
.Y(n_2388)
);

AO31x2_ASAP7_75t_L g2389 ( 
.A1(n_2011),
.A2(n_2014),
.A3(n_1705),
.B(n_1640),
.Y(n_2389)
);

AOI221xp5_ASAP7_75t_L g2390 ( 
.A1(n_1689),
.A2(n_2096),
.B1(n_2191),
.B2(n_2162),
.C(n_2084),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_2116),
.Y(n_2391)
);

AOI21xp5_ASAP7_75t_L g2392 ( 
.A1(n_1627),
.A2(n_2070),
.B(n_2079),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2116),
.Y(n_2393)
);

BUFx3_ASAP7_75t_L g2394 ( 
.A(n_1798),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2116),
.Y(n_2395)
);

AOI21xp5_ASAP7_75t_L g2396 ( 
.A1(n_1627),
.A2(n_2070),
.B(n_2308),
.Y(n_2396)
);

AOI21xp5_ASAP7_75t_L g2397 ( 
.A1(n_2308),
.A2(n_1713),
.B(n_1670),
.Y(n_2397)
);

BUFx12f_ASAP7_75t_L g2398 ( 
.A(n_1745),
.Y(n_2398)
);

OAI21xp5_ASAP7_75t_L g2399 ( 
.A1(n_1630),
.A2(n_2206),
.B(n_2198),
.Y(n_2399)
);

NAND3xp33_ASAP7_75t_L g2400 ( 
.A(n_1630),
.B(n_2245),
.C(n_2224),
.Y(n_2400)
);

AOI21xp33_ASAP7_75t_L g2401 ( 
.A1(n_1696),
.A2(n_1763),
.B(n_1682),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2131),
.Y(n_2402)
);

OAI21xp33_ASAP7_75t_L g2403 ( 
.A1(n_1704),
.A2(n_1782),
.B(n_1657),
.Y(n_2403)
);

OAI21xp5_ASAP7_75t_L g2404 ( 
.A1(n_1650),
.A2(n_1705),
.B(n_1657),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_2131),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2131),
.Y(n_2406)
);

O2A1O1Ixp33_ASAP7_75t_L g2407 ( 
.A1(n_1803),
.A2(n_2073),
.B(n_2080),
.C(n_2077),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2137),
.Y(n_2408)
);

INVx11_ASAP7_75t_L g2409 ( 
.A(n_1745),
.Y(n_2409)
);

INVxp67_ASAP7_75t_L g2410 ( 
.A(n_1885),
.Y(n_2410)
);

CKINVDCx5p33_ASAP7_75t_R g2411 ( 
.A(n_2071),
.Y(n_2411)
);

NOR2x1_ASAP7_75t_L g2412 ( 
.A(n_1651),
.B(n_1832),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_1775),
.B(n_1800),
.Y(n_2413)
);

AOI21x1_ASAP7_75t_L g2414 ( 
.A1(n_1700),
.A2(n_1833),
.B(n_2044),
.Y(n_2414)
);

AOI21xp5_ASAP7_75t_L g2415 ( 
.A1(n_1670),
.A2(n_1714),
.B(n_1713),
.Y(n_2415)
);

OAI21x1_ASAP7_75t_L g2416 ( 
.A1(n_1990),
.A2(n_1980),
.B(n_1962),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_SL g2417 ( 
.A(n_2073),
.B(n_2077),
.Y(n_2417)
);

NOR2xp33_ASAP7_75t_L g2418 ( 
.A(n_1784),
.B(n_1695),
.Y(n_2418)
);

AOI21xp5_ASAP7_75t_L g2419 ( 
.A1(n_1714),
.A2(n_1716),
.B(n_1715),
.Y(n_2419)
);

BUFx12f_ASAP7_75t_L g2420 ( 
.A(n_1745),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2080),
.B(n_2090),
.Y(n_2421)
);

NAND3xp33_ASAP7_75t_L g2422 ( 
.A(n_1809),
.B(n_1650),
.C(n_1649),
.Y(n_2422)
);

BUFx6f_ASAP7_75t_L g2423 ( 
.A(n_1623),
.Y(n_2423)
);

NOR3xp33_ASAP7_75t_L g2424 ( 
.A(n_1757),
.B(n_1700),
.C(n_2090),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2200),
.B(n_2249),
.Y(n_2425)
);

INVx5_ASAP7_75t_L g2426 ( 
.A(n_2082),
.Y(n_2426)
);

AOI21xp5_ASAP7_75t_L g2427 ( 
.A1(n_1715),
.A2(n_1730),
.B(n_1716),
.Y(n_2427)
);

OAI22xp5_ASAP7_75t_L g2428 ( 
.A1(n_2197),
.A2(n_2275),
.B1(n_2238),
.B2(n_1646),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_2103),
.B(n_2104),
.Y(n_2429)
);

AOI21xp5_ASAP7_75t_L g2430 ( 
.A1(n_1730),
.A2(n_1732),
.B(n_1663),
.Y(n_2430)
);

O2A1O1Ixp33_ASAP7_75t_L g2431 ( 
.A1(n_2103),
.A2(n_2107),
.B(n_2113),
.C(n_2104),
.Y(n_2431)
);

AOI21xp5_ASAP7_75t_L g2432 ( 
.A1(n_1732),
.A2(n_1734),
.B(n_1694),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2107),
.B(n_2113),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2137),
.Y(n_2434)
);

AOI21xp5_ASAP7_75t_L g2435 ( 
.A1(n_1694),
.A2(n_1734),
.B(n_1629),
.Y(n_2435)
);

OAI21xp5_ASAP7_75t_L g2436 ( 
.A1(n_1649),
.A2(n_1797),
.B(n_1725),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2137),
.Y(n_2437)
);

INVxp67_ASAP7_75t_L g2438 ( 
.A(n_1616),
.Y(n_2438)
);

AOI21xp5_ASAP7_75t_L g2439 ( 
.A1(n_1694),
.A2(n_1734),
.B(n_1629),
.Y(n_2439)
);

NAND3xp33_ASAP7_75t_L g2440 ( 
.A(n_1725),
.B(n_1797),
.C(n_1761),
.Y(n_2440)
);

A2O1A1Ixp33_ASAP7_75t_L g2441 ( 
.A1(n_1884),
.A2(n_2065),
.B(n_2109),
.C(n_2078),
.Y(n_2441)
);

OAI22xp5_ASAP7_75t_L g2442 ( 
.A1(n_2197),
.A2(n_2238),
.B1(n_2275),
.B2(n_1646),
.Y(n_2442)
);

OAI21xp5_ASAP7_75t_L g2443 ( 
.A1(n_1776),
.A2(n_2119),
.B(n_2115),
.Y(n_2443)
);

O2A1O1Ixp5_ASAP7_75t_L g2444 ( 
.A1(n_1847),
.A2(n_1998),
.B(n_2020),
.C(n_1766),
.Y(n_2444)
);

OAI22xp5_ASAP7_75t_L g2445 ( 
.A1(n_2129),
.A2(n_2175),
.B1(n_1743),
.B2(n_2142),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2115),
.B(n_2121),
.Y(n_2446)
);

AOI21xp5_ASAP7_75t_L g2447 ( 
.A1(n_2082),
.A2(n_2122),
.B(n_2121),
.Y(n_2447)
);

NOR2x1_ASAP7_75t_L g2448 ( 
.A(n_1651),
.B(n_2298),
.Y(n_2448)
);

INVxp67_ASAP7_75t_L g2449 ( 
.A(n_2063),
.Y(n_2449)
);

OR2x2_ASAP7_75t_L g2450 ( 
.A(n_1656),
.B(n_1740),
.Y(n_2450)
);

O2A1O1Ixp5_ASAP7_75t_L g2451 ( 
.A1(n_2020),
.A2(n_2047),
.B(n_2033),
.C(n_2054),
.Y(n_2451)
);

AOI22xp5_ASAP7_75t_L g2452 ( 
.A1(n_2176),
.A2(n_2221),
.B1(n_2225),
.B2(n_2216),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2145),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_SL g2454 ( 
.A(n_2122),
.B(n_2132),
.Y(n_2454)
);

AOI22xp33_ASAP7_75t_L g2455 ( 
.A1(n_2283),
.A2(n_1676),
.B1(n_2175),
.B2(n_2129),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2298),
.B(n_2132),
.Y(n_2456)
);

AOI21xp5_ASAP7_75t_L g2457 ( 
.A1(n_2134),
.A2(n_2150),
.B(n_2149),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2134),
.B(n_2149),
.Y(n_2458)
);

NOR2xp33_ASAP7_75t_L g2459 ( 
.A(n_1695),
.B(n_1839),
.Y(n_2459)
);

AOI21xp5_ASAP7_75t_L g2460 ( 
.A1(n_2150),
.A2(n_2160),
.B(n_2157),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_SL g2461 ( 
.A(n_2157),
.B(n_2160),
.Y(n_2461)
);

NOR2xp33_ASAP7_75t_L g2462 ( 
.A(n_1757),
.B(n_1743),
.Y(n_2462)
);

NAND2xp33_ASAP7_75t_L g2463 ( 
.A(n_1641),
.B(n_2161),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_2161),
.B(n_2183),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_L g2465 ( 
.A(n_2183),
.B(n_2186),
.Y(n_2465)
);

INVx3_ASAP7_75t_L g2466 ( 
.A(n_1878),
.Y(n_2466)
);

AOI21xp5_ASAP7_75t_L g2467 ( 
.A1(n_2186),
.A2(n_2222),
.B(n_2189),
.Y(n_2467)
);

AOI21xp5_ASAP7_75t_L g2468 ( 
.A1(n_2189),
.A2(n_2223),
.B(n_2222),
.Y(n_2468)
);

INVx2_ASAP7_75t_L g2469 ( 
.A(n_2145),
.Y(n_2469)
);

AOI21xp5_ASAP7_75t_L g2470 ( 
.A1(n_2223),
.A2(n_2240),
.B(n_2227),
.Y(n_2470)
);

INVx11_ASAP7_75t_L g2471 ( 
.A(n_1745),
.Y(n_2471)
);

INVx2_ASAP7_75t_SL g2472 ( 
.A(n_1900),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_SL g2473 ( 
.A(n_2227),
.B(n_2240),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_SL g2474 ( 
.A(n_2246),
.B(n_2259),
.Y(n_2474)
);

AOI21xp5_ASAP7_75t_L g2475 ( 
.A1(n_2246),
.A2(n_2276),
.B(n_2259),
.Y(n_2475)
);

AOI21xp5_ASAP7_75t_L g2476 ( 
.A1(n_2276),
.A2(n_2290),
.B(n_2284),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2284),
.B(n_2290),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2295),
.B(n_2303),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2295),
.B(n_2303),
.Y(n_2479)
);

AND2x2_ASAP7_75t_L g2480 ( 
.A(n_1697),
.B(n_1818),
.Y(n_2480)
);

CKINVDCx10_ASAP7_75t_R g2481 ( 
.A(n_2129),
.Y(n_2481)
);

AOI21xp5_ASAP7_75t_L g2482 ( 
.A1(n_2306),
.A2(n_2311),
.B(n_2261),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_SL g2483 ( 
.A(n_2306),
.B(n_2311),
.Y(n_2483)
);

AOI21xp5_ASAP7_75t_L g2484 ( 
.A1(n_1788),
.A2(n_1802),
.B(n_2013),
.Y(n_2484)
);

OAI321xp33_ASAP7_75t_L g2485 ( 
.A1(n_1884),
.A2(n_1819),
.A3(n_1735),
.B1(n_1804),
.B2(n_1959),
.C(n_1796),
.Y(n_2485)
);

AND2x4_ASAP7_75t_L g2486 ( 
.A(n_1625),
.B(n_1688),
.Y(n_2486)
);

O2A1O1Ixp33_ASAP7_75t_L g2487 ( 
.A1(n_1834),
.A2(n_1852),
.B(n_1816),
.C(n_1991),
.Y(n_2487)
);

AOI33xp33_ASAP7_75t_L g2488 ( 
.A1(n_2105),
.A2(n_2120),
.A3(n_2182),
.B1(n_2279),
.B2(n_2241),
.B3(n_2127),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2146),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_1620),
.B(n_1626),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_1654),
.B(n_1662),
.Y(n_2491)
);

BUFx6f_ASAP7_75t_L g2492 ( 
.A(n_1623),
.Y(n_2492)
);

A2O1A1Ixp33_ASAP7_75t_L g2493 ( 
.A1(n_1655),
.A2(n_1804),
.B(n_1740),
.C(n_1735),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_2146),
.Y(n_2494)
);

AOI21xp5_ASAP7_75t_L g2495 ( 
.A1(n_2024),
.A2(n_2017),
.B(n_1718),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_1665),
.B(n_1687),
.Y(n_2496)
);

INVx4_ASAP7_75t_L g2497 ( 
.A(n_2175),
.Y(n_2497)
);

AOI22xp5_ASAP7_75t_L g2498 ( 
.A1(n_2175),
.A2(n_2105),
.B1(n_2127),
.B2(n_2120),
.Y(n_2498)
);

INVxp67_ASAP7_75t_L g2499 ( 
.A(n_2067),
.Y(n_2499)
);

AOI21xp5_ASAP7_75t_L g2500 ( 
.A1(n_2017),
.A2(n_1718),
.B(n_1712),
.Y(n_2500)
);

OR2x6_ASAP7_75t_L g2501 ( 
.A(n_1787),
.B(n_1796),
.Y(n_2501)
);

NOR2xp33_ASAP7_75t_L g2502 ( 
.A(n_2182),
.B(n_2241),
.Y(n_2502)
);

INVx3_ASAP7_75t_L g2503 ( 
.A(n_1878),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_1702),
.B(n_1736),
.Y(n_2504)
);

AOI21x1_ASAP7_75t_L g2505 ( 
.A1(n_2054),
.A2(n_2021),
.B(n_1841),
.Y(n_2505)
);

OAI22xp33_ASAP7_75t_L g2506 ( 
.A1(n_1930),
.A2(n_1806),
.B1(n_1796),
.B2(n_1787),
.Y(n_2506)
);

BUFx4f_ASAP7_75t_L g2507 ( 
.A(n_1631),
.Y(n_2507)
);

NOR2xp33_ASAP7_75t_L g2508 ( 
.A(n_2279),
.B(n_2280),
.Y(n_2508)
);

A2O1A1Ixp33_ASAP7_75t_L g2509 ( 
.A1(n_1676),
.A2(n_1873),
.B(n_1899),
.C(n_1718),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_L g2510 ( 
.A(n_1741),
.B(n_1752),
.Y(n_2510)
);

AOI21xp5_ASAP7_75t_L g2511 ( 
.A1(n_2017),
.A2(n_1718),
.B(n_1712),
.Y(n_2511)
);

CKINVDCx5p33_ASAP7_75t_R g2512 ( 
.A(n_1739),
.Y(n_2512)
);

HB1xp67_ASAP7_75t_L g2513 ( 
.A(n_2108),
.Y(n_2513)
);

AND2x2_ASAP7_75t_L g2514 ( 
.A(n_1697),
.B(n_1818),
.Y(n_2514)
);

INVx2_ASAP7_75t_L g2515 ( 
.A(n_2164),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2164),
.Y(n_2516)
);

NOR2xp33_ASAP7_75t_L g2517 ( 
.A(n_2280),
.B(n_2294),
.Y(n_2517)
);

INVxp67_ASAP7_75t_L g2518 ( 
.A(n_2152),
.Y(n_2518)
);

BUFx2_ASAP7_75t_SL g2519 ( 
.A(n_1635),
.Y(n_2519)
);

O2A1O1Ixp33_ASAP7_75t_L g2520 ( 
.A1(n_1760),
.A2(n_1777),
.B(n_1762),
.C(n_2226),
.Y(n_2520)
);

BUFx6f_ASAP7_75t_L g2521 ( 
.A(n_1631),
.Y(n_2521)
);

NOR2xp33_ASAP7_75t_L g2522 ( 
.A(n_2294),
.B(n_2310),
.Y(n_2522)
);

AOI22xp5_ASAP7_75t_L g2523 ( 
.A1(n_2310),
.A2(n_2312),
.B1(n_2166),
.B2(n_1908),
.Y(n_2523)
);

INVx3_ASAP7_75t_L g2524 ( 
.A(n_1878),
.Y(n_2524)
);

O2A1O1Ixp33_ASAP7_75t_L g2525 ( 
.A1(n_2230),
.A2(n_2248),
.B(n_2288),
.C(n_2264),
.Y(n_2525)
);

OAI21x1_ASAP7_75t_L g2526 ( 
.A1(n_1962),
.A2(n_2003),
.B(n_1980),
.Y(n_2526)
);

NOR2xp33_ASAP7_75t_L g2527 ( 
.A(n_2312),
.B(n_1748),
.Y(n_2527)
);

BUFx8_ASAP7_75t_L g2528 ( 
.A(n_2118),
.Y(n_2528)
);

AOI21xp5_ASAP7_75t_L g2529 ( 
.A1(n_1712),
.A2(n_2016),
.B(n_1635),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_1634),
.B(n_1843),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2169),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_SL g2532 ( 
.A(n_1625),
.B(n_1688),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2169),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2169),
.Y(n_2534)
);

NAND3xp33_ASAP7_75t_L g2535 ( 
.A(n_1888),
.B(n_1903),
.C(n_2015),
.Y(n_2535)
);

INVx2_ASAP7_75t_SL g2536 ( 
.A(n_1900),
.Y(n_2536)
);

OAI21xp5_ASAP7_75t_L g2537 ( 
.A1(n_1903),
.A2(n_1841),
.B(n_2018),
.Y(n_2537)
);

AOI22xp5_ASAP7_75t_L g2538 ( 
.A1(n_2166),
.A2(n_1908),
.B1(n_1807),
.B2(n_1930),
.Y(n_2538)
);

INVx6_ASAP7_75t_L g2539 ( 
.A(n_1900),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_1634),
.B(n_1843),
.Y(n_2540)
);

AND2x4_ASAP7_75t_L g2541 ( 
.A(n_1688),
.B(n_1710),
.Y(n_2541)
);

NOR3xp33_ASAP7_75t_L g2542 ( 
.A(n_1993),
.B(n_2056),
.C(n_2037),
.Y(n_2542)
);

AND2x2_ASAP7_75t_L g2543 ( 
.A(n_1664),
.B(n_1996),
.Y(n_2543)
);

AOI22xp5_ASAP7_75t_L g2544 ( 
.A1(n_2166),
.A2(n_1822),
.B1(n_2095),
.B2(n_1710),
.Y(n_2544)
);

O2A1O1Ixp5_ASAP7_75t_L g2545 ( 
.A1(n_1892),
.A2(n_1893),
.B(n_1914),
.C(n_1898),
.Y(n_2545)
);

OAI21xp5_ASAP7_75t_L g2546 ( 
.A1(n_2057),
.A2(n_1883),
.B(n_1822),
.Y(n_2546)
);

INVx4_ASAP7_75t_L g2547 ( 
.A(n_1635),
.Y(n_2547)
);

AOI33xp33_ASAP7_75t_L g2548 ( 
.A1(n_1653),
.A2(n_1709),
.A3(n_2299),
.B1(n_2066),
.B2(n_1972),
.B3(n_1955),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_1724),
.B(n_1667),
.Y(n_2549)
);

INVx2_ASAP7_75t_SL g2550 ( 
.A(n_1900),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_1667),
.B(n_1668),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_1668),
.B(n_1674),
.Y(n_2552)
);

AO32x1_ASAP7_75t_L g2553 ( 
.A1(n_2171),
.A2(n_2213),
.A3(n_2239),
.B1(n_2199),
.B2(n_2174),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_SL g2554 ( 
.A(n_1710),
.B(n_2095),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_SL g2555 ( 
.A(n_1710),
.B(n_2095),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_1674),
.B(n_1675),
.Y(n_2556)
);

CKINVDCx10_ASAP7_75t_R g2557 ( 
.A(n_1669),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2171),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_2174),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_SL g2560 ( 
.A(n_2095),
.B(n_2110),
.Y(n_2560)
);

NOR2xp33_ASAP7_75t_L g2561 ( 
.A(n_1795),
.B(n_2317),
.Y(n_2561)
);

OAI22xp5_ASAP7_75t_L g2562 ( 
.A1(n_1791),
.A2(n_1737),
.B1(n_1796),
.B2(n_1787),
.Y(n_2562)
);

O2A1O1Ixp33_ASAP7_75t_L g2563 ( 
.A1(n_1939),
.A2(n_1643),
.B(n_1896),
.C(n_1891),
.Y(n_2563)
);

NOR2xp33_ASAP7_75t_L g2564 ( 
.A(n_1795),
.B(n_1982),
.Y(n_2564)
);

INVxp67_ASAP7_75t_SL g2565 ( 
.A(n_1883),
.Y(n_2565)
);

NAND3xp33_ASAP7_75t_L g2566 ( 
.A(n_2049),
.B(n_1656),
.C(n_2036),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_SL g2567 ( 
.A(n_2110),
.B(n_2123),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_1675),
.B(n_1678),
.Y(n_2568)
);

O2A1O1Ixp33_ASAP7_75t_L g2569 ( 
.A1(n_1939),
.A2(n_1891),
.B(n_1901),
.C(n_1896),
.Y(n_2569)
);

A2O1A1Ixp33_ASAP7_75t_L g2570 ( 
.A1(n_1899),
.A2(n_1999),
.B(n_1678),
.C(n_1854),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_1978),
.B(n_1988),
.Y(n_2571)
);

OAI22xp5_ASAP7_75t_L g2572 ( 
.A1(n_1791),
.A2(n_1737),
.B1(n_1796),
.B2(n_1787),
.Y(n_2572)
);

AOI22xp5_ASAP7_75t_L g2573 ( 
.A1(n_2166),
.A2(n_2123),
.B1(n_2184),
.B2(n_2110),
.Y(n_2573)
);

OR2x6_ASAP7_75t_L g2574 ( 
.A(n_1787),
.B(n_1669),
.Y(n_2574)
);

O2A1O1Ixp33_ASAP7_75t_L g2575 ( 
.A1(n_1901),
.A2(n_1904),
.B(n_1928),
.C(n_1927),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2174),
.Y(n_2576)
);

INVx1_ASAP7_75t_SL g2577 ( 
.A(n_1653),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_2199),
.Y(n_2578)
);

OR2x6_ASAP7_75t_L g2579 ( 
.A(n_1669),
.B(n_1723),
.Y(n_2579)
);

OR2x2_ASAP7_75t_L g2580 ( 
.A(n_2199),
.B(n_2320),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2213),
.Y(n_2581)
);

AOI21xp5_ASAP7_75t_L g2582 ( 
.A1(n_2260),
.A2(n_1938),
.B(n_1957),
.Y(n_2582)
);

AOI21xp5_ASAP7_75t_L g2583 ( 
.A1(n_2260),
.A2(n_1938),
.B(n_1957),
.Y(n_2583)
);

NAND2x1_ASAP7_75t_L g2584 ( 
.A(n_2166),
.B(n_1962),
.Y(n_2584)
);

AOI22x1_ASAP7_75t_L g2585 ( 
.A1(n_1867),
.A2(n_1881),
.B1(n_1875),
.B2(n_2019),
.Y(n_2585)
);

AOI21x1_ASAP7_75t_L g2586 ( 
.A1(n_2021),
.A2(n_2031),
.B(n_2029),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_1979),
.B(n_2066),
.Y(n_2587)
);

OR2x2_ASAP7_75t_L g2588 ( 
.A(n_2213),
.B(n_2320),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2239),
.Y(n_2589)
);

A2O1A1Ixp33_ASAP7_75t_L g2590 ( 
.A1(n_1912),
.A2(n_1904),
.B(n_1928),
.C(n_1927),
.Y(n_2590)
);

OR2x6_ASAP7_75t_L g2591 ( 
.A(n_1669),
.B(n_1723),
.Y(n_2591)
);

OAI22xp5_ASAP7_75t_L g2592 ( 
.A1(n_1944),
.A2(n_1949),
.B1(n_1954),
.B2(n_1945),
.Y(n_2592)
);

AND2x2_ASAP7_75t_L g2593 ( 
.A(n_1664),
.B(n_1996),
.Y(n_2593)
);

AOI21xp33_ASAP7_75t_L g2594 ( 
.A1(n_1709),
.A2(n_2299),
.B(n_2038),
.Y(n_2594)
);

O2A1O1Ixp33_ASAP7_75t_L g2595 ( 
.A1(n_1944),
.A2(n_1949),
.B(n_1954),
.C(n_1945),
.Y(n_2595)
);

OA22x2_ASAP7_75t_L g2596 ( 
.A1(n_1912),
.A2(n_2123),
.B1(n_2184),
.B2(n_2110),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_1882),
.B(n_1952),
.Y(n_2597)
);

INVx2_ASAP7_75t_L g2598 ( 
.A(n_2250),
.Y(n_2598)
);

NAND3xp33_ASAP7_75t_L g2599 ( 
.A(n_2036),
.B(n_2042),
.C(n_2038),
.Y(n_2599)
);

INVx3_ASAP7_75t_L g2600 ( 
.A(n_1878),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_1882),
.B(n_1952),
.Y(n_2601)
);

AO22x1_ASAP7_75t_L g2602 ( 
.A1(n_2166),
.A2(n_1856),
.B1(n_2184),
.B2(n_2123),
.Y(n_2602)
);

BUFx2_ASAP7_75t_L g2603 ( 
.A(n_2166),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_L g2604 ( 
.A(n_1955),
.B(n_1972),
.Y(n_2604)
);

HB1xp67_ASAP7_75t_L g2605 ( 
.A(n_1850),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2250),
.Y(n_2606)
);

OR2x2_ASAP7_75t_L g2607 ( 
.A(n_2250),
.B(n_2320),
.Y(n_2607)
);

O2A1O1Ixp33_ASAP7_75t_L g2608 ( 
.A1(n_1963),
.A2(n_1983),
.B(n_1992),
.C(n_1977),
.Y(n_2608)
);

AOI33xp33_ASAP7_75t_L g2609 ( 
.A1(n_1621),
.A2(n_1622),
.A3(n_1624),
.B1(n_1659),
.B2(n_1652),
.B3(n_1637),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_1845),
.B(n_1907),
.Y(n_2610)
);

OAI21xp33_ASAP7_75t_L g2611 ( 
.A1(n_1679),
.A2(n_1977),
.B(n_1963),
.Y(n_2611)
);

NOR3xp33_ASAP7_75t_L g2612 ( 
.A(n_2037),
.B(n_2056),
.C(n_1974),
.Y(n_2612)
);

AND2x2_ASAP7_75t_L g2613 ( 
.A(n_1978),
.B(n_1988),
.Y(n_2613)
);

NAND3xp33_ASAP7_75t_L g2614 ( 
.A(n_2045),
.B(n_2050),
.C(n_2046),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_SL g2615 ( 
.A(n_2184),
.B(n_2214),
.Y(n_2615)
);

AOI21xp5_ASAP7_75t_L g2616 ( 
.A1(n_1931),
.A2(n_1994),
.B(n_1961),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_1845),
.B(n_1759),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_L g2618 ( 
.A(n_1759),
.B(n_1925),
.Y(n_2618)
);

NAND2x1p5_ASAP7_75t_L g2619 ( 
.A(n_1631),
.B(n_2136),
.Y(n_2619)
);

INVx2_ASAP7_75t_L g2620 ( 
.A(n_2254),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_1915),
.B(n_1872),
.Y(n_2621)
);

NOR2xp33_ASAP7_75t_L g2622 ( 
.A(n_1814),
.B(n_1981),
.Y(n_2622)
);

O2A1O1Ixp33_ASAP7_75t_L g2623 ( 
.A1(n_1983),
.A2(n_1992),
.B(n_1849),
.C(n_1848),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_1853),
.B(n_1859),
.Y(n_2624)
);

NAND2xp33_ASAP7_75t_L g2625 ( 
.A(n_1948),
.B(n_1875),
.Y(n_2625)
);

A2O1A1Ixp33_ASAP7_75t_L g2626 ( 
.A1(n_1857),
.A2(n_1997),
.B(n_1624),
.C(n_1621),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_1853),
.B(n_1859),
.Y(n_2627)
);

AOI22x1_ASAP7_75t_L g2628 ( 
.A1(n_1875),
.A2(n_2019),
.B1(n_2006),
.B2(n_1994),
.Y(n_2628)
);

NOR2xp33_ASAP7_75t_L g2629 ( 
.A(n_1814),
.B(n_1750),
.Y(n_2629)
);

O2A1O1Ixp33_ASAP7_75t_L g2630 ( 
.A1(n_1789),
.A2(n_1837),
.B(n_1810),
.C(n_1886),
.Y(n_2630)
);

BUFx6f_ASAP7_75t_L g2631 ( 
.A(n_1631),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2254),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_1868),
.B(n_1876),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_1868),
.B(n_1876),
.Y(n_2634)
);

NOR2xp33_ASAP7_75t_L g2635 ( 
.A(n_1750),
.B(n_1785),
.Y(n_2635)
);

HB1xp67_ASAP7_75t_L g2636 ( 
.A(n_2025),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2262),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_L g2638 ( 
.A(n_1879),
.B(n_1622),
.Y(n_2638)
);

AND2x2_ASAP7_75t_L g2639 ( 
.A(n_1637),
.B(n_1652),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_1879),
.B(n_1659),
.Y(n_2640)
);

AOI21xp5_ASAP7_75t_L g2641 ( 
.A1(n_2006),
.A2(n_1723),
.B(n_1669),
.Y(n_2641)
);

CKINVDCx20_ASAP7_75t_R g2642 ( 
.A(n_1786),
.Y(n_2642)
);

NOR2xp33_ASAP7_75t_L g2643 ( 
.A(n_1785),
.B(n_1793),
.Y(n_2643)
);

AOI21xp5_ASAP7_75t_L g2644 ( 
.A1(n_2006),
.A2(n_2185),
.B(n_1723),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_1661),
.B(n_2059),
.Y(n_2645)
);

NOR2xp33_ASAP7_75t_R g2646 ( 
.A(n_2074),
.B(n_2128),
.Y(n_2646)
);

INVxp67_ASAP7_75t_L g2647 ( 
.A(n_1789),
.Y(n_2647)
);

AOI21xp5_ASAP7_75t_L g2648 ( 
.A1(n_1723),
.A2(n_2229),
.B(n_2185),
.Y(n_2648)
);

INVx2_ASAP7_75t_SL g2649 ( 
.A(n_1900),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_1661),
.B(n_2059),
.Y(n_2650)
);

A2O1A1Ixp33_ASAP7_75t_L g2651 ( 
.A1(n_2060),
.A2(n_2075),
.B(n_2083),
.C(n_2061),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_L g2652 ( 
.A(n_2060),
.B(n_2061),
.Y(n_2652)
);

O2A1O1Ixp5_ASAP7_75t_L g2653 ( 
.A1(n_1933),
.A2(n_1921),
.B(n_2008),
.C(n_2043),
.Y(n_2653)
);

OAI22xp5_ASAP7_75t_L g2654 ( 
.A1(n_1793),
.A2(n_2215),
.B1(n_2219),
.B2(n_2214),
.Y(n_2654)
);

A2O1A1Ixp33_ASAP7_75t_L g2655 ( 
.A1(n_2075),
.A2(n_2086),
.B(n_2087),
.C(n_2083),
.Y(n_2655)
);

O2A1O1Ixp33_ASAP7_75t_L g2656 ( 
.A1(n_1810),
.A2(n_1837),
.B(n_1913),
.C(n_1886),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_SL g2657 ( 
.A(n_2214),
.B(n_2215),
.Y(n_2657)
);

AOI22xp5_ASAP7_75t_L g2658 ( 
.A1(n_2166),
.A2(n_2215),
.B1(n_2219),
.B2(n_2214),
.Y(n_2658)
);

AOI21xp5_ASAP7_75t_L g2659 ( 
.A1(n_2185),
.A2(n_2229),
.B(n_2027),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_SL g2660 ( 
.A(n_2215),
.B(n_2219),
.Y(n_2660)
);

O2A1O1Ixp33_ASAP7_75t_SL g2661 ( 
.A1(n_1632),
.A2(n_1642),
.B(n_2098),
.C(n_1749),
.Y(n_2661)
);

AND2x2_ASAP7_75t_L g2662 ( 
.A(n_2086),
.B(n_2087),
.Y(n_2662)
);

OAI22xp5_ASAP7_75t_L g2663 ( 
.A1(n_2219),
.A2(n_2251),
.B1(n_2287),
.B2(n_2247),
.Y(n_2663)
);

NOR2xp33_ASAP7_75t_L g2664 ( 
.A(n_1913),
.B(n_2005),
.Y(n_2664)
);

AOI21xp5_ASAP7_75t_L g2665 ( 
.A1(n_2185),
.A2(n_2229),
.B(n_2027),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_2088),
.B(n_2089),
.Y(n_2666)
);

AOI22xp33_ASAP7_75t_L g2667 ( 
.A1(n_1870),
.A2(n_1842),
.B1(n_1758),
.B2(n_1864),
.Y(n_2667)
);

O2A1O1Ixp33_ASAP7_75t_SL g2668 ( 
.A1(n_1632),
.A2(n_1642),
.B(n_2098),
.C(n_1749),
.Y(n_2668)
);

NOR2xp33_ASAP7_75t_L g2669 ( 
.A(n_2318),
.B(n_1794),
.Y(n_2669)
);

AOI22xp5_ASAP7_75t_L g2670 ( 
.A1(n_2247),
.A2(n_2287),
.B1(n_2313),
.B2(n_2251),
.Y(n_2670)
);

AO32x2_ASAP7_75t_L g2671 ( 
.A1(n_1679),
.A2(n_1958),
.A3(n_1836),
.B1(n_1986),
.B2(n_1936),
.Y(n_2671)
);

A2O1A1Ixp33_ASAP7_75t_L g2672 ( 
.A1(n_2088),
.A2(n_2089),
.B(n_2099),
.C(n_2093),
.Y(n_2672)
);

INVx3_ASAP7_75t_L g2673 ( 
.A(n_1878),
.Y(n_2673)
);

NOR3xp33_ASAP7_75t_L g2674 ( 
.A(n_2144),
.B(n_2188),
.C(n_2170),
.Y(n_2674)
);

INVx3_ASAP7_75t_SL g2675 ( 
.A(n_1727),
.Y(n_2675)
);

OAI22xp5_ASAP7_75t_L g2676 ( 
.A1(n_2247),
.A2(n_2287),
.B1(n_2313),
.B2(n_2251),
.Y(n_2676)
);

A2O1A1Ixp33_ASAP7_75t_L g2677 ( 
.A1(n_2093),
.A2(n_2099),
.B(n_2114),
.C(n_2111),
.Y(n_2677)
);

OAI22xp5_ASAP7_75t_L g2678 ( 
.A1(n_2251),
.A2(n_2287),
.B1(n_2313),
.B2(n_2272),
.Y(n_2678)
);

OAI21x1_ASAP7_75t_L g2679 ( 
.A1(n_1962),
.A2(n_2003),
.B(n_1980),
.Y(n_2679)
);

BUFx3_ASAP7_75t_L g2680 ( 
.A(n_1798),
.Y(n_2680)
);

BUFx6f_ASAP7_75t_L g2681 ( 
.A(n_1631),
.Y(n_2681)
);

O2A1O1Ixp33_ASAP7_75t_L g2682 ( 
.A1(n_2035),
.A2(n_2039),
.B(n_2052),
.C(n_2050),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2267),
.Y(n_2683)
);

BUFx12f_ASAP7_75t_L g2684 ( 
.A(n_2244),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2111),
.B(n_2114),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_SL g2686 ( 
.A(n_2313),
.B(n_2023),
.Y(n_2686)
);

AOI21x1_ASAP7_75t_L g2687 ( 
.A1(n_2034),
.A2(n_2055),
.B(n_2032),
.Y(n_2687)
);

AOI22xp33_ASAP7_75t_L g2688 ( 
.A1(n_1864),
.A2(n_1677),
.B1(n_1690),
.B2(n_1684),
.Y(n_2688)
);

INVxp67_ASAP7_75t_L g2689 ( 
.A(n_1836),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_SL g2690 ( 
.A(n_2023),
.B(n_1738),
.Y(n_2690)
);

OAI22xp5_ASAP7_75t_L g2691 ( 
.A1(n_2272),
.A2(n_1738),
.B1(n_2139),
.B2(n_2138),
.Y(n_2691)
);

AOI21xp5_ASAP7_75t_L g2692 ( 
.A1(n_1633),
.A2(n_1666),
.B(n_1647),
.Y(n_2692)
);

OAI21xp5_ASAP7_75t_L g2693 ( 
.A1(n_2051),
.A2(n_2032),
.B(n_2010),
.Y(n_2693)
);

NOR2xp33_ASAP7_75t_L g2694 ( 
.A(n_1894),
.B(n_1880),
.Y(n_2694)
);

AOI21x1_ASAP7_75t_L g2695 ( 
.A1(n_2051),
.A2(n_2010),
.B(n_2138),
.Y(n_2695)
);

AO21x2_ASAP7_75t_L g2696 ( 
.A1(n_2267),
.A2(n_2273),
.B(n_2271),
.Y(n_2696)
);

OAI22xp5_ASAP7_75t_L g2697 ( 
.A1(n_1738),
.A2(n_2141),
.B1(n_2151),
.B2(n_2139),
.Y(n_2697)
);

AOI21xp5_ASAP7_75t_L g2698 ( 
.A1(n_1633),
.A2(n_1666),
.B(n_1647),
.Y(n_2698)
);

CKINVDCx10_ASAP7_75t_R g2699 ( 
.A(n_2118),
.Y(n_2699)
);

NOR2xp33_ASAP7_75t_L g2700 ( 
.A(n_1894),
.B(n_1880),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_2141),
.B(n_2151),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_2154),
.B(n_2156),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_2271),
.Y(n_2703)
);

HB1xp67_ASAP7_75t_L g2704 ( 
.A(n_2048),
.Y(n_2704)
);

A2O1A1Ixp33_ASAP7_75t_L g2705 ( 
.A1(n_2154),
.A2(n_2156),
.B(n_2163),
.C(n_2158),
.Y(n_2705)
);

AOI22xp33_ASAP7_75t_L g2706 ( 
.A1(n_1864),
.A2(n_1677),
.B1(n_1690),
.B2(n_1684),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2158),
.B(n_2163),
.Y(n_2707)
);

A2O1A1Ixp33_ASAP7_75t_L g2708 ( 
.A1(n_2167),
.A2(n_2168),
.B(n_2196),
.C(n_2172),
.Y(n_2708)
);

BUFx6f_ASAP7_75t_L g2709 ( 
.A(n_1631),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2167),
.B(n_2168),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2172),
.B(n_2196),
.Y(n_2711)
);

OAI21xp5_ASAP7_75t_L g2712 ( 
.A1(n_1846),
.A2(n_2022),
.B(n_2204),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2204),
.B(n_2209),
.Y(n_2713)
);

AO21x1_ASAP7_75t_L g2714 ( 
.A1(n_1677),
.A2(n_1679),
.B(n_2209),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2210),
.B(n_2232),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_L g2716 ( 
.A(n_2210),
.B(n_2232),
.Y(n_2716)
);

OR2x2_ASAP7_75t_L g2717 ( 
.A(n_2271),
.B(n_2273),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_SL g2718 ( 
.A(n_1738),
.B(n_1856),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2233),
.B(n_2234),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_2233),
.B(n_2234),
.Y(n_2720)
);

BUFx3_ASAP7_75t_L g2721 ( 
.A(n_1798),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2236),
.B(n_2237),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2273),
.Y(n_2723)
);

OAI321xp33_ASAP7_75t_L g2724 ( 
.A1(n_1638),
.A2(n_2069),
.A3(n_1672),
.B1(n_2201),
.B2(n_2228),
.C(n_2236),
.Y(n_2724)
);

AOI22xp5_ASAP7_75t_L g2725 ( 
.A1(n_1806),
.A2(n_1871),
.B1(n_1768),
.B2(n_2237),
.Y(n_2725)
);

OAI21xp5_ASAP7_75t_L g2726 ( 
.A1(n_1846),
.A2(n_2022),
.B(n_2242),
.Y(n_2726)
);

O2A1O1Ixp33_ASAP7_75t_L g2727 ( 
.A1(n_2242),
.A2(n_2255),
.B(n_2256),
.C(n_2252),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2291),
.Y(n_2728)
);

A2O1A1Ixp33_ASAP7_75t_L g2729 ( 
.A1(n_2252),
.A2(n_2256),
.B(n_2266),
.C(n_2255),
.Y(n_2729)
);

BUFx8_ASAP7_75t_L g2730 ( 
.A(n_2118),
.Y(n_2730)
);

AND2x4_ASAP7_75t_L g2731 ( 
.A(n_2040),
.B(n_1768),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2266),
.B(n_2270),
.Y(n_2732)
);

INVx2_ASAP7_75t_L g2733 ( 
.A(n_2291),
.Y(n_2733)
);

AOI21x1_ASAP7_75t_L g2734 ( 
.A1(n_2270),
.A2(n_2278),
.B(n_2277),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2291),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2301),
.Y(n_2736)
);

OAI22xp5_ASAP7_75t_L g2737 ( 
.A1(n_2277),
.A2(n_2282),
.B1(n_2289),
.B2(n_2278),
.Y(n_2737)
);

A2O1A1Ixp33_ASAP7_75t_L g2738 ( 
.A1(n_2282),
.A2(n_2305),
.B(n_2309),
.C(n_2289),
.Y(n_2738)
);

O2A1O1Ixp33_ASAP7_75t_SL g2739 ( 
.A1(n_2144),
.A2(n_2170),
.B(n_2194),
.C(n_2188),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2301),
.Y(n_2740)
);

OAI22xp5_ASAP7_75t_L g2741 ( 
.A1(n_2305),
.A2(n_2316),
.B1(n_2309),
.B2(n_1790),
.Y(n_2741)
);

OAI21xp5_ASAP7_75t_L g2742 ( 
.A1(n_1846),
.A2(n_2316),
.B(n_2030),
.Y(n_2742)
);

NOR2xp33_ASAP7_75t_L g2743 ( 
.A(n_1894),
.B(n_1880),
.Y(n_2743)
);

BUFx8_ASAP7_75t_L g2744 ( 
.A(n_2126),
.Y(n_2744)
);

AO32x2_ASAP7_75t_L g2745 ( 
.A1(n_1958),
.A2(n_1986),
.A3(n_1936),
.B1(n_1864),
.B2(n_1769),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_1744),
.B(n_1780),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2301),
.Y(n_2747)
);

HB1xp67_ASAP7_75t_L g2748 ( 
.A(n_2048),
.Y(n_2748)
);

NOR2xp67_ASAP7_75t_L g2749 ( 
.A(n_1900),
.B(n_2043),
.Y(n_2749)
);

AOI22xp33_ASAP7_75t_L g2750 ( 
.A1(n_1864),
.A2(n_1824),
.B1(n_1964),
.B2(n_1947),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2304),
.Y(n_2751)
);

NAND3xp33_ASAP7_75t_L g2752 ( 
.A(n_2053),
.B(n_2048),
.C(n_2244),
.Y(n_2752)
);

NOR2xp33_ASAP7_75t_L g2753 ( 
.A(n_2085),
.B(n_2268),
.Y(n_2753)
);

AOI22xp5_ASAP7_75t_L g2754 ( 
.A1(n_1871),
.A2(n_1768),
.B1(n_1856),
.B2(n_1769),
.Y(n_2754)
);

BUFx8_ASAP7_75t_L g2755 ( 
.A(n_2126),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2304),
.Y(n_2756)
);

CKINVDCx5p33_ASAP7_75t_R g2757 ( 
.A(n_2126),
.Y(n_2757)
);

NOR2xp33_ASAP7_75t_L g2758 ( 
.A(n_1744),
.B(n_1780),
.Y(n_2758)
);

NAND2x1p5_ASAP7_75t_L g2759 ( 
.A(n_2136),
.B(n_2140),
.Y(n_2759)
);

O2A1O1Ixp33_ASAP7_75t_L g2760 ( 
.A1(n_2194),
.A2(n_2319),
.B(n_2207),
.C(n_2243),
.Y(n_2760)
);

AOI22xp33_ASAP7_75t_L g2761 ( 
.A1(n_1691),
.A2(n_1905),
.B1(n_1910),
.B2(n_1906),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_1744),
.B(n_1780),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_1744),
.B(n_1790),
.Y(n_2763)
);

O2A1O1Ixp33_ASAP7_75t_L g2764 ( 
.A1(n_2207),
.A2(n_2319),
.B(n_2243),
.C(n_2269),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_1790),
.B(n_1779),
.Y(n_2765)
);

AOI22xp33_ASAP7_75t_L g2766 ( 
.A1(n_1691),
.A2(n_1905),
.B1(n_1910),
.B2(n_1917),
.Y(n_2766)
);

BUFx6f_ASAP7_75t_L g2767 ( 
.A(n_2136),
.Y(n_2767)
);

AND2x4_ASAP7_75t_L g2768 ( 
.A(n_2040),
.B(n_1768),
.Y(n_2768)
);

AND2x4_ASAP7_75t_L g2769 ( 
.A(n_2040),
.B(n_2041),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_1706),
.Y(n_2770)
);

AO22x1_ASAP7_75t_L g2771 ( 
.A1(n_1871),
.A2(n_2314),
.B1(n_2136),
.B2(n_2140),
.Y(n_2771)
);

BUFx12f_ASAP7_75t_L g2772 ( 
.A(n_2244),
.Y(n_2772)
);

BUFx4f_ASAP7_75t_L g2773 ( 
.A(n_2136),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_1692),
.Y(n_2774)
);

AOI22xp33_ASAP7_75t_SL g2775 ( 
.A1(n_2140),
.A2(n_2187),
.B1(n_2177),
.B2(n_2314),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_SL g2776 ( 
.A(n_1887),
.B(n_2041),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_1779),
.B(n_2203),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_SL g2778 ( 
.A(n_1887),
.B(n_2041),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_1692),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_L g2780 ( 
.A(n_2007),
.B(n_1851),
.Y(n_2780)
);

AOI22xp5_ASAP7_75t_L g2781 ( 
.A1(n_1861),
.A2(n_1909),
.B1(n_1946),
.B2(n_2202),
.Y(n_2781)
);

AND2x2_ASAP7_75t_L g2782 ( 
.A(n_2007),
.B(n_2041),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_1703),
.Y(n_2783)
);

INVx1_ASAP7_75t_SL g2784 ( 
.A(n_1953),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_L g2785 ( 
.A(n_1858),
.B(n_1897),
.Y(n_2785)
);

OAI21xp5_ASAP7_75t_L g2786 ( 
.A1(n_2106),
.A2(n_2148),
.B(n_1887),
.Y(n_2786)
);

INVx4_ASAP7_75t_L g2787 ( 
.A(n_2177),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_SL g2788 ( 
.A(n_1887),
.B(n_1874),
.Y(n_2788)
);

AOI22xp5_ASAP7_75t_L g2789 ( 
.A1(n_2202),
.A2(n_2302),
.B1(n_1773),
.B2(n_1874),
.Y(n_2789)
);

AO21x1_ASAP7_75t_L g2790 ( 
.A1(n_1638),
.A2(n_2069),
.B(n_1672),
.Y(n_2790)
);

AOI22xp5_ASAP7_75t_L g2791 ( 
.A1(n_2302),
.A2(n_1773),
.B1(n_1874),
.B2(n_1671),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_1703),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_1711),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_1897),
.B(n_1711),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_1719),
.B(n_1722),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_SL g2796 ( 
.A(n_1874),
.B(n_2028),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_1719),
.B(n_1722),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_1726),
.B(n_1729),
.Y(n_2798)
);

O2A1O1Ixp33_ASAP7_75t_SL g2799 ( 
.A1(n_2269),
.A2(n_1987),
.B(n_1671),
.C(n_1683),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_1726),
.Y(n_2800)
);

HB1xp67_ASAP7_75t_L g2801 ( 
.A(n_1951),
.Y(n_2801)
);

O2A1O1Ixp33_ASAP7_75t_L g2802 ( 
.A1(n_2004),
.A2(n_2012),
.B(n_2220),
.C(n_2217),
.Y(n_2802)
);

INVx4_ASAP7_75t_L g2803 ( 
.A(n_2187),
.Y(n_2803)
);

INVx3_ASAP7_75t_L g2804 ( 
.A(n_1951),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2053),
.B(n_2004),
.Y(n_2805)
);

INVx1_ASAP7_75t_SL g2806 ( 
.A(n_2004),
.Y(n_2806)
);

OAI22xp5_ASAP7_75t_L g2807 ( 
.A1(n_1728),
.A2(n_2179),
.B1(n_2097),
.B2(n_2285),
.Y(n_2807)
);

O2A1O1Ixp33_ASAP7_75t_SL g2808 ( 
.A1(n_1671),
.A2(n_1708),
.B(n_1721),
.C(n_1683),
.Y(n_2808)
);

HB1xp67_ASAP7_75t_L g2809 ( 
.A(n_1951),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_SL g2810 ( 
.A(n_2028),
.B(n_1936),
.Y(n_2810)
);

OAI22xp5_ASAP7_75t_L g2811 ( 
.A1(n_1728),
.A2(n_2220),
.B1(n_2217),
.B2(n_2285),
.Y(n_2811)
);

BUFx12f_ASAP7_75t_L g2812 ( 
.A(n_2244),
.Y(n_2812)
);

AOI22xp5_ASAP7_75t_L g2813 ( 
.A1(n_1773),
.A2(n_1708),
.B1(n_1721),
.B2(n_1683),
.Y(n_2813)
);

AOI22xp5_ASAP7_75t_L g2814 ( 
.A1(n_1683),
.A2(n_1708),
.B1(n_1721),
.B2(n_1733),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_L g2815 ( 
.A(n_1753),
.B(n_1765),
.Y(n_2815)
);

AND2x2_ASAP7_75t_L g2816 ( 
.A(n_2053),
.B(n_2012),
.Y(n_2816)
);

OAI21xp5_ASAP7_75t_L g2817 ( 
.A1(n_2106),
.A2(n_2148),
.B(n_2026),
.Y(n_2817)
);

BUFx2_ASAP7_75t_L g2818 ( 
.A(n_2053),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_1771),
.B(n_1774),
.Y(n_2819)
);

AOI21xp5_ASAP7_75t_L g2820 ( 
.A1(n_2026),
.A2(n_2000),
.B(n_2012),
.Y(n_2820)
);

AOI21xp5_ASAP7_75t_L g2821 ( 
.A1(n_2026),
.A2(n_2002),
.B(n_1984),
.Y(n_2821)
);

AND2x4_ASAP7_75t_L g2822 ( 
.A(n_2028),
.B(n_1733),
.Y(n_2822)
);

NOR2xp33_ASAP7_75t_L g2823 ( 
.A(n_2296),
.B(n_1728),
.Y(n_2823)
);

AOI21x1_ASAP7_75t_L g2824 ( 
.A1(n_1778),
.A2(n_1965),
.B(n_1942),
.Y(n_2824)
);

O2A1O1Ixp33_ASAP7_75t_L g2825 ( 
.A1(n_2097),
.A2(n_2220),
.B(n_2179),
.C(n_2285),
.Y(n_2825)
);

NAND2x1p5_ASAP7_75t_L g2826 ( 
.A(n_1733),
.B(n_2028),
.Y(n_2826)
);

NOR2xp33_ASAP7_75t_L g2827 ( 
.A(n_2296),
.B(n_2097),
.Y(n_2827)
);

AOI22xp5_ASAP7_75t_L g2828 ( 
.A1(n_1686),
.A2(n_1693),
.B1(n_1783),
.B2(n_2296),
.Y(n_2828)
);

OAI22xp5_ASAP7_75t_L g2829 ( 
.A1(n_2179),
.A2(n_2217),
.B1(n_1937),
.B2(n_1902),
.Y(n_2829)
);

AOI21x1_ASAP7_75t_L g2830 ( 
.A1(n_1799),
.A2(n_1890),
.B(n_1971),
.Y(n_2830)
);

AOI21xp5_ASAP7_75t_L g2831 ( 
.A1(n_1970),
.A2(n_1973),
.B(n_1984),
.Y(n_2831)
);

OR2x6_ASAP7_75t_L g2832 ( 
.A(n_1638),
.B(n_1672),
.Y(n_2832)
);

OAI22xp5_ASAP7_75t_L g2833 ( 
.A1(n_1902),
.A2(n_1937),
.B1(n_2228),
.B2(n_2201),
.Y(n_2833)
);

BUFx3_ASAP7_75t_L g2834 ( 
.A(n_1829),
.Y(n_2834)
);

NOR2xp33_ASAP7_75t_L g2835 ( 
.A(n_2296),
.B(n_1801),
.Y(n_2835)
);

BUFx12f_ASAP7_75t_L g2836 ( 
.A(n_1829),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_L g2837 ( 
.A(n_1808),
.B(n_1812),
.Y(n_2837)
);

A2O1A1Ixp33_ASAP7_75t_SL g2838 ( 
.A1(n_1801),
.A2(n_1830),
.B(n_1828),
.C(n_1717),
.Y(n_2838)
);

NOR2xp33_ASAP7_75t_L g2839 ( 
.A(n_1801),
.B(n_1828),
.Y(n_2839)
);

AOI21xp5_ASAP7_75t_L g2840 ( 
.A1(n_1970),
.A2(n_1973),
.B(n_1984),
.Y(n_2840)
);

NAND3xp33_ASAP7_75t_L g2841 ( 
.A(n_2053),
.B(n_1860),
.C(n_1829),
.Y(n_2841)
);

OAI22xp5_ASAP7_75t_L g2842 ( 
.A1(n_2069),
.A2(n_2201),
.B1(n_2228),
.B2(n_1686),
.Y(n_2842)
);

AND2x2_ASAP7_75t_L g2843 ( 
.A(n_2053),
.B(n_1812),
.Y(n_2843)
);

BUFx4f_ASAP7_75t_L g2844 ( 
.A(n_1686),
.Y(n_2844)
);

AOI22xp5_ASAP7_75t_L g2845 ( 
.A1(n_1686),
.A2(n_1693),
.B1(n_1783),
.B2(n_1920),
.Y(n_2845)
);

NOR2xp33_ASAP7_75t_L g2846 ( 
.A(n_1801),
.B(n_1828),
.Y(n_2846)
);

AOI221xp5_ASAP7_75t_L g2847 ( 
.A1(n_1889),
.A2(n_2001),
.B1(n_1995),
.B2(n_1989),
.C(n_1976),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_1717),
.Y(n_2848)
);

OAI21xp5_ASAP7_75t_L g2849 ( 
.A1(n_1828),
.A2(n_1830),
.B(n_1911),
.Y(n_2849)
);

CKINVDCx20_ASAP7_75t_R g2850 ( 
.A(n_1968),
.Y(n_2850)
);

CKINVDCx20_ASAP7_75t_R g2851 ( 
.A(n_1968),
.Y(n_2851)
);

AOI22xp5_ASAP7_75t_L g2852 ( 
.A1(n_1686),
.A2(n_1693),
.B1(n_1783),
.B2(n_1920),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_1813),
.B(n_1815),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_1815),
.B(n_1820),
.Y(n_2854)
);

AOI21xp5_ASAP7_75t_L g2855 ( 
.A1(n_1970),
.A2(n_2002),
.B(n_1984),
.Y(n_2855)
);

AND2x2_ASAP7_75t_SL g2856 ( 
.A(n_1693),
.B(n_1783),
.Y(n_2856)
);

NOR2xp67_ASAP7_75t_L g2857 ( 
.A(n_1830),
.B(n_1970),
.Y(n_2857)
);

AND2x2_ASAP7_75t_L g2858 ( 
.A(n_1820),
.B(n_1824),
.Y(n_2858)
);

AOI21xp5_ASAP7_75t_L g2859 ( 
.A1(n_1970),
.A2(n_2002),
.B(n_1973),
.Y(n_2859)
);

INVx1_ASAP7_75t_SL g2860 ( 
.A(n_1973),
.Y(n_2860)
);

AOI21x1_ASAP7_75t_L g2861 ( 
.A1(n_1825),
.A2(n_1906),
.B(n_1995),
.Y(n_2861)
);

NOR2x1p5_ASAP7_75t_SL g2862 ( 
.A(n_1720),
.B(n_1731),
.Y(n_2862)
);

INVx2_ASAP7_75t_L g2863 ( 
.A(n_1720),
.Y(n_2863)
);

NOR2xp33_ASAP7_75t_R g2864 ( 
.A(n_1830),
.B(n_1968),
.Y(n_2864)
);

AOI21xp5_ASAP7_75t_L g2865 ( 
.A1(n_1860),
.A2(n_1862),
.B(n_1920),
.Y(n_2865)
);

OAI21xp5_ASAP7_75t_L g2866 ( 
.A1(n_1934),
.A2(n_1940),
.B(n_1976),
.Y(n_2866)
);

BUFx6f_ASAP7_75t_L g2867 ( 
.A(n_1693),
.Y(n_2867)
);

AOI21xp5_ASAP7_75t_L g2868 ( 
.A1(n_1862),
.A2(n_1693),
.B(n_1783),
.Y(n_2868)
);

BUFx4f_ASAP7_75t_L g2869 ( 
.A(n_1783),
.Y(n_2869)
);

AO21x1_ASAP7_75t_L g2870 ( 
.A1(n_1825),
.A2(n_1989),
.B(n_1975),
.Y(n_2870)
);

CKINVDCx11_ASAP7_75t_R g2871 ( 
.A(n_1862),
.Y(n_2871)
);

INVx3_ASAP7_75t_L g2872 ( 
.A(n_1969),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_1826),
.B(n_1966),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_SL g2874 ( 
.A(n_1969),
.B(n_1929),
.Y(n_2874)
);

INVx5_ASAP7_75t_L g2875 ( 
.A(n_1747),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_SL g2876 ( 
.A(n_1827),
.B(n_1926),
.Y(n_2876)
);

OAI22xp5_ASAP7_75t_L g2877 ( 
.A1(n_1835),
.A2(n_1965),
.B1(n_1964),
.B2(n_1947),
.Y(n_2877)
);

INVx1_ASAP7_75t_SL g2878 ( 
.A(n_1835),
.Y(n_2878)
);

INVxp67_ASAP7_75t_L g2879 ( 
.A(n_1865),
.Y(n_2879)
);

BUFx6f_ASAP7_75t_L g2880 ( 
.A(n_1770),
.Y(n_2880)
);

AOI33xp33_ASAP7_75t_L g2881 ( 
.A1(n_1866),
.A2(n_1926),
.A3(n_1943),
.B1(n_1942),
.B2(n_1941),
.B3(n_1869),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_SL g2882 ( 
.A(n_1866),
.B(n_1943),
.Y(n_2882)
);

NOR2xp33_ASAP7_75t_L g2883 ( 
.A(n_1869),
.B(n_1919),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_1917),
.Y(n_2884)
);

NAND2x1p5_ASAP7_75t_L g2885 ( 
.A(n_1919),
.B(n_1772),
.Y(n_2885)
);

NOR2xp67_ASAP7_75t_SL g2886 ( 
.A(n_1781),
.B(n_1792),
.Y(n_2886)
);

NOR3xp33_ASAP7_75t_L g2887 ( 
.A(n_1792),
.B(n_1805),
.C(n_1811),
.Y(n_2887)
);

OAI22xp5_ASAP7_75t_L g2888 ( 
.A1(n_1805),
.A2(n_1811),
.B1(n_1817),
.B2(n_1821),
.Y(n_2888)
);

NOR3xp33_ASAP7_75t_L g2889 ( 
.A(n_1805),
.B(n_1811),
.C(n_1817),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2009),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_L g2891 ( 
.A(n_1817),
.B(n_1821),
.Y(n_2891)
);

OAI22xp5_ASAP7_75t_L g2892 ( 
.A1(n_1823),
.A2(n_1831),
.B1(n_1855),
.B2(n_1863),
.Y(n_2892)
);

BUFx2_ASAP7_75t_L g2893 ( 
.A(n_1823),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_1831),
.B(n_1855),
.Y(n_2894)
);

BUFx3_ASAP7_75t_L g2895 ( 
.A(n_1855),
.Y(n_2895)
);

BUFx3_ASAP7_75t_L g2896 ( 
.A(n_1863),
.Y(n_2896)
);

BUFx6f_ASAP7_75t_L g2897 ( 
.A(n_1877),
.Y(n_2897)
);

NOR2xp33_ASAP7_75t_L g2898 ( 
.A(n_1916),
.B(n_1918),
.Y(n_2898)
);

AND2x2_ASAP7_75t_L g2899 ( 
.A(n_1922),
.B(n_1923),
.Y(n_2899)
);

A2O1A1Ixp33_ASAP7_75t_L g2900 ( 
.A1(n_1924),
.A2(n_1935),
.B(n_1950),
.C(n_1956),
.Y(n_2900)
);

A2O1A1Ixp33_ASAP7_75t_L g2901 ( 
.A1(n_1960),
.A2(n_1967),
.B(n_1985),
.C(n_2009),
.Y(n_2901)
);

AND2x2_ASAP7_75t_L g2902 ( 
.A(n_1960),
.B(n_1967),
.Y(n_2902)
);

AOI21xp5_ASAP7_75t_L g2903 ( 
.A1(n_1960),
.A2(n_1967),
.B(n_1985),
.Y(n_2903)
);

INVx3_ASAP7_75t_L g2904 ( 
.A(n_1985),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_1658),
.B(n_1660),
.Y(n_2905)
);

OAI21xp5_ASAP7_75t_L g2906 ( 
.A1(n_2211),
.A2(n_1107),
.B(n_1437),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_1645),
.Y(n_2907)
);

INVxp67_ASAP7_75t_SL g2908 ( 
.A(n_2286),
.Y(n_2908)
);

A2O1A1Ixp33_ASAP7_75t_L g2909 ( 
.A1(n_2211),
.A2(n_1552),
.B(n_1492),
.C(n_1107),
.Y(n_2909)
);

AND2x4_ASAP7_75t_L g2910 ( 
.A(n_2068),
.B(n_1625),
.Y(n_2910)
);

OAI22xp5_ASAP7_75t_L g2911 ( 
.A1(n_1615),
.A2(n_2102),
.B1(n_2124),
.B2(n_2094),
.Y(n_2911)
);

AND2x2_ASAP7_75t_SL g2912 ( 
.A(n_1627),
.B(n_2070),
.Y(n_2912)
);

AOI21xp5_ASAP7_75t_L g2913 ( 
.A1(n_2058),
.A2(n_1107),
.B(n_2117),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_1658),
.B(n_1660),
.Y(n_2914)
);

NOR2xp33_ASAP7_75t_L g2915 ( 
.A(n_1636),
.B(n_1639),
.Y(n_2915)
);

AOI21xp5_ASAP7_75t_L g2916 ( 
.A1(n_2058),
.A2(n_1107),
.B(n_2117),
.Y(n_2916)
);

O2A1O1Ixp33_ASAP7_75t_L g2917 ( 
.A1(n_2212),
.A2(n_1107),
.B(n_1439),
.C(n_1437),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_1658),
.B(n_1660),
.Y(n_2918)
);

NOR2xp33_ASAP7_75t_L g2919 ( 
.A(n_1636),
.B(n_1639),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_SL g2920 ( 
.A(n_2076),
.B(n_1107),
.Y(n_2920)
);

NOR2x1_ASAP7_75t_L g2921 ( 
.A(n_1651),
.B(n_1832),
.Y(n_2921)
);

AOI21xp5_ASAP7_75t_L g2922 ( 
.A1(n_2058),
.A2(n_1107),
.B(n_2117),
.Y(n_2922)
);

AOI21x1_ASAP7_75t_L g2923 ( 
.A1(n_1673),
.A2(n_1932),
.B(n_1101),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_1645),
.Y(n_2924)
);

NAND2xp5_ASAP7_75t_SL g2925 ( 
.A(n_2076),
.B(n_1107),
.Y(n_2925)
);

CKINVDCx10_ASAP7_75t_R g2926 ( 
.A(n_2180),
.Y(n_2926)
);

AND2x4_ASAP7_75t_L g2927 ( 
.A(n_2068),
.B(n_1625),
.Y(n_2927)
);

AOI33xp33_ASAP7_75t_L g2928 ( 
.A1(n_2212),
.A2(n_2257),
.A3(n_762),
.B1(n_1552),
.B2(n_1492),
.B3(n_2211),
.Y(n_2928)
);

AOI21x1_ASAP7_75t_L g2929 ( 
.A1(n_1673),
.A2(n_1932),
.B(n_1101),
.Y(n_2929)
);

A2O1A1Ixp33_ASAP7_75t_L g2930 ( 
.A1(n_2211),
.A2(n_1552),
.B(n_1492),
.C(n_1107),
.Y(n_2930)
);

NAND3xp33_ASAP7_75t_L g2931 ( 
.A(n_2211),
.B(n_1107),
.C(n_1437),
.Y(n_2931)
);

AOI22xp5_ASAP7_75t_L g2932 ( 
.A1(n_2079),
.A2(n_1568),
.B1(n_1437),
.B2(n_1439),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_SL g2933 ( 
.A(n_2076),
.B(n_1107),
.Y(n_2933)
);

INVx2_ASAP7_75t_L g2934 ( 
.A(n_1645),
.Y(n_2934)
);

CKINVDCx5p33_ASAP7_75t_R g2935 ( 
.A(n_2071),
.Y(n_2935)
);

OAI21x1_ASAP7_75t_L g2936 ( 
.A1(n_1932),
.A2(n_1673),
.B(n_1895),
.Y(n_2936)
);

AOI22xp5_ASAP7_75t_L g2937 ( 
.A1(n_2079),
.A2(n_1568),
.B1(n_1437),
.B2(n_1439),
.Y(n_2937)
);

AOI21xp5_ASAP7_75t_L g2938 ( 
.A1(n_2058),
.A2(n_1107),
.B(n_2117),
.Y(n_2938)
);

AOI21xp5_ASAP7_75t_L g2939 ( 
.A1(n_2058),
.A2(n_1107),
.B(n_2117),
.Y(n_2939)
);

AOI21xp5_ASAP7_75t_L g2940 ( 
.A1(n_2058),
.A2(n_1107),
.B(n_2117),
.Y(n_2940)
);

NOR2xp67_ASAP7_75t_L g2941 ( 
.A(n_1635),
.B(n_2062),
.Y(n_2941)
);

AOI21xp5_ASAP7_75t_L g2942 ( 
.A1(n_2058),
.A2(n_1107),
.B(n_2117),
.Y(n_2942)
);

OAI22xp5_ASAP7_75t_L g2943 ( 
.A1(n_1615),
.A2(n_2102),
.B1(n_2124),
.B2(n_2094),
.Y(n_2943)
);

AOI21xp5_ASAP7_75t_L g2944 ( 
.A1(n_2058),
.A2(n_1107),
.B(n_2117),
.Y(n_2944)
);

NAND2xp5_ASAP7_75t_L g2945 ( 
.A(n_1658),
.B(n_1660),
.Y(n_2945)
);

OA21x2_ASAP7_75t_L g2946 ( 
.A1(n_1673),
.A2(n_1932),
.B(n_1701),
.Y(n_2946)
);

AND2x2_ASAP7_75t_L g2947 ( 
.A(n_2143),
.B(n_2068),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_1658),
.B(n_1660),
.Y(n_2948)
);

AOI22xp5_ASAP7_75t_L g2949 ( 
.A1(n_2079),
.A2(n_1568),
.B1(n_1437),
.B2(n_1439),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_L g2950 ( 
.A(n_1658),
.B(n_1660),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_L g2951 ( 
.A(n_1658),
.B(n_1660),
.Y(n_2951)
);

AND2x4_ASAP7_75t_L g2952 ( 
.A(n_2068),
.B(n_1625),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_L g2953 ( 
.A(n_1658),
.B(n_1660),
.Y(n_2953)
);

OAI21xp5_ASAP7_75t_L g2954 ( 
.A1(n_2211),
.A2(n_1107),
.B(n_1437),
.Y(n_2954)
);

INVx2_ASAP7_75t_L g2955 ( 
.A(n_1645),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_1658),
.B(n_1660),
.Y(n_2956)
);

BUFx12f_ASAP7_75t_L g2957 ( 
.A(n_2180),
.Y(n_2957)
);

AOI22xp33_ASAP7_75t_L g2958 ( 
.A1(n_2079),
.A2(n_1568),
.B1(n_1414),
.B2(n_1534),
.Y(n_2958)
);

A2O1A1Ixp33_ASAP7_75t_SL g2959 ( 
.A1(n_2084),
.A2(n_757),
.B(n_1461),
.C(n_1407),
.Y(n_2959)
);

OAI21xp5_ASAP7_75t_L g2960 ( 
.A1(n_2211),
.A2(n_1107),
.B(n_1437),
.Y(n_2960)
);

OAI21x1_ASAP7_75t_L g2961 ( 
.A1(n_1932),
.A2(n_1673),
.B(n_1895),
.Y(n_2961)
);

AOI21xp5_ASAP7_75t_L g2962 ( 
.A1(n_2058),
.A2(n_1107),
.B(n_2117),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_L g2963 ( 
.A(n_1658),
.B(n_1660),
.Y(n_2963)
);

O2A1O1Ixp5_ASAP7_75t_L g2964 ( 
.A1(n_2092),
.A2(n_1107),
.B(n_1439),
.C(n_1437),
.Y(n_2964)
);

A2O1A1Ixp33_ASAP7_75t_L g2965 ( 
.A1(n_2211),
.A2(n_1552),
.B(n_1492),
.C(n_1107),
.Y(n_2965)
);

AOI22xp5_ASAP7_75t_L g2966 ( 
.A1(n_2079),
.A2(n_1568),
.B1(n_1437),
.B2(n_1439),
.Y(n_2966)
);

AND2x2_ASAP7_75t_SL g2967 ( 
.A(n_1627),
.B(n_2070),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_L g2968 ( 
.A(n_1658),
.B(n_1660),
.Y(n_2968)
);

NAND2xp5_ASAP7_75t_L g2969 ( 
.A(n_1658),
.B(n_1660),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_1645),
.Y(n_2970)
);

AOI21xp5_ASAP7_75t_L g2971 ( 
.A1(n_2058),
.A2(n_1107),
.B(n_2117),
.Y(n_2971)
);

NOR3xp33_ASAP7_75t_L g2972 ( 
.A(n_2112),
.B(n_1539),
.C(n_1453),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_1658),
.B(n_1660),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_1658),
.B(n_1660),
.Y(n_2974)
);

AOI21xp5_ASAP7_75t_L g2975 ( 
.A1(n_2058),
.A2(n_1107),
.B(n_2117),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_L g2976 ( 
.A(n_1658),
.B(n_1660),
.Y(n_2976)
);

NAND2xp33_ASAP7_75t_SL g2977 ( 
.A(n_2129),
.B(n_1437),
.Y(n_2977)
);

BUFx6f_ASAP7_75t_L g2978 ( 
.A(n_1623),
.Y(n_2978)
);

CKINVDCx16_ASAP7_75t_R g2979 ( 
.A(n_2071),
.Y(n_2979)
);

AOI21xp5_ASAP7_75t_L g2980 ( 
.A1(n_2058),
.A2(n_1107),
.B(n_2117),
.Y(n_2980)
);

NAND2x1p5_ASAP7_75t_L g2981 ( 
.A(n_1627),
.B(n_2070),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_1645),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_SL g2983 ( 
.A(n_2076),
.B(n_1107),
.Y(n_2983)
);

OR2x2_ASAP7_75t_L g2984 ( 
.A(n_1682),
.B(n_1640),
.Y(n_2984)
);

AOI21xp5_ASAP7_75t_L g2985 ( 
.A1(n_2058),
.A2(n_1107),
.B(n_2117),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_L g2986 ( 
.A(n_1618),
.B(n_1685),
.Y(n_2986)
);

BUFx4f_ASAP7_75t_L g2987 ( 
.A(n_1623),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_L g2988 ( 
.A(n_1618),
.B(n_1685),
.Y(n_2988)
);

INVx2_ASAP7_75t_L g2989 ( 
.A(n_1645),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_1645),
.Y(n_2990)
);

INVx3_ASAP7_75t_L g2991 ( 
.A(n_2584),
.Y(n_2991)
);

NOR2x1_ASAP7_75t_SL g2992 ( 
.A(n_2579),
.B(n_2591),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_SL g2993 ( 
.A(n_2390),
.B(n_2321),
.Y(n_2993)
);

AND2x4_ASAP7_75t_L g2994 ( 
.A(n_2603),
.B(n_2769),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_SL g2995 ( 
.A(n_2321),
.B(n_2399),
.Y(n_2995)
);

OAI21xp5_ASAP7_75t_L g2996 ( 
.A1(n_2400),
.A2(n_2369),
.B(n_2350),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2351),
.B(n_2357),
.Y(n_2997)
);

NOR2x1_ASAP7_75t_SL g2998 ( 
.A(n_2579),
.B(n_2591),
.Y(n_2998)
);

AOI22xp5_ASAP7_75t_L g2999 ( 
.A1(n_2388),
.A2(n_2937),
.B1(n_2949),
.B2(n_2932),
.Y(n_2999)
);

AOI21xp5_ASAP7_75t_L g3000 ( 
.A1(n_2350),
.A2(n_2917),
.B(n_2386),
.Y(n_3000)
);

AOI21xp5_ASAP7_75t_L g3001 ( 
.A1(n_2913),
.A2(n_2922),
.B(n_2916),
.Y(n_3001)
);

BUFx6f_ASAP7_75t_L g3002 ( 
.A(n_2912),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3003)
);

AOI21xp33_ASAP7_75t_L g3004 ( 
.A1(n_2428),
.A2(n_2442),
.B(n_2932),
.Y(n_3004)
);

CKINVDCx5p33_ASAP7_75t_R g3005 ( 
.A(n_2322),
.Y(n_3005)
);

AND2x2_ASAP7_75t_L g3006 ( 
.A(n_2480),
.B(n_2514),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2986),
.B(n_2988),
.Y(n_3007)
);

AOI21xp5_ASAP7_75t_L g3008 ( 
.A1(n_2938),
.A2(n_2940),
.B(n_2939),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2986),
.B(n_2988),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2397),
.B(n_2592),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_2592),
.B(n_2456),
.Y(n_3011)
);

OAI21x1_ASAP7_75t_L g3012 ( 
.A1(n_2923),
.A2(n_2929),
.B(n_2416),
.Y(n_3012)
);

OAI22xp5_ASAP7_75t_L g3013 ( 
.A1(n_2937),
.A2(n_2949),
.B1(n_2966),
.B2(n_2388),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_2456),
.B(n_2415),
.Y(n_3014)
);

A2O1A1Ixp33_ASAP7_75t_L g3015 ( 
.A1(n_2462),
.A2(n_2966),
.B(n_2964),
.C(n_2399),
.Y(n_3015)
);

OAI21xp5_ASAP7_75t_L g3016 ( 
.A1(n_2400),
.A2(n_2370),
.B(n_2375),
.Y(n_3016)
);

AO21x1_ASAP7_75t_L g3017 ( 
.A1(n_2428),
.A2(n_2442),
.B(n_2920),
.Y(n_3017)
);

AND2x2_ASAP7_75t_L g3018 ( 
.A(n_2480),
.B(n_2514),
.Y(n_3018)
);

INVx5_ASAP7_75t_L g3019 ( 
.A(n_2579),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_L g3020 ( 
.A(n_2419),
.B(n_2427),
.Y(n_3020)
);

OAI21xp5_ASAP7_75t_L g3021 ( 
.A1(n_2370),
.A2(n_2375),
.B(n_2931),
.Y(n_3021)
);

OA22x2_ASAP7_75t_L g3022 ( 
.A1(n_2498),
.A2(n_2538),
.B1(n_2523),
.B2(n_2452),
.Y(n_3022)
);

OAI21xp5_ASAP7_75t_L g3023 ( 
.A1(n_2931),
.A2(n_2346),
.B(n_2344),
.Y(n_3023)
);

AOI22xp5_ASAP7_75t_L g3024 ( 
.A1(n_2958),
.A2(n_2340),
.B1(n_2933),
.B2(n_2925),
.Y(n_3024)
);

AOI21xp5_ASAP7_75t_L g3025 ( 
.A1(n_2942),
.A2(n_2962),
.B(n_2944),
.Y(n_3025)
);

AO31x2_ASAP7_75t_L g3026 ( 
.A1(n_2714),
.A2(n_2352),
.A3(n_2911),
.B(n_2342),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_2908),
.B(n_2457),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2460),
.B(n_2467),
.Y(n_3028)
);

OR2x2_ASAP7_75t_L g3029 ( 
.A(n_2450),
.B(n_2385),
.Y(n_3029)
);

INVx2_ASAP7_75t_L g3030 ( 
.A(n_2696),
.Y(n_3030)
);

AO31x2_ASAP7_75t_L g3031 ( 
.A1(n_2714),
.A2(n_2352),
.A3(n_2911),
.B(n_2342),
.Y(n_3031)
);

OAI21x1_ASAP7_75t_SL g3032 ( 
.A1(n_2346),
.A2(n_2954),
.B(n_2906),
.Y(n_3032)
);

AOI21xp33_ASAP7_75t_L g3033 ( 
.A1(n_2403),
.A2(n_2954),
.B(n_2906),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_L g3034 ( 
.A(n_2468),
.B(n_2470),
.Y(n_3034)
);

INVx1_ASAP7_75t_SL g3035 ( 
.A(n_2577),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2475),
.B(n_2476),
.Y(n_3036)
);

AOI21x1_ASAP7_75t_L g3037 ( 
.A1(n_2354),
.A2(n_2339),
.B(n_2687),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_L g3038 ( 
.A(n_2379),
.B(n_2380),
.Y(n_3038)
);

OAI21x1_ASAP7_75t_L g3039 ( 
.A1(n_2529),
.A2(n_2698),
.B(n_2692),
.Y(n_3039)
);

AOI21xp5_ASAP7_75t_L g3040 ( 
.A1(n_2971),
.A2(n_2980),
.B(n_2975),
.Y(n_3040)
);

AOI21xp5_ASAP7_75t_L g3041 ( 
.A1(n_2985),
.A2(n_2334),
.B(n_2960),
.Y(n_3041)
);

NAND3xp33_ASAP7_75t_L g3042 ( 
.A(n_2330),
.B(n_2919),
.C(n_2915),
.Y(n_3042)
);

AND2x4_ASAP7_75t_L g3043 ( 
.A(n_2603),
.B(n_2769),
.Y(n_3043)
);

INVx5_ASAP7_75t_L g3044 ( 
.A(n_2579),
.Y(n_3044)
);

O2A1O1Ixp5_ASAP7_75t_L g3045 ( 
.A1(n_2960),
.A2(n_2983),
.B(n_2930),
.C(n_2965),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_L g3046 ( 
.A(n_2493),
.B(n_2360),
.Y(n_3046)
);

AND2x2_ASAP7_75t_L g3047 ( 
.A(n_2326),
.B(n_2947),
.Y(n_3047)
);

AND2x2_ASAP7_75t_L g3048 ( 
.A(n_2326),
.B(n_2947),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2695),
.Y(n_3049)
);

O2A1O1Ixp5_ASAP7_75t_L g3050 ( 
.A1(n_2909),
.A2(n_2338),
.B(n_2436),
.C(n_2354),
.Y(n_3050)
);

XNOR2xp5_ASAP7_75t_L g3051 ( 
.A(n_2523),
.B(n_2642),
.Y(n_3051)
);

OAI21xp5_ASAP7_75t_L g3052 ( 
.A1(n_2332),
.A2(n_2403),
.B(n_2348),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_2425),
.B(n_2424),
.Y(n_3053)
);

OAI21xp33_ASAP7_75t_SL g3054 ( 
.A1(n_2928),
.A2(n_2371),
.B(n_2345),
.Y(n_3054)
);

AOI221xp5_ASAP7_75t_SL g3055 ( 
.A1(n_2341),
.A2(n_2359),
.B1(n_2358),
.B2(n_2338),
.C(n_2407),
.Y(n_3055)
);

AOI21xp5_ASAP7_75t_L g3056 ( 
.A1(n_2430),
.A2(n_2495),
.B(n_2943),
.Y(n_3056)
);

OAI21xp5_ASAP7_75t_L g3057 ( 
.A1(n_2349),
.A2(n_2972),
.B(n_2444),
.Y(n_3057)
);

BUFx2_ASAP7_75t_L g3058 ( 
.A(n_2448),
.Y(n_3058)
);

A2O1A1Ixp33_ASAP7_75t_L g3059 ( 
.A1(n_2441),
.A2(n_2977),
.B(n_2452),
.C(n_2436),
.Y(n_3059)
);

OAI21xp5_ASAP7_75t_L g3060 ( 
.A1(n_2943),
.A2(n_2440),
.B(n_2959),
.Y(n_3060)
);

AO31x2_ASAP7_75t_L g3061 ( 
.A1(n_2870),
.A2(n_2888),
.A3(n_2892),
.B(n_2877),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_2611),
.B(n_2443),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2329),
.Y(n_3063)
);

INVx2_ASAP7_75t_L g3064 ( 
.A(n_2696),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_L g3065 ( 
.A(n_2611),
.B(n_2443),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_2549),
.B(n_2537),
.Y(n_3066)
);

INVx1_ASAP7_75t_SL g3067 ( 
.A(n_2577),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_2549),
.B(n_2537),
.Y(n_3068)
);

NAND2xp33_ASAP7_75t_L g3069 ( 
.A(n_2542),
.B(n_2612),
.Y(n_3069)
);

OAI21x1_ASAP7_75t_SL g3070 ( 
.A1(n_2392),
.A2(n_2569),
.B(n_2432),
.Y(n_3070)
);

NOR2x1_ASAP7_75t_L g3071 ( 
.A(n_2412),
.B(n_2921),
.Y(n_3071)
);

AO31x2_ASAP7_75t_L g3072 ( 
.A1(n_2870),
.A2(n_2888),
.A3(n_2892),
.B(n_2877),
.Y(n_3072)
);

NOR4xp25_ASAP7_75t_L g3073 ( 
.A(n_2440),
.B(n_2485),
.C(n_2590),
.D(n_2404),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_L g3074 ( 
.A(n_2458),
.B(n_2479),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_L g3075 ( 
.A(n_2458),
.B(n_2479),
.Y(n_3075)
);

AOI21x1_ASAP7_75t_L g3076 ( 
.A1(n_2687),
.A2(n_2505),
.B(n_2414),
.Y(n_3076)
);

OAI21x1_ASAP7_75t_L g3077 ( 
.A1(n_2526),
.A2(n_2679),
.B(n_2821),
.Y(n_3077)
);

AOI21xp5_ASAP7_75t_L g3078 ( 
.A1(n_2946),
.A2(n_2484),
.B(n_2396),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2329),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_2551),
.B(n_2552),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2551),
.B(n_2552),
.Y(n_3081)
);

OA21x2_ASAP7_75t_L g3082 ( 
.A1(n_2404),
.A2(n_2482),
.B(n_2599),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2337),
.Y(n_3083)
);

AOI21x1_ASAP7_75t_L g3084 ( 
.A1(n_2414),
.A2(n_2840),
.B(n_2831),
.Y(n_3084)
);

AOI21x1_ASAP7_75t_L g3085 ( 
.A1(n_2855),
.A2(n_2859),
.B(n_2868),
.Y(n_3085)
);

NAND2x1p5_ASAP7_75t_L g3086 ( 
.A(n_2497),
.B(n_2426),
.Y(n_3086)
);

AOI21xp5_ASAP7_75t_L g3087 ( 
.A1(n_2628),
.A2(n_2808),
.B(n_2431),
.Y(n_3087)
);

NOR2xp33_ASAP7_75t_L g3088 ( 
.A(n_2410),
.B(n_2378),
.Y(n_3088)
);

BUFx2_ASAP7_75t_L g3089 ( 
.A(n_2448),
.Y(n_3089)
);

BUFx2_ASAP7_75t_SL g3090 ( 
.A(n_2331),
.Y(n_3090)
);

AOI21xp5_ASAP7_75t_L g3091 ( 
.A1(n_2628),
.A2(n_2585),
.B(n_2447),
.Y(n_3091)
);

AOI21xp5_ASAP7_75t_L g3092 ( 
.A1(n_2435),
.A2(n_2439),
.B(n_2368),
.Y(n_3092)
);

BUFx6f_ASAP7_75t_L g3093 ( 
.A(n_2912),
.Y(n_3093)
);

AND2x2_ASAP7_75t_L g3094 ( 
.A(n_2639),
.B(n_2662),
.Y(n_3094)
);

OAI21xp5_ASAP7_75t_L g3095 ( 
.A1(n_2422),
.A2(n_2535),
.B(n_2451),
.Y(n_3095)
);

BUFx6f_ASAP7_75t_L g3096 ( 
.A(n_2967),
.Y(n_3096)
);

O2A1O1Ixp5_ASAP7_75t_L g3097 ( 
.A1(n_2365),
.A2(n_2366),
.B(n_2422),
.C(n_2829),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_2556),
.B(n_2568),
.Y(n_3098)
);

NOR2xp33_ASAP7_75t_L g3099 ( 
.A(n_2463),
.B(n_2372),
.Y(n_3099)
);

AOI21xp33_ASAP7_75t_L g3100 ( 
.A1(n_2485),
.A2(n_2445),
.B(n_2371),
.Y(n_3100)
);

NAND2xp5_ASAP7_75t_L g3101 ( 
.A(n_2556),
.B(n_2568),
.Y(n_3101)
);

AOI22xp5_ASAP7_75t_L g3102 ( 
.A1(n_2345),
.A2(n_2445),
.B1(n_2367),
.B2(n_2401),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2624),
.B(n_2627),
.Y(n_3103)
);

BUFx6f_ASAP7_75t_L g3104 ( 
.A(n_2967),
.Y(n_3104)
);

OAI21x1_ASAP7_75t_SL g3105 ( 
.A1(n_2802),
.A2(n_2563),
.B(n_2825),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_2633),
.B(n_2634),
.Y(n_3106)
);

A2O1A1Ixp33_ASAP7_75t_L g3107 ( 
.A1(n_2548),
.A2(n_2487),
.B(n_2401),
.C(n_2535),
.Y(n_3107)
);

NOR2xp33_ASAP7_75t_L g3108 ( 
.A(n_2411),
.B(n_2935),
.Y(n_3108)
);

AOI21xp5_ASAP7_75t_L g3109 ( 
.A1(n_2838),
.A2(n_2820),
.B(n_2585),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_2373),
.Y(n_3110)
);

AND2x2_ASAP7_75t_L g3111 ( 
.A(n_2639),
.B(n_2662),
.Y(n_3111)
);

INVxp67_ASAP7_75t_L g3112 ( 
.A(n_2502),
.Y(n_3112)
);

AOI21xp5_ASAP7_75t_SL g3113 ( 
.A1(n_2500),
.A2(n_2511),
.B(n_2663),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_2575),
.B(n_2595),
.Y(n_3114)
);

AND2x4_ASAP7_75t_L g3115 ( 
.A(n_2769),
.B(n_2584),
.Y(n_3115)
);

AOI21xp33_ASAP7_75t_L g3116 ( 
.A1(n_2566),
.A2(n_2572),
.B(n_2562),
.Y(n_3116)
);

OAI21x1_ASAP7_75t_L g3117 ( 
.A1(n_2648),
.A2(n_2665),
.B(n_2659),
.Y(n_3117)
);

OAI21xp5_ASAP7_75t_L g3118 ( 
.A1(n_2566),
.A2(n_2921),
.B(n_2412),
.Y(n_3118)
);

AOI21xp5_ASAP7_75t_L g3119 ( 
.A1(n_2616),
.A2(n_2806),
.B(n_2454),
.Y(n_3119)
);

OR2x6_ASAP7_75t_L g3120 ( 
.A(n_2602),
.B(n_2574),
.Y(n_3120)
);

AOI21x1_ASAP7_75t_L g3121 ( 
.A1(n_2362),
.A2(n_2865),
.B(n_2586),
.Y(n_3121)
);

INVx2_ASAP7_75t_SL g3122 ( 
.A(n_2704),
.Y(n_3122)
);

AOI21xp5_ASAP7_75t_L g3123 ( 
.A1(n_2806),
.A2(n_2461),
.B(n_2417),
.Y(n_3123)
);

NOR2xp33_ASAP7_75t_L g3124 ( 
.A(n_2411),
.B(n_2935),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_L g3125 ( 
.A(n_2608),
.B(n_2421),
.Y(n_3125)
);

OAI22xp5_ASAP7_75t_L g3126 ( 
.A1(n_2429),
.A2(n_2446),
.B1(n_2464),
.B2(n_2433),
.Y(n_3126)
);

INVx2_ASAP7_75t_L g3127 ( 
.A(n_2377),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_2465),
.B(n_2477),
.Y(n_3128)
);

AOI21xp5_ASAP7_75t_L g3129 ( 
.A1(n_2473),
.A2(n_2483),
.B(n_2474),
.Y(n_3129)
);

AOI21xp5_ASAP7_75t_L g3130 ( 
.A1(n_2582),
.A2(n_2583),
.B(n_2841),
.Y(n_3130)
);

OAI21xp5_ASAP7_75t_L g3131 ( 
.A1(n_2599),
.A2(n_2614),
.B(n_2520),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_L g3132 ( 
.A(n_2478),
.B(n_2609),
.Y(n_3132)
);

OR2x6_ASAP7_75t_L g3133 ( 
.A(n_2602),
.B(n_2574),
.Y(n_3133)
);

AOI21x1_ASAP7_75t_L g3134 ( 
.A1(n_2586),
.A2(n_2811),
.B(n_2807),
.Y(n_3134)
);

OAI21xp33_ASAP7_75t_L g3135 ( 
.A1(n_2488),
.A2(n_2546),
.B(n_2562),
.Y(n_3135)
);

BUFx4f_ASAP7_75t_SL g3136 ( 
.A(n_2957),
.Y(n_3136)
);

NOR2x1_ASAP7_75t_L g3137 ( 
.A(n_2614),
.B(n_2752),
.Y(n_3137)
);

A2O1A1Ixp33_ASAP7_75t_L g3138 ( 
.A1(n_2626),
.A2(n_2509),
.B(n_2572),
.C(n_2538),
.Y(n_3138)
);

NOR2xp33_ASAP7_75t_L g3139 ( 
.A(n_2364),
.B(n_2979),
.Y(n_3139)
);

OAI21x1_ASAP7_75t_L g3140 ( 
.A1(n_2817),
.A2(n_2644),
.B(n_2641),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_SL g3141 ( 
.A(n_2829),
.B(n_2725),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_2546),
.B(n_2333),
.Y(n_3142)
);

AND2x2_ASAP7_75t_L g3143 ( 
.A(n_2543),
.B(n_2593),
.Y(n_3143)
);

NAND2x1p5_ASAP7_75t_L g3144 ( 
.A(n_2497),
.B(n_2426),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2337),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_L g3146 ( 
.A(n_2343),
.B(n_2347),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2355),
.Y(n_3147)
);

INVx2_ASAP7_75t_L g3148 ( 
.A(n_2377),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_SL g3149 ( 
.A(n_2725),
.B(n_2570),
.Y(n_3149)
);

OAI21x1_ASAP7_75t_L g3150 ( 
.A1(n_2826),
.A2(n_2842),
.B(n_2734),
.Y(n_3150)
);

CKINVDCx20_ASAP7_75t_R g3151 ( 
.A(n_2979),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2355),
.Y(n_3152)
);

OAI22xp5_ASAP7_75t_L g3153 ( 
.A1(n_2573),
.A2(n_2658),
.B1(n_2517),
.B2(n_2522),
.Y(n_3153)
);

OAI22xp5_ASAP7_75t_L g3154 ( 
.A1(n_2573),
.A2(n_2658),
.B1(n_2508),
.B2(n_2544),
.Y(n_3154)
);

BUFx2_ASAP7_75t_L g3155 ( 
.A(n_2745),
.Y(n_3155)
);

AOI21x1_ASAP7_75t_L g3156 ( 
.A1(n_2807),
.A2(n_2811),
.B(n_2857),
.Y(n_3156)
);

A2O1A1Ixp33_ASAP7_75t_L g3157 ( 
.A1(n_2667),
.A2(n_2623),
.B(n_2691),
.C(n_2561),
.Y(n_3157)
);

AND3x2_ASAP7_75t_L g3158 ( 
.A(n_2564),
.B(n_2700),
.C(n_2694),
.Y(n_3158)
);

AOI21xp5_ASAP7_75t_L g3159 ( 
.A1(n_2712),
.A2(n_2726),
.B(n_2625),
.Y(n_3159)
);

AND2x2_ASAP7_75t_L g3160 ( 
.A(n_2543),
.B(n_2593),
.Y(n_3160)
);

AOI21x1_ASAP7_75t_L g3161 ( 
.A1(n_2857),
.A2(n_2749),
.B(n_2771),
.Y(n_3161)
);

INVx5_ASAP7_75t_L g3162 ( 
.A(n_2591),
.Y(n_3162)
);

INVx2_ASAP7_75t_L g3163 ( 
.A(n_2391),
.Y(n_3163)
);

NAND2x1p5_ASAP7_75t_L g3164 ( 
.A(n_2497),
.B(n_2426),
.Y(n_3164)
);

AOI21x1_ASAP7_75t_L g3165 ( 
.A1(n_2749),
.A2(n_2771),
.B(n_2810),
.Y(n_3165)
);

NAND2x1_ASAP7_75t_L g3166 ( 
.A(n_2814),
.B(n_2539),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2391),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_2374),
.B(n_2376),
.Y(n_3168)
);

OAI21x1_ASAP7_75t_L g3169 ( 
.A1(n_2824),
.A2(n_2861),
.B(n_2830),
.Y(n_3169)
);

AOI22xp33_ASAP7_75t_L g3170 ( 
.A1(n_2784),
.A2(n_2596),
.B1(n_2455),
.B2(n_2794),
.Y(n_3170)
);

INVxp67_ASAP7_75t_SL g3171 ( 
.A(n_2571),
.Y(n_3171)
);

AOI21xp5_ASAP7_75t_L g3172 ( 
.A1(n_2712),
.A2(n_2726),
.B(n_2724),
.Y(n_3172)
);

OAI22xp5_ASAP7_75t_L g3173 ( 
.A1(n_2544),
.A2(n_2450),
.B1(n_2984),
.B2(n_2385),
.Y(n_3173)
);

BUFx2_ASAP7_75t_L g3174 ( 
.A(n_2745),
.Y(n_3174)
);

OAI21xp5_ASAP7_75t_L g3175 ( 
.A1(n_2741),
.A2(n_2682),
.B(n_2653),
.Y(n_3175)
);

BUFx8_ASAP7_75t_SL g3176 ( 
.A(n_2957),
.Y(n_3176)
);

AND2x2_ASAP7_75t_L g3177 ( 
.A(n_2984),
.B(n_2613),
.Y(n_3177)
);

AO31x2_ASAP7_75t_L g3178 ( 
.A1(n_2790),
.A2(n_2741),
.A3(n_2901),
.B(n_2900),
.Y(n_3178)
);

OR2x2_ASAP7_75t_L g3179 ( 
.A(n_2389),
.B(n_2571),
.Y(n_3179)
);

OAI21x1_ASAP7_75t_L g3180 ( 
.A1(n_2824),
.A2(n_2861),
.B(n_2830),
.Y(n_3180)
);

OR2x2_ASAP7_75t_L g3181 ( 
.A(n_2389),
.B(n_2604),
.Y(n_3181)
);

AND2x2_ASAP7_75t_L g3182 ( 
.A(n_2613),
.B(n_2782),
.Y(n_3182)
);

INVx1_ASAP7_75t_SL g3183 ( 
.A(n_2587),
.Y(n_3183)
);

A2O1A1Ixp33_ASAP7_75t_L g3184 ( 
.A1(n_2691),
.A2(n_2784),
.B(n_2498),
.C(n_2689),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_SL g3185 ( 
.A(n_2833),
.B(n_2791),
.Y(n_3185)
);

AOI21xp5_ASAP7_75t_L g3186 ( 
.A1(n_2724),
.A2(n_2668),
.B(n_2661),
.Y(n_3186)
);

OR2x6_ASAP7_75t_L g3187 ( 
.A(n_2574),
.B(n_2501),
.Y(n_3187)
);

A2O1A1Ixp33_ASAP7_75t_L g3188 ( 
.A1(n_2381),
.A2(n_2413),
.B(n_2387),
.C(n_2418),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_2638),
.B(n_2640),
.Y(n_3189)
);

OAI22xp5_ASAP7_75t_L g3190 ( 
.A1(n_2670),
.A2(n_2527),
.B1(n_2449),
.B2(n_2499),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2393),
.Y(n_3191)
);

AOI21xp5_ASAP7_75t_L g3192 ( 
.A1(n_2739),
.A2(n_2676),
.B(n_2663),
.Y(n_3192)
);

OAI21x1_ASAP7_75t_L g3193 ( 
.A1(n_2619),
.A2(n_2759),
.B(n_2814),
.Y(n_3193)
);

INVx1_ASAP7_75t_SL g3194 ( 
.A(n_2871),
.Y(n_3194)
);

AOI21x1_ASAP7_75t_L g3195 ( 
.A1(n_2886),
.A2(n_2941),
.B(n_2809),
.Y(n_3195)
);

OAI21x1_ASAP7_75t_L g3196 ( 
.A1(n_2619),
.A2(n_2849),
.B(n_2813),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_2393),
.Y(n_3197)
);

OAI21x1_ASAP7_75t_L g3198 ( 
.A1(n_2619),
.A2(n_2849),
.B(n_2813),
.Y(n_3198)
);

INVxp67_ASAP7_75t_SL g3199 ( 
.A(n_2885),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_2402),
.Y(n_3200)
);

OAI21xp5_ASAP7_75t_L g3201 ( 
.A1(n_2525),
.A2(n_2697),
.B(n_2545),
.Y(n_3201)
);

AOI21xp5_ASAP7_75t_L g3202 ( 
.A1(n_2676),
.A2(n_2799),
.B(n_2967),
.Y(n_3202)
);

A2O1A1Ixp33_ASAP7_75t_L g3203 ( 
.A1(n_2833),
.A2(n_2328),
.B(n_2914),
.C(n_2905),
.Y(n_3203)
);

OAI22xp33_ASAP7_75t_L g3204 ( 
.A1(n_2675),
.A2(n_2754),
.B1(n_2670),
.B2(n_2596),
.Y(n_3204)
);

A2O1A1Ixp33_ASAP7_75t_L g3205 ( 
.A1(n_2918),
.A2(n_2945),
.B(n_2950),
.C(n_2948),
.Y(n_3205)
);

NOR2xp33_ASAP7_75t_L g3206 ( 
.A(n_2664),
.B(n_2635),
.Y(n_3206)
);

INVxp67_ASAP7_75t_L g3207 ( 
.A(n_2324),
.Y(n_3207)
);

INVx1_ASAP7_75t_SL g3208 ( 
.A(n_2818),
.Y(n_3208)
);

AND2x2_ASAP7_75t_L g3209 ( 
.A(n_2782),
.B(n_2805),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_SL g3210 ( 
.A(n_2791),
.B(n_2754),
.Y(n_3210)
);

NOR2xp33_ASAP7_75t_SL g3211 ( 
.A(n_2497),
.B(n_2361),
.Y(n_3211)
);

OR2x2_ASAP7_75t_L g3212 ( 
.A(n_2389),
.B(n_2580),
.Y(n_3212)
);

OR2x6_ASAP7_75t_L g3213 ( 
.A(n_2574),
.B(n_2501),
.Y(n_3213)
);

INVx3_ASAP7_75t_L g3214 ( 
.A(n_2336),
.Y(n_3214)
);

A2O1A1Ixp33_ASAP7_75t_L g3215 ( 
.A1(n_2951),
.A2(n_2953),
.B(n_2963),
.C(n_2956),
.Y(n_3215)
);

OAI22xp5_ASAP7_75t_L g3216 ( 
.A1(n_2438),
.A2(n_2518),
.B1(n_2617),
.B2(n_2605),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_2402),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_2597),
.B(n_2601),
.Y(n_3218)
);

OAI21x1_ASAP7_75t_L g3219 ( 
.A1(n_2941),
.A2(n_2503),
.B(n_2466),
.Y(n_3219)
);

OAI22xp5_ASAP7_75t_L g3220 ( 
.A1(n_2654),
.A2(n_2675),
.B1(n_2513),
.B2(n_2789),
.Y(n_3220)
);

OA22x2_ASAP7_75t_L g3221 ( 
.A1(n_2675),
.A2(n_2654),
.B1(n_2678),
.B2(n_2501),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_2737),
.B(n_2651),
.Y(n_3222)
);

OAI21xp5_ASAP7_75t_L g3223 ( 
.A1(n_2697),
.A2(n_2594),
.B(n_2656),
.Y(n_3223)
);

OAI21xp33_ASAP7_75t_L g3224 ( 
.A1(n_2596),
.A2(n_2969),
.B(n_2968),
.Y(n_3224)
);

INVx3_ASAP7_75t_L g3225 ( 
.A(n_2466),
.Y(n_3225)
);

OAI21x1_ASAP7_75t_L g3226 ( 
.A1(n_2466),
.A2(n_2524),
.B(n_2503),
.Y(n_3226)
);

AO31x2_ASAP7_75t_L g3227 ( 
.A1(n_2790),
.A2(n_2737),
.A3(n_2893),
.B(n_2898),
.Y(n_3227)
);

OAI21x1_ASAP7_75t_L g3228 ( 
.A1(n_2503),
.A2(n_2600),
.B(n_2524),
.Y(n_3228)
);

OAI21x1_ASAP7_75t_L g3229 ( 
.A1(n_2524),
.A2(n_2673),
.B(n_2600),
.Y(n_3229)
);

OAI21xp5_ASAP7_75t_L g3230 ( 
.A1(n_2594),
.A2(n_2491),
.B(n_2490),
.Y(n_3230)
);

BUFx3_ASAP7_75t_L g3231 ( 
.A(n_2818),
.Y(n_3231)
);

NAND2xp5_ASAP7_75t_L g3232 ( 
.A(n_2655),
.B(n_2672),
.Y(n_3232)
);

OAI21x1_ASAP7_75t_L g3233 ( 
.A1(n_2600),
.A2(n_2804),
.B(n_2673),
.Y(n_3233)
);

AOI21xp5_ASAP7_75t_L g3234 ( 
.A1(n_2507),
.A2(n_2987),
.B(n_2773),
.Y(n_3234)
);

AOI21xp5_ASAP7_75t_L g3235 ( 
.A1(n_2507),
.A2(n_2987),
.B(n_2773),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_2406),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_2677),
.B(n_2705),
.Y(n_3237)
);

AOI21xp5_ASAP7_75t_L g3238 ( 
.A1(n_2507),
.A2(n_2987),
.B(n_2773),
.Y(n_3238)
);

AND2x2_ASAP7_75t_L g3239 ( 
.A(n_2805),
.B(n_2816),
.Y(n_3239)
);

AO31x2_ASAP7_75t_L g3240 ( 
.A1(n_2893),
.A2(n_2395),
.A3(n_2453),
.B(n_2405),
.Y(n_3240)
);

AOI21xp5_ASAP7_75t_L g3241 ( 
.A1(n_2844),
.A2(n_2869),
.B(n_2742),
.Y(n_3241)
);

OAI21xp5_ASAP7_75t_L g3242 ( 
.A1(n_2496),
.A2(n_2510),
.B(n_2504),
.Y(n_3242)
);

AOI21xp5_ASAP7_75t_L g3243 ( 
.A1(n_2844),
.A2(n_2869),
.B(n_2742),
.Y(n_3243)
);

BUFx2_ASAP7_75t_L g3244 ( 
.A(n_2745),
.Y(n_3244)
);

OAI21xp5_ASAP7_75t_L g3245 ( 
.A1(n_2630),
.A2(n_2974),
.B(n_2973),
.Y(n_3245)
);

AOI21x1_ASAP7_75t_L g3246 ( 
.A1(n_2801),
.A2(n_2796),
.B(n_2690),
.Y(n_3246)
);

NOR2xp33_ASAP7_75t_L g3247 ( 
.A(n_2643),
.B(n_2753),
.Y(n_3247)
);

AOI21xp33_ASAP7_75t_L g3248 ( 
.A1(n_2335),
.A2(n_2727),
.B(n_2636),
.Y(n_3248)
);

AOI22xp33_ASAP7_75t_L g3249 ( 
.A1(n_2501),
.A2(n_2506),
.B1(n_2706),
.B2(n_2688),
.Y(n_3249)
);

AOI21xp5_ASAP7_75t_SL g3250 ( 
.A1(n_2981),
.A2(n_2591),
.B(n_2678),
.Y(n_3250)
);

A2O1A1Ixp33_ASAP7_75t_L g3251 ( 
.A1(n_2976),
.A2(n_2785),
.B(n_2459),
.C(n_2789),
.Y(n_3251)
);

BUFx2_ASAP7_75t_L g3252 ( 
.A(n_2745),
.Y(n_3252)
);

AOI21xp5_ASAP7_75t_L g3253 ( 
.A1(n_2844),
.A2(n_2869),
.B(n_2788),
.Y(n_3253)
);

AOI21xp5_ASAP7_75t_L g3254 ( 
.A1(n_2532),
.A2(n_2555),
.B(n_2554),
.Y(n_3254)
);

AND2x4_ASAP7_75t_L g3255 ( 
.A(n_2731),
.B(n_2768),
.Y(n_3255)
);

INVx2_ASAP7_75t_SL g3256 ( 
.A(n_2748),
.Y(n_3256)
);

BUFx2_ASAP7_75t_SL g3257 ( 
.A(n_2426),
.Y(n_3257)
);

AOI21xp5_ASAP7_75t_L g3258 ( 
.A1(n_2560),
.A2(n_2615),
.B(n_2567),
.Y(n_3258)
);

OAI21xp5_ASAP7_75t_L g3259 ( 
.A1(n_2693),
.A2(n_2621),
.B(n_2708),
.Y(n_3259)
);

AOI21xp5_ASAP7_75t_L g3260 ( 
.A1(n_2657),
.A2(n_2660),
.B(n_2686),
.Y(n_3260)
);

A2O1A1Ixp33_ASAP7_75t_L g3261 ( 
.A1(n_2780),
.A2(n_2752),
.B(n_2610),
.C(n_2743),
.Y(n_3261)
);

AOI21xp5_ASAP7_75t_L g3262 ( 
.A1(n_2472),
.A2(n_2550),
.B(n_2536),
.Y(n_3262)
);

AND2x4_ASAP7_75t_L g3263 ( 
.A(n_2731),
.B(n_2768),
.Y(n_3263)
);

AOI21xp5_ASAP7_75t_L g3264 ( 
.A1(n_2550),
.A2(n_2649),
.B(n_2860),
.Y(n_3264)
);

INVx3_ASAP7_75t_L g3265 ( 
.A(n_2804),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_L g3266 ( 
.A(n_2729),
.B(n_2738),
.Y(n_3266)
);

INVxp67_ASAP7_75t_SL g3267 ( 
.A(n_2885),
.Y(n_3267)
);

INVx4_ASAP7_75t_L g3268 ( 
.A(n_2426),
.Y(n_3268)
);

AOI21xp5_ASAP7_75t_L g3269 ( 
.A1(n_2875),
.A2(n_2764),
.B(n_2760),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_2406),
.Y(n_3270)
);

NAND2xp5_ASAP7_75t_L g3271 ( 
.A(n_2701),
.B(n_2702),
.Y(n_3271)
);

NAND2xp5_ASAP7_75t_L g3272 ( 
.A(n_2701),
.B(n_2702),
.Y(n_3272)
);

NAND2xp5_ASAP7_75t_L g3273 ( 
.A(n_2707),
.B(n_2710),
.Y(n_3273)
);

CKINVDCx6p67_ASAP7_75t_R g3274 ( 
.A(n_2322),
.Y(n_3274)
);

AND2x2_ASAP7_75t_L g3275 ( 
.A(n_2816),
.B(n_2843),
.Y(n_3275)
);

AOI21x1_ASAP7_75t_L g3276 ( 
.A1(n_2822),
.A2(n_2777),
.B(n_2765),
.Y(n_3276)
);

BUFx6f_ASAP7_75t_L g3277 ( 
.A(n_2327),
.Y(n_3277)
);

AOI21xp5_ASAP7_75t_L g3278 ( 
.A1(n_2875),
.A2(n_2786),
.B(n_2778),
.Y(n_3278)
);

OAI21xp5_ASAP7_75t_L g3279 ( 
.A1(n_2693),
.A2(n_2647),
.B(n_2674),
.Y(n_3279)
);

A2O1A1Ixp33_ASAP7_75t_L g3280 ( 
.A1(n_2835),
.A2(n_2828),
.B(n_2629),
.C(n_2862),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_2707),
.B(n_2710),
.Y(n_3281)
);

INVxp67_ASAP7_75t_SL g3282 ( 
.A(n_2904),
.Y(n_3282)
);

INVx2_ASAP7_75t_SL g3283 ( 
.A(n_2834),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_2408),
.Y(n_3284)
);

NAND2xp5_ASAP7_75t_L g3285 ( 
.A(n_2645),
.B(n_2650),
.Y(n_3285)
);

OAI21xp5_ASAP7_75t_L g3286 ( 
.A1(n_2828),
.A2(n_2666),
.B(n_2652),
.Y(n_3286)
);

AOI21x1_ASAP7_75t_L g3287 ( 
.A1(n_2822),
.A2(n_2882),
.B(n_2876),
.Y(n_3287)
);

OAI21xp5_ASAP7_75t_L g3288 ( 
.A1(n_2685),
.A2(n_2713),
.B(n_2711),
.Y(n_3288)
);

AOI22xp5_ASAP7_75t_L g3289 ( 
.A1(n_2618),
.A2(n_2718),
.B1(n_2776),
.B2(n_2758),
.Y(n_3289)
);

INVx1_ASAP7_75t_SL g3290 ( 
.A(n_2864),
.Y(n_3290)
);

AO31x2_ASAP7_75t_L g3291 ( 
.A1(n_2395),
.A2(n_2453),
.A3(n_2469),
.B(n_2405),
.Y(n_3291)
);

INVx2_ASAP7_75t_L g3292 ( 
.A(n_2469),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_2715),
.B(n_2716),
.Y(n_3293)
);

INVx2_ASAP7_75t_L g3294 ( 
.A(n_2494),
.Y(n_3294)
);

AND2x4_ASAP7_75t_L g3295 ( 
.A(n_2731),
.B(n_2768),
.Y(n_3295)
);

AOI21xp5_ASAP7_75t_L g3296 ( 
.A1(n_2574),
.A2(n_2878),
.B(n_2832),
.Y(n_3296)
);

CKINVDCx5p33_ASAP7_75t_R g3297 ( 
.A(n_2926),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_L g3298 ( 
.A(n_2719),
.B(n_2720),
.Y(n_3298)
);

AOI21xp5_ASAP7_75t_L g3299 ( 
.A1(n_2832),
.A2(n_2335),
.B(n_2383),
.Y(n_3299)
);

AND2x2_ASAP7_75t_L g3300 ( 
.A(n_2843),
.B(n_2731),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_L g3301 ( 
.A(n_2722),
.B(n_2732),
.Y(n_3301)
);

INVx5_ASAP7_75t_L g3302 ( 
.A(n_2832),
.Y(n_3302)
);

AOI21xp5_ASAP7_75t_L g3303 ( 
.A1(n_2547),
.A2(n_2846),
.B(n_2839),
.Y(n_3303)
);

INVx2_ASAP7_75t_L g3304 ( 
.A(n_2494),
.Y(n_3304)
);

INVx2_ASAP7_75t_L g3305 ( 
.A(n_2515),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_2408),
.Y(n_3306)
);

AO221x2_ASAP7_75t_L g3307 ( 
.A1(n_2671),
.A2(n_2745),
.B1(n_2382),
.B2(n_2501),
.C(n_2763),
.Y(n_3307)
);

AND2x2_ASAP7_75t_L g3308 ( 
.A(n_2768),
.B(n_2389),
.Y(n_3308)
);

OAI21xp5_ASAP7_75t_L g3309 ( 
.A1(n_2847),
.A2(n_2879),
.B(n_2866),
.Y(n_3309)
);

OAI21xp5_ASAP7_75t_L g3310 ( 
.A1(n_2866),
.A2(n_2852),
.B(n_2845),
.Y(n_3310)
);

AO31x2_ASAP7_75t_L g3311 ( 
.A1(n_2515),
.A2(n_2733),
.A3(n_2598),
.B(n_2989),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_2774),
.B(n_2779),
.Y(n_3312)
);

OAI21xp5_ASAP7_75t_L g3313 ( 
.A1(n_2845),
.A2(n_2852),
.B(n_2827),
.Y(n_3313)
);

INVx2_ASAP7_75t_L g3314 ( 
.A(n_2531),
.Y(n_3314)
);

AOI221xp5_ASAP7_75t_L g3315 ( 
.A1(n_2530),
.A2(n_2540),
.B1(n_2622),
.B2(n_2750),
.C(n_2823),
.Y(n_3315)
);

CKINVDCx20_ASAP7_75t_R g3316 ( 
.A(n_2646),
.Y(n_3316)
);

AND2x2_ASAP7_75t_L g3317 ( 
.A(n_2389),
.B(n_2323),
.Y(n_3317)
);

OR2x2_ASAP7_75t_L g3318 ( 
.A(n_2580),
.B(n_2588),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_L g3319 ( 
.A(n_2774),
.B(n_2779),
.Y(n_3319)
);

OAI21x1_ASAP7_75t_L g3320 ( 
.A1(n_2903),
.A2(n_2872),
.B(n_2837),
.Y(n_3320)
);

AOI21xp5_ASAP7_75t_L g3321 ( 
.A1(n_2547),
.A2(n_2553),
.B(n_2856),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_2783),
.B(n_2792),
.Y(n_3322)
);

AOI21xp5_ASAP7_75t_L g3323 ( 
.A1(n_2553),
.A2(n_2856),
.B(n_2887),
.Y(n_3323)
);

AND2x2_ASAP7_75t_L g3324 ( 
.A(n_2323),
.B(n_2910),
.Y(n_3324)
);

AOI21xp5_ASAP7_75t_L g3325 ( 
.A1(n_2553),
.A2(n_2856),
.B(n_2889),
.Y(n_3325)
);

AOI21xp5_ASAP7_75t_L g3326 ( 
.A1(n_2553),
.A2(n_2822),
.B(n_2356),
.Y(n_3326)
);

NAND2xp5_ASAP7_75t_L g3327 ( 
.A(n_2783),
.B(n_2792),
.Y(n_3327)
);

OAI21x1_ASAP7_75t_L g3328 ( 
.A1(n_2872),
.A2(n_2837),
.B(n_2797),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_SL g3329 ( 
.A(n_2867),
.B(n_2382),
.Y(n_3329)
);

INVx2_ASAP7_75t_L g3330 ( 
.A(n_2531),
.Y(n_3330)
);

OAI21x1_ASAP7_75t_L g3331 ( 
.A1(n_2872),
.A2(n_2853),
.B(n_2797),
.Y(n_3331)
);

INVx3_ASAP7_75t_L g3332 ( 
.A(n_2822),
.Y(n_3332)
);

INVx2_ASAP7_75t_L g3333 ( 
.A(n_2533),
.Y(n_3333)
);

OR2x6_ASAP7_75t_L g3334 ( 
.A(n_2519),
.B(n_2862),
.Y(n_3334)
);

BUFx10_ASAP7_75t_L g3335 ( 
.A(n_2867),
.Y(n_3335)
);

OAI21x1_ASAP7_75t_L g3336 ( 
.A1(n_2854),
.A2(n_2873),
.B(n_2904),
.Y(n_3336)
);

AND2x4_ASAP7_75t_L g3337 ( 
.A(n_2323),
.B(n_2910),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_2434),
.Y(n_3338)
);

OAI21x1_ASAP7_75t_L g3339 ( 
.A1(n_2904),
.A2(n_2800),
.B(n_2793),
.Y(n_3339)
);

HB1xp67_ASAP7_75t_L g3340 ( 
.A(n_2588),
.Y(n_3340)
);

CKINVDCx8_ASAP7_75t_R g3341 ( 
.A(n_2926),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_SL g3342 ( 
.A(n_2867),
.B(n_2383),
.Y(n_3342)
);

OAI21xp5_ASAP7_75t_L g3343 ( 
.A1(n_2883),
.A2(n_2874),
.B(n_2781),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_2434),
.Y(n_3344)
);

AND2x4_ASAP7_75t_L g3345 ( 
.A(n_2323),
.B(n_2910),
.Y(n_3345)
);

NOR2xp33_ASAP7_75t_L g3346 ( 
.A(n_2669),
.B(n_2512),
.Y(n_3346)
);

OAI21x1_ASAP7_75t_L g3347 ( 
.A1(n_2884),
.A2(n_2798),
.B(n_2795),
.Y(n_3347)
);

AOI21xp5_ASAP7_75t_L g3348 ( 
.A1(n_2383),
.A2(n_2541),
.B(n_2486),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_2884),
.B(n_2858),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_2437),
.Y(n_3350)
);

BUFx2_ASAP7_75t_L g3351 ( 
.A(n_2671),
.Y(n_3351)
);

AOI21xp33_ASAP7_75t_L g3352 ( 
.A1(n_2361),
.A2(n_2819),
.B(n_2815),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_L g3353 ( 
.A(n_2858),
.B(n_2881),
.Y(n_3353)
);

INVx2_ASAP7_75t_L g3354 ( 
.A(n_2533),
.Y(n_3354)
);

A2O1A1Ixp33_ASAP7_75t_L g3355 ( 
.A1(n_2781),
.A2(n_2952),
.B(n_2927),
.C(n_2910),
.Y(n_3355)
);

AND2x4_ASAP7_75t_L g3356 ( 
.A(n_2927),
.B(n_2952),
.Y(n_3356)
);

AND2x2_ASAP7_75t_L g3357 ( 
.A(n_2927),
.B(n_2952),
.Y(n_3357)
);

NOR2xp33_ASAP7_75t_L g3358 ( 
.A(n_2512),
.B(n_2757),
.Y(n_3358)
);

AND2x2_ASAP7_75t_L g3359 ( 
.A(n_2927),
.B(n_2952),
.Y(n_3359)
);

AND2x2_ASAP7_75t_L g3360 ( 
.A(n_2353),
.B(n_2394),
.Y(n_3360)
);

AOI21xp5_ASAP7_75t_L g3361 ( 
.A1(n_2553),
.A2(n_2327),
.B(n_2978),
.Y(n_3361)
);

NOR2xp33_ASAP7_75t_L g3362 ( 
.A(n_2757),
.B(n_2699),
.Y(n_3362)
);

AOI211x1_ASAP7_75t_L g3363 ( 
.A1(n_2746),
.A2(n_2762),
.B(n_2990),
.C(n_2728),
.Y(n_3363)
);

AOI21x1_ASAP7_75t_L g3364 ( 
.A1(n_2891),
.A2(n_2894),
.B(n_2890),
.Y(n_3364)
);

INVx2_ASAP7_75t_L g3365 ( 
.A(n_2559),
.Y(n_3365)
);

INVx3_ASAP7_75t_SL g3366 ( 
.A(n_2867),
.Y(n_3366)
);

INVx2_ASAP7_75t_SL g3367 ( 
.A(n_2353),
.Y(n_3367)
);

AOI21xp5_ASAP7_75t_L g3368 ( 
.A1(n_2383),
.A2(n_2541),
.B(n_2486),
.Y(n_3368)
);

OAI21xp5_ASAP7_75t_L g3369 ( 
.A1(n_2761),
.A2(n_2766),
.B(n_2924),
.Y(n_3369)
);

AOI21xp5_ASAP7_75t_L g3370 ( 
.A1(n_2486),
.A2(n_2541),
.B(n_2775),
.Y(n_3370)
);

AO31x2_ASAP7_75t_L g3371 ( 
.A1(n_2559),
.A2(n_2989),
.A3(n_2982),
.B(n_2970),
.Y(n_3371)
);

AO31x2_ASAP7_75t_L g3372 ( 
.A1(n_2578),
.A2(n_2982),
.A3(n_2970),
.B(n_2955),
.Y(n_3372)
);

AND2x2_ASAP7_75t_L g3373 ( 
.A(n_2394),
.B(n_2680),
.Y(n_3373)
);

AOI21x1_ASAP7_75t_L g3374 ( 
.A1(n_2489),
.A2(n_2747),
.B(n_2751),
.Y(n_3374)
);

AND2x2_ASAP7_75t_L g3375 ( 
.A(n_2680),
.B(n_2721),
.Y(n_3375)
);

AO31x2_ASAP7_75t_L g3376 ( 
.A1(n_2578),
.A2(n_2955),
.A3(n_2934),
.B(n_2736),
.Y(n_3376)
);

OAI21x1_ASAP7_75t_L g3377 ( 
.A1(n_2516),
.A2(n_2589),
.B(n_2924),
.Y(n_3377)
);

OAI21x1_ASAP7_75t_L g3378 ( 
.A1(n_2516),
.A2(n_2723),
.B(n_2735),
.Y(n_3378)
);

NOR2xp67_ASAP7_75t_L g3379 ( 
.A(n_2607),
.B(n_2717),
.Y(n_3379)
);

AND2x2_ASAP7_75t_L g3380 ( 
.A(n_2680),
.B(n_2721),
.Y(n_3380)
);

OAI21x1_ASAP7_75t_L g3381 ( 
.A1(n_2534),
.A2(n_2589),
.B(n_2907),
.Y(n_3381)
);

INVx2_ASAP7_75t_L g3382 ( 
.A(n_2581),
.Y(n_3382)
);

AOI21xp5_ASAP7_75t_L g3383 ( 
.A1(n_2486),
.A2(n_2541),
.B(n_2721),
.Y(n_3383)
);

BUFx3_ASAP7_75t_L g3384 ( 
.A(n_2361),
.Y(n_3384)
);

CKINVDCx5p33_ASAP7_75t_R g3385 ( 
.A(n_2699),
.Y(n_3385)
);

OAI21x1_ASAP7_75t_L g3386 ( 
.A1(n_2558),
.A2(n_2606),
.B(n_2907),
.Y(n_3386)
);

BUFx3_ASAP7_75t_L g3387 ( 
.A(n_2361),
.Y(n_3387)
);

BUFx6f_ASAP7_75t_L g3388 ( 
.A(n_2356),
.Y(n_3388)
);

HB1xp67_ASAP7_75t_L g3389 ( 
.A(n_2607),
.Y(n_3389)
);

HB1xp67_ASAP7_75t_L g3390 ( 
.A(n_2717),
.Y(n_3390)
);

INVxp67_ASAP7_75t_SL g3391 ( 
.A(n_2895),
.Y(n_3391)
);

BUFx2_ASAP7_75t_L g3392 ( 
.A(n_2671),
.Y(n_3392)
);

INVx1_ASAP7_75t_SL g3393 ( 
.A(n_2836),
.Y(n_3393)
);

OAI21x1_ASAP7_75t_L g3394 ( 
.A1(n_2576),
.A2(n_2740),
.B(n_2751),
.Y(n_3394)
);

OAI21x1_ASAP7_75t_L g3395 ( 
.A1(n_2606),
.A2(n_2756),
.B(n_2632),
.Y(n_3395)
);

BUFx4f_ASAP7_75t_L g3396 ( 
.A(n_2539),
.Y(n_3396)
);

BUFx10_ASAP7_75t_L g3397 ( 
.A(n_2363),
.Y(n_3397)
);

NAND2xp33_ASAP7_75t_L g3398 ( 
.A(n_2363),
.B(n_2978),
.Y(n_3398)
);

BUFx8_ASAP7_75t_L g3399 ( 
.A(n_2398),
.Y(n_3399)
);

INVxp67_ASAP7_75t_L g3400 ( 
.A(n_2899),
.Y(n_3400)
);

INVx2_ASAP7_75t_L g3401 ( 
.A(n_2581),
.Y(n_3401)
);

NOR2xp67_ASAP7_75t_L g3402 ( 
.A(n_2787),
.B(n_2803),
.Y(n_3402)
);

OR2x2_ASAP7_75t_L g3403 ( 
.A(n_2620),
.B(n_2637),
.Y(n_3403)
);

INVx2_ASAP7_75t_SL g3404 ( 
.A(n_2384),
.Y(n_3404)
);

INVx1_ASAP7_75t_SL g3405 ( 
.A(n_2836),
.Y(n_3405)
);

AND2x2_ASAP7_75t_L g3406 ( 
.A(n_2671),
.B(n_2683),
.Y(n_3406)
);

OR2x6_ASAP7_75t_L g3407 ( 
.A(n_2895),
.B(n_2896),
.Y(n_3407)
);

CKINVDCx5p33_ASAP7_75t_R g3408 ( 
.A(n_2398),
.Y(n_3408)
);

INVx1_ASAP7_75t_L g3409 ( 
.A(n_2683),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_2703),
.Y(n_3410)
);

INVx2_ASAP7_75t_L g3411 ( 
.A(n_2703),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_2770),
.Y(n_3412)
);

AND3x4_ASAP7_75t_L g3413 ( 
.A(n_2557),
.B(n_2409),
.C(n_2471),
.Y(n_3413)
);

NOR2xp33_ASAP7_75t_SL g3414 ( 
.A(n_2420),
.B(n_2812),
.Y(n_3414)
);

INVx2_ASAP7_75t_SL g3415 ( 
.A(n_2423),
.Y(n_3415)
);

AND2x2_ASAP7_75t_L g3416 ( 
.A(n_2896),
.B(n_2902),
.Y(n_3416)
);

NOR2xp33_ASAP7_75t_L g3417 ( 
.A(n_2409),
.B(n_2471),
.Y(n_3417)
);

INVx2_ASAP7_75t_L g3418 ( 
.A(n_2848),
.Y(n_3418)
);

OA22x2_ASAP7_75t_L g3419 ( 
.A1(n_2803),
.A2(n_2481),
.B1(n_2899),
.B2(n_2902),
.Y(n_3419)
);

A2O1A1Ixp33_ASAP7_75t_L g3420 ( 
.A1(n_2481),
.A2(n_2681),
.B(n_2423),
.C(n_2492),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_2880),
.B(n_2897),
.Y(n_3421)
);

AO31x2_ASAP7_75t_L g3422 ( 
.A1(n_2863),
.A2(n_2897),
.A3(n_2880),
.B(n_2521),
.Y(n_3422)
);

OAI22xp5_ASAP7_75t_L g3423 ( 
.A1(n_2850),
.A2(n_2851),
.B1(n_2772),
.B2(n_2812),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_L g3424 ( 
.A(n_2880),
.B(n_2897),
.Y(n_3424)
);

A2O1A1Ixp33_ASAP7_75t_L g3425 ( 
.A1(n_2492),
.A2(n_2709),
.B(n_2521),
.C(n_2767),
.Y(n_3425)
);

INVx1_ASAP7_75t_SL g3426 ( 
.A(n_2631),
.Y(n_3426)
);

INVx3_ASAP7_75t_L g3427 ( 
.A(n_2681),
.Y(n_3427)
);

A2O1A1Ixp33_ASAP7_75t_L g3428 ( 
.A1(n_2557),
.A2(n_2897),
.B(n_2420),
.C(n_2684),
.Y(n_3428)
);

OAI22xp5_ASAP7_75t_L g3429 ( 
.A1(n_2684),
.A2(n_2772),
.B1(n_2730),
.B2(n_2744),
.Y(n_3429)
);

INVx2_ASAP7_75t_L g3430 ( 
.A(n_2528),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_2528),
.Y(n_3431)
);

A2O1A1Ixp33_ASAP7_75t_L g3432 ( 
.A1(n_2528),
.A2(n_2730),
.B(n_2744),
.C(n_2755),
.Y(n_3432)
);

OAI21x1_ASAP7_75t_L g3433 ( 
.A1(n_2528),
.A2(n_2730),
.B(n_2744),
.Y(n_3433)
);

O2A1O1Ixp5_ASAP7_75t_L g3434 ( 
.A1(n_2730),
.A2(n_1107),
.B(n_2350),
.C(n_1439),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_2744),
.Y(n_3435)
);

OAI21x1_ASAP7_75t_SL g3436 ( 
.A1(n_2755),
.A2(n_2350),
.B(n_2932),
.Y(n_3436)
);

AOI21xp5_ASAP7_75t_L g3437 ( 
.A1(n_2755),
.A2(n_1107),
.B(n_2058),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_L g3438 ( 
.A(n_2755),
.B(n_2351),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_L g3439 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_2695),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3441)
);

OAI21x1_ASAP7_75t_SL g3442 ( 
.A1(n_2350),
.A2(n_2937),
.B(n_2932),
.Y(n_3442)
);

AO21x1_ASAP7_75t_L g3443 ( 
.A1(n_2428),
.A2(n_2135),
.B(n_2442),
.Y(n_3443)
);

OAI21xp5_ASAP7_75t_L g3444 ( 
.A1(n_2400),
.A2(n_1107),
.B(n_1437),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_L g3445 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3446)
);

OAI22x1_ASAP7_75t_L g3447 ( 
.A1(n_2388),
.A2(n_2937),
.B1(n_2949),
.B2(n_2932),
.Y(n_3447)
);

OAI21xp5_ASAP7_75t_L g3448 ( 
.A1(n_2400),
.A2(n_1107),
.B(n_1437),
.Y(n_3448)
);

AOI22xp5_ASAP7_75t_L g3449 ( 
.A1(n_2321),
.A2(n_2079),
.B1(n_2388),
.B2(n_1568),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3450)
);

OR2x2_ASAP7_75t_L g3451 ( 
.A(n_2450),
.B(n_2385),
.Y(n_3451)
);

INVxp67_ASAP7_75t_SL g3452 ( 
.A(n_2908),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3453)
);

AOI21xp5_ASAP7_75t_L g3454 ( 
.A1(n_2369),
.A2(n_1107),
.B(n_2058),
.Y(n_3454)
);

NAND2xp5_ASAP7_75t_L g3455 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3455)
);

AOI22xp5_ASAP7_75t_L g3456 ( 
.A1(n_2321),
.A2(n_2079),
.B1(n_2388),
.B2(n_1568),
.Y(n_3456)
);

OAI21xp5_ASAP7_75t_L g3457 ( 
.A1(n_2400),
.A2(n_1107),
.B(n_1437),
.Y(n_3457)
);

AND2x2_ASAP7_75t_L g3458 ( 
.A(n_2480),
.B(n_2514),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_L g3459 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3459)
);

A2O1A1Ixp33_ASAP7_75t_L g3460 ( 
.A1(n_2321),
.A2(n_1552),
.B(n_1492),
.C(n_2462),
.Y(n_3460)
);

AOI21xp5_ASAP7_75t_L g3461 ( 
.A1(n_2369),
.A2(n_1107),
.B(n_2058),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3462)
);

AOI21xp5_ASAP7_75t_L g3463 ( 
.A1(n_2369),
.A2(n_1107),
.B(n_2058),
.Y(n_3463)
);

AO21x1_ASAP7_75t_L g3464 ( 
.A1(n_2428),
.A2(n_2135),
.B(n_2442),
.Y(n_3464)
);

INVx4_ASAP7_75t_L g3465 ( 
.A(n_2579),
.Y(n_3465)
);

O2A1O1Ixp5_ASAP7_75t_L g3466 ( 
.A1(n_2350),
.A2(n_1107),
.B(n_1439),
.C(n_1437),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_L g3467 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3467)
);

BUFx6f_ASAP7_75t_L g3468 ( 
.A(n_2912),
.Y(n_3468)
);

AOI21xp33_ASAP7_75t_L g3469 ( 
.A1(n_2917),
.A2(n_1107),
.B(n_2211),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_L g3470 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3470)
);

AOI21xp5_ASAP7_75t_L g3471 ( 
.A1(n_2369),
.A2(n_1107),
.B(n_2058),
.Y(n_3471)
);

NAND3xp33_ASAP7_75t_SL g3472 ( 
.A(n_2390),
.B(n_1461),
.C(n_1407),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_2695),
.Y(n_3473)
);

AOI21xp5_ASAP7_75t_L g3474 ( 
.A1(n_2369),
.A2(n_1107),
.B(n_2058),
.Y(n_3474)
);

OAI22xp5_ASAP7_75t_L g3475 ( 
.A1(n_2932),
.A2(n_2937),
.B1(n_2966),
.B2(n_2949),
.Y(n_3475)
);

CKINVDCx11_ASAP7_75t_R g3476 ( 
.A(n_2957),
.Y(n_3476)
);

AOI21xp33_ASAP7_75t_L g3477 ( 
.A1(n_2917),
.A2(n_1107),
.B(n_2211),
.Y(n_3477)
);

OAI21xp5_ASAP7_75t_L g3478 ( 
.A1(n_2400),
.A2(n_1107),
.B(n_1437),
.Y(n_3478)
);

O2A1O1Ixp5_ASAP7_75t_L g3479 ( 
.A1(n_2350),
.A2(n_1107),
.B(n_1439),
.C(n_1437),
.Y(n_3479)
);

AND2x2_ASAP7_75t_L g3480 ( 
.A(n_2480),
.B(n_2514),
.Y(n_3480)
);

OAI21xp5_ASAP7_75t_L g3481 ( 
.A1(n_2400),
.A2(n_1107),
.B(n_1437),
.Y(n_3481)
);

AO21x2_ASAP7_75t_L g3482 ( 
.A1(n_2404),
.A2(n_2143),
.B(n_1101),
.Y(n_3482)
);

OAI21x1_ASAP7_75t_SL g3483 ( 
.A1(n_2350),
.A2(n_2937),
.B(n_2932),
.Y(n_3483)
);

A2O1A1Ixp33_ASAP7_75t_L g3484 ( 
.A1(n_2321),
.A2(n_1552),
.B(n_1492),
.C(n_2462),
.Y(n_3484)
);

A2O1A1Ixp33_ASAP7_75t_L g3485 ( 
.A1(n_2321),
.A2(n_1552),
.B(n_1492),
.C(n_2462),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_L g3486 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_2695),
.Y(n_3487)
);

BUFx5_ASAP7_75t_L g3488 ( 
.A(n_2912),
.Y(n_3488)
);

OAI22x1_ASAP7_75t_L g3489 ( 
.A1(n_2388),
.A2(n_2937),
.B1(n_2949),
.B2(n_2932),
.Y(n_3489)
);

OAI21xp5_ASAP7_75t_L g3490 ( 
.A1(n_2400),
.A2(n_1107),
.B(n_1437),
.Y(n_3490)
);

OAI21x1_ASAP7_75t_SL g3491 ( 
.A1(n_2350),
.A2(n_2937),
.B(n_2932),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_2695),
.Y(n_3492)
);

AOI21xp5_ASAP7_75t_L g3493 ( 
.A1(n_2369),
.A2(n_1107),
.B(n_2058),
.Y(n_3493)
);

NAND3xp33_ASAP7_75t_L g3494 ( 
.A(n_2390),
.B(n_1107),
.C(n_2369),
.Y(n_3494)
);

NOR2x1_ASAP7_75t_SL g3495 ( 
.A(n_2579),
.B(n_2591),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_L g3496 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3496)
);

INVx1_ASAP7_75t_SL g3497 ( 
.A(n_2577),
.Y(n_3497)
);

AOI22xp5_ASAP7_75t_L g3498 ( 
.A1(n_2321),
.A2(n_2079),
.B1(n_2388),
.B2(n_1568),
.Y(n_3498)
);

INVx2_ASAP7_75t_L g3499 ( 
.A(n_2696),
.Y(n_3499)
);

NOR2xp33_ASAP7_75t_L g3500 ( 
.A(n_2330),
.B(n_2344),
.Y(n_3500)
);

AOI21xp5_ASAP7_75t_L g3501 ( 
.A1(n_2913),
.A2(n_1107),
.B(n_2058),
.Y(n_3501)
);

INVx3_ASAP7_75t_L g3502 ( 
.A(n_2584),
.Y(n_3502)
);

AND2x2_ASAP7_75t_SL g3503 ( 
.A(n_2603),
.B(n_1627),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3504)
);

AOI21xp5_ASAP7_75t_L g3505 ( 
.A1(n_2913),
.A2(n_1107),
.B(n_2058),
.Y(n_3505)
);

AOI21xp5_ASAP7_75t_L g3506 ( 
.A1(n_2913),
.A2(n_1107),
.B(n_2058),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3507)
);

BUFx2_ASAP7_75t_L g3508 ( 
.A(n_2565),
.Y(n_3508)
);

OAI21xp5_ASAP7_75t_L g3509 ( 
.A1(n_2400),
.A2(n_1107),
.B(n_1437),
.Y(n_3509)
);

O2A1O1Ixp5_ASAP7_75t_L g3510 ( 
.A1(n_2350),
.A2(n_1107),
.B(n_1439),
.C(n_1437),
.Y(n_3510)
);

AOI21xp5_ASAP7_75t_L g3511 ( 
.A1(n_2913),
.A2(n_1107),
.B(n_2058),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_L g3512 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3512)
);

INVx5_ASAP7_75t_L g3513 ( 
.A(n_2579),
.Y(n_3513)
);

OAI21x1_ASAP7_75t_SL g3514 ( 
.A1(n_2350),
.A2(n_2937),
.B(n_2932),
.Y(n_3514)
);

INVxp67_ASAP7_75t_L g3515 ( 
.A(n_2330),
.Y(n_3515)
);

A2O1A1Ixp33_ASAP7_75t_L g3516 ( 
.A1(n_2321),
.A2(n_1552),
.B(n_1492),
.C(n_2462),
.Y(n_3516)
);

A2O1A1Ixp33_ASAP7_75t_L g3517 ( 
.A1(n_2321),
.A2(n_1552),
.B(n_1492),
.C(n_2462),
.Y(n_3517)
);

OR2x2_ASAP7_75t_L g3518 ( 
.A(n_2450),
.B(n_2385),
.Y(n_3518)
);

BUFx3_ASAP7_75t_L g3519 ( 
.A(n_2818),
.Y(n_3519)
);

OAI22xp5_ASAP7_75t_L g3520 ( 
.A1(n_2932),
.A2(n_2937),
.B1(n_2966),
.B2(n_2949),
.Y(n_3520)
);

OAI21xp5_ASAP7_75t_SL g3521 ( 
.A1(n_2932),
.A2(n_2949),
.B(n_2937),
.Y(n_3521)
);

AOI21xp5_ASAP7_75t_L g3522 ( 
.A1(n_2913),
.A2(n_1107),
.B(n_2058),
.Y(n_3522)
);

AO31x2_ASAP7_75t_L g3523 ( 
.A1(n_2714),
.A2(n_2352),
.A3(n_2911),
.B(n_2342),
.Y(n_3523)
);

INVx2_ASAP7_75t_SL g3524 ( 
.A(n_2704),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3525)
);

NOR2xp33_ASAP7_75t_L g3526 ( 
.A(n_2330),
.B(n_2344),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_L g3527 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3527)
);

INVx3_ASAP7_75t_L g3528 ( 
.A(n_2584),
.Y(n_3528)
);

OAI22x1_ASAP7_75t_L g3529 ( 
.A1(n_2388),
.A2(n_2937),
.B1(n_2949),
.B2(n_2932),
.Y(n_3529)
);

INVx2_ASAP7_75t_L g3530 ( 
.A(n_2696),
.Y(n_3530)
);

A2O1A1Ixp33_ASAP7_75t_L g3531 ( 
.A1(n_2321),
.A2(n_1552),
.B(n_1492),
.C(n_2462),
.Y(n_3531)
);

INVx2_ASAP7_75t_SL g3532 ( 
.A(n_2704),
.Y(n_3532)
);

INVx3_ASAP7_75t_L g3533 ( 
.A(n_2584),
.Y(n_3533)
);

A2O1A1Ixp33_ASAP7_75t_L g3534 ( 
.A1(n_2321),
.A2(n_1552),
.B(n_1492),
.C(n_2462),
.Y(n_3534)
);

AOI21xp5_ASAP7_75t_L g3535 ( 
.A1(n_2369),
.A2(n_1107),
.B(n_2058),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3536)
);

INVx3_ASAP7_75t_L g3537 ( 
.A(n_2584),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_2695),
.Y(n_3538)
);

OAI21xp5_ASAP7_75t_L g3539 ( 
.A1(n_2400),
.A2(n_1107),
.B(n_1437),
.Y(n_3539)
);

AO31x2_ASAP7_75t_L g3540 ( 
.A1(n_2714),
.A2(n_2352),
.A3(n_2911),
.B(n_2342),
.Y(n_3540)
);

OAI21xp5_ASAP7_75t_L g3541 ( 
.A1(n_2400),
.A2(n_1107),
.B(n_1437),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_2695),
.Y(n_3542)
);

AOI221xp5_ASAP7_75t_SL g3543 ( 
.A1(n_2321),
.A2(n_2369),
.B1(n_2386),
.B2(n_2442),
.C(n_2428),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_SL g3544 ( 
.A(n_2390),
.B(n_2321),
.Y(n_3544)
);

OAI22xp5_ASAP7_75t_L g3545 ( 
.A1(n_2932),
.A2(n_2937),
.B1(n_2966),
.B2(n_2949),
.Y(n_3545)
);

INVx2_ASAP7_75t_SL g3546 ( 
.A(n_2704),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3547)
);

NAND2xp5_ASAP7_75t_SL g3548 ( 
.A(n_2390),
.B(n_2321),
.Y(n_3548)
);

AOI21xp5_ASAP7_75t_L g3549 ( 
.A1(n_2369),
.A2(n_1107),
.B(n_2058),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_2695),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_L g3551 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3551)
);

INVx2_ASAP7_75t_SL g3552 ( 
.A(n_2704),
.Y(n_3552)
);

AO21x1_ASAP7_75t_L g3553 ( 
.A1(n_2428),
.A2(n_2135),
.B(n_2442),
.Y(n_3553)
);

AOI21xp5_ASAP7_75t_L g3554 ( 
.A1(n_2369),
.A2(n_1107),
.B(n_2058),
.Y(n_3554)
);

BUFx12f_ASAP7_75t_L g3555 ( 
.A(n_2957),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_L g3556 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3556)
);

NOR2x1_ASAP7_75t_L g3557 ( 
.A(n_2375),
.B(n_2412),
.Y(n_3557)
);

AOI21xp5_ASAP7_75t_L g3558 ( 
.A1(n_2369),
.A2(n_1107),
.B(n_2058),
.Y(n_3558)
);

AOI21x1_ASAP7_75t_L g3559 ( 
.A1(n_2923),
.A2(n_1673),
.B(n_2929),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_L g3560 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3560)
);

BUFx4f_ASAP7_75t_SL g3561 ( 
.A(n_2957),
.Y(n_3561)
);

BUFx5_ASAP7_75t_L g3562 ( 
.A(n_2912),
.Y(n_3562)
);

AOI221xp5_ASAP7_75t_SL g3563 ( 
.A1(n_2321),
.A2(n_2369),
.B1(n_2386),
.B2(n_2442),
.C(n_2428),
.Y(n_3563)
);

AOI21xp5_ASAP7_75t_L g3564 ( 
.A1(n_2369),
.A2(n_1107),
.B(n_2058),
.Y(n_3564)
);

OAI21xp5_ASAP7_75t_L g3565 ( 
.A1(n_2400),
.A2(n_1107),
.B(n_1437),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3566)
);

AOI21xp5_ASAP7_75t_SL g3567 ( 
.A1(n_2932),
.A2(n_2175),
.B(n_2129),
.Y(n_3567)
);

OAI21x1_ASAP7_75t_L g3568 ( 
.A1(n_2325),
.A2(n_2961),
.B(n_2936),
.Y(n_3568)
);

INVx3_ASAP7_75t_L g3569 ( 
.A(n_2584),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3570)
);

AOI21xp5_ASAP7_75t_L g3571 ( 
.A1(n_2369),
.A2(n_1107),
.B(n_2058),
.Y(n_3571)
);

A2O1A1Ixp33_ASAP7_75t_L g3572 ( 
.A1(n_2321),
.A2(n_1552),
.B(n_1492),
.C(n_2462),
.Y(n_3572)
);

OAI21x1_ASAP7_75t_L g3573 ( 
.A1(n_2325),
.A2(n_2961),
.B(n_2936),
.Y(n_3573)
);

INVxp67_ASAP7_75t_SL g3574 ( 
.A(n_2908),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_L g3575 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3575)
);

OAI22xp5_ASAP7_75t_L g3576 ( 
.A1(n_2932),
.A2(n_2937),
.B1(n_2966),
.B2(n_2949),
.Y(n_3576)
);

NOR2xp33_ASAP7_75t_L g3577 ( 
.A(n_2330),
.B(n_2344),
.Y(n_3577)
);

AND2x4_ASAP7_75t_L g3578 ( 
.A(n_2603),
.B(n_2769),
.Y(n_3578)
);

AOI222xp33_ASAP7_75t_L g3579 ( 
.A1(n_2321),
.A2(n_2079),
.B1(n_2390),
.B2(n_2340),
.C1(n_1689),
.C2(n_2958),
.Y(n_3579)
);

OAI22xp5_ASAP7_75t_L g3580 ( 
.A1(n_2932),
.A2(n_2937),
.B1(n_2966),
.B2(n_2949),
.Y(n_3580)
);

INVx2_ASAP7_75t_L g3581 ( 
.A(n_2696),
.Y(n_3581)
);

CKINVDCx20_ASAP7_75t_R g3582 ( 
.A(n_2642),
.Y(n_3582)
);

CKINVDCx20_ASAP7_75t_R g3583 ( 
.A(n_2642),
.Y(n_3583)
);

OAI21xp5_ASAP7_75t_L g3584 ( 
.A1(n_2400),
.A2(n_1107),
.B(n_1437),
.Y(n_3584)
);

OAI21x1_ASAP7_75t_L g3585 ( 
.A1(n_2325),
.A2(n_2961),
.B(n_2936),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3586)
);

AND2x2_ASAP7_75t_L g3587 ( 
.A(n_2480),
.B(n_2514),
.Y(n_3587)
);

AOI21xp5_ASAP7_75t_L g3588 ( 
.A1(n_2369),
.A2(n_1107),
.B(n_2058),
.Y(n_3588)
);

INVxp67_ASAP7_75t_SL g3589 ( 
.A(n_2908),
.Y(n_3589)
);

AO31x2_ASAP7_75t_L g3590 ( 
.A1(n_2714),
.A2(n_2352),
.A3(n_2911),
.B(n_2342),
.Y(n_3590)
);

AOI211x1_ASAP7_75t_L g3591 ( 
.A1(n_2399),
.A2(n_2321),
.B(n_2400),
.C(n_2428),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3592)
);

A2O1A1Ixp33_ASAP7_75t_L g3593 ( 
.A1(n_2321),
.A2(n_1552),
.B(n_1492),
.C(n_2462),
.Y(n_3593)
);

OAI21xp5_ASAP7_75t_L g3594 ( 
.A1(n_2400),
.A2(n_1107),
.B(n_1437),
.Y(n_3594)
);

INVx1_ASAP7_75t_SL g3595 ( 
.A(n_2577),
.Y(n_3595)
);

INVx3_ASAP7_75t_L g3596 ( 
.A(n_2584),
.Y(n_3596)
);

AOI21xp5_ASAP7_75t_L g3597 ( 
.A1(n_2369),
.A2(n_1107),
.B(n_2058),
.Y(n_3597)
);

AOI21x1_ASAP7_75t_L g3598 ( 
.A1(n_2923),
.A2(n_1673),
.B(n_2929),
.Y(n_3598)
);

AOI21x1_ASAP7_75t_SL g3599 ( 
.A1(n_2421),
.A2(n_1704),
.B(n_1700),
.Y(n_3599)
);

OR2x2_ASAP7_75t_L g3600 ( 
.A(n_2450),
.B(n_2385),
.Y(n_3600)
);

O2A1O1Ixp33_ASAP7_75t_L g3601 ( 
.A1(n_2959),
.A2(n_1107),
.B(n_1439),
.C(n_1437),
.Y(n_3601)
);

AOI21xp33_ASAP7_75t_L g3602 ( 
.A1(n_2917),
.A2(n_1107),
.B(n_2211),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3603)
);

A2O1A1Ixp33_ASAP7_75t_L g3604 ( 
.A1(n_2321),
.A2(n_1552),
.B(n_1492),
.C(n_2462),
.Y(n_3604)
);

AOI21xp5_ASAP7_75t_L g3605 ( 
.A1(n_2913),
.A2(n_1107),
.B(n_2058),
.Y(n_3605)
);

OAI21xp33_ASAP7_75t_L g3606 ( 
.A1(n_2321),
.A2(n_2079),
.B(n_2350),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_SL g3607 ( 
.A(n_2390),
.B(n_2321),
.Y(n_3607)
);

AOI21xp5_ASAP7_75t_L g3608 ( 
.A1(n_2913),
.A2(n_1107),
.B(n_2058),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_L g3609 ( 
.A(n_2351),
.B(n_2357),
.Y(n_3609)
);

A2O1A1Ixp33_ASAP7_75t_L g3610 ( 
.A1(n_2321),
.A2(n_1552),
.B(n_1492),
.C(n_2462),
.Y(n_3610)
);

BUFx6f_ASAP7_75t_L g3611 ( 
.A(n_3277),
.Y(n_3611)
);

BUFx2_ASAP7_75t_L g3612 ( 
.A(n_3452),
.Y(n_3612)
);

BUFx4_ASAP7_75t_SL g3613 ( 
.A(n_3316),
.Y(n_3613)
);

BUFx5_ASAP7_75t_L g3614 ( 
.A(n_3503),
.Y(n_3614)
);

AOI22xp33_ASAP7_75t_L g3615 ( 
.A1(n_3606),
.A2(n_3579),
.B1(n_2993),
.B2(n_3548),
.Y(n_3615)
);

BUFx12f_ASAP7_75t_L g3616 ( 
.A(n_3476),
.Y(n_3616)
);

INVx1_ASAP7_75t_SL g3617 ( 
.A(n_3035),
.Y(n_3617)
);

BUFx2_ASAP7_75t_L g3618 ( 
.A(n_3574),
.Y(n_3618)
);

AND2x4_ASAP7_75t_L g3619 ( 
.A(n_3115),
.B(n_2991),
.Y(n_3619)
);

INVx1_ASAP7_75t_SL g3620 ( 
.A(n_3035),
.Y(n_3620)
);

INVxp67_ASAP7_75t_SL g3621 ( 
.A(n_3028),
.Y(n_3621)
);

CKINVDCx5p33_ASAP7_75t_R g3622 ( 
.A(n_3176),
.Y(n_3622)
);

CKINVDCx14_ASAP7_75t_R g3623 ( 
.A(n_3274),
.Y(n_3623)
);

INVx1_ASAP7_75t_SL g3624 ( 
.A(n_3067),
.Y(n_3624)
);

OR2x6_ASAP7_75t_SL g3625 ( 
.A(n_3013),
.B(n_3475),
.Y(n_3625)
);

INVx2_ASAP7_75t_L g3626 ( 
.A(n_3374),
.Y(n_3626)
);

BUFx8_ASAP7_75t_L g3627 ( 
.A(n_3555),
.Y(n_3627)
);

CKINVDCx20_ASAP7_75t_R g3628 ( 
.A(n_3582),
.Y(n_3628)
);

INVx5_ASAP7_75t_L g3629 ( 
.A(n_3334),
.Y(n_3629)
);

BUFx2_ASAP7_75t_L g3630 ( 
.A(n_3589),
.Y(n_3630)
);

BUFx2_ASAP7_75t_L g3631 ( 
.A(n_3508),
.Y(n_3631)
);

INVx5_ASAP7_75t_L g3632 ( 
.A(n_3334),
.Y(n_3632)
);

INVx2_ASAP7_75t_SL g3633 ( 
.A(n_3231),
.Y(n_3633)
);

CKINVDCx5p33_ASAP7_75t_R g3634 ( 
.A(n_3555),
.Y(n_3634)
);

INVx4_ASAP7_75t_L g3635 ( 
.A(n_3384),
.Y(n_3635)
);

INVx4_ASAP7_75t_L g3636 ( 
.A(n_3384),
.Y(n_3636)
);

INVx2_ASAP7_75t_L g3637 ( 
.A(n_3374),
.Y(n_3637)
);

INVx3_ASAP7_75t_L g3638 ( 
.A(n_2991),
.Y(n_3638)
);

CKINVDCx20_ASAP7_75t_R g3639 ( 
.A(n_3583),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_L g3640 ( 
.A(n_3014),
.B(n_3011),
.Y(n_3640)
);

NAND2xp5_ASAP7_75t_L g3641 ( 
.A(n_3014),
.B(n_3011),
.Y(n_3641)
);

INVx4_ASAP7_75t_L g3642 ( 
.A(n_3384),
.Y(n_3642)
);

BUFx4f_ASAP7_75t_L g3643 ( 
.A(n_3503),
.Y(n_3643)
);

CKINVDCx6p67_ASAP7_75t_R g3644 ( 
.A(n_3387),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_SL g3645 ( 
.A(n_3023),
.B(n_3443),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3063),
.Y(n_3646)
);

AND2x4_ASAP7_75t_L g3647 ( 
.A(n_3115),
.B(n_3502),
.Y(n_3647)
);

INVxp67_ASAP7_75t_SL g3648 ( 
.A(n_3028),
.Y(n_3648)
);

NAND2x1p5_ASAP7_75t_L g3649 ( 
.A(n_3019),
.B(n_3044),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_L g3650 ( 
.A(n_3010),
.B(n_3125),
.Y(n_3650)
);

INVx2_ASAP7_75t_L g3651 ( 
.A(n_3377),
.Y(n_3651)
);

INVx6_ASAP7_75t_L g3652 ( 
.A(n_3019),
.Y(n_3652)
);

NAND2x1p5_ASAP7_75t_L g3653 ( 
.A(n_3019),
.B(n_3044),
.Y(n_3653)
);

CKINVDCx5p33_ASAP7_75t_R g3654 ( 
.A(n_3555),
.Y(n_3654)
);

INVx5_ASAP7_75t_SL g3655 ( 
.A(n_3002),
.Y(n_3655)
);

INVxp67_ASAP7_75t_SL g3656 ( 
.A(n_3034),
.Y(n_3656)
);

HB1xp67_ASAP7_75t_L g3657 ( 
.A(n_3328),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_3010),
.B(n_3125),
.Y(n_3658)
);

BUFx12f_ASAP7_75t_L g3659 ( 
.A(n_3005),
.Y(n_3659)
);

OR2x6_ASAP7_75t_SL g3660 ( 
.A(n_3013),
.B(n_3475),
.Y(n_3660)
);

INVx1_ASAP7_75t_SL g3661 ( 
.A(n_3067),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3063),
.Y(n_3662)
);

NAND2x1p5_ASAP7_75t_L g3663 ( 
.A(n_3019),
.B(n_3044),
.Y(n_3663)
);

NAND2x1p5_ASAP7_75t_L g3664 ( 
.A(n_3019),
.B(n_3044),
.Y(n_3664)
);

INVx5_ASAP7_75t_L g3665 ( 
.A(n_3334),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3079),
.Y(n_3666)
);

INVx1_ASAP7_75t_SL g3667 ( 
.A(n_3497),
.Y(n_3667)
);

INVx1_ASAP7_75t_L g3668 ( 
.A(n_3079),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_L g3669 ( 
.A(n_3020),
.B(n_3126),
.Y(n_3669)
);

INVx6_ASAP7_75t_L g3670 ( 
.A(n_3019),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3083),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_3020),
.B(n_3126),
.Y(n_3672)
);

INVx1_ASAP7_75t_SL g3673 ( 
.A(n_3497),
.Y(n_3673)
);

INVx2_ASAP7_75t_L g3674 ( 
.A(n_3378),
.Y(n_3674)
);

BUFx6f_ASAP7_75t_SL g3675 ( 
.A(n_3268),
.Y(n_3675)
);

INVx4_ASAP7_75t_L g3676 ( 
.A(n_3387),
.Y(n_3676)
);

HB1xp67_ASAP7_75t_L g3677 ( 
.A(n_3328),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3083),
.Y(n_3678)
);

BUFx4f_ASAP7_75t_L g3679 ( 
.A(n_3503),
.Y(n_3679)
);

AND2x4_ASAP7_75t_L g3680 ( 
.A(n_3115),
.B(n_3502),
.Y(n_3680)
);

NAND2xp5_ASAP7_75t_L g3681 ( 
.A(n_2997),
.B(n_3003),
.Y(n_3681)
);

CKINVDCx11_ASAP7_75t_R g3682 ( 
.A(n_3341),
.Y(n_3682)
);

INVx2_ASAP7_75t_L g3683 ( 
.A(n_3378),
.Y(n_3683)
);

INVx1_ASAP7_75t_L g3684 ( 
.A(n_3145),
.Y(n_3684)
);

BUFx2_ASAP7_75t_L g3685 ( 
.A(n_3519),
.Y(n_3685)
);

INVx6_ASAP7_75t_L g3686 ( 
.A(n_3044),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_3145),
.Y(n_3687)
);

CKINVDCx16_ASAP7_75t_R g3688 ( 
.A(n_3414),
.Y(n_3688)
);

NOR2xp33_ASAP7_75t_L g3689 ( 
.A(n_3500),
.B(n_3526),
.Y(n_3689)
);

BUFx10_ASAP7_75t_L g3690 ( 
.A(n_3417),
.Y(n_3690)
);

BUFx12f_ASAP7_75t_L g3691 ( 
.A(n_3297),
.Y(n_3691)
);

INVx1_ASAP7_75t_SL g3692 ( 
.A(n_3595),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3147),
.Y(n_3693)
);

BUFx12f_ASAP7_75t_L g3694 ( 
.A(n_3399),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3147),
.Y(n_3695)
);

BUFx8_ASAP7_75t_L g3696 ( 
.A(n_3430),
.Y(n_3696)
);

BUFx3_ASAP7_75t_L g3697 ( 
.A(n_3433),
.Y(n_3697)
);

INVx4_ASAP7_75t_L g3698 ( 
.A(n_3387),
.Y(n_3698)
);

CKINVDCx16_ASAP7_75t_R g3699 ( 
.A(n_3414),
.Y(n_3699)
);

INVx2_ASAP7_75t_L g3700 ( 
.A(n_3381),
.Y(n_3700)
);

INVx1_ASAP7_75t_SL g3701 ( 
.A(n_3595),
.Y(n_3701)
);

INVx3_ASAP7_75t_L g3702 ( 
.A(n_3502),
.Y(n_3702)
);

INVx1_ASAP7_75t_SL g3703 ( 
.A(n_3183),
.Y(n_3703)
);

INVxp67_ASAP7_75t_SL g3704 ( 
.A(n_3034),
.Y(n_3704)
);

INVx2_ASAP7_75t_L g3705 ( 
.A(n_3381),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3152),
.Y(n_3706)
);

BUFx3_ASAP7_75t_L g3707 ( 
.A(n_3433),
.Y(n_3707)
);

AOI22xp5_ASAP7_75t_L g3708 ( 
.A1(n_3606),
.A2(n_3456),
.B1(n_3498),
.B2(n_3449),
.Y(n_3708)
);

INVx4_ASAP7_75t_L g3709 ( 
.A(n_3268),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3152),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_L g3711 ( 
.A(n_2997),
.B(n_3003),
.Y(n_3711)
);

BUFx12f_ASAP7_75t_L g3712 ( 
.A(n_3399),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_3007),
.B(n_3009),
.Y(n_3713)
);

NAND2x1p5_ASAP7_75t_L g3714 ( 
.A(n_3044),
.B(n_3162),
.Y(n_3714)
);

CKINVDCx14_ASAP7_75t_R g3715 ( 
.A(n_3274),
.Y(n_3715)
);

CKINVDCx5p33_ASAP7_75t_R g3716 ( 
.A(n_3341),
.Y(n_3716)
);

BUFx2_ASAP7_75t_L g3717 ( 
.A(n_3058),
.Y(n_3717)
);

INVx1_ASAP7_75t_SL g3718 ( 
.A(n_3183),
.Y(n_3718)
);

INVx4_ASAP7_75t_L g3719 ( 
.A(n_3268),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_L g3720 ( 
.A(n_3007),
.B(n_3009),
.Y(n_3720)
);

NAND2x1p5_ASAP7_75t_L g3721 ( 
.A(n_3162),
.B(n_3513),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_3191),
.Y(n_3722)
);

INVx3_ASAP7_75t_L g3723 ( 
.A(n_3502),
.Y(n_3723)
);

BUFx12f_ASAP7_75t_L g3724 ( 
.A(n_3399),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3191),
.Y(n_3725)
);

AND2x4_ASAP7_75t_L g3726 ( 
.A(n_3115),
.B(n_3528),
.Y(n_3726)
);

BUFx4f_ASAP7_75t_SL g3727 ( 
.A(n_3151),
.Y(n_3727)
);

BUFx3_ASAP7_75t_L g3728 ( 
.A(n_3166),
.Y(n_3728)
);

AOI22xp5_ASAP7_75t_L g3729 ( 
.A1(n_3449),
.A2(n_3498),
.B1(n_3456),
.B2(n_3544),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_3197),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3197),
.Y(n_3731)
);

BUFx4f_ASAP7_75t_L g3732 ( 
.A(n_3086),
.Y(n_3732)
);

INVx4_ASAP7_75t_L g3733 ( 
.A(n_3413),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3200),
.Y(n_3734)
);

NAND2xp5_ASAP7_75t_L g3735 ( 
.A(n_3439),
.B(n_3441),
.Y(n_3735)
);

BUFx12f_ASAP7_75t_L g3736 ( 
.A(n_3399),
.Y(n_3736)
);

INVx3_ASAP7_75t_L g3737 ( 
.A(n_3528),
.Y(n_3737)
);

HB1xp67_ASAP7_75t_L g3738 ( 
.A(n_3331),
.Y(n_3738)
);

BUFx3_ASAP7_75t_L g3739 ( 
.A(n_3166),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3200),
.Y(n_3740)
);

INVx3_ASAP7_75t_L g3741 ( 
.A(n_3528),
.Y(n_3741)
);

INVx1_ASAP7_75t_SL g3742 ( 
.A(n_3208),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3217),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3217),
.Y(n_3744)
);

BUFx12f_ASAP7_75t_L g3745 ( 
.A(n_3385),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3236),
.Y(n_3746)
);

NAND2xp5_ASAP7_75t_L g3747 ( 
.A(n_3439),
.B(n_3441),
.Y(n_3747)
);

BUFx2_ASAP7_75t_L g3748 ( 
.A(n_3058),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3236),
.Y(n_3749)
);

BUFx12f_ASAP7_75t_L g3750 ( 
.A(n_3408),
.Y(n_3750)
);

INVx2_ASAP7_75t_L g3751 ( 
.A(n_3386),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3270),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3270),
.Y(n_3753)
);

BUFx3_ASAP7_75t_L g3754 ( 
.A(n_3431),
.Y(n_3754)
);

BUFx3_ASAP7_75t_L g3755 ( 
.A(n_3431),
.Y(n_3755)
);

BUFx3_ASAP7_75t_L g3756 ( 
.A(n_3435),
.Y(n_3756)
);

BUFx3_ASAP7_75t_L g3757 ( 
.A(n_3435),
.Y(n_3757)
);

INVx6_ASAP7_75t_SL g3758 ( 
.A(n_3120),
.Y(n_3758)
);

BUFx12f_ASAP7_75t_L g3759 ( 
.A(n_3335),
.Y(n_3759)
);

BUFx12f_ASAP7_75t_L g3760 ( 
.A(n_3335),
.Y(n_3760)
);

BUFx3_ASAP7_75t_L g3761 ( 
.A(n_3089),
.Y(n_3761)
);

NAND2xp5_ASAP7_75t_L g3762 ( 
.A(n_3445),
.B(n_3446),
.Y(n_3762)
);

BUFx12f_ASAP7_75t_L g3763 ( 
.A(n_3335),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3284),
.Y(n_3764)
);

AND2x4_ASAP7_75t_L g3765 ( 
.A(n_3528),
.B(n_3533),
.Y(n_3765)
);

BUFx6f_ASAP7_75t_SL g3766 ( 
.A(n_3334),
.Y(n_3766)
);

BUFx3_ASAP7_75t_L g3767 ( 
.A(n_3089),
.Y(n_3767)
);

CKINVDCx5p33_ASAP7_75t_R g3768 ( 
.A(n_3136),
.Y(n_3768)
);

NAND2x1p5_ASAP7_75t_L g3769 ( 
.A(n_3162),
.B(n_3513),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_3284),
.Y(n_3770)
);

BUFx2_ASAP7_75t_SL g3771 ( 
.A(n_3443),
.Y(n_3771)
);

INVxp67_ASAP7_75t_SL g3772 ( 
.A(n_3036),
.Y(n_3772)
);

NAND2xp5_ASAP7_75t_L g3773 ( 
.A(n_3445),
.B(n_3446),
.Y(n_3773)
);

BUFx2_ASAP7_75t_SL g3774 ( 
.A(n_3464),
.Y(n_3774)
);

AND2x2_ASAP7_75t_L g3775 ( 
.A(n_3094),
.B(n_3111),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_L g3776 ( 
.A(n_3450),
.B(n_3453),
.Y(n_3776)
);

INVx1_ASAP7_75t_SL g3777 ( 
.A(n_3208),
.Y(n_3777)
);

INVx3_ASAP7_75t_L g3778 ( 
.A(n_3533),
.Y(n_3778)
);

CKINVDCx5p33_ASAP7_75t_R g3779 ( 
.A(n_3561),
.Y(n_3779)
);

INVx1_ASAP7_75t_L g3780 ( 
.A(n_3306),
.Y(n_3780)
);

INVx6_ASAP7_75t_SL g3781 ( 
.A(n_3120),
.Y(n_3781)
);

BUFx4f_ASAP7_75t_SL g3782 ( 
.A(n_3194),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3306),
.Y(n_3783)
);

BUFx12f_ASAP7_75t_L g3784 ( 
.A(n_3335),
.Y(n_3784)
);

INVx3_ASAP7_75t_L g3785 ( 
.A(n_3533),
.Y(n_3785)
);

CKINVDCx6p67_ASAP7_75t_R g3786 ( 
.A(n_3366),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3338),
.Y(n_3787)
);

INVx3_ASAP7_75t_L g3788 ( 
.A(n_3537),
.Y(n_3788)
);

INVx1_ASAP7_75t_SL g3789 ( 
.A(n_3366),
.Y(n_3789)
);

NOR2x1_ASAP7_75t_R g3790 ( 
.A(n_3607),
.B(n_2995),
.Y(n_3790)
);

AOI22xp5_ASAP7_75t_L g3791 ( 
.A1(n_3579),
.A2(n_2999),
.B1(n_3489),
.B2(n_3447),
.Y(n_3791)
);

BUFx2_ASAP7_75t_L g3792 ( 
.A(n_3122),
.Y(n_3792)
);

INVx3_ASAP7_75t_SL g3793 ( 
.A(n_3366),
.Y(n_3793)
);

OAI22xp5_ASAP7_75t_L g3794 ( 
.A1(n_2999),
.A2(n_3494),
.B1(n_3521),
.B2(n_3484),
.Y(n_3794)
);

NAND2xp5_ASAP7_75t_L g3795 ( 
.A(n_3450),
.B(n_3453),
.Y(n_3795)
);

AOI22xp5_ASAP7_75t_L g3796 ( 
.A1(n_3447),
.A2(n_3529),
.B1(n_3489),
.B2(n_3520),
.Y(n_3796)
);

INVx5_ASAP7_75t_L g3797 ( 
.A(n_3334),
.Y(n_3797)
);

CKINVDCx5p33_ASAP7_75t_R g3798 ( 
.A(n_3362),
.Y(n_3798)
);

NOR2xp33_ASAP7_75t_L g3799 ( 
.A(n_3577),
.B(n_3042),
.Y(n_3799)
);

CKINVDCx8_ASAP7_75t_R g3800 ( 
.A(n_3257),
.Y(n_3800)
);

AND2x2_ASAP7_75t_L g3801 ( 
.A(n_3094),
.B(n_3111),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3338),
.Y(n_3802)
);

INVx8_ASAP7_75t_L g3803 ( 
.A(n_3162),
.Y(n_3803)
);

CKINVDCx20_ASAP7_75t_R g3804 ( 
.A(n_3194),
.Y(n_3804)
);

INVx2_ASAP7_75t_L g3805 ( 
.A(n_3386),
.Y(n_3805)
);

INVx3_ASAP7_75t_L g3806 ( 
.A(n_3537),
.Y(n_3806)
);

BUFx3_ASAP7_75t_L g3807 ( 
.A(n_3193),
.Y(n_3807)
);

INVx4_ASAP7_75t_L g3808 ( 
.A(n_3413),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_3344),
.Y(n_3809)
);

BUFx12f_ASAP7_75t_L g3810 ( 
.A(n_3397),
.Y(n_3810)
);

CKINVDCx5p33_ASAP7_75t_R g3811 ( 
.A(n_3108),
.Y(n_3811)
);

BUFx12f_ASAP7_75t_L g3812 ( 
.A(n_3397),
.Y(n_3812)
);

INVx2_ASAP7_75t_L g3813 ( 
.A(n_3394),
.Y(n_3813)
);

INVx3_ASAP7_75t_L g3814 ( 
.A(n_3537),
.Y(n_3814)
);

INVx4_ASAP7_75t_L g3815 ( 
.A(n_3413),
.Y(n_3815)
);

NAND2xp5_ASAP7_75t_L g3816 ( 
.A(n_3455),
.B(n_3459),
.Y(n_3816)
);

INVx1_ASAP7_75t_SL g3817 ( 
.A(n_3290),
.Y(n_3817)
);

INVx6_ASAP7_75t_L g3818 ( 
.A(n_3513),
.Y(n_3818)
);

BUFx10_ASAP7_75t_L g3819 ( 
.A(n_3099),
.Y(n_3819)
);

AOI22xp33_ASAP7_75t_L g3820 ( 
.A1(n_3024),
.A2(n_3529),
.B1(n_3017),
.B2(n_3520),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3344),
.Y(n_3821)
);

AND2x2_ASAP7_75t_SL g3822 ( 
.A(n_3155),
.B(n_3174),
.Y(n_3822)
);

BUFx2_ASAP7_75t_L g3823 ( 
.A(n_3122),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_L g3824 ( 
.A(n_3455),
.B(n_3459),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_L g3825 ( 
.A(n_3462),
.B(n_3467),
.Y(n_3825)
);

NAND2x1p5_ASAP7_75t_L g3826 ( 
.A(n_3513),
.B(n_3302),
.Y(n_3826)
);

INVx5_ASAP7_75t_L g3827 ( 
.A(n_3120),
.Y(n_3827)
);

INVx6_ASAP7_75t_L g3828 ( 
.A(n_3120),
.Y(n_3828)
);

INVx2_ASAP7_75t_L g3829 ( 
.A(n_3394),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_L g3830 ( 
.A(n_3462),
.B(n_3467),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_L g3831 ( 
.A(n_3470),
.B(n_3486),
.Y(n_3831)
);

AND2x2_ASAP7_75t_L g3832 ( 
.A(n_3047),
.B(n_3048),
.Y(n_3832)
);

BUFx2_ASAP7_75t_L g3833 ( 
.A(n_3256),
.Y(n_3833)
);

BUFx3_ASAP7_75t_L g3834 ( 
.A(n_3193),
.Y(n_3834)
);

HB1xp67_ASAP7_75t_L g3835 ( 
.A(n_3331),
.Y(n_3835)
);

INVx1_ASAP7_75t_L g3836 ( 
.A(n_3350),
.Y(n_3836)
);

AO21x2_ASAP7_75t_L g3837 ( 
.A1(n_3076),
.A2(n_3180),
.B(n_3169),
.Y(n_3837)
);

HB1xp67_ASAP7_75t_L g3838 ( 
.A(n_3027),
.Y(n_3838)
);

BUFx4f_ASAP7_75t_L g3839 ( 
.A(n_3086),
.Y(n_3839)
);

INVxp67_ASAP7_75t_SL g3840 ( 
.A(n_3036),
.Y(n_3840)
);

INVx6_ASAP7_75t_L g3841 ( 
.A(n_3133),
.Y(n_3841)
);

BUFx10_ASAP7_75t_L g3842 ( 
.A(n_3139),
.Y(n_3842)
);

INVx1_ASAP7_75t_SL g3843 ( 
.A(n_3290),
.Y(n_3843)
);

INVx3_ASAP7_75t_SL g3844 ( 
.A(n_3388),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_L g3845 ( 
.A(n_3470),
.B(n_3486),
.Y(n_3845)
);

INVx3_ASAP7_75t_L g3846 ( 
.A(n_3537),
.Y(n_3846)
);

BUFx3_ASAP7_75t_L g3847 ( 
.A(n_3105),
.Y(n_3847)
);

AND2x2_ASAP7_75t_L g3848 ( 
.A(n_3047),
.B(n_3048),
.Y(n_3848)
);

BUFx4f_ASAP7_75t_L g3849 ( 
.A(n_3086),
.Y(n_3849)
);

INVx3_ASAP7_75t_L g3850 ( 
.A(n_3569),
.Y(n_3850)
);

INVxp67_ASAP7_75t_SL g3851 ( 
.A(n_3027),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_3395),
.Y(n_3852)
);

OR2x2_ASAP7_75t_L g3853 ( 
.A(n_3181),
.B(n_3029),
.Y(n_3853)
);

NAND2xp5_ASAP7_75t_L g3854 ( 
.A(n_3496),
.B(n_3504),
.Y(n_3854)
);

INVx3_ASAP7_75t_L g3855 ( 
.A(n_3569),
.Y(n_3855)
);

HB1xp67_ASAP7_75t_L g3856 ( 
.A(n_3336),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_L g3857 ( 
.A(n_3496),
.B(n_3504),
.Y(n_3857)
);

AND2x4_ASAP7_75t_L g3858 ( 
.A(n_3569),
.B(n_3596),
.Y(n_3858)
);

BUFx2_ASAP7_75t_SL g3859 ( 
.A(n_3464),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_3312),
.Y(n_3860)
);

BUFx2_ASAP7_75t_SL g3861 ( 
.A(n_3553),
.Y(n_3861)
);

INVx8_ASAP7_75t_L g3862 ( 
.A(n_3133),
.Y(n_3862)
);

CKINVDCx5p33_ASAP7_75t_R g3863 ( 
.A(n_3124),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_3312),
.Y(n_3864)
);

INVx3_ASAP7_75t_L g3865 ( 
.A(n_3569),
.Y(n_3865)
);

BUFx4f_ASAP7_75t_SL g3866 ( 
.A(n_3393),
.Y(n_3866)
);

CKINVDCx14_ASAP7_75t_R g3867 ( 
.A(n_3423),
.Y(n_3867)
);

BUFx3_ASAP7_75t_L g3868 ( 
.A(n_3105),
.Y(n_3868)
);

BUFx2_ASAP7_75t_R g3869 ( 
.A(n_3051),
.Y(n_3869)
);

AND2x2_ASAP7_75t_L g3870 ( 
.A(n_3275),
.B(n_3317),
.Y(n_3870)
);

AND2x2_ASAP7_75t_L g3871 ( 
.A(n_3275),
.B(n_3317),
.Y(n_3871)
);

INVx3_ASAP7_75t_L g3872 ( 
.A(n_3596),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_3507),
.B(n_3512),
.Y(n_3873)
);

BUFx6f_ASAP7_75t_L g3874 ( 
.A(n_3121),
.Y(n_3874)
);

CKINVDCx11_ASAP7_75t_R g3875 ( 
.A(n_3423),
.Y(n_3875)
);

INVx6_ASAP7_75t_SL g3876 ( 
.A(n_3133),
.Y(n_3876)
);

BUFx2_ASAP7_75t_L g3877 ( 
.A(n_3256),
.Y(n_3877)
);

AND2x2_ASAP7_75t_L g3878 ( 
.A(n_3239),
.B(n_3308),
.Y(n_3878)
);

INVx8_ASAP7_75t_L g3879 ( 
.A(n_3133),
.Y(n_3879)
);

INVx3_ASAP7_75t_SL g3880 ( 
.A(n_3149),
.Y(n_3880)
);

INVx3_ASAP7_75t_SL g3881 ( 
.A(n_3419),
.Y(n_3881)
);

INVx3_ASAP7_75t_L g3882 ( 
.A(n_3596),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3319),
.Y(n_3883)
);

NOR2xp33_ASAP7_75t_L g3884 ( 
.A(n_3042),
.B(n_3515),
.Y(n_3884)
);

INVx5_ASAP7_75t_L g3885 ( 
.A(n_3133),
.Y(n_3885)
);

BUFx4f_ASAP7_75t_SL g3886 ( 
.A(n_3393),
.Y(n_3886)
);

BUFx4f_ASAP7_75t_L g3887 ( 
.A(n_3144),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_L g3888 ( 
.A(n_3507),
.B(n_3512),
.Y(n_3888)
);

CKINVDCx8_ASAP7_75t_R g3889 ( 
.A(n_3257),
.Y(n_3889)
);

INVx1_ASAP7_75t_SL g3890 ( 
.A(n_3524),
.Y(n_3890)
);

BUFx6f_ASAP7_75t_L g3891 ( 
.A(n_3121),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_L g3892 ( 
.A(n_3525),
.B(n_3527),
.Y(n_3892)
);

INVx6_ASAP7_75t_L g3893 ( 
.A(n_3302),
.Y(n_3893)
);

INVxp67_ASAP7_75t_SL g3894 ( 
.A(n_3062),
.Y(n_3894)
);

INVx1_ASAP7_75t_L g3895 ( 
.A(n_3319),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3322),
.Y(n_3896)
);

INVx2_ASAP7_75t_SL g3897 ( 
.A(n_3071),
.Y(n_3897)
);

BUFx2_ASAP7_75t_L g3898 ( 
.A(n_3524),
.Y(n_3898)
);

HB1xp67_ASAP7_75t_L g3899 ( 
.A(n_3336),
.Y(n_3899)
);

CKINVDCx5p33_ASAP7_75t_R g3900 ( 
.A(n_3346),
.Y(n_3900)
);

INVx1_ASAP7_75t_SL g3901 ( 
.A(n_3532),
.Y(n_3901)
);

AND2x2_ASAP7_75t_L g3902 ( 
.A(n_3239),
.B(n_3308),
.Y(n_3902)
);

INVx2_ASAP7_75t_SL g3903 ( 
.A(n_3071),
.Y(n_3903)
);

INVx1_ASAP7_75t_L g3904 ( 
.A(n_3322),
.Y(n_3904)
);

INVx3_ASAP7_75t_L g3905 ( 
.A(n_3596),
.Y(n_3905)
);

CKINVDCx20_ASAP7_75t_R g3906 ( 
.A(n_3429),
.Y(n_3906)
);

INVx5_ASAP7_75t_L g3907 ( 
.A(n_3407),
.Y(n_3907)
);

AND2x2_ASAP7_75t_L g3908 ( 
.A(n_3182),
.B(n_3006),
.Y(n_3908)
);

INVx2_ASAP7_75t_SL g3909 ( 
.A(n_3337),
.Y(n_3909)
);

INVx5_ASAP7_75t_L g3910 ( 
.A(n_3407),
.Y(n_3910)
);

BUFx2_ASAP7_75t_L g3911 ( 
.A(n_3532),
.Y(n_3911)
);

INVx1_ASAP7_75t_L g3912 ( 
.A(n_3327),
.Y(n_3912)
);

AND2x4_ASAP7_75t_L g3913 ( 
.A(n_3337),
.B(n_3345),
.Y(n_3913)
);

BUFx4_ASAP7_75t_SL g3914 ( 
.A(n_3494),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3327),
.Y(n_3915)
);

INVx8_ASAP7_75t_L g3916 ( 
.A(n_3093),
.Y(n_3916)
);

INVx3_ASAP7_75t_L g3917 ( 
.A(n_3077),
.Y(n_3917)
);

OR2x2_ASAP7_75t_L g3918 ( 
.A(n_3451),
.B(n_3518),
.Y(n_3918)
);

INVx5_ASAP7_75t_L g3919 ( 
.A(n_3407),
.Y(n_3919)
);

NAND2xp5_ASAP7_75t_SL g3920 ( 
.A(n_3023),
.B(n_3553),
.Y(n_3920)
);

OR2x6_ASAP7_75t_L g3921 ( 
.A(n_3567),
.B(n_3187),
.Y(n_3921)
);

AND2x2_ASAP7_75t_L g3922 ( 
.A(n_3182),
.B(n_3006),
.Y(n_3922)
);

BUFx2_ASAP7_75t_SL g3923 ( 
.A(n_3017),
.Y(n_3923)
);

BUFx2_ASAP7_75t_L g3924 ( 
.A(n_3546),
.Y(n_3924)
);

INVx1_ASAP7_75t_SL g3925 ( 
.A(n_3546),
.Y(n_3925)
);

INVx6_ASAP7_75t_L g3926 ( 
.A(n_3093),
.Y(n_3926)
);

NOR2x1_ASAP7_75t_L g3927 ( 
.A(n_3557),
.B(n_3131),
.Y(n_3927)
);

AND2x2_ASAP7_75t_L g3928 ( 
.A(n_3018),
.B(n_3458),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_L g3929 ( 
.A(n_3525),
.B(n_3527),
.Y(n_3929)
);

BUFx2_ASAP7_75t_SL g3930 ( 
.A(n_3429),
.Y(n_3930)
);

INVx2_ASAP7_75t_SL g3931 ( 
.A(n_3337),
.Y(n_3931)
);

AOI22xp33_ASAP7_75t_L g3932 ( 
.A1(n_3024),
.A2(n_3576),
.B1(n_3580),
.B2(n_3545),
.Y(n_3932)
);

CKINVDCx20_ASAP7_75t_R g3933 ( 
.A(n_3358),
.Y(n_3933)
);

CKINVDCx5p33_ASAP7_75t_R g3934 ( 
.A(n_3206),
.Y(n_3934)
);

AND2x2_ASAP7_75t_L g3935 ( 
.A(n_3018),
.B(n_3458),
.Y(n_3935)
);

INVxp67_ASAP7_75t_SL g3936 ( 
.A(n_3062),
.Y(n_3936)
);

INVx6_ASAP7_75t_L g3937 ( 
.A(n_3096),
.Y(n_3937)
);

CKINVDCx14_ASAP7_75t_R g3938 ( 
.A(n_3247),
.Y(n_3938)
);

INVx1_ASAP7_75t_SL g3939 ( 
.A(n_3552),
.Y(n_3939)
);

INVxp67_ASAP7_75t_SL g3940 ( 
.A(n_3065),
.Y(n_3940)
);

AOI22xp33_ASAP7_75t_L g3941 ( 
.A1(n_3545),
.A2(n_3580),
.B1(n_3576),
.B2(n_3442),
.Y(n_3941)
);

BUFx3_ASAP7_75t_L g3942 ( 
.A(n_3407),
.Y(n_3942)
);

INVx3_ASAP7_75t_SL g3943 ( 
.A(n_3419),
.Y(n_3943)
);

INVx3_ASAP7_75t_L g3944 ( 
.A(n_3085),
.Y(n_3944)
);

INVx3_ASAP7_75t_L g3945 ( 
.A(n_3085),
.Y(n_3945)
);

BUFx10_ASAP7_75t_L g3946 ( 
.A(n_3158),
.Y(n_3946)
);

HB1xp67_ASAP7_75t_L g3947 ( 
.A(n_3339),
.Y(n_3947)
);

INVx2_ASAP7_75t_L g3948 ( 
.A(n_3110),
.Y(n_3948)
);

CKINVDCx16_ASAP7_75t_R g3949 ( 
.A(n_3337),
.Y(n_3949)
);

CKINVDCx5p33_ASAP7_75t_R g3950 ( 
.A(n_3088),
.Y(n_3950)
);

BUFx8_ASAP7_75t_SL g3951 ( 
.A(n_3438),
.Y(n_3951)
);

INVx8_ASAP7_75t_L g3952 ( 
.A(n_3104),
.Y(n_3952)
);

INVx2_ASAP7_75t_SL g3953 ( 
.A(n_3345),
.Y(n_3953)
);

BUFx4f_ASAP7_75t_SL g3954 ( 
.A(n_3405),
.Y(n_3954)
);

BUFx4f_ASAP7_75t_SL g3955 ( 
.A(n_3405),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3536),
.B(n_3547),
.Y(n_3956)
);

BUFx4f_ASAP7_75t_L g3957 ( 
.A(n_3144),
.Y(n_3957)
);

INVx2_ASAP7_75t_L g3958 ( 
.A(n_3110),
.Y(n_3958)
);

INVxp67_ASAP7_75t_SL g3959 ( 
.A(n_3065),
.Y(n_3959)
);

AND2x2_ASAP7_75t_L g3960 ( 
.A(n_3480),
.B(n_3587),
.Y(n_3960)
);

INVx1_ASAP7_75t_SL g3961 ( 
.A(n_3438),
.Y(n_3961)
);

CKINVDCx5p33_ASAP7_75t_R g3962 ( 
.A(n_3207),
.Y(n_3962)
);

INVx2_ASAP7_75t_SL g3963 ( 
.A(n_3345),
.Y(n_3963)
);

BUFx4f_ASAP7_75t_SL g3964 ( 
.A(n_3329),
.Y(n_3964)
);

INVx2_ASAP7_75t_L g3965 ( 
.A(n_3110),
.Y(n_3965)
);

BUFx4f_ASAP7_75t_SL g3966 ( 
.A(n_3342),
.Y(n_3966)
);

BUFx3_ASAP7_75t_L g3967 ( 
.A(n_3407),
.Y(n_3967)
);

INVx2_ASAP7_75t_SL g3968 ( 
.A(n_3345),
.Y(n_3968)
);

BUFx2_ASAP7_75t_L g3969 ( 
.A(n_3332),
.Y(n_3969)
);

BUFx2_ASAP7_75t_L g3970 ( 
.A(n_3332),
.Y(n_3970)
);

AOI22xp33_ASAP7_75t_L g3971 ( 
.A1(n_3483),
.A2(n_3442),
.B1(n_3514),
.B2(n_3491),
.Y(n_3971)
);

BUFx2_ASAP7_75t_L g3972 ( 
.A(n_3332),
.Y(n_3972)
);

OR2x6_ASAP7_75t_L g3973 ( 
.A(n_3567),
.B(n_3187),
.Y(n_3973)
);

CKINVDCx14_ASAP7_75t_R g3974 ( 
.A(n_3051),
.Y(n_3974)
);

INVxp67_ASAP7_75t_SL g3975 ( 
.A(n_3222),
.Y(n_3975)
);

INVx2_ASAP7_75t_SL g3976 ( 
.A(n_3356),
.Y(n_3976)
);

BUFx4_ASAP7_75t_SL g3977 ( 
.A(n_3432),
.Y(n_3977)
);

NOR2xp33_ASAP7_75t_L g3978 ( 
.A(n_3128),
.B(n_3112),
.Y(n_3978)
);

INVx6_ASAP7_75t_SL g3979 ( 
.A(n_3187),
.Y(n_3979)
);

BUFx2_ASAP7_75t_L g3980 ( 
.A(n_3283),
.Y(n_3980)
);

BUFx2_ASAP7_75t_SL g3981 ( 
.A(n_3402),
.Y(n_3981)
);

CKINVDCx8_ASAP7_75t_R g3982 ( 
.A(n_3090),
.Y(n_3982)
);

INVx2_ASAP7_75t_SL g3983 ( 
.A(n_3356),
.Y(n_3983)
);

INVx1_ASAP7_75t_L g3984 ( 
.A(n_3339),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3409),
.Y(n_3985)
);

BUFx2_ASAP7_75t_L g3986 ( 
.A(n_3283),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3409),
.Y(n_3987)
);

BUFx3_ASAP7_75t_L g3988 ( 
.A(n_3117),
.Y(n_3988)
);

INVx6_ASAP7_75t_L g3989 ( 
.A(n_3468),
.Y(n_3989)
);

OR2x6_ASAP7_75t_L g3990 ( 
.A(n_3187),
.B(n_3213),
.Y(n_3990)
);

NOR2x1_ASAP7_75t_R g3991 ( 
.A(n_3185),
.B(n_3210),
.Y(n_3991)
);

NAND2xp5_ASAP7_75t_L g3992 ( 
.A(n_3536),
.B(n_3547),
.Y(n_3992)
);

CKINVDCx11_ASAP7_75t_R g3993 ( 
.A(n_3216),
.Y(n_3993)
);

INVx5_ASAP7_75t_L g3994 ( 
.A(n_3187),
.Y(n_3994)
);

INVx1_ASAP7_75t_L g3995 ( 
.A(n_3410),
.Y(n_3995)
);

BUFx2_ASAP7_75t_L g3996 ( 
.A(n_3171),
.Y(n_3996)
);

AND2x2_ASAP7_75t_L g3997 ( 
.A(n_3480),
.B(n_3587),
.Y(n_3997)
);

INVx2_ASAP7_75t_L g3998 ( 
.A(n_3127),
.Y(n_3998)
);

BUFx3_ASAP7_75t_L g3999 ( 
.A(n_3117),
.Y(n_3999)
);

BUFx3_ASAP7_75t_L g4000 ( 
.A(n_3196),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_3349),
.Y(n_4001)
);

BUFx4_ASAP7_75t_SL g4002 ( 
.A(n_3069),
.Y(n_4002)
);

INVx2_ASAP7_75t_L g4003 ( 
.A(n_3127),
.Y(n_4003)
);

INVxp67_ASAP7_75t_L g4004 ( 
.A(n_3557),
.Y(n_4004)
);

INVx2_ASAP7_75t_L g4005 ( 
.A(n_3127),
.Y(n_4005)
);

BUFx2_ASAP7_75t_L g4006 ( 
.A(n_3223),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3349),
.Y(n_4007)
);

BUFx2_ASAP7_75t_SL g4008 ( 
.A(n_3202),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_L g4009 ( 
.A(n_3551),
.B(n_3556),
.Y(n_4009)
);

NAND2xp5_ASAP7_75t_L g4010 ( 
.A(n_3551),
.B(n_3556),
.Y(n_4010)
);

INVx2_ASAP7_75t_SL g4011 ( 
.A(n_3356),
.Y(n_4011)
);

AND2x2_ASAP7_75t_L g4012 ( 
.A(n_3209),
.B(n_3177),
.Y(n_4012)
);

BUFx2_ASAP7_75t_L g4013 ( 
.A(n_3223),
.Y(n_4013)
);

BUFx3_ASAP7_75t_L g4014 ( 
.A(n_3196),
.Y(n_4014)
);

BUFx4_ASAP7_75t_SL g4015 ( 
.A(n_3451),
.Y(n_4015)
);

BUFx3_ASAP7_75t_L g4016 ( 
.A(n_3198),
.Y(n_4016)
);

INVx4_ASAP7_75t_L g4017 ( 
.A(n_3396),
.Y(n_4017)
);

BUFx3_ASAP7_75t_L g4018 ( 
.A(n_3198),
.Y(n_4018)
);

INVx2_ASAP7_75t_L g4019 ( 
.A(n_3148),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_3212),
.Y(n_4020)
);

INVx4_ASAP7_75t_L g4021 ( 
.A(n_3396),
.Y(n_4021)
);

CKINVDCx16_ASAP7_75t_R g4022 ( 
.A(n_3356),
.Y(n_4022)
);

NAND2xp5_ASAP7_75t_L g4023 ( 
.A(n_3560),
.B(n_3566),
.Y(n_4023)
);

AOI22xp33_ASAP7_75t_L g4024 ( 
.A1(n_3483),
.A2(n_3514),
.B1(n_3491),
.B2(n_2996),
.Y(n_4024)
);

NOR2xp33_ASAP7_75t_L g4025 ( 
.A(n_3128),
.B(n_3188),
.Y(n_4025)
);

NOR2xp33_ASAP7_75t_L g4026 ( 
.A(n_3146),
.B(n_3168),
.Y(n_4026)
);

INVx5_ASAP7_75t_L g4027 ( 
.A(n_3213),
.Y(n_4027)
);

INVx1_ASAP7_75t_SL g4028 ( 
.A(n_3137),
.Y(n_4028)
);

INVx2_ASAP7_75t_L g4029 ( 
.A(n_3148),
.Y(n_4029)
);

AO22x2_ASAP7_75t_L g4030 ( 
.A1(n_3591),
.A2(n_3521),
.B1(n_3154),
.B2(n_3173),
.Y(n_4030)
);

BUFx2_ASAP7_75t_L g4031 ( 
.A(n_3118),
.Y(n_4031)
);

INVx2_ASAP7_75t_L g4032 ( 
.A(n_3148),
.Y(n_4032)
);

OR2x6_ASAP7_75t_L g4033 ( 
.A(n_3213),
.B(n_3250),
.Y(n_4033)
);

BUFx2_ASAP7_75t_L g4034 ( 
.A(n_3118),
.Y(n_4034)
);

INVx1_ASAP7_75t_L g4035 ( 
.A(n_3347),
.Y(n_4035)
);

INVx8_ASAP7_75t_L g4036 ( 
.A(n_3213),
.Y(n_4036)
);

INVx1_ASAP7_75t_L g4037 ( 
.A(n_3347),
.Y(n_4037)
);

INVx4_ASAP7_75t_L g4038 ( 
.A(n_3396),
.Y(n_4038)
);

AOI22xp5_ASAP7_75t_L g4039 ( 
.A1(n_3543),
.A2(n_3563),
.B1(n_3054),
.B2(n_2996),
.Y(n_4039)
);

INVx1_ASAP7_75t_SL g4040 ( 
.A(n_3137),
.Y(n_4040)
);

NOR2xp33_ASAP7_75t_L g4041 ( 
.A(n_3146),
.B(n_3168),
.Y(n_4041)
);

BUFx2_ASAP7_75t_L g4042 ( 
.A(n_3214),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_L g4043 ( 
.A(n_3560),
.B(n_3566),
.Y(n_4043)
);

INVx8_ASAP7_75t_L g4044 ( 
.A(n_3213),
.Y(n_4044)
);

INVx1_ASAP7_75t_L g4045 ( 
.A(n_3364),
.Y(n_4045)
);

INVx1_ASAP7_75t_SL g4046 ( 
.A(n_3179),
.Y(n_4046)
);

INVx2_ASAP7_75t_SL g4047 ( 
.A(n_3324),
.Y(n_4047)
);

NAND2xp5_ASAP7_75t_L g4048 ( 
.A(n_3570),
.B(n_3575),
.Y(n_4048)
);

INVx2_ASAP7_75t_SL g4049 ( 
.A(n_3324),
.Y(n_4049)
);

INVx2_ASAP7_75t_SL g4050 ( 
.A(n_3357),
.Y(n_4050)
);

BUFx4f_ASAP7_75t_L g4051 ( 
.A(n_3164),
.Y(n_4051)
);

INVx1_ASAP7_75t_SL g4052 ( 
.A(n_3179),
.Y(n_4052)
);

INVx1_ASAP7_75t_L g4053 ( 
.A(n_3364),
.Y(n_4053)
);

HB1xp67_ASAP7_75t_L g4054 ( 
.A(n_3082),
.Y(n_4054)
);

INVx3_ASAP7_75t_SL g4055 ( 
.A(n_3419),
.Y(n_4055)
);

INVx8_ASAP7_75t_L g4056 ( 
.A(n_3255),
.Y(n_4056)
);

INVx6_ASAP7_75t_SL g4057 ( 
.A(n_2994),
.Y(n_4057)
);

BUFx2_ASAP7_75t_L g4058 ( 
.A(n_3214),
.Y(n_4058)
);

CKINVDCx5p33_ASAP7_75t_R g4059 ( 
.A(n_3216),
.Y(n_4059)
);

NAND2x1p5_ASAP7_75t_L g4060 ( 
.A(n_3465),
.B(n_3156),
.Y(n_4060)
);

INVx2_ASAP7_75t_L g4061 ( 
.A(n_3163),
.Y(n_4061)
);

NOR2xp33_ASAP7_75t_L g4062 ( 
.A(n_3472),
.B(n_3074),
.Y(n_4062)
);

INVx5_ASAP7_75t_L g4063 ( 
.A(n_3465),
.Y(n_4063)
);

INVx5_ASAP7_75t_L g4064 ( 
.A(n_3465),
.Y(n_4064)
);

AOI22xp33_ASAP7_75t_L g4065 ( 
.A1(n_3004),
.A2(n_3060),
.B1(n_3057),
.B2(n_3033),
.Y(n_4065)
);

BUFx3_ASAP7_75t_L g4066 ( 
.A(n_3488),
.Y(n_4066)
);

INVx2_ASAP7_75t_L g4067 ( 
.A(n_3163),
.Y(n_4067)
);

INVx6_ASAP7_75t_L g4068 ( 
.A(n_3255),
.Y(n_4068)
);

BUFx3_ASAP7_75t_L g4069 ( 
.A(n_3488),
.Y(n_4069)
);

INVx2_ASAP7_75t_L g4070 ( 
.A(n_3163),
.Y(n_4070)
);

BUFx4f_ASAP7_75t_SL g4071 ( 
.A(n_3426),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_L g4072 ( 
.A(n_3570),
.B(n_3575),
.Y(n_4072)
);

INVx2_ASAP7_75t_SL g4073 ( 
.A(n_3357),
.Y(n_4073)
);

AOI22xp33_ASAP7_75t_L g4074 ( 
.A1(n_3004),
.A2(n_3060),
.B1(n_3057),
.B2(n_3033),
.Y(n_4074)
);

INVx2_ASAP7_75t_SL g4075 ( 
.A(n_3359),
.Y(n_4075)
);

NAND2xp5_ASAP7_75t_L g4076 ( 
.A(n_3586),
.B(n_3592),
.Y(n_4076)
);

AND2x2_ASAP7_75t_L g4077 ( 
.A(n_3209),
.B(n_3177),
.Y(n_4077)
);

BUFx2_ASAP7_75t_L g4078 ( 
.A(n_3225),
.Y(n_4078)
);

AND2x2_ASAP7_75t_L g4079 ( 
.A(n_3143),
.B(n_3160),
.Y(n_4079)
);

AOI22xp33_ASAP7_75t_L g4080 ( 
.A1(n_3032),
.A2(n_3100),
.B1(n_3000),
.B2(n_3444),
.Y(n_4080)
);

INVx2_ASAP7_75t_L g4081 ( 
.A(n_3167),
.Y(n_4081)
);

BUFx2_ASAP7_75t_L g4082 ( 
.A(n_3225),
.Y(n_4082)
);

BUFx2_ASAP7_75t_R g4083 ( 
.A(n_3141),
.Y(n_4083)
);

NAND2xp5_ASAP7_75t_SL g4084 ( 
.A(n_3543),
.B(n_3563),
.Y(n_4084)
);

BUFx3_ASAP7_75t_L g4085 ( 
.A(n_3488),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_L g4086 ( 
.A(n_3586),
.B(n_3592),
.Y(n_4086)
);

INVx5_ASAP7_75t_SL g4087 ( 
.A(n_3482),
.Y(n_4087)
);

NAND2x1p5_ASAP7_75t_L g4088 ( 
.A(n_3156),
.B(n_3140),
.Y(n_4088)
);

INVx1_ASAP7_75t_SL g4089 ( 
.A(n_3518),
.Y(n_4089)
);

BUFx4f_ASAP7_75t_SL g4090 ( 
.A(n_3426),
.Y(n_4090)
);

BUFx3_ASAP7_75t_L g4091 ( 
.A(n_3488),
.Y(n_4091)
);

INVx1_ASAP7_75t_SL g4092 ( 
.A(n_3600),
.Y(n_4092)
);

BUFx3_ASAP7_75t_L g4093 ( 
.A(n_3562),
.Y(n_4093)
);

OR2x2_ASAP7_75t_L g4094 ( 
.A(n_3600),
.B(n_3318),
.Y(n_4094)
);

BUFx2_ASAP7_75t_SL g4095 ( 
.A(n_3186),
.Y(n_4095)
);

BUFx3_ASAP7_75t_L g4096 ( 
.A(n_3562),
.Y(n_4096)
);

BUFx3_ASAP7_75t_L g4097 ( 
.A(n_3562),
.Y(n_4097)
);

INVxp67_ASAP7_75t_SL g4098 ( 
.A(n_3222),
.Y(n_4098)
);

CKINVDCx20_ASAP7_75t_R g4099 ( 
.A(n_3218),
.Y(n_4099)
);

INVx1_ASAP7_75t_SL g4100 ( 
.A(n_3318),
.Y(n_4100)
);

BUFx2_ASAP7_75t_SL g4101 ( 
.A(n_3192),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_3403),
.Y(n_4102)
);

BUFx2_ASAP7_75t_R g4103 ( 
.A(n_3053),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_3403),
.Y(n_4104)
);

INVxp67_ASAP7_75t_SL g4105 ( 
.A(n_3049),
.Y(n_4105)
);

BUFx2_ASAP7_75t_L g4106 ( 
.A(n_3265),
.Y(n_4106)
);

INVx3_ASAP7_75t_SL g4107 ( 
.A(n_3404),
.Y(n_4107)
);

INVx1_ASAP7_75t_L g4108 ( 
.A(n_3240),
.Y(n_4108)
);

AND2x2_ASAP7_75t_L g4109 ( 
.A(n_3143),
.B(n_3160),
.Y(n_4109)
);

NAND2x1p5_ASAP7_75t_L g4110 ( 
.A(n_3140),
.B(n_3161),
.Y(n_4110)
);

INVx3_ASAP7_75t_SL g4111 ( 
.A(n_3415),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_3603),
.B(n_3609),
.Y(n_4112)
);

INVx2_ASAP7_75t_SL g4113 ( 
.A(n_3359),
.Y(n_4113)
);

INVx8_ASAP7_75t_L g4114 ( 
.A(n_3255),
.Y(n_4114)
);

CKINVDCx20_ASAP7_75t_R g4115 ( 
.A(n_3218),
.Y(n_4115)
);

BUFx2_ASAP7_75t_L g4116 ( 
.A(n_3265),
.Y(n_4116)
);

AND2x2_ASAP7_75t_L g4117 ( 
.A(n_3300),
.B(n_3416),
.Y(n_4117)
);

INVx3_ASAP7_75t_L g4118 ( 
.A(n_3219),
.Y(n_4118)
);

AND2x2_ASAP7_75t_L g4119 ( 
.A(n_3300),
.B(n_3416),
.Y(n_4119)
);

INVx2_ASAP7_75t_SL g4120 ( 
.A(n_3263),
.Y(n_4120)
);

AOI22xp33_ASAP7_75t_L g4121 ( 
.A1(n_3032),
.A2(n_3100),
.B1(n_3448),
.B2(n_3444),
.Y(n_4121)
);

BUFx3_ASAP7_75t_L g4122 ( 
.A(n_3562),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_3240),
.Y(n_4123)
);

BUFx3_ASAP7_75t_L g4124 ( 
.A(n_3562),
.Y(n_4124)
);

NAND2xp5_ASAP7_75t_L g4125 ( 
.A(n_3603),
.B(n_3609),
.Y(n_4125)
);

INVx2_ASAP7_75t_L g4126 ( 
.A(n_3167),
.Y(n_4126)
);

INVx1_ASAP7_75t_L g4127 ( 
.A(n_3240),
.Y(n_4127)
);

CKINVDCx20_ASAP7_75t_R g4128 ( 
.A(n_3340),
.Y(n_4128)
);

INVx1_ASAP7_75t_L g4129 ( 
.A(n_3240),
.Y(n_4129)
);

AOI21xp5_ASAP7_75t_L g4130 ( 
.A1(n_3645),
.A2(n_3041),
.B(n_3008),
.Y(n_4130)
);

OAI22xp5_ASAP7_75t_L g4131 ( 
.A1(n_3932),
.A2(n_3015),
.B1(n_3485),
.B2(n_3460),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_3646),
.Y(n_4132)
);

OR2x2_ASAP7_75t_L g4133 ( 
.A(n_3853),
.B(n_3351),
.Y(n_4133)
);

OAI21xp5_ASAP7_75t_L g4134 ( 
.A1(n_3794),
.A2(n_3045),
.B(n_3016),
.Y(n_4134)
);

OAI21xp5_ASAP7_75t_L g4135 ( 
.A1(n_3794),
.A2(n_3016),
.B(n_3516),
.Y(n_4135)
);

AND2x2_ASAP7_75t_L g4136 ( 
.A(n_3870),
.B(n_3155),
.Y(n_4136)
);

INVx1_ASAP7_75t_L g4137 ( 
.A(n_3646),
.Y(n_4137)
);

AOI22xp33_ASAP7_75t_L g4138 ( 
.A1(n_3615),
.A2(n_3307),
.B1(n_3022),
.B2(n_3224),
.Y(n_4138)
);

BUFx6f_ASAP7_75t_L g4139 ( 
.A(n_3611),
.Y(n_4139)
);

NAND2xp5_ASAP7_75t_L g4140 ( 
.A(n_3650),
.B(n_3114),
.Y(n_4140)
);

NOR3xp33_ASAP7_75t_SL g4141 ( 
.A(n_3634),
.B(n_3531),
.C(n_3517),
.Y(n_4141)
);

AOI21xp5_ASAP7_75t_SL g4142 ( 
.A1(n_3920),
.A2(n_3052),
.B(n_3448),
.Y(n_4142)
);

NOR2xp67_ASAP7_75t_L g4143 ( 
.A(n_3838),
.B(n_3078),
.Y(n_4143)
);

AOI22xp33_ASAP7_75t_SL g4144 ( 
.A1(n_3923),
.A2(n_3307),
.B1(n_3022),
.B2(n_3221),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_3662),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_3662),
.Y(n_4146)
);

INVx1_ASAP7_75t_SL g4147 ( 
.A(n_4015),
.Y(n_4147)
);

NAND3x1_ASAP7_75t_L g4148 ( 
.A(n_3927),
.B(n_3478),
.C(n_3457),
.Y(n_4148)
);

AOI21x1_ASAP7_75t_L g4149 ( 
.A1(n_4006),
.A2(n_3084),
.B(n_3037),
.Y(n_4149)
);

AOI21xp5_ASAP7_75t_L g4150 ( 
.A1(n_3927),
.A2(n_3025),
.B(n_3001),
.Y(n_4150)
);

OAI21x1_ASAP7_75t_L g4151 ( 
.A1(n_4110),
.A2(n_4088),
.B(n_3945),
.Y(n_4151)
);

OAI21xp5_ASAP7_75t_L g4152 ( 
.A1(n_4039),
.A2(n_3572),
.B(n_3534),
.Y(n_4152)
);

OAI21xp5_ASAP7_75t_L g4153 ( 
.A1(n_4039),
.A2(n_3604),
.B(n_3593),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_L g4154 ( 
.A(n_3650),
.B(n_3114),
.Y(n_4154)
);

OR2x2_ASAP7_75t_L g4155 ( 
.A(n_3853),
.B(n_3392),
.Y(n_4155)
);

AOI21xp5_ASAP7_75t_L g4156 ( 
.A1(n_3669),
.A2(n_3040),
.B(n_3501),
.Y(n_4156)
);

AOI21xp5_ASAP7_75t_L g4157 ( 
.A1(n_3669),
.A2(n_3505),
.B(n_3501),
.Y(n_4157)
);

AND2x4_ASAP7_75t_L g4158 ( 
.A(n_3629),
.B(n_3263),
.Y(n_4158)
);

AND2x2_ASAP7_75t_L g4159 ( 
.A(n_3870),
.B(n_3174),
.Y(n_4159)
);

OR2x6_ASAP7_75t_L g4160 ( 
.A(n_3862),
.B(n_3250),
.Y(n_4160)
);

INVx4_ASAP7_75t_SL g4161 ( 
.A(n_3881),
.Y(n_4161)
);

INVxp67_ASAP7_75t_L g4162 ( 
.A(n_3884),
.Y(n_4162)
);

OAI21x1_ASAP7_75t_L g4163 ( 
.A1(n_4088),
.A2(n_3945),
.B(n_3944),
.Y(n_4163)
);

OAI21xp5_ASAP7_75t_L g4164 ( 
.A1(n_4084),
.A2(n_3610),
.B(n_3073),
.Y(n_4164)
);

OAI22xp5_ASAP7_75t_L g4165 ( 
.A1(n_3932),
.A2(n_3591),
.B1(n_3457),
.B2(n_3481),
.Y(n_4165)
);

AOI22xp33_ASAP7_75t_L g4166 ( 
.A1(n_3615),
.A2(n_3307),
.B1(n_3923),
.B2(n_4030),
.Y(n_4166)
);

OAI21xp5_ASAP7_75t_L g4167 ( 
.A1(n_4065),
.A2(n_3073),
.B(n_3454),
.Y(n_4167)
);

NAND2x1p5_ASAP7_75t_L g4168 ( 
.A(n_3643),
.B(n_3165),
.Y(n_4168)
);

AOI21xp5_ASAP7_75t_L g4169 ( 
.A1(n_3672),
.A2(n_3506),
.B(n_3505),
.Y(n_4169)
);

INVx3_ASAP7_75t_L g4170 ( 
.A(n_3765),
.Y(n_4170)
);

AND2x2_ASAP7_75t_L g4171 ( 
.A(n_3870),
.B(n_3244),
.Y(n_4171)
);

INVx1_ASAP7_75t_L g4172 ( 
.A(n_3666),
.Y(n_4172)
);

INVx3_ASAP7_75t_L g4173 ( 
.A(n_3765),
.Y(n_4173)
);

OAI21x1_ASAP7_75t_SL g4174 ( 
.A1(n_3733),
.A2(n_3481),
.B(n_3478),
.Y(n_4174)
);

AOI22xp33_ASAP7_75t_L g4175 ( 
.A1(n_4030),
.A2(n_3307),
.B1(n_3022),
.B2(n_3224),
.Y(n_4175)
);

A2O1A1Ixp33_ASAP7_75t_SL g4176 ( 
.A1(n_3799),
.A2(n_3095),
.B(n_3021),
.C(n_3490),
.Y(n_4176)
);

HB1xp67_ASAP7_75t_L g4177 ( 
.A(n_3631),
.Y(n_4177)
);

AND2x4_ASAP7_75t_L g4178 ( 
.A(n_3629),
.B(n_3632),
.Y(n_4178)
);

AND2x2_ASAP7_75t_L g4179 ( 
.A(n_3871),
.B(n_3252),
.Y(n_4179)
);

OA21x2_ASAP7_75t_L g4180 ( 
.A1(n_3626),
.A2(n_3361),
.B(n_3095),
.Y(n_4180)
);

NAND2x1p5_ASAP7_75t_L g4181 ( 
.A(n_3643),
.B(n_3165),
.Y(n_4181)
);

NAND2x1p5_ASAP7_75t_L g4182 ( 
.A(n_3643),
.B(n_3269),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_3666),
.Y(n_4183)
);

NAND2xp5_ASAP7_75t_L g4184 ( 
.A(n_3658),
.B(n_3066),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_L g4185 ( 
.A(n_3658),
.B(n_3066),
.Y(n_4185)
);

BUFx2_ASAP7_75t_L g4186 ( 
.A(n_4057),
.Y(n_4186)
);

OA21x2_ASAP7_75t_L g4187 ( 
.A1(n_3626),
.A2(n_3361),
.B(n_3321),
.Y(n_4187)
);

AOI22xp33_ASAP7_75t_SL g4188 ( 
.A1(n_3771),
.A2(n_3221),
.B1(n_3509),
.B2(n_3490),
.Y(n_4188)
);

INVx1_ASAP7_75t_L g4189 ( 
.A(n_3668),
.Y(n_4189)
);

AOI21x1_ASAP7_75t_L g4190 ( 
.A1(n_4013),
.A2(n_3084),
.B(n_3037),
.Y(n_4190)
);

AO31x2_ASAP7_75t_L g4191 ( 
.A1(n_4108),
.A2(n_3172),
.A3(n_3325),
.B(n_3323),
.Y(n_4191)
);

NOR2xp33_ASAP7_75t_L g4192 ( 
.A(n_3689),
.B(n_3053),
.Y(n_4192)
);

AND2x4_ASAP7_75t_L g4193 ( 
.A(n_3629),
.B(n_3295),
.Y(n_4193)
);

AOI21xp5_ASAP7_75t_L g4194 ( 
.A1(n_3672),
.A2(n_3511),
.B(n_3506),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_L g4195 ( 
.A(n_3838),
.B(n_3068),
.Y(n_4195)
);

OAI22xp5_ASAP7_75t_L g4196 ( 
.A1(n_3941),
.A2(n_3539),
.B1(n_3541),
.B2(n_3509),
.Y(n_4196)
);

OAI21x1_ASAP7_75t_L g4197 ( 
.A1(n_3917),
.A2(n_3573),
.B(n_3568),
.Y(n_4197)
);

OA21x2_ASAP7_75t_L g4198 ( 
.A1(n_3637),
.A2(n_3321),
.B(n_3323),
.Y(n_4198)
);

A2O1A1Ixp33_ASAP7_75t_L g4199 ( 
.A1(n_3791),
.A2(n_3157),
.B(n_3107),
.C(n_3054),
.Y(n_4199)
);

OAI21x1_ASAP7_75t_L g4200 ( 
.A1(n_3917),
.A2(n_3585),
.B(n_3573),
.Y(n_4200)
);

AO21x1_ASAP7_75t_L g4201 ( 
.A1(n_4062),
.A2(n_3541),
.B(n_3539),
.Y(n_4201)
);

INVx1_ASAP7_75t_L g4202 ( 
.A(n_3668),
.Y(n_4202)
);

OAI21xp5_ASAP7_75t_L g4203 ( 
.A1(n_4065),
.A2(n_3463),
.B(n_3461),
.Y(n_4203)
);

OAI21xp5_ASAP7_75t_L g4204 ( 
.A1(n_4074),
.A2(n_3474),
.B(n_3471),
.Y(n_4204)
);

OA21x2_ASAP7_75t_L g4205 ( 
.A1(n_3637),
.A2(n_3325),
.B(n_3092),
.Y(n_4205)
);

INVxp67_ASAP7_75t_L g4206 ( 
.A(n_4025),
.Y(n_4206)
);

INVx1_ASAP7_75t_SL g4207 ( 
.A(n_4015),
.Y(n_4207)
);

AND2x2_ASAP7_75t_L g4208 ( 
.A(n_3871),
.B(n_2994),
.Y(n_4208)
);

INVx1_ASAP7_75t_SL g4209 ( 
.A(n_3890),
.Y(n_4209)
);

NOR2xp33_ASAP7_75t_L g4210 ( 
.A(n_3938),
.B(n_3074),
.Y(n_4210)
);

OAI21xp33_ASAP7_75t_L g4211 ( 
.A1(n_4074),
.A2(n_3021),
.B(n_3565),
.Y(n_4211)
);

INVxp67_ASAP7_75t_L g4212 ( 
.A(n_3792),
.Y(n_4212)
);

NOR2xp33_ASAP7_75t_L g4213 ( 
.A(n_3934),
.B(n_3075),
.Y(n_4213)
);

AOI222xp33_ASAP7_75t_L g4214 ( 
.A1(n_3790),
.A2(n_3059),
.B1(n_3052),
.B2(n_3584),
.C1(n_3594),
.C2(n_3565),
.Y(n_4214)
);

NAND3xp33_ASAP7_75t_L g4215 ( 
.A(n_4080),
.B(n_3594),
.C(n_3584),
.Y(n_4215)
);

BUFx3_ASAP7_75t_L g4216 ( 
.A(n_3694),
.Y(n_4216)
);

INVx2_ASAP7_75t_L g4217 ( 
.A(n_3651),
.Y(n_4217)
);

INVx2_ASAP7_75t_L g4218 ( 
.A(n_3651),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_3671),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_3671),
.Y(n_4220)
);

HB1xp67_ASAP7_75t_L g4221 ( 
.A(n_3631),
.Y(n_4221)
);

BUFx12f_ASAP7_75t_L g4222 ( 
.A(n_3616),
.Y(n_4222)
);

INVx1_ASAP7_75t_L g4223 ( 
.A(n_3678),
.Y(n_4223)
);

INVx1_ASAP7_75t_L g4224 ( 
.A(n_3678),
.Y(n_4224)
);

OA21x2_ASAP7_75t_L g4225 ( 
.A1(n_3637),
.A2(n_3092),
.B(n_3326),
.Y(n_4225)
);

NOR2xp67_ASAP7_75t_L g4226 ( 
.A(n_4004),
.B(n_3109),
.Y(n_4226)
);

HB1xp67_ASAP7_75t_L g4227 ( 
.A(n_3996),
.Y(n_4227)
);

OR2x6_ASAP7_75t_L g4228 ( 
.A(n_3862),
.B(n_3296),
.Y(n_4228)
);

NAND2xp5_ASAP7_75t_L g4229 ( 
.A(n_3640),
.B(n_3068),
.Y(n_4229)
);

OAI21xp5_ASAP7_75t_L g4230 ( 
.A1(n_4080),
.A2(n_3535),
.B(n_3493),
.Y(n_4230)
);

INVx3_ASAP7_75t_L g4231 ( 
.A(n_3765),
.Y(n_4231)
);

INVx8_ASAP7_75t_L g4232 ( 
.A(n_3694),
.Y(n_4232)
);

AO21x2_ASAP7_75t_L g4233 ( 
.A1(n_4045),
.A2(n_4053),
.B(n_3473),
.Y(n_4233)
);

NOR2xp33_ASAP7_75t_SL g4234 ( 
.A(n_3771),
.B(n_3138),
.Y(n_4234)
);

INVx2_ASAP7_75t_L g4235 ( 
.A(n_3651),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_3684),
.Y(n_4236)
);

AO21x2_ASAP7_75t_L g4237 ( 
.A1(n_4045),
.A2(n_4053),
.B(n_3473),
.Y(n_4237)
);

BUFx2_ASAP7_75t_SL g4238 ( 
.A(n_3982),
.Y(n_4238)
);

CKINVDCx5p33_ASAP7_75t_R g4239 ( 
.A(n_3613),
.Y(n_4239)
);

OAI21x1_ASAP7_75t_L g4240 ( 
.A1(n_4118),
.A2(n_3598),
.B(n_3559),
.Y(n_4240)
);

NAND2xp5_ASAP7_75t_L g4241 ( 
.A(n_3640),
.B(n_3641),
.Y(n_4241)
);

OR2x2_ASAP7_75t_L g4242 ( 
.A(n_4089),
.B(n_4092),
.Y(n_4242)
);

NAND2xp5_ASAP7_75t_L g4243 ( 
.A(n_3641),
.B(n_3482),
.Y(n_4243)
);

CKINVDCx5p33_ASAP7_75t_R g4244 ( 
.A(n_3613),
.Y(n_4244)
);

O2A1O1Ixp33_ASAP7_75t_L g4245 ( 
.A1(n_3941),
.A2(n_3601),
.B(n_3479),
.C(n_3510),
.Y(n_4245)
);

OAI21x1_ASAP7_75t_L g4246 ( 
.A1(n_4118),
.A2(n_3012),
.B(n_3091),
.Y(n_4246)
);

AOI22xp33_ASAP7_75t_L g4247 ( 
.A1(n_4030),
.A2(n_3135),
.B1(n_3482),
.B2(n_3170),
.Y(n_4247)
);

A2O1A1Ixp33_ASAP7_75t_L g4248 ( 
.A1(n_3791),
.A2(n_3097),
.B(n_3466),
.C(n_3135),
.Y(n_4248)
);

CKINVDCx11_ASAP7_75t_R g4249 ( 
.A(n_3628),
.Y(n_4249)
);

AOI21xp33_ASAP7_75t_L g4250 ( 
.A1(n_3790),
.A2(n_3050),
.B(n_3131),
.Y(n_4250)
);

INVx1_ASAP7_75t_L g4251 ( 
.A(n_3684),
.Y(n_4251)
);

CKINVDCx5p33_ASAP7_75t_R g4252 ( 
.A(n_3682),
.Y(n_4252)
);

INVx1_ASAP7_75t_SL g4253 ( 
.A(n_3890),
.Y(n_4253)
);

OA21x2_ASAP7_75t_L g4254 ( 
.A1(n_4054),
.A2(n_4127),
.B(n_4123),
.Y(n_4254)
);

HB1xp67_ASAP7_75t_L g4255 ( 
.A(n_3996),
.Y(n_4255)
);

BUFx2_ASAP7_75t_L g4256 ( 
.A(n_4057),
.Y(n_4256)
);

AOI22xp5_ASAP7_75t_L g4257 ( 
.A1(n_3708),
.A2(n_3102),
.B1(n_3554),
.B2(n_3549),
.Y(n_4257)
);

INVx1_ASAP7_75t_SL g4258 ( 
.A(n_3901),
.Y(n_4258)
);

INVx1_ASAP7_75t_SL g4259 ( 
.A(n_3901),
.Y(n_4259)
);

INVx4_ASAP7_75t_SL g4260 ( 
.A(n_3881),
.Y(n_4260)
);

AND2x2_ASAP7_75t_L g4261 ( 
.A(n_3871),
.B(n_2994),
.Y(n_4261)
);

CKINVDCx16_ASAP7_75t_R g4262 ( 
.A(n_3949),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_3687),
.Y(n_4263)
);

AOI222xp33_ASAP7_75t_L g4264 ( 
.A1(n_3820),
.A2(n_3309),
.B1(n_3259),
.B2(n_3153),
.C1(n_3237),
.C2(n_3266),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_3687),
.Y(n_4265)
);

OR2x2_ASAP7_75t_L g4266 ( 
.A(n_4089),
.B(n_3227),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_3693),
.Y(n_4267)
);

OAI22xp33_ASAP7_75t_L g4268 ( 
.A1(n_3708),
.A2(n_3102),
.B1(n_3564),
.B2(n_3558),
.Y(n_4268)
);

AO21x2_ASAP7_75t_L g4269 ( 
.A1(n_3837),
.A2(n_3487),
.B(n_3440),
.Y(n_4269)
);

OAI21x1_ASAP7_75t_L g4270 ( 
.A1(n_4060),
.A2(n_3039),
.B(n_3134),
.Y(n_4270)
);

AO31x2_ASAP7_75t_L g4271 ( 
.A1(n_4129),
.A2(n_3237),
.A3(n_3266),
.B(n_3232),
.Y(n_4271)
);

BUFx3_ASAP7_75t_L g4272 ( 
.A(n_3694),
.Y(n_4272)
);

OAI21xp5_ASAP7_75t_L g4273 ( 
.A1(n_4121),
.A2(n_3588),
.B(n_3571),
.Y(n_4273)
);

INVx1_ASAP7_75t_L g4274 ( 
.A(n_3693),
.Y(n_4274)
);

INVx3_ASAP7_75t_L g4275 ( 
.A(n_3765),
.Y(n_4275)
);

INVx1_ASAP7_75t_SL g4276 ( 
.A(n_3925),
.Y(n_4276)
);

INVx4_ASAP7_75t_L g4277 ( 
.A(n_3712),
.Y(n_4277)
);

INVx1_ASAP7_75t_L g4278 ( 
.A(n_3695),
.Y(n_4278)
);

HB1xp67_ASAP7_75t_L g4279 ( 
.A(n_3612),
.Y(n_4279)
);

INVx1_ASAP7_75t_L g4280 ( 
.A(n_3695),
.Y(n_4280)
);

OAI21x1_ASAP7_75t_SL g4281 ( 
.A1(n_3733),
.A2(n_3201),
.B(n_3608),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_3706),
.Y(n_4282)
);

INVx1_ASAP7_75t_L g4283 ( 
.A(n_3706),
.Y(n_4283)
);

OAI22xp5_ASAP7_75t_L g4284 ( 
.A1(n_3625),
.A2(n_3597),
.B1(n_3522),
.B2(n_3511),
.Y(n_4284)
);

INVx1_ASAP7_75t_SL g4285 ( 
.A(n_3925),
.Y(n_4285)
);

OAI22xp5_ASAP7_75t_L g4286 ( 
.A1(n_3625),
.A2(n_3605),
.B1(n_3608),
.B2(n_3522),
.Y(n_4286)
);

BUFx6f_ASAP7_75t_L g4287 ( 
.A(n_3611),
.Y(n_4287)
);

INVx6_ASAP7_75t_L g4288 ( 
.A(n_3627),
.Y(n_4288)
);

NOR2xp33_ASAP7_75t_SL g4289 ( 
.A(n_3774),
.B(n_3056),
.Y(n_4289)
);

CKINVDCx6p67_ASAP7_75t_R g4290 ( 
.A(n_3712),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_3710),
.Y(n_4291)
);

AOI22xp33_ASAP7_75t_L g4292 ( 
.A1(n_4030),
.A2(n_3482),
.B1(n_3221),
.B2(n_3309),
.Y(n_4292)
);

AOI21xp5_ASAP7_75t_L g4293 ( 
.A1(n_3621),
.A2(n_3605),
.B(n_3477),
.Y(n_4293)
);

NAND2xp5_ASAP7_75t_L g4294 ( 
.A(n_3851),
.B(n_3142),
.Y(n_4294)
);

INVxp67_ASAP7_75t_L g4295 ( 
.A(n_3792),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_3710),
.Y(n_4296)
);

O2A1O1Ixp5_ASAP7_75t_L g4297 ( 
.A1(n_3975),
.A2(n_3434),
.B(n_3201),
.C(n_3230),
.Y(n_4297)
);

NAND3xp33_ASAP7_75t_SL g4298 ( 
.A(n_4059),
.B(n_3437),
.C(n_3245),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_3722),
.Y(n_4299)
);

OAI22xp5_ASAP7_75t_L g4300 ( 
.A1(n_3625),
.A2(n_3469),
.B1(n_3602),
.B2(n_3477),
.Y(n_4300)
);

AO21x2_ASAP7_75t_L g4301 ( 
.A1(n_3837),
.A2(n_3487),
.B(n_3440),
.Y(n_4301)
);

CKINVDCx20_ASAP7_75t_R g4302 ( 
.A(n_3639),
.Y(n_4302)
);

OAI22xp33_ASAP7_75t_L g4303 ( 
.A1(n_3660),
.A2(n_3154),
.B1(n_3232),
.B2(n_3153),
.Y(n_4303)
);

AO31x2_ASAP7_75t_L g4304 ( 
.A1(n_3674),
.A2(n_3700),
.A3(n_3705),
.B(n_3683),
.Y(n_4304)
);

AOI22x1_ASAP7_75t_L g4305 ( 
.A1(n_3774),
.A2(n_3070),
.B1(n_3087),
.B2(n_3129),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_3722),
.Y(n_4306)
);

AOI221xp5_ASAP7_75t_L g4307 ( 
.A1(n_4030),
.A2(n_3602),
.B1(n_3469),
.B2(n_3132),
.C(n_3203),
.Y(n_4307)
);

NOR2xp33_ASAP7_75t_L g4308 ( 
.A(n_3900),
.B(n_3075),
.Y(n_4308)
);

O2A1O1Ixp33_ASAP7_75t_SL g4309 ( 
.A1(n_4002),
.A2(n_3428),
.B(n_3355),
.C(n_3251),
.Y(n_4309)
);

NOR2xp33_ASAP7_75t_L g4310 ( 
.A(n_3950),
.B(n_3190),
.Y(n_4310)
);

INVx1_ASAP7_75t_L g4311 ( 
.A(n_3725),
.Y(n_4311)
);

AOI21xp5_ASAP7_75t_SL g4312 ( 
.A1(n_3991),
.A2(n_3175),
.B(n_3420),
.Y(n_4312)
);

INVx1_ASAP7_75t_SL g4313 ( 
.A(n_3939),
.Y(n_4313)
);

OR2x6_ASAP7_75t_L g4314 ( 
.A(n_3862),
.B(n_3299),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_3725),
.Y(n_4315)
);

NAND2xp5_ASAP7_75t_L g4316 ( 
.A(n_3851),
.B(n_3142),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_3730),
.Y(n_4317)
);

BUFx4_ASAP7_75t_SL g4318 ( 
.A(n_3804),
.Y(n_4318)
);

AOI21x1_ASAP7_75t_L g4319 ( 
.A1(n_3657),
.A2(n_3538),
.B(n_3492),
.Y(n_4319)
);

OA21x2_ASAP7_75t_L g4320 ( 
.A1(n_3648),
.A2(n_3248),
.B(n_3150),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_3730),
.Y(n_4321)
);

INVx3_ASAP7_75t_L g4322 ( 
.A(n_3765),
.Y(n_4322)
);

INVx3_ASAP7_75t_L g4323 ( 
.A(n_3858),
.Y(n_4323)
);

OAI21xp5_ASAP7_75t_L g4324 ( 
.A1(n_4121),
.A2(n_3175),
.B(n_3055),
.Y(n_4324)
);

A2O1A1Ixp33_ASAP7_75t_L g4325 ( 
.A1(n_3729),
.A2(n_3184),
.B(n_3315),
.C(n_3259),
.Y(n_4325)
);

AOI22xp33_ASAP7_75t_L g4326 ( 
.A1(n_3820),
.A2(n_3116),
.B1(n_3249),
.B2(n_3204),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_3731),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_3731),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_3734),
.Y(n_4329)
);

OAI21xp5_ASAP7_75t_L g4330 ( 
.A1(n_3729),
.A2(n_3055),
.B(n_3159),
.Y(n_4330)
);

INVx3_ASAP7_75t_L g4331 ( 
.A(n_3858),
.Y(n_4331)
);

OAI211xp5_ASAP7_75t_L g4332 ( 
.A1(n_3796),
.A2(n_3132),
.B(n_3343),
.C(n_3315),
.Y(n_4332)
);

INVx1_ASAP7_75t_L g4333 ( 
.A(n_3734),
.Y(n_4333)
);

OAI21x1_ASAP7_75t_SL g4334 ( 
.A1(n_3733),
.A2(n_3436),
.B(n_3070),
.Y(n_4334)
);

CKINVDCx5p33_ASAP7_75t_R g4335 ( 
.A(n_3616),
.Y(n_4335)
);

BUFx2_ASAP7_75t_L g4336 ( 
.A(n_4057),
.Y(n_4336)
);

NAND2xp5_ASAP7_75t_L g4337 ( 
.A(n_3656),
.B(n_3271),
.Y(n_4337)
);

INVx1_ASAP7_75t_SL g4338 ( 
.A(n_3939),
.Y(n_4338)
);

OAI221xp5_ASAP7_75t_L g4339 ( 
.A1(n_3859),
.A2(n_3245),
.B1(n_3343),
.B2(n_3116),
.C(n_3205),
.Y(n_4339)
);

OAI21xp5_ASAP7_75t_L g4340 ( 
.A1(n_3796),
.A2(n_3123),
.B(n_3129),
.Y(n_4340)
);

OAI21xp5_ASAP7_75t_L g4341 ( 
.A1(n_4024),
.A2(n_4098),
.B(n_3975),
.Y(n_4341)
);

BUFx3_ASAP7_75t_L g4342 ( 
.A(n_3712),
.Y(n_4342)
);

OR2x2_ASAP7_75t_L g4343 ( 
.A(n_4092),
.B(n_3227),
.Y(n_4343)
);

OA21x2_ASAP7_75t_L g4344 ( 
.A1(n_3656),
.A2(n_3248),
.B(n_3130),
.Y(n_4344)
);

INVx1_ASAP7_75t_L g4345 ( 
.A(n_3740),
.Y(n_4345)
);

AO32x2_ASAP7_75t_L g4346 ( 
.A1(n_4047),
.A2(n_3173),
.A3(n_3190),
.B1(n_3220),
.B2(n_3367),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_3740),
.Y(n_4347)
);

INVx1_ASAP7_75t_L g4348 ( 
.A(n_3743),
.Y(n_4348)
);

OAI21xp5_ASAP7_75t_L g4349 ( 
.A1(n_4024),
.A2(n_3123),
.B(n_3119),
.Y(n_4349)
);

OAI21xp33_ASAP7_75t_SL g4350 ( 
.A1(n_3822),
.A2(n_3279),
.B(n_3113),
.Y(n_4350)
);

AO31x2_ASAP7_75t_L g4351 ( 
.A1(n_3751),
.A2(n_3813),
.A3(n_3829),
.B(n_3805),
.Y(n_4351)
);

AOI22xp33_ASAP7_75t_L g4352 ( 
.A1(n_3859),
.A2(n_3310),
.B1(n_3562),
.B2(n_3406),
.Y(n_4352)
);

INVx1_ASAP7_75t_L g4353 ( 
.A(n_3743),
.Y(n_4353)
);

CKINVDCx20_ASAP7_75t_R g4354 ( 
.A(n_3727),
.Y(n_4354)
);

INVx1_ASAP7_75t_L g4355 ( 
.A(n_3744),
.Y(n_4355)
);

AOI22xp33_ASAP7_75t_L g4356 ( 
.A1(n_3861),
.A2(n_3310),
.B1(n_3562),
.B2(n_3406),
.Y(n_4356)
);

INVx1_ASAP7_75t_L g4357 ( 
.A(n_3744),
.Y(n_4357)
);

INVxp67_ASAP7_75t_L g4358 ( 
.A(n_3823),
.Y(n_4358)
);

INVx1_ASAP7_75t_L g4359 ( 
.A(n_3746),
.Y(n_4359)
);

NOR2xp33_ASAP7_75t_L g4360 ( 
.A(n_3811),
.B(n_3261),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_3746),
.Y(n_4361)
);

NAND2xp5_ASAP7_75t_L g4362 ( 
.A(n_3704),
.B(n_3271),
.Y(n_4362)
);

OR2x2_ASAP7_75t_L g4363 ( 
.A(n_3918),
.B(n_3227),
.Y(n_4363)
);

AOI22xp33_ASAP7_75t_L g4364 ( 
.A1(n_3861),
.A2(n_3562),
.B1(n_3220),
.B2(n_3353),
.Y(n_4364)
);

AND2x2_ASAP7_75t_L g4365 ( 
.A(n_3878),
.B(n_3043),
.Y(n_4365)
);

CKINVDCx5p33_ASAP7_75t_R g4366 ( 
.A(n_3616),
.Y(n_4366)
);

CKINVDCx12_ASAP7_75t_R g4367 ( 
.A(n_3991),
.Y(n_4367)
);

BUFx2_ASAP7_75t_L g4368 ( 
.A(n_4057),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_3749),
.Y(n_4369)
);

NAND2xp5_ASAP7_75t_L g4370 ( 
.A(n_3704),
.B(n_3272),
.Y(n_4370)
);

OR2x6_ASAP7_75t_L g4371 ( 
.A(n_3862),
.B(n_3113),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_3749),
.Y(n_4372)
);

OAI22x1_ASAP7_75t_L g4373 ( 
.A1(n_3881),
.A2(n_3943),
.B1(n_4055),
.B2(n_4034),
.Y(n_4373)
);

OAI21xp5_ASAP7_75t_L g4374 ( 
.A1(n_4098),
.A2(n_3119),
.B(n_3046),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_3752),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_3752),
.Y(n_4376)
);

OAI21xp5_ASAP7_75t_L g4377 ( 
.A1(n_3971),
.A2(n_3046),
.B(n_3279),
.Y(n_4377)
);

CKINVDCx5p33_ASAP7_75t_R g4378 ( 
.A(n_3768),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_3753),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_3753),
.Y(n_4380)
);

AND2x2_ASAP7_75t_L g4381 ( 
.A(n_3878),
.B(n_3043),
.Y(n_4381)
);

AOI22xp33_ASAP7_75t_L g4382 ( 
.A1(n_3993),
.A2(n_3562),
.B1(n_3353),
.B2(n_3436),
.Y(n_4382)
);

CKINVDCx5p33_ASAP7_75t_R g4383 ( 
.A(n_3779),
.Y(n_4383)
);

AOI22xp33_ASAP7_75t_L g4384 ( 
.A1(n_3880),
.A2(n_3369),
.B1(n_3313),
.B2(n_3352),
.Y(n_4384)
);

CKINVDCx11_ASAP7_75t_R g4385 ( 
.A(n_3659),
.Y(n_4385)
);

AO32x2_ASAP7_75t_L g4386 ( 
.A1(n_4047),
.A2(n_4073),
.A3(n_4075),
.B1(n_4050),
.B2(n_4049),
.Y(n_4386)
);

AND2x2_ASAP7_75t_L g4387 ( 
.A(n_3878),
.B(n_3578),
.Y(n_4387)
);

AOI22xp33_ASAP7_75t_L g4388 ( 
.A1(n_3880),
.A2(n_3369),
.B1(n_3313),
.B2(n_3352),
.Y(n_4388)
);

OA21x2_ASAP7_75t_L g4389 ( 
.A1(n_3772),
.A2(n_3550),
.B(n_3542),
.Y(n_4389)
);

INVxp67_ASAP7_75t_SL g4390 ( 
.A(n_4004),
.Y(n_4390)
);

AOI21x1_ASAP7_75t_L g4391 ( 
.A1(n_3657),
.A2(n_3550),
.B(n_3542),
.Y(n_4391)
);

BUFx3_ASAP7_75t_L g4392 ( 
.A(n_3724),
.Y(n_4392)
);

AOI22xp33_ASAP7_75t_SL g4393 ( 
.A1(n_3867),
.A2(n_2992),
.B1(n_2998),
.B2(n_3495),
.Y(n_4393)
);

BUFx2_ASAP7_75t_L g4394 ( 
.A(n_4057),
.Y(n_4394)
);

INVx5_ASAP7_75t_L g4395 ( 
.A(n_3921),
.Y(n_4395)
);

A2O1A1Ixp33_ASAP7_75t_L g4396 ( 
.A1(n_4031),
.A2(n_3280),
.B(n_3289),
.C(n_3215),
.Y(n_4396)
);

OAI21xp5_ASAP7_75t_L g4397 ( 
.A1(n_3971),
.A2(n_3082),
.B(n_3230),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_3764),
.Y(n_4398)
);

OR2x6_ASAP7_75t_L g4399 ( 
.A(n_3862),
.B(n_3363),
.Y(n_4399)
);

OAI21x1_ASAP7_75t_L g4400 ( 
.A1(n_3984),
.A2(n_3276),
.B(n_3195),
.Y(n_4400)
);

OR2x6_ASAP7_75t_L g4401 ( 
.A(n_3879),
.B(n_3363),
.Y(n_4401)
);

BUFx6f_ASAP7_75t_L g4402 ( 
.A(n_3611),
.Y(n_4402)
);

OAI22xp33_ASAP7_75t_L g4403 ( 
.A1(n_3660),
.A2(n_3289),
.B1(n_3260),
.B2(n_3258),
.Y(n_4403)
);

OA21x2_ASAP7_75t_L g4404 ( 
.A1(n_3772),
.A2(n_3840),
.B(n_3984),
.Y(n_4404)
);

O2A1O1Ixp33_ASAP7_75t_SL g4405 ( 
.A1(n_4002),
.A2(n_3038),
.B(n_3106),
.C(n_3103),
.Y(n_4405)
);

OAI21x1_ASAP7_75t_SL g4406 ( 
.A1(n_3733),
.A2(n_3038),
.B(n_3241),
.Y(n_4406)
);

NAND2xp5_ASAP7_75t_L g4407 ( 
.A(n_3840),
.B(n_3272),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_3764),
.Y(n_4408)
);

OAI21x1_ASAP7_75t_L g4409 ( 
.A1(n_3852),
.A2(n_3276),
.B(n_3195),
.Y(n_4409)
);

AOI221xp5_ASAP7_75t_L g4410 ( 
.A1(n_3894),
.A2(n_3242),
.B1(n_3106),
.B2(n_3103),
.C(n_3286),
.Y(n_4410)
);

CKINVDCx6p67_ASAP7_75t_R g4411 ( 
.A(n_3724),
.Y(n_4411)
);

BUFx2_ASAP7_75t_R g4412 ( 
.A(n_3660),
.Y(n_4412)
);

AOI21xp5_ASAP7_75t_L g4413 ( 
.A1(n_3643),
.A2(n_3082),
.B(n_3398),
.Y(n_4413)
);

A2O1A1Ixp33_ASAP7_75t_L g4414 ( 
.A1(n_4031),
.A2(n_3243),
.B(n_3286),
.C(n_3278),
.Y(n_4414)
);

BUFx3_ASAP7_75t_L g4415 ( 
.A(n_3724),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_3770),
.Y(n_4416)
);

A2O1A1Ixp33_ASAP7_75t_L g4417 ( 
.A1(n_4034),
.A2(n_3370),
.B(n_3254),
.C(n_3523),
.Y(n_4417)
);

AND2x2_ASAP7_75t_L g4418 ( 
.A(n_3902),
.B(n_3360),
.Y(n_4418)
);

OAI21xp5_ASAP7_75t_L g4419 ( 
.A1(n_4028),
.A2(n_3082),
.B(n_3242),
.Y(n_4419)
);

NAND2xp5_ASAP7_75t_SL g4420 ( 
.A(n_3819),
.B(n_3189),
.Y(n_4420)
);

BUFx2_ASAP7_75t_L g4421 ( 
.A(n_3949),
.Y(n_4421)
);

AND2x4_ASAP7_75t_L g4422 ( 
.A(n_3665),
.B(n_3797),
.Y(n_4422)
);

OAI21xp5_ASAP7_75t_L g4423 ( 
.A1(n_4028),
.A2(n_3264),
.B(n_3287),
.Y(n_4423)
);

OAI21xp5_ASAP7_75t_L g4424 ( 
.A1(n_4040),
.A2(n_3287),
.B(n_3253),
.Y(n_4424)
);

OAI221xp5_ASAP7_75t_L g4425 ( 
.A1(n_3880),
.A2(n_3026),
.B1(n_3540),
.B2(n_3031),
.C(n_3523),
.Y(n_4425)
);

AOI21xp5_ASAP7_75t_L g4426 ( 
.A1(n_3679),
.A2(n_3936),
.B(n_3894),
.Y(n_4426)
);

OAI21xp5_ASAP7_75t_L g4427 ( 
.A1(n_4040),
.A2(n_3320),
.B(n_3262),
.Y(n_4427)
);

OR2x2_ASAP7_75t_L g4428 ( 
.A(n_3918),
.B(n_3227),
.Y(n_4428)
);

BUFx3_ASAP7_75t_L g4429 ( 
.A(n_3736),
.Y(n_4429)
);

CKINVDCx5p33_ASAP7_75t_R g4430 ( 
.A(n_3659),
.Y(n_4430)
);

NOR2xp67_ASAP7_75t_L g4431 ( 
.A(n_3808),
.B(n_3030),
.Y(n_4431)
);

NAND2xp5_ASAP7_75t_L g4432 ( 
.A(n_3936),
.B(n_3273),
.Y(n_4432)
);

AND2x2_ASAP7_75t_L g4433 ( 
.A(n_3902),
.B(n_3360),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_L g4434 ( 
.A(n_3940),
.B(n_3273),
.Y(n_4434)
);

OAI22xp5_ASAP7_75t_L g4435 ( 
.A1(n_4083),
.A2(n_3368),
.B1(n_3348),
.B2(n_3281),
.Y(n_4435)
);

NAND3xp33_ASAP7_75t_L g4436 ( 
.A(n_3868),
.B(n_3288),
.C(n_3101),
.Y(n_4436)
);

BUFx2_ASAP7_75t_L g4437 ( 
.A(n_4022),
.Y(n_4437)
);

O2A1O1Ixp33_ASAP7_75t_SL g4438 ( 
.A1(n_3933),
.A2(n_3189),
.B(n_3281),
.C(n_3599),
.Y(n_4438)
);

INVxp67_ASAP7_75t_SL g4439 ( 
.A(n_3612),
.Y(n_4439)
);

OAI21xp5_ASAP7_75t_L g4440 ( 
.A1(n_3914),
.A2(n_3959),
.B(n_3940),
.Y(n_4440)
);

AND2x2_ASAP7_75t_L g4441 ( 
.A(n_3902),
.B(n_3373),
.Y(n_4441)
);

INVx2_ASAP7_75t_SL g4442 ( 
.A(n_4022),
.Y(n_4442)
);

BUFx3_ASAP7_75t_L g4443 ( 
.A(n_3736),
.Y(n_4443)
);

NOR2x1_ASAP7_75t_SL g4444 ( 
.A(n_3930),
.B(n_3090),
.Y(n_4444)
);

OAI21xp5_ASAP7_75t_L g4445 ( 
.A1(n_3914),
.A2(n_3246),
.B(n_3288),
.Y(n_4445)
);

AOI21xp5_ASAP7_75t_L g4446 ( 
.A1(n_3679),
.A2(n_3282),
.B(n_3391),
.Y(n_4446)
);

INVx1_ASAP7_75t_L g4447 ( 
.A(n_3770),
.Y(n_4447)
);

OAI21xp5_ASAP7_75t_L g4448 ( 
.A1(n_3959),
.A2(n_3246),
.B(n_3303),
.Y(n_4448)
);

INVx1_ASAP7_75t_L g4449 ( 
.A(n_3780),
.Y(n_4449)
);

INVx1_ASAP7_75t_L g4450 ( 
.A(n_3780),
.Y(n_4450)
);

OA21x2_ASAP7_75t_L g4451 ( 
.A1(n_4035),
.A2(n_4037),
.B(n_3947),
.Y(n_4451)
);

AOI222xp33_ASAP7_75t_L g4452 ( 
.A1(n_3875),
.A2(n_3026),
.B1(n_3031),
.B2(n_3540),
.C1(n_3523),
.C2(n_3590),
.Y(n_4452)
);

AND2x2_ASAP7_75t_L g4453 ( 
.A(n_3832),
.B(n_3848),
.Y(n_4453)
);

INVx1_ASAP7_75t_L g4454 ( 
.A(n_3783),
.Y(n_4454)
);

NAND2xp5_ASAP7_75t_L g4455 ( 
.A(n_3618),
.B(n_3080),
.Y(n_4455)
);

OAI21xp5_ASAP7_75t_L g4456 ( 
.A1(n_3847),
.A2(n_3868),
.B(n_3630),
.Y(n_4456)
);

AND2x2_ASAP7_75t_L g4457 ( 
.A(n_3832),
.B(n_3375),
.Y(n_4457)
);

NAND2x1p5_ASAP7_75t_L g4458 ( 
.A(n_3679),
.B(n_3427),
.Y(n_4458)
);

OAI21x1_ASAP7_75t_L g4459 ( 
.A1(n_3638),
.A2(n_3228),
.B(n_3226),
.Y(n_4459)
);

INVx5_ASAP7_75t_L g4460 ( 
.A(n_3921),
.Y(n_4460)
);

AOI21xp5_ASAP7_75t_L g4461 ( 
.A1(n_3679),
.A2(n_3839),
.B(n_3732),
.Y(n_4461)
);

OAI21x1_ASAP7_75t_L g4462 ( 
.A1(n_3702),
.A2(n_3228),
.B(n_3226),
.Y(n_4462)
);

AND2x2_ASAP7_75t_L g4463 ( 
.A(n_3832),
.B(n_3375),
.Y(n_4463)
);

O2A1O1Ixp33_ASAP7_75t_L g4464 ( 
.A1(n_3847),
.A2(n_3101),
.B(n_3098),
.C(n_3081),
.Y(n_4464)
);

OAI22xp33_ASAP7_75t_L g4465 ( 
.A1(n_3943),
.A2(n_4055),
.B1(n_3688),
.B2(n_3699),
.Y(n_4465)
);

OA21x2_ASAP7_75t_L g4466 ( 
.A1(n_3947),
.A2(n_3499),
.B(n_3581),
.Y(n_4466)
);

HB1xp67_ASAP7_75t_L g4467 ( 
.A(n_3618),
.Y(n_4467)
);

NOR2xp33_ASAP7_75t_L g4468 ( 
.A(n_3863),
.B(n_3285),
.Y(n_4468)
);

OAI21xp5_ASAP7_75t_L g4469 ( 
.A1(n_3847),
.A2(n_3303),
.B(n_3031),
.Y(n_4469)
);

AOI22xp33_ASAP7_75t_L g4470 ( 
.A1(n_3822),
.A2(n_3379),
.B1(n_3400),
.B2(n_3389),
.Y(n_4470)
);

OAI22xp5_ASAP7_75t_L g4471 ( 
.A1(n_4083),
.A2(n_3383),
.B1(n_3081),
.B2(n_3098),
.Y(n_4471)
);

INVxp67_ASAP7_75t_SL g4472 ( 
.A(n_3630),
.Y(n_4472)
);

BUFx6f_ASAP7_75t_L g4473 ( 
.A(n_3611),
.Y(n_4473)
);

OAI21x1_ASAP7_75t_L g4474 ( 
.A1(n_3702),
.A2(n_3233),
.B(n_3229),
.Y(n_4474)
);

HB1xp67_ASAP7_75t_L g4475 ( 
.A(n_3742),
.Y(n_4475)
);

OAI21x1_ASAP7_75t_L g4476 ( 
.A1(n_3702),
.A2(n_3233),
.B(n_3229),
.Y(n_4476)
);

AOI22xp33_ASAP7_75t_L g4477 ( 
.A1(n_3822),
.A2(n_3390),
.B1(n_3080),
.B2(n_3380),
.Y(n_4477)
);

NAND2xp5_ASAP7_75t_L g4478 ( 
.A(n_4026),
.B(n_3301),
.Y(n_4478)
);

OAI21xp5_ASAP7_75t_L g4479 ( 
.A1(n_3868),
.A2(n_3026),
.B(n_3031),
.Y(n_4479)
);

AND2x4_ASAP7_75t_L g4480 ( 
.A(n_3665),
.B(n_3227),
.Y(n_4480)
);

A2O1A1Ixp33_ASAP7_75t_L g4481 ( 
.A1(n_3974),
.A2(n_3026),
.B(n_3031),
.C(n_3540),
.Y(n_4481)
);

CKINVDCx5p33_ASAP7_75t_R g4482 ( 
.A(n_3659),
.Y(n_4482)
);

AND2x2_ASAP7_75t_L g4483 ( 
.A(n_3848),
.B(n_3227),
.Y(n_4483)
);

INVx6_ASAP7_75t_L g4484 ( 
.A(n_3627),
.Y(n_4484)
);

AND2x2_ASAP7_75t_L g4485 ( 
.A(n_3848),
.B(n_3072),
.Y(n_4485)
);

AND2x2_ASAP7_75t_L g4486 ( 
.A(n_3775),
.B(n_3072),
.Y(n_4486)
);

INVx2_ASAP7_75t_SL g4487 ( 
.A(n_4068),
.Y(n_4487)
);

CKINVDCx5p33_ASAP7_75t_R g4488 ( 
.A(n_3691),
.Y(n_4488)
);

AOI21xp5_ASAP7_75t_L g4489 ( 
.A1(n_3732),
.A2(n_3425),
.B(n_3199),
.Y(n_4489)
);

CKINVDCx6p67_ASAP7_75t_R g4490 ( 
.A(n_3736),
.Y(n_4490)
);

OAI21x1_ASAP7_75t_L g4491 ( 
.A1(n_3723),
.A2(n_3741),
.B(n_3737),
.Y(n_4491)
);

INVx1_ASAP7_75t_L g4492 ( 
.A(n_3783),
.Y(n_4492)
);

INVx1_ASAP7_75t_L g4493 ( 
.A(n_3787),
.Y(n_4493)
);

A2O1A1Ixp33_ASAP7_75t_L g4494 ( 
.A1(n_4095),
.A2(n_3026),
.B(n_3031),
.C(n_3540),
.Y(n_4494)
);

AOI22xp33_ASAP7_75t_L g4495 ( 
.A1(n_4095),
.A2(n_3354),
.B1(n_3333),
.B2(n_3330),
.Y(n_4495)
);

INVx1_ASAP7_75t_L g4496 ( 
.A(n_3787),
.Y(n_4496)
);

CKINVDCx5p33_ASAP7_75t_R g4497 ( 
.A(n_3691),
.Y(n_4497)
);

INVx1_ASAP7_75t_L g4498 ( 
.A(n_3802),
.Y(n_4498)
);

NAND2xp5_ASAP7_75t_L g4499 ( 
.A(n_4041),
.B(n_3301),
.Y(n_4499)
);

BUFx2_ASAP7_75t_L g4500 ( 
.A(n_3761),
.Y(n_4500)
);

NAND2xp5_ASAP7_75t_L g4501 ( 
.A(n_3681),
.B(n_3298),
.Y(n_4501)
);

AOI22xp33_ASAP7_75t_L g4502 ( 
.A1(n_4087),
.A2(n_3292),
.B1(n_3333),
.B2(n_3330),
.Y(n_4502)
);

NAND2x1p5_ASAP7_75t_L g4503 ( 
.A(n_3732),
.B(n_3234),
.Y(n_4503)
);

BUFx2_ASAP7_75t_L g4504 ( 
.A(n_3761),
.Y(n_4504)
);

OAI221xp5_ASAP7_75t_L g4505 ( 
.A1(n_4101),
.A2(n_3026),
.B1(n_3540),
.B2(n_3523),
.C(n_3590),
.Y(n_4505)
);

BUFx10_ASAP7_75t_L g4506 ( 
.A(n_3675),
.Y(n_4506)
);

NOR2xp67_ASAP7_75t_L g4507 ( 
.A(n_3808),
.B(n_3815),
.Y(n_4507)
);

NAND2xp5_ASAP7_75t_L g4508 ( 
.A(n_3681),
.B(n_3298),
.Y(n_4508)
);

BUFx12f_ASAP7_75t_L g4509 ( 
.A(n_3622),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_3802),
.Y(n_4510)
);

AND2x4_ASAP7_75t_L g4511 ( 
.A(n_3665),
.B(n_3590),
.Y(n_4511)
);

AO21x2_ASAP7_75t_L g4512 ( 
.A1(n_4105),
.A2(n_3530),
.B(n_3064),
.Y(n_4512)
);

HB1xp67_ASAP7_75t_L g4513 ( 
.A(n_3742),
.Y(n_4513)
);

BUFx2_ASAP7_75t_L g4514 ( 
.A(n_3761),
.Y(n_4514)
);

NAND2xp5_ASAP7_75t_L g4515 ( 
.A(n_3711),
.B(n_3293),
.Y(n_4515)
);

HB1xp67_ASAP7_75t_L g4516 ( 
.A(n_3777),
.Y(n_4516)
);

XOR2xp5_ASAP7_75t_L g4517 ( 
.A(n_3869),
.B(n_3293),
.Y(n_4517)
);

INVx1_ASAP7_75t_L g4518 ( 
.A(n_3809),
.Y(n_4518)
);

AND2x2_ASAP7_75t_L g4519 ( 
.A(n_3775),
.B(n_3061),
.Y(n_4519)
);

AOI22xp5_ASAP7_75t_L g4520 ( 
.A1(n_4099),
.A2(n_3211),
.B1(n_3285),
.B2(n_3523),
.Y(n_4520)
);

NAND3xp33_ASAP7_75t_L g4521 ( 
.A(n_3677),
.B(n_3267),
.C(n_3421),
.Y(n_4521)
);

BUFx2_ASAP7_75t_L g4522 ( 
.A(n_3767),
.Y(n_4522)
);

HB1xp67_ASAP7_75t_L g4523 ( 
.A(n_3777),
.Y(n_4523)
);

BUFx3_ASAP7_75t_L g4524 ( 
.A(n_3627),
.Y(n_4524)
);

BUFx4_ASAP7_75t_SL g4525 ( 
.A(n_3716),
.Y(n_4525)
);

AOI21xp5_ASAP7_75t_L g4526 ( 
.A1(n_3839),
.A2(n_3424),
.B(n_3235),
.Y(n_4526)
);

NAND2xp5_ASAP7_75t_L g4527 ( 
.A(n_3711),
.B(n_3590),
.Y(n_4527)
);

OAI22xp33_ASAP7_75t_L g4528 ( 
.A1(n_3943),
.A2(n_4055),
.B1(n_3688),
.B2(n_3699),
.Y(n_4528)
);

AND2x4_ASAP7_75t_L g4529 ( 
.A(n_3797),
.B(n_3590),
.Y(n_4529)
);

OAI21x1_ASAP7_75t_SL g4530 ( 
.A1(n_3808),
.A2(n_3238),
.B(n_3424),
.Y(n_4530)
);

AOI21xp33_ASAP7_75t_SL g4531 ( 
.A1(n_3654),
.A2(n_3590),
.B(n_3540),
.Y(n_4531)
);

CKINVDCx5p33_ASAP7_75t_R g4532 ( 
.A(n_3691),
.Y(n_4532)
);

CKINVDCx16_ASAP7_75t_R g4533 ( 
.A(n_3808),
.Y(n_4533)
);

OAI21x1_ASAP7_75t_L g4534 ( 
.A1(n_3778),
.A2(n_3333),
.B(n_3354),
.Y(n_4534)
);

AND2x2_ASAP7_75t_L g4535 ( 
.A(n_3775),
.B(n_3061),
.Y(n_4535)
);

NOR2xp33_ASAP7_75t_L g4536 ( 
.A(n_3782),
.B(n_3211),
.Y(n_4536)
);

INVx2_ASAP7_75t_SL g4537 ( 
.A(n_4068),
.Y(n_4537)
);

CKINVDCx5p33_ASAP7_75t_R g4538 ( 
.A(n_3745),
.Y(n_4538)
);

OAI21xp5_ASAP7_75t_L g4539 ( 
.A1(n_3617),
.A2(n_3523),
.B(n_3072),
.Y(n_4539)
);

OAI22xp33_ASAP7_75t_L g4540 ( 
.A1(n_4115),
.A2(n_3061),
.B1(n_3072),
.B2(n_3330),
.Y(n_4540)
);

OAI21x1_ASAP7_75t_L g4541 ( 
.A1(n_3778),
.A2(n_3788),
.B(n_3785),
.Y(n_4541)
);

OAI221xp5_ASAP7_75t_L g4542 ( 
.A1(n_4101),
.A2(n_3061),
.B1(n_3072),
.B2(n_3314),
.C(n_3382),
.Y(n_4542)
);

BUFx6f_ASAP7_75t_L g4543 ( 
.A(n_3611),
.Y(n_4543)
);

NAND2xp5_ASAP7_75t_L g4544 ( 
.A(n_3713),
.B(n_3061),
.Y(n_4544)
);

AOI21x1_ASAP7_75t_L g4545 ( 
.A1(n_3677),
.A2(n_3314),
.B(n_3365),
.Y(n_4545)
);

AND2x4_ASAP7_75t_L g4546 ( 
.A(n_3797),
.B(n_3061),
.Y(n_4546)
);

INVx1_ASAP7_75t_L g4547 ( 
.A(n_3809),
.Y(n_4547)
);

HB1xp67_ASAP7_75t_L g4548 ( 
.A(n_3823),
.Y(n_4548)
);

NAND2xp5_ASAP7_75t_L g4549 ( 
.A(n_3713),
.B(n_3072),
.Y(n_4549)
);

NOR2xp33_ASAP7_75t_L g4550 ( 
.A(n_3782),
.B(n_3365),
.Y(n_4550)
);

A2O1A1Ixp33_ASAP7_75t_L g4551 ( 
.A1(n_4008),
.A2(n_3365),
.B(n_3382),
.C(n_3401),
.Y(n_4551)
);

INVx4_ASAP7_75t_SL g4552 ( 
.A(n_3828),
.Y(n_4552)
);

OAI21x1_ASAP7_75t_L g4553 ( 
.A1(n_3778),
.A2(n_3304),
.B(n_3401),
.Y(n_4553)
);

AND2x2_ASAP7_75t_L g4554 ( 
.A(n_3801),
.B(n_3422),
.Y(n_4554)
);

NAND2x1_ASAP7_75t_L g4555 ( 
.A(n_3619),
.B(n_3304),
.Y(n_4555)
);

AO21x2_ASAP7_75t_L g4556 ( 
.A1(n_4105),
.A2(n_3304),
.B(n_3401),
.Y(n_4556)
);

OAI21x1_ASAP7_75t_L g4557 ( 
.A1(n_3785),
.A2(n_3294),
.B(n_3314),
.Y(n_4557)
);

HB1xp67_ASAP7_75t_L g4558 ( 
.A(n_3833),
.Y(n_4558)
);

INVx2_ASAP7_75t_SL g4559 ( 
.A(n_4068),
.Y(n_4559)
);

OAI21x1_ASAP7_75t_L g4560 ( 
.A1(n_3785),
.A2(n_3294),
.B(n_3411),
.Y(n_4560)
);

OAI22xp5_ASAP7_75t_L g4561 ( 
.A1(n_4103),
.A2(n_3294),
.B1(n_3411),
.B2(n_3305),
.Y(n_4561)
);

INVx1_ASAP7_75t_L g4562 ( 
.A(n_3821),
.Y(n_4562)
);

INVx1_ASAP7_75t_L g4563 ( 
.A(n_3821),
.Y(n_4563)
);

OAI21x1_ASAP7_75t_L g4564 ( 
.A1(n_3785),
.A2(n_3292),
.B(n_3305),
.Y(n_4564)
);

OR2x2_ASAP7_75t_L g4565 ( 
.A(n_4094),
.B(n_3240),
.Y(n_4565)
);

OAI22xp5_ASAP7_75t_L g4566 ( 
.A1(n_4103),
.A2(n_3305),
.B1(n_3411),
.B2(n_3382),
.Y(n_4566)
);

INVx1_ASAP7_75t_SL g4567 ( 
.A(n_3817),
.Y(n_4567)
);

OAI21x1_ASAP7_75t_L g4568 ( 
.A1(n_3788),
.A2(n_3418),
.B(n_3412),
.Y(n_4568)
);

NAND2xp33_ASAP7_75t_SL g4569 ( 
.A(n_3815),
.B(n_3178),
.Y(n_4569)
);

NOR2xp67_ASAP7_75t_L g4570 ( 
.A(n_3815),
.B(n_3178),
.Y(n_4570)
);

NAND3xp33_ASAP7_75t_L g4571 ( 
.A(n_3738),
.B(n_3178),
.C(n_3422),
.Y(n_4571)
);

INVx1_ASAP7_75t_L g4572 ( 
.A(n_3836),
.Y(n_4572)
);

HB1xp67_ASAP7_75t_L g4573 ( 
.A(n_3833),
.Y(n_4573)
);

INVx1_ASAP7_75t_SL g4574 ( 
.A(n_3817),
.Y(n_4574)
);

AND2x4_ASAP7_75t_L g4575 ( 
.A(n_3797),
.B(n_3913),
.Y(n_4575)
);

O2A1O1Ixp33_ASAP7_75t_SL g4576 ( 
.A1(n_3623),
.A2(n_3178),
.B(n_3422),
.C(n_3240),
.Y(n_4576)
);

INVx4_ASAP7_75t_L g4577 ( 
.A(n_3815),
.Y(n_4577)
);

HB1xp67_ASAP7_75t_L g4578 ( 
.A(n_3877),
.Y(n_4578)
);

AND2x6_ASAP7_75t_L g4579 ( 
.A(n_3655),
.B(n_3291),
.Y(n_4579)
);

AND2x2_ASAP7_75t_L g4580 ( 
.A(n_3801),
.B(n_3291),
.Y(n_4580)
);

OAI21x1_ASAP7_75t_L g4581 ( 
.A1(n_3788),
.A2(n_3291),
.B(n_3311),
.Y(n_4581)
);

OAI21xp5_ASAP7_75t_L g4582 ( 
.A1(n_3620),
.A2(n_3291),
.B(n_3311),
.Y(n_4582)
);

AOI21x1_ASAP7_75t_L g4583 ( 
.A1(n_3738),
.A2(n_3291),
.B(n_3311),
.Y(n_4583)
);

OAI21x1_ASAP7_75t_L g4584 ( 
.A1(n_3788),
.A2(n_3371),
.B(n_3372),
.Y(n_4584)
);

OAI21x1_ASAP7_75t_L g4585 ( 
.A1(n_3806),
.A2(n_3371),
.B(n_3372),
.Y(n_4585)
);

CKINVDCx5p33_ASAP7_75t_R g4586 ( 
.A(n_3745),
.Y(n_4586)
);

OA21x2_ASAP7_75t_L g4587 ( 
.A1(n_3835),
.A2(n_3371),
.B(n_3372),
.Y(n_4587)
);

OAI21x1_ASAP7_75t_L g4588 ( 
.A1(n_3806),
.A2(n_3371),
.B(n_3372),
.Y(n_4588)
);

NAND2xp5_ASAP7_75t_L g4589 ( 
.A(n_3720),
.B(n_3371),
.Y(n_4589)
);

NAND2xp5_ASAP7_75t_L g4590 ( 
.A(n_3720),
.B(n_3371),
.Y(n_4590)
);

OAI21x1_ASAP7_75t_L g4591 ( 
.A1(n_3806),
.A2(n_3372),
.B(n_3376),
.Y(n_4591)
);

OAI21x1_ASAP7_75t_SL g4592 ( 
.A1(n_3635),
.A2(n_3642),
.B(n_3636),
.Y(n_4592)
);

OAI21x1_ASAP7_75t_L g4593 ( 
.A1(n_3806),
.A2(n_3372),
.B(n_3376),
.Y(n_4593)
);

OA21x2_ASAP7_75t_L g4594 ( 
.A1(n_3835),
.A2(n_3376),
.B(n_3856),
.Y(n_4594)
);

A2O1A1Ixp33_ASAP7_75t_L g4595 ( 
.A1(n_4008),
.A2(n_3376),
.B(n_3739),
.C(n_3728),
.Y(n_4595)
);

OAI221xp5_ASAP7_75t_L g4596 ( 
.A1(n_3930),
.A2(n_3376),
.B1(n_4046),
.B2(n_4052),
.C(n_3978),
.Y(n_4596)
);

CKINVDCx8_ASAP7_75t_R g4597 ( 
.A(n_3981),
.Y(n_4597)
);

OAI21x1_ASAP7_75t_L g4598 ( 
.A1(n_3814),
.A2(n_3376),
.B(n_3846),
.Y(n_4598)
);

OAI21x1_ASAP7_75t_L g4599 ( 
.A1(n_3814),
.A2(n_3850),
.B(n_3846),
.Y(n_4599)
);

OAI21x1_ASAP7_75t_L g4600 ( 
.A1(n_3814),
.A2(n_3850),
.B(n_3846),
.Y(n_4600)
);

O2A1O1Ixp33_ASAP7_75t_L g4601 ( 
.A1(n_3843),
.A2(n_3624),
.B(n_3661),
.C(n_3620),
.Y(n_4601)
);

CKINVDCx5p33_ASAP7_75t_R g4602 ( 
.A(n_3745),
.Y(n_4602)
);

OAI21x1_ASAP7_75t_L g4603 ( 
.A1(n_3814),
.A2(n_3850),
.B(n_3846),
.Y(n_4603)
);

OAI21x1_ASAP7_75t_SL g4604 ( 
.A1(n_3635),
.A2(n_3642),
.B(n_3636),
.Y(n_4604)
);

OAI22xp5_ASAP7_75t_L g4605 ( 
.A1(n_4128),
.A2(n_3869),
.B1(n_3935),
.B2(n_3928),
.Y(n_4605)
);

NAND2x1p5_ASAP7_75t_L g4606 ( 
.A(n_3839),
.B(n_3849),
.Y(n_4606)
);

HB1xp67_ASAP7_75t_L g4607 ( 
.A(n_3877),
.Y(n_4607)
);

INVxp67_ASAP7_75t_L g4608 ( 
.A(n_3898),
.Y(n_4608)
);

NAND2xp5_ASAP7_75t_L g4609 ( 
.A(n_3735),
.B(n_3747),
.Y(n_4609)
);

OAI21x1_ASAP7_75t_L g4610 ( 
.A1(n_3850),
.A2(n_3865),
.B(n_3855),
.Y(n_4610)
);

INVxp33_ASAP7_75t_L g4611 ( 
.A(n_3951),
.Y(n_4611)
);

OAI22xp5_ASAP7_75t_L g4612 ( 
.A1(n_3928),
.A2(n_3935),
.B1(n_3997),
.B2(n_3960),
.Y(n_4612)
);

INVx3_ASAP7_75t_L g4613 ( 
.A(n_3619),
.Y(n_4613)
);

NOR2xp67_ASAP7_75t_L g4614 ( 
.A(n_3797),
.B(n_3907),
.Y(n_4614)
);

OAI21x1_ASAP7_75t_L g4615 ( 
.A1(n_3855),
.A2(n_3872),
.B(n_3865),
.Y(n_4615)
);

AOI21xp5_ASAP7_75t_L g4616 ( 
.A1(n_3849),
.A2(n_3957),
.B(n_3887),
.Y(n_4616)
);

OAI21x1_ASAP7_75t_L g4617 ( 
.A1(n_3855),
.A2(n_3872),
.B(n_3865),
.Y(n_4617)
);

OAI21x1_ASAP7_75t_L g4618 ( 
.A1(n_3855),
.A2(n_3872),
.B(n_3865),
.Y(n_4618)
);

OAI21xp33_ASAP7_75t_L g4619 ( 
.A1(n_4046),
.A2(n_4052),
.B(n_4007),
.Y(n_4619)
);

AND2x2_ASAP7_75t_SL g4620 ( 
.A(n_3913),
.B(n_3849),
.Y(n_4620)
);

O2A1O1Ixp33_ASAP7_75t_SL g4621 ( 
.A1(n_3715),
.A2(n_3906),
.B(n_3627),
.C(n_3843),
.Y(n_4621)
);

NAND2xp5_ASAP7_75t_L g4622 ( 
.A(n_3735),
.B(n_3747),
.Y(n_4622)
);

AO21x2_ASAP7_75t_L g4623 ( 
.A1(n_3856),
.A2(n_3899),
.B(n_4020),
.Y(n_4623)
);

A2O1A1Ixp33_ASAP7_75t_L g4624 ( 
.A1(n_3728),
.A2(n_3739),
.B(n_4014),
.C(n_4000),
.Y(n_4624)
);

HB1xp67_ASAP7_75t_L g4625 ( 
.A(n_3898),
.Y(n_4625)
);

O2A1O1Ixp33_ASAP7_75t_SL g4626 ( 
.A1(n_3727),
.A2(n_3977),
.B(n_3789),
.C(n_3633),
.Y(n_4626)
);

OAI21x1_ASAP7_75t_L g4627 ( 
.A1(n_3872),
.A2(n_3905),
.B(n_3882),
.Y(n_4627)
);

AOI221xp5_ASAP7_75t_L g4628 ( 
.A1(n_3762),
.A2(n_3773),
.B1(n_3816),
.B2(n_3795),
.C(n_3776),
.Y(n_4628)
);

AO31x2_ASAP7_75t_L g4629 ( 
.A1(n_4020),
.A2(n_3987),
.A3(n_3995),
.B(n_3985),
.Y(n_4629)
);

OAI22xp5_ASAP7_75t_L g4630 ( 
.A1(n_3928),
.A2(n_3935),
.B1(n_3997),
.B2(n_3960),
.Y(n_4630)
);

HB1xp67_ASAP7_75t_L g4631 ( 
.A(n_3911),
.Y(n_4631)
);

NAND2xp5_ASAP7_75t_L g4632 ( 
.A(n_3762),
.B(n_3773),
.Y(n_4632)
);

OA21x2_ASAP7_75t_L g4633 ( 
.A1(n_3899),
.A2(n_3958),
.B(n_3948),
.Y(n_4633)
);

OR2x2_ASAP7_75t_L g4634 ( 
.A(n_4094),
.B(n_4100),
.Y(n_4634)
);

HB1xp67_ASAP7_75t_L g4635 ( 
.A(n_3911),
.Y(n_4635)
);

O2A1O1Ixp33_ASAP7_75t_L g4636 ( 
.A1(n_3624),
.A2(n_3667),
.B(n_3673),
.C(n_3661),
.Y(n_4636)
);

AND2x2_ASAP7_75t_L g4637 ( 
.A(n_3801),
.B(n_4012),
.Y(n_4637)
);

O2A1O1Ixp33_ASAP7_75t_L g4638 ( 
.A1(n_3667),
.A2(n_3692),
.B(n_3701),
.C(n_3673),
.Y(n_4638)
);

NAND2x1p5_ASAP7_75t_L g4639 ( 
.A(n_3849),
.B(n_3887),
.Y(n_4639)
);

OAI22xp33_ASAP7_75t_L g4640 ( 
.A1(n_3964),
.A2(n_3966),
.B1(n_3973),
.B2(n_3921),
.Y(n_4640)
);

BUFx2_ASAP7_75t_L g4641 ( 
.A(n_3767),
.Y(n_4641)
);

OAI22xp5_ASAP7_75t_L g4642 ( 
.A1(n_3960),
.A2(n_3997),
.B1(n_4109),
.B2(n_4079),
.Y(n_4642)
);

BUFx2_ASAP7_75t_L g4643 ( 
.A(n_3767),
.Y(n_4643)
);

CKINVDCx16_ASAP7_75t_R g4644 ( 
.A(n_3750),
.Y(n_4644)
);

OAI21x1_ASAP7_75t_L g4645 ( 
.A1(n_3826),
.A2(n_3653),
.B(n_3649),
.Y(n_4645)
);

AND2x4_ASAP7_75t_L g4646 ( 
.A(n_3913),
.B(n_3619),
.Y(n_4646)
);

OAI21x1_ASAP7_75t_L g4647 ( 
.A1(n_3826),
.A2(n_3653),
.B(n_3649),
.Y(n_4647)
);

OAI22xp33_ASAP7_75t_L g4648 ( 
.A1(n_3964),
.A2(n_3966),
.B1(n_3973),
.B2(n_3921),
.Y(n_4648)
);

NAND2xp5_ASAP7_75t_L g4649 ( 
.A(n_3776),
.B(n_3795),
.Y(n_4649)
);

AO21x1_ASAP7_75t_L g4650 ( 
.A1(n_3816),
.A2(n_3825),
.B(n_3824),
.Y(n_4650)
);

INVx1_ASAP7_75t_L g4651 ( 
.A(n_3985),
.Y(n_4651)
);

INVx1_ASAP7_75t_L g4652 ( 
.A(n_3987),
.Y(n_4652)
);

INVx1_ASAP7_75t_L g4653 ( 
.A(n_3995),
.Y(n_4653)
);

AOI21xp5_ASAP7_75t_SL g4654 ( 
.A1(n_3973),
.A2(n_3707),
.B(n_3697),
.Y(n_4654)
);

AOI22xp33_ASAP7_75t_L g4655 ( 
.A1(n_4087),
.A2(n_3614),
.B1(n_4044),
.B2(n_4036),
.Y(n_4655)
);

AO21x2_ASAP7_75t_L g4656 ( 
.A1(n_3958),
.A2(n_3998),
.B(n_3965),
.Y(n_4656)
);

HB1xp67_ASAP7_75t_L g4657 ( 
.A(n_3924),
.Y(n_4657)
);

OAI22xp5_ASAP7_75t_L g4658 ( 
.A1(n_4079),
.A2(n_4109),
.B1(n_3908),
.B2(n_3922),
.Y(n_4658)
);

OAI21xp5_ASAP7_75t_L g4659 ( 
.A1(n_3692),
.A2(n_3701),
.B(n_3703),
.Y(n_4659)
);

AND2x4_ASAP7_75t_L g4660 ( 
.A(n_3913),
.B(n_3619),
.Y(n_4660)
);

OA21x2_ASAP7_75t_L g4661 ( 
.A1(n_3958),
.A2(n_3998),
.B(n_3965),
.Y(n_4661)
);

HB1xp67_ASAP7_75t_L g4662 ( 
.A(n_3924),
.Y(n_4662)
);

OAI21xp5_ASAP7_75t_L g4663 ( 
.A1(n_3703),
.A2(n_3718),
.B(n_3887),
.Y(n_4663)
);

OR2x6_ASAP7_75t_L g4664 ( 
.A(n_3973),
.B(n_4033),
.Y(n_4664)
);

NAND2xp5_ASAP7_75t_L g4665 ( 
.A(n_3824),
.B(n_3825),
.Y(n_4665)
);

AOI22xp33_ASAP7_75t_L g4666 ( 
.A1(n_4087),
.A2(n_3614),
.B1(n_4044),
.B2(n_4036),
.Y(n_4666)
);

OR2x2_ASAP7_75t_L g4667 ( 
.A(n_4100),
.B(n_3908),
.Y(n_4667)
);

NAND2xp5_ASAP7_75t_L g4668 ( 
.A(n_3830),
.B(n_3831),
.Y(n_4668)
);

NAND2xp5_ASAP7_75t_L g4669 ( 
.A(n_3830),
.B(n_3831),
.Y(n_4669)
);

CKINVDCx20_ASAP7_75t_R g4670 ( 
.A(n_4249),
.Y(n_4670)
);

AOI222xp33_ASAP7_75t_L g4671 ( 
.A1(n_4152),
.A2(n_4087),
.B1(n_3718),
.B2(n_3946),
.C1(n_3854),
.C2(n_3873),
.Y(n_4671)
);

NAND2xp5_ASAP7_75t_L g4672 ( 
.A(n_4650),
.B(n_4001),
.Y(n_4672)
);

AND2x4_ASAP7_75t_L g4673 ( 
.A(n_4646),
.B(n_3619),
.Y(n_4673)
);

INVx2_ASAP7_75t_L g4674 ( 
.A(n_4633),
.Y(n_4674)
);

INVx6_ASAP7_75t_L g4675 ( 
.A(n_4222),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_4629),
.Y(n_4676)
);

INVx1_ASAP7_75t_L g4677 ( 
.A(n_4629),
.Y(n_4677)
);

INVx2_ASAP7_75t_L g4678 ( 
.A(n_4633),
.Y(n_4678)
);

AND2x2_ASAP7_75t_L g4679 ( 
.A(n_4386),
.B(n_3908),
.Y(n_4679)
);

CKINVDCx6p67_ASAP7_75t_R g4680 ( 
.A(n_4222),
.Y(n_4680)
);

BUFx3_ASAP7_75t_L g4681 ( 
.A(n_4222),
.Y(n_4681)
);

HB1xp67_ASAP7_75t_L g4682 ( 
.A(n_4227),
.Y(n_4682)
);

AO21x1_ASAP7_75t_SL g4683 ( 
.A1(n_4469),
.A2(n_4330),
.B(n_4349),
.Y(n_4683)
);

INVx1_ASAP7_75t_SL g4684 ( 
.A(n_4318),
.Y(n_4684)
);

CKINVDCx11_ASAP7_75t_R g4685 ( 
.A(n_4302),
.Y(n_4685)
);

INVx1_ASAP7_75t_L g4686 ( 
.A(n_4629),
.Y(n_4686)
);

INVx2_ASAP7_75t_L g4687 ( 
.A(n_4633),
.Y(n_4687)
);

AOI22xp33_ASAP7_75t_SL g4688 ( 
.A1(n_4425),
.A2(n_4087),
.B1(n_4000),
.B2(n_4016),
.Y(n_4688)
);

OA21x2_ASAP7_75t_L g4689 ( 
.A1(n_4163),
.A2(n_3748),
.B(n_3717),
.Y(n_4689)
);

AO21x2_ASAP7_75t_L g4690 ( 
.A1(n_4540),
.A2(n_3998),
.B(n_3965),
.Y(n_4690)
);

AOI22xp33_ASAP7_75t_L g4691 ( 
.A1(n_4452),
.A2(n_4087),
.B1(n_3614),
.B2(n_4044),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_4629),
.Y(n_4692)
);

AND2x2_ASAP7_75t_L g4693 ( 
.A(n_4386),
.B(n_3922),
.Y(n_4693)
);

INVx1_ASAP7_75t_L g4694 ( 
.A(n_4629),
.Y(n_4694)
);

HB1xp67_ASAP7_75t_L g4695 ( 
.A(n_4255),
.Y(n_4695)
);

INVx2_ASAP7_75t_L g4696 ( 
.A(n_4633),
.Y(n_4696)
);

CKINVDCx20_ASAP7_75t_R g4697 ( 
.A(n_4354),
.Y(n_4697)
);

INVx2_ASAP7_75t_L g4698 ( 
.A(n_4633),
.Y(n_4698)
);

BUFx2_ASAP7_75t_L g4699 ( 
.A(n_4386),
.Y(n_4699)
);

AO21x1_ASAP7_75t_L g4700 ( 
.A1(n_4167),
.A2(n_3854),
.B(n_3845),
.Y(n_4700)
);

INVx1_ASAP7_75t_L g4701 ( 
.A(n_4629),
.Y(n_4701)
);

INVx2_ASAP7_75t_L g4702 ( 
.A(n_4545),
.Y(n_4702)
);

INVx2_ASAP7_75t_L g4703 ( 
.A(n_4545),
.Y(n_4703)
);

INVx1_ASAP7_75t_L g4704 ( 
.A(n_4132),
.Y(n_4704)
);

BUFx2_ASAP7_75t_L g4705 ( 
.A(n_4386),
.Y(n_4705)
);

CKINVDCx5p33_ASAP7_75t_R g4706 ( 
.A(n_4378),
.Y(n_4706)
);

BUFx2_ASAP7_75t_L g4707 ( 
.A(n_4386),
.Y(n_4707)
);

AND2x4_ASAP7_75t_L g4708 ( 
.A(n_4646),
.B(n_3647),
.Y(n_4708)
);

HB1xp67_ASAP7_75t_L g4709 ( 
.A(n_4279),
.Y(n_4709)
);

INVx1_ASAP7_75t_L g4710 ( 
.A(n_4132),
.Y(n_4710)
);

NAND2x1p5_ASAP7_75t_L g4711 ( 
.A(n_4620),
.B(n_3907),
.Y(n_4711)
);

OAI22xp33_ASAP7_75t_L g4712 ( 
.A1(n_4234),
.A2(n_3973),
.B1(n_3739),
.B2(n_3728),
.Y(n_4712)
);

CKINVDCx11_ASAP7_75t_R g4713 ( 
.A(n_4509),
.Y(n_4713)
);

INVx2_ASAP7_75t_L g4714 ( 
.A(n_4556),
.Y(n_4714)
);

BUFx6f_ASAP7_75t_L g4715 ( 
.A(n_4386),
.Y(n_4715)
);

INVx2_ASAP7_75t_L g4716 ( 
.A(n_4556),
.Y(n_4716)
);

INVx2_ASAP7_75t_L g4717 ( 
.A(n_4556),
.Y(n_4717)
);

AND2x2_ASAP7_75t_L g4718 ( 
.A(n_4386),
.B(n_3922),
.Y(n_4718)
);

INVx1_ASAP7_75t_L g4719 ( 
.A(n_4137),
.Y(n_4719)
);

INVx3_ASAP7_75t_L g4720 ( 
.A(n_4646),
.Y(n_4720)
);

INVx2_ASAP7_75t_L g4721 ( 
.A(n_4556),
.Y(n_4721)
);

AND2x4_ASAP7_75t_L g4722 ( 
.A(n_4646),
.B(n_3647),
.Y(n_4722)
);

INVx2_ASAP7_75t_L g4723 ( 
.A(n_4661),
.Y(n_4723)
);

INVx3_ASAP7_75t_L g4724 ( 
.A(n_4660),
.Y(n_4724)
);

AOI22xp33_ASAP7_75t_SL g4725 ( 
.A1(n_4425),
.A2(n_4000),
.B1(n_4016),
.B2(n_4014),
.Y(n_4725)
);

NAND2x1p5_ASAP7_75t_L g4726 ( 
.A(n_4620),
.B(n_3907),
.Y(n_4726)
);

INVx1_ASAP7_75t_L g4727 ( 
.A(n_4137),
.Y(n_4727)
);

INVx2_ASAP7_75t_L g4728 ( 
.A(n_4661),
.Y(n_4728)
);

AOI22xp33_ASAP7_75t_L g4729 ( 
.A1(n_4452),
.A2(n_3614),
.B1(n_4044),
.B2(n_4036),
.Y(n_4729)
);

INVx1_ASAP7_75t_L g4730 ( 
.A(n_4145),
.Y(n_4730)
);

HB1xp67_ASAP7_75t_L g4731 ( 
.A(n_4467),
.Y(n_4731)
);

BUFx3_ASAP7_75t_L g4732 ( 
.A(n_4385),
.Y(n_4732)
);

HB1xp67_ASAP7_75t_L g4733 ( 
.A(n_4177),
.Y(n_4733)
);

INVx2_ASAP7_75t_L g4734 ( 
.A(n_4661),
.Y(n_4734)
);

BUFx8_ASAP7_75t_L g4735 ( 
.A(n_4509),
.Y(n_4735)
);

OA21x2_ASAP7_75t_L g4736 ( 
.A1(n_4163),
.A2(n_3748),
.B(n_3717),
.Y(n_4736)
);

OAI22xp5_ASAP7_75t_L g4737 ( 
.A1(n_4215),
.A2(n_4079),
.B1(n_4109),
.B2(n_3982),
.Y(n_4737)
);

AOI222xp33_ASAP7_75t_L g4738 ( 
.A1(n_4152),
.A2(n_3946),
.B1(n_3845),
.B2(n_3857),
.C1(n_3892),
.C2(n_3888),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_4145),
.Y(n_4739)
);

OA21x2_ASAP7_75t_L g4740 ( 
.A1(n_4163),
.A2(n_3970),
.B(n_3969),
.Y(n_4740)
);

AOI22xp33_ASAP7_75t_L g4741 ( 
.A1(n_4138),
.A2(n_3614),
.B1(n_4044),
.B2(n_4036),
.Y(n_4741)
);

AOI22xp33_ASAP7_75t_L g4742 ( 
.A1(n_4175),
.A2(n_3614),
.B1(n_4044),
.B2(n_4036),
.Y(n_4742)
);

AOI21x1_ASAP7_75t_L g4743 ( 
.A1(n_4226),
.A2(n_4058),
.B(n_4042),
.Y(n_4743)
);

NAND2x1p5_ASAP7_75t_L g4744 ( 
.A(n_4620),
.B(n_3907),
.Y(n_4744)
);

INVx2_ASAP7_75t_L g4745 ( 
.A(n_4661),
.Y(n_4745)
);

BUFx2_ASAP7_75t_L g4746 ( 
.A(n_4262),
.Y(n_4746)
);

CKINVDCx20_ASAP7_75t_R g4747 ( 
.A(n_4252),
.Y(n_4747)
);

BUFx8_ASAP7_75t_L g4748 ( 
.A(n_4509),
.Y(n_4748)
);

OAI21x1_ASAP7_75t_L g4749 ( 
.A1(n_4270),
.A2(n_3663),
.B(n_3649),
.Y(n_4749)
);

BUFx3_ASAP7_75t_L g4750 ( 
.A(n_4335),
.Y(n_4750)
);

AOI22xp33_ASAP7_75t_L g4751 ( 
.A1(n_4144),
.A2(n_3614),
.B1(n_4036),
.B2(n_3841),
.Y(n_4751)
);

BUFx4f_ASAP7_75t_SL g4752 ( 
.A(n_4290),
.Y(n_4752)
);

BUFx12f_ASAP7_75t_L g4753 ( 
.A(n_4366),
.Y(n_4753)
);

INVx2_ASAP7_75t_L g4754 ( 
.A(n_4661),
.Y(n_4754)
);

BUFx3_ASAP7_75t_L g4755 ( 
.A(n_4524),
.Y(n_4755)
);

AOI22xp33_ASAP7_75t_L g4756 ( 
.A1(n_4166),
.A2(n_3614),
.B1(n_3841),
.B2(n_3828),
.Y(n_4756)
);

AOI22xp33_ASAP7_75t_L g4757 ( 
.A1(n_4167),
.A2(n_3614),
.B1(n_3841),
.B2(n_3828),
.Y(n_4757)
);

INVx1_ASAP7_75t_L g4758 ( 
.A(n_4146),
.Y(n_4758)
);

INVx2_ASAP7_75t_L g4759 ( 
.A(n_4656),
.Y(n_4759)
);

INVx1_ASAP7_75t_L g4760 ( 
.A(n_4146),
.Y(n_4760)
);

BUFx3_ASAP7_75t_L g4761 ( 
.A(n_4524),
.Y(n_4761)
);

OAI21x1_ASAP7_75t_L g4762 ( 
.A1(n_4270),
.A2(n_3664),
.B(n_3663),
.Y(n_4762)
);

INVx2_ASAP7_75t_L g4763 ( 
.A(n_4656),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4172),
.Y(n_4764)
);

BUFx2_ASAP7_75t_L g4765 ( 
.A(n_4262),
.Y(n_4765)
);

AO21x1_ASAP7_75t_L g4766 ( 
.A1(n_4153),
.A2(n_4234),
.B(n_4300),
.Y(n_4766)
);

INVx1_ASAP7_75t_L g4767 ( 
.A(n_4172),
.Y(n_4767)
);

HB1xp67_ASAP7_75t_L g4768 ( 
.A(n_4221),
.Y(n_4768)
);

AND2x2_ASAP7_75t_L g4769 ( 
.A(n_4485),
.B(n_4012),
.Y(n_4769)
);

AOI22xp33_ASAP7_75t_L g4770 ( 
.A1(n_4247),
.A2(n_3614),
.B1(n_3841),
.B2(n_3828),
.Y(n_4770)
);

OAI22xp33_ASAP7_75t_L g4771 ( 
.A1(n_4257),
.A2(n_3973),
.B1(n_4033),
.B2(n_3885),
.Y(n_4771)
);

INVx1_ASAP7_75t_SL g4772 ( 
.A(n_4567),
.Y(n_4772)
);

BUFx2_ASAP7_75t_R g4773 ( 
.A(n_4239),
.Y(n_4773)
);

CKINVDCx5p33_ASAP7_75t_R g4774 ( 
.A(n_4383),
.Y(n_4774)
);

INVx1_ASAP7_75t_L g4775 ( 
.A(n_4183),
.Y(n_4775)
);

INVx2_ASAP7_75t_L g4776 ( 
.A(n_4656),
.Y(n_4776)
);

INVx3_ASAP7_75t_L g4777 ( 
.A(n_4660),
.Y(n_4777)
);

INVx1_ASAP7_75t_SL g4778 ( 
.A(n_4567),
.Y(n_4778)
);

AOI21x1_ASAP7_75t_L g4779 ( 
.A1(n_4226),
.A2(n_4058),
.B(n_4042),
.Y(n_4779)
);

INVx6_ASAP7_75t_L g4780 ( 
.A(n_4506),
.Y(n_4780)
);

BUFx10_ASAP7_75t_L g4781 ( 
.A(n_4288),
.Y(n_4781)
);

BUFx2_ASAP7_75t_L g4782 ( 
.A(n_4660),
.Y(n_4782)
);

INVx1_ASAP7_75t_L g4783 ( 
.A(n_4183),
.Y(n_4783)
);

AO21x1_ASAP7_75t_L g4784 ( 
.A1(n_4153),
.A2(n_3873),
.B(n_3857),
.Y(n_4784)
);

AND2x2_ASAP7_75t_L g4785 ( 
.A(n_4485),
.B(n_4486),
.Y(n_4785)
);

INVx1_ASAP7_75t_L g4786 ( 
.A(n_4189),
.Y(n_4786)
);

NAND2xp5_ASAP7_75t_L g4787 ( 
.A(n_4650),
.B(n_4001),
.Y(n_4787)
);

INVx2_ASAP7_75t_L g4788 ( 
.A(n_4656),
.Y(n_4788)
);

AOI21x1_ASAP7_75t_L g4789 ( 
.A1(n_4149),
.A2(n_4082),
.B(n_4078),
.Y(n_4789)
);

BUFx2_ASAP7_75t_L g4790 ( 
.A(n_4660),
.Y(n_4790)
);

AOI22xp33_ASAP7_75t_L g4791 ( 
.A1(n_4211),
.A2(n_4505),
.B1(n_4201),
.B2(n_4164),
.Y(n_4791)
);

NAND2xp5_ASAP7_75t_L g4792 ( 
.A(n_4544),
.B(n_4007),
.Y(n_4792)
);

INVx2_ASAP7_75t_L g4793 ( 
.A(n_4587),
.Y(n_4793)
);

BUFx4f_ASAP7_75t_L g4794 ( 
.A(n_4290),
.Y(n_4794)
);

AND2x4_ASAP7_75t_L g4795 ( 
.A(n_4575),
.B(n_3647),
.Y(n_4795)
);

CKINVDCx5p33_ASAP7_75t_R g4796 ( 
.A(n_4525),
.Y(n_4796)
);

AOI22xp33_ASAP7_75t_L g4797 ( 
.A1(n_4211),
.A2(n_3614),
.B1(n_3841),
.B2(n_3828),
.Y(n_4797)
);

BUFx3_ASAP7_75t_L g4798 ( 
.A(n_4524),
.Y(n_4798)
);

INVx1_ASAP7_75t_L g4799 ( 
.A(n_4189),
.Y(n_4799)
);

AND2x2_ASAP7_75t_L g4800 ( 
.A(n_4486),
.B(n_4519),
.Y(n_4800)
);

CKINVDCx11_ASAP7_75t_R g4801 ( 
.A(n_4644),
.Y(n_4801)
);

INVx2_ASAP7_75t_L g4802 ( 
.A(n_4587),
.Y(n_4802)
);

INVx1_ASAP7_75t_L g4803 ( 
.A(n_4202),
.Y(n_4803)
);

AND2x2_ASAP7_75t_L g4804 ( 
.A(n_4519),
.B(n_4535),
.Y(n_4804)
);

INVx11_ASAP7_75t_L g4805 ( 
.A(n_4244),
.Y(n_4805)
);

INVx1_ASAP7_75t_L g4806 ( 
.A(n_4202),
.Y(n_4806)
);

INVx6_ASAP7_75t_L g4807 ( 
.A(n_4506),
.Y(n_4807)
);

AOI22xp33_ASAP7_75t_L g4808 ( 
.A1(n_4505),
.A2(n_3990),
.B1(n_4033),
.B2(n_3979),
.Y(n_4808)
);

AOI22xp33_ASAP7_75t_L g4809 ( 
.A1(n_4201),
.A2(n_3990),
.B1(n_4033),
.B2(n_3979),
.Y(n_4809)
);

BUFx3_ASAP7_75t_L g4810 ( 
.A(n_4232),
.Y(n_4810)
);

INVx1_ASAP7_75t_L g4811 ( 
.A(n_4219),
.Y(n_4811)
);

BUFx2_ASAP7_75t_L g4812 ( 
.A(n_4421),
.Y(n_4812)
);

AOI22xp33_ASAP7_75t_L g4813 ( 
.A1(n_4164),
.A2(n_3990),
.B1(n_4033),
.B2(n_3979),
.Y(n_4813)
);

AND2x4_ASAP7_75t_L g4814 ( 
.A(n_4575),
.B(n_3647),
.Y(n_4814)
);

AOI22xp33_ASAP7_75t_L g4815 ( 
.A1(n_4135),
.A2(n_3990),
.B1(n_4033),
.B2(n_3979),
.Y(n_4815)
);

INVx2_ASAP7_75t_L g4816 ( 
.A(n_4587),
.Y(n_4816)
);

AOI22xp33_ASAP7_75t_L g4817 ( 
.A1(n_4135),
.A2(n_3990),
.B1(n_3979),
.B2(n_3781),
.Y(n_4817)
);

NAND2xp5_ASAP7_75t_L g4818 ( 
.A(n_4544),
.B(n_3860),
.Y(n_4818)
);

AOI22xp33_ASAP7_75t_L g4819 ( 
.A1(n_4292),
.A2(n_3990),
.B1(n_3781),
.B2(n_3876),
.Y(n_4819)
);

OAI22xp5_ASAP7_75t_L g4820 ( 
.A1(n_4215),
.A2(n_3982),
.B1(n_4049),
.B2(n_4047),
.Y(n_4820)
);

AND2x2_ASAP7_75t_L g4821 ( 
.A(n_4535),
.B(n_4483),
.Y(n_4821)
);

OAI22xp5_ASAP7_75t_L g4822 ( 
.A1(n_4257),
.A2(n_4050),
.B1(n_4073),
.B2(n_4049),
.Y(n_4822)
);

AND2x2_ASAP7_75t_L g4823 ( 
.A(n_4483),
.B(n_4012),
.Y(n_4823)
);

INVx1_ASAP7_75t_L g4824 ( 
.A(n_4219),
.Y(n_4824)
);

HB1xp67_ASAP7_75t_L g4825 ( 
.A(n_4475),
.Y(n_4825)
);

INVx2_ASAP7_75t_SL g4826 ( 
.A(n_4421),
.Y(n_4826)
);

NAND2x1p5_ASAP7_75t_L g4827 ( 
.A(n_4395),
.B(n_3907),
.Y(n_4827)
);

INVx2_ASAP7_75t_L g4828 ( 
.A(n_4587),
.Y(n_4828)
);

INVx1_ASAP7_75t_L g4829 ( 
.A(n_4220),
.Y(n_4829)
);

INVx1_ASAP7_75t_L g4830 ( 
.A(n_4220),
.Y(n_4830)
);

OAI22xp5_ASAP7_75t_L g4831 ( 
.A1(n_4286),
.A2(n_4073),
.B1(n_4075),
.B2(n_4050),
.Y(n_4831)
);

INVx2_ASAP7_75t_L g4832 ( 
.A(n_4587),
.Y(n_4832)
);

INVx6_ASAP7_75t_L g4833 ( 
.A(n_4506),
.Y(n_4833)
);

AOI22xp33_ASAP7_75t_L g4834 ( 
.A1(n_4188),
.A2(n_3781),
.B1(n_3876),
.B2(n_3758),
.Y(n_4834)
);

INVx1_ASAP7_75t_L g4835 ( 
.A(n_4223),
.Y(n_4835)
);

INVx4_ASAP7_75t_L g4836 ( 
.A(n_4288),
.Y(n_4836)
);

AND2x2_ASAP7_75t_L g4837 ( 
.A(n_4554),
.B(n_4077),
.Y(n_4837)
);

BUFx5_ASAP7_75t_L g4838 ( 
.A(n_4579),
.Y(n_4838)
);

OR2x6_ASAP7_75t_L g4839 ( 
.A(n_4654),
.B(n_3803),
.Y(n_4839)
);

INVx1_ASAP7_75t_L g4840 ( 
.A(n_4223),
.Y(n_4840)
);

INVx1_ASAP7_75t_L g4841 ( 
.A(n_4224),
.Y(n_4841)
);

INVx2_ASAP7_75t_L g4842 ( 
.A(n_4581),
.Y(n_4842)
);

AND2x2_ASAP7_75t_L g4843 ( 
.A(n_4554),
.B(n_4077),
.Y(n_4843)
);

AOI22xp33_ASAP7_75t_SL g4844 ( 
.A1(n_4332),
.A2(n_4016),
.B1(n_4018),
.B2(n_4014),
.Y(n_4844)
);

AO21x2_ASAP7_75t_L g4845 ( 
.A1(n_4539),
.A2(n_4005),
.B(n_4003),
.Y(n_4845)
);

INVx2_ASAP7_75t_SL g4846 ( 
.A(n_4437),
.Y(n_4846)
);

NAND2x1p5_ASAP7_75t_L g4847 ( 
.A(n_4395),
.B(n_3907),
.Y(n_4847)
);

CKINVDCx5p33_ASAP7_75t_R g4848 ( 
.A(n_4430),
.Y(n_4848)
);

INVx4_ASAP7_75t_L g4849 ( 
.A(n_4288),
.Y(n_4849)
);

INVx2_ASAP7_75t_L g4850 ( 
.A(n_4581),
.Y(n_4850)
);

INVx2_ASAP7_75t_L g4851 ( 
.A(n_4581),
.Y(n_4851)
);

INVx5_ASAP7_75t_L g4852 ( 
.A(n_4579),
.Y(n_4852)
);

CKINVDCx20_ASAP7_75t_R g4853 ( 
.A(n_4644),
.Y(n_4853)
);

NAND2x1p5_ASAP7_75t_L g4854 ( 
.A(n_4395),
.B(n_3910),
.Y(n_4854)
);

NAND2x1p5_ASAP7_75t_L g4855 ( 
.A(n_4395),
.B(n_3910),
.Y(n_4855)
);

AOI22xp33_ASAP7_75t_L g4856 ( 
.A1(n_4264),
.A2(n_3781),
.B1(n_3876),
.B2(n_3758),
.Y(n_4856)
);

INVx1_ASAP7_75t_L g4857 ( 
.A(n_4224),
.Y(n_4857)
);

INVx2_ASAP7_75t_L g4858 ( 
.A(n_4584),
.Y(n_4858)
);

BUFx6f_ASAP7_75t_L g4859 ( 
.A(n_4139),
.Y(n_4859)
);

BUFx6f_ASAP7_75t_L g4860 ( 
.A(n_4139),
.Y(n_4860)
);

AOI22xp33_ASAP7_75t_SL g4861 ( 
.A1(n_4332),
.A2(n_4286),
.B1(n_4284),
.B2(n_4300),
.Y(n_4861)
);

NAND2x1p5_ASAP7_75t_L g4862 ( 
.A(n_4395),
.B(n_3910),
.Y(n_4862)
);

OR2x2_ASAP7_75t_L g4863 ( 
.A(n_4133),
.B(n_4077),
.Y(n_4863)
);

CKINVDCx5p33_ASAP7_75t_R g4864 ( 
.A(n_4482),
.Y(n_4864)
);

AND2x4_ASAP7_75t_L g4865 ( 
.A(n_4575),
.B(n_4161),
.Y(n_4865)
);

INVx1_ASAP7_75t_L g4866 ( 
.A(n_4236),
.Y(n_4866)
);

HB1xp67_ASAP7_75t_L g4867 ( 
.A(n_4513),
.Y(n_4867)
);

BUFx6f_ASAP7_75t_L g4868 ( 
.A(n_4139),
.Y(n_4868)
);

BUFx6f_ASAP7_75t_L g4869 ( 
.A(n_4139),
.Y(n_4869)
);

INVx1_ASAP7_75t_L g4870 ( 
.A(n_4236),
.Y(n_4870)
);

AO21x2_ASAP7_75t_L g4871 ( 
.A1(n_4539),
.A2(n_4005),
.B(n_4003),
.Y(n_4871)
);

INVx1_ASAP7_75t_SL g4872 ( 
.A(n_4574),
.Y(n_4872)
);

AND2x2_ASAP7_75t_L g4873 ( 
.A(n_4453),
.B(n_4117),
.Y(n_4873)
);

CKINVDCx5p33_ASAP7_75t_R g4874 ( 
.A(n_4488),
.Y(n_4874)
);

INVx1_ASAP7_75t_L g4875 ( 
.A(n_4251),
.Y(n_4875)
);

AO21x2_ASAP7_75t_L g4876 ( 
.A1(n_4542),
.A2(n_4005),
.B(n_4003),
.Y(n_4876)
);

INVx1_ASAP7_75t_L g4877 ( 
.A(n_4251),
.Y(n_4877)
);

INVx1_ASAP7_75t_L g4878 ( 
.A(n_4263),
.Y(n_4878)
);

INVx3_ASAP7_75t_L g4879 ( 
.A(n_4613),
.Y(n_4879)
);

INVx2_ASAP7_75t_L g4880 ( 
.A(n_4584),
.Y(n_4880)
);

INVx2_ASAP7_75t_L g4881 ( 
.A(n_4584),
.Y(n_4881)
);

BUFx3_ASAP7_75t_L g4882 ( 
.A(n_4232),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4263),
.Y(n_4883)
);

BUFx12f_ASAP7_75t_L g4884 ( 
.A(n_4497),
.Y(n_4884)
);

OA21x2_ASAP7_75t_L g4885 ( 
.A1(n_4151),
.A2(n_3970),
.B(n_3969),
.Y(n_4885)
);

HB1xp67_ASAP7_75t_L g4886 ( 
.A(n_4516),
.Y(n_4886)
);

CKINVDCx5p33_ASAP7_75t_R g4887 ( 
.A(n_4532),
.Y(n_4887)
);

NAND2xp5_ASAP7_75t_L g4888 ( 
.A(n_4549),
.B(n_3860),
.Y(n_4888)
);

INVx4_ASAP7_75t_L g4889 ( 
.A(n_4288),
.Y(n_4889)
);

HB1xp67_ASAP7_75t_L g4890 ( 
.A(n_4523),
.Y(n_4890)
);

BUFx12f_ASAP7_75t_L g4891 ( 
.A(n_4538),
.Y(n_4891)
);

AOI22xp33_ASAP7_75t_L g4892 ( 
.A1(n_4264),
.A2(n_3781),
.B1(n_3876),
.B2(n_3758),
.Y(n_4892)
);

INVx2_ASAP7_75t_L g4893 ( 
.A(n_4585),
.Y(n_4893)
);

BUFx3_ASAP7_75t_L g4894 ( 
.A(n_4232),
.Y(n_4894)
);

INVxp33_ASAP7_75t_L g4895 ( 
.A(n_4611),
.Y(n_4895)
);

AOI22xp33_ASAP7_75t_L g4896 ( 
.A1(n_4307),
.A2(n_3876),
.B1(n_3758),
.B2(n_3961),
.Y(n_4896)
);

AND2x2_ASAP7_75t_L g4897 ( 
.A(n_4453),
.B(n_4117),
.Y(n_4897)
);

INVx2_ASAP7_75t_L g4898 ( 
.A(n_4585),
.Y(n_4898)
);

OAI22xp33_ASAP7_75t_L g4899 ( 
.A1(n_4520),
.A2(n_4203),
.B1(n_4204),
.B2(n_4284),
.Y(n_4899)
);

INVx1_ASAP7_75t_L g4900 ( 
.A(n_4265),
.Y(n_4900)
);

BUFx12f_ASAP7_75t_L g4901 ( 
.A(n_4586),
.Y(n_4901)
);

AND2x4_ASAP7_75t_L g4902 ( 
.A(n_4575),
.B(n_3647),
.Y(n_4902)
);

INVx1_ASAP7_75t_L g4903 ( 
.A(n_4265),
.Y(n_4903)
);

OA21x2_ASAP7_75t_L g4904 ( 
.A1(n_4151),
.A2(n_3972),
.B(n_4019),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4267),
.Y(n_4905)
);

INVx3_ASAP7_75t_L g4906 ( 
.A(n_4613),
.Y(n_4906)
);

INVx8_ASAP7_75t_L g4907 ( 
.A(n_4232),
.Y(n_4907)
);

INVx1_ASAP7_75t_L g4908 ( 
.A(n_4267),
.Y(n_4908)
);

NAND2xp5_ASAP7_75t_L g4909 ( 
.A(n_4549),
.B(n_3864),
.Y(n_4909)
);

OAI21xp5_ASAP7_75t_L g4910 ( 
.A1(n_4148),
.A2(n_3961),
.B(n_3903),
.Y(n_4910)
);

AND2x2_ASAP7_75t_L g4911 ( 
.A(n_4637),
.B(n_4117),
.Y(n_4911)
);

NAND2xp5_ASAP7_75t_L g4912 ( 
.A(n_4140),
.B(n_3864),
.Y(n_4912)
);

OAI22xp5_ASAP7_75t_L g4913 ( 
.A1(n_4196),
.A2(n_4113),
.B1(n_4075),
.B2(n_3931),
.Y(n_4913)
);

INVx2_ASAP7_75t_L g4914 ( 
.A(n_4585),
.Y(n_4914)
);

INVx1_ASAP7_75t_L g4915 ( 
.A(n_4274),
.Y(n_4915)
);

INVx1_ASAP7_75t_L g4916 ( 
.A(n_4274),
.Y(n_4916)
);

CKINVDCx5p33_ASAP7_75t_R g4917 ( 
.A(n_4602),
.Y(n_4917)
);

AOI22xp33_ASAP7_75t_SL g4918 ( 
.A1(n_4131),
.A2(n_4018),
.B1(n_3827),
.B2(n_3885),
.Y(n_4918)
);

INVx1_ASAP7_75t_L g4919 ( 
.A(n_4278),
.Y(n_4919)
);

OAI22xp5_ASAP7_75t_L g4920 ( 
.A1(n_4196),
.A2(n_4113),
.B1(n_3931),
.B2(n_3953),
.Y(n_4920)
);

NAND2xp5_ASAP7_75t_L g4921 ( 
.A(n_4140),
.B(n_3883),
.Y(n_4921)
);

INVx2_ASAP7_75t_SL g4922 ( 
.A(n_4437),
.Y(n_4922)
);

CKINVDCx5p33_ASAP7_75t_R g4923 ( 
.A(n_4290),
.Y(n_4923)
);

INVx2_ASAP7_75t_L g4924 ( 
.A(n_4588),
.Y(n_4924)
);

INVx2_ASAP7_75t_L g4925 ( 
.A(n_4588),
.Y(n_4925)
);

NAND2x1p5_ASAP7_75t_L g4926 ( 
.A(n_4395),
.B(n_3910),
.Y(n_4926)
);

AO21x1_ASAP7_75t_L g4927 ( 
.A1(n_4531),
.A2(n_4569),
.B(n_4131),
.Y(n_4927)
);

INVx2_ASAP7_75t_SL g4928 ( 
.A(n_4500),
.Y(n_4928)
);

OR2x2_ASAP7_75t_L g4929 ( 
.A(n_4133),
.B(n_3888),
.Y(n_4929)
);

INVx1_ASAP7_75t_L g4930 ( 
.A(n_4278),
.Y(n_4930)
);

BUFx3_ASAP7_75t_L g4931 ( 
.A(n_4232),
.Y(n_4931)
);

CKINVDCx16_ASAP7_75t_R g4932 ( 
.A(n_4533),
.Y(n_4932)
);

INVx1_ASAP7_75t_L g4933 ( 
.A(n_4280),
.Y(n_4933)
);

INVx3_ASAP7_75t_L g4934 ( 
.A(n_4613),
.Y(n_4934)
);

OAI22xp5_ASAP7_75t_L g4935 ( 
.A1(n_4148),
.A2(n_4113),
.B1(n_3931),
.B2(n_3953),
.Y(n_4935)
);

AO21x1_ASAP7_75t_L g4936 ( 
.A1(n_4531),
.A2(n_3929),
.B(n_3892),
.Y(n_4936)
);

AND2x4_ASAP7_75t_L g4937 ( 
.A(n_4161),
.B(n_3680),
.Y(n_4937)
);

CKINVDCx20_ASAP7_75t_R g4938 ( 
.A(n_4411),
.Y(n_4938)
);

AOI22xp33_ASAP7_75t_L g4939 ( 
.A1(n_4307),
.A2(n_3758),
.B1(n_4027),
.B2(n_3994),
.Y(n_4939)
);

AOI22xp33_ASAP7_75t_L g4940 ( 
.A1(n_4203),
.A2(n_4027),
.B1(n_3994),
.B2(n_3707),
.Y(n_4940)
);

NAND2xp5_ASAP7_75t_L g4941 ( 
.A(n_4154),
.B(n_3883),
.Y(n_4941)
);

INVx4_ASAP7_75t_L g4942 ( 
.A(n_4288),
.Y(n_4942)
);

HB1xp67_ASAP7_75t_L g4943 ( 
.A(n_4548),
.Y(n_4943)
);

AOI22xp5_ASAP7_75t_L g4944 ( 
.A1(n_4214),
.A2(n_3819),
.B1(n_3946),
.B2(n_3929),
.Y(n_4944)
);

NAND2xp5_ASAP7_75t_L g4945 ( 
.A(n_4154),
.B(n_3895),
.Y(n_4945)
);

AND2x4_ASAP7_75t_L g4946 ( 
.A(n_4161),
.B(n_3680),
.Y(n_4946)
);

INVx1_ASAP7_75t_SL g4947 ( 
.A(n_4574),
.Y(n_4947)
);

INVx4_ASAP7_75t_L g4948 ( 
.A(n_4484),
.Y(n_4948)
);

INVx1_ASAP7_75t_SL g4949 ( 
.A(n_4412),
.Y(n_4949)
);

INVx1_ASAP7_75t_L g4950 ( 
.A(n_4280),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_4282),
.Y(n_4951)
);

AOI21x1_ASAP7_75t_L g4952 ( 
.A1(n_4149),
.A2(n_4082),
.B(n_4078),
.Y(n_4952)
);

INVx6_ASAP7_75t_L g4953 ( 
.A(n_4506),
.Y(n_4953)
);

INVxp67_ASAP7_75t_SL g4954 ( 
.A(n_4148),
.Y(n_4954)
);

INVx1_ASAP7_75t_L g4955 ( 
.A(n_4282),
.Y(n_4955)
);

INVx1_ASAP7_75t_L g4956 ( 
.A(n_4283),
.Y(n_4956)
);

INVx2_ASAP7_75t_L g4957 ( 
.A(n_4588),
.Y(n_4957)
);

BUFx12f_ASAP7_75t_L g4958 ( 
.A(n_4277),
.Y(n_4958)
);

OAI22xp5_ASAP7_75t_L g4959 ( 
.A1(n_4303),
.A2(n_3953),
.B1(n_3963),
.B2(n_3909),
.Y(n_4959)
);

OAI22xp5_ASAP7_75t_L g4960 ( 
.A1(n_4165),
.A2(n_3963),
.B1(n_3968),
.B2(n_3909),
.Y(n_4960)
);

BUFx6f_ASAP7_75t_L g4961 ( 
.A(n_4139),
.Y(n_4961)
);

INVx2_ASAP7_75t_L g4962 ( 
.A(n_4591),
.Y(n_4962)
);

AOI22xp33_ASAP7_75t_L g4963 ( 
.A1(n_4204),
.A2(n_4027),
.B1(n_3994),
.B2(n_3707),
.Y(n_4963)
);

INVx1_ASAP7_75t_L g4964 ( 
.A(n_4283),
.Y(n_4964)
);

BUFx10_ASAP7_75t_L g4965 ( 
.A(n_4484),
.Y(n_4965)
);

AND2x2_ASAP7_75t_L g4966 ( 
.A(n_4637),
.B(n_4119),
.Y(n_4966)
);

HB1xp67_ASAP7_75t_L g4967 ( 
.A(n_4558),
.Y(n_4967)
);

INVx1_ASAP7_75t_L g4968 ( 
.A(n_4291),
.Y(n_4968)
);

INVx6_ASAP7_75t_L g4969 ( 
.A(n_4161),
.Y(n_4969)
);

INVx1_ASAP7_75t_L g4970 ( 
.A(n_4291),
.Y(n_4970)
);

INVx2_ASAP7_75t_L g4971 ( 
.A(n_4591),
.Y(n_4971)
);

BUFx3_ASAP7_75t_L g4972 ( 
.A(n_4232),
.Y(n_4972)
);

BUFx2_ASAP7_75t_L g4973 ( 
.A(n_4456),
.Y(n_4973)
);

INVx2_ASAP7_75t_L g4974 ( 
.A(n_4591),
.Y(n_4974)
);

AOI22xp33_ASAP7_75t_SL g4975 ( 
.A1(n_4479),
.A2(n_4018),
.B1(n_3885),
.B2(n_3827),
.Y(n_4975)
);

OR2x6_ASAP7_75t_L g4976 ( 
.A(n_4654),
.B(n_3803),
.Y(n_4976)
);

INVx1_ASAP7_75t_L g4977 ( 
.A(n_4296),
.Y(n_4977)
);

INVx2_ASAP7_75t_L g4978 ( 
.A(n_4593),
.Y(n_4978)
);

INVx1_ASAP7_75t_L g4979 ( 
.A(n_4296),
.Y(n_4979)
);

INVx1_ASAP7_75t_L g4980 ( 
.A(n_4299),
.Y(n_4980)
);

AOI22xp33_ASAP7_75t_SL g4981 ( 
.A1(n_4542),
.A2(n_3807),
.B1(n_3834),
.B2(n_3827),
.Y(n_4981)
);

INVx2_ASAP7_75t_L g4982 ( 
.A(n_4593),
.Y(n_4982)
);

INVx2_ASAP7_75t_L g4983 ( 
.A(n_4593),
.Y(n_4983)
);

INVx1_ASAP7_75t_L g4984 ( 
.A(n_4299),
.Y(n_4984)
);

INVx2_ASAP7_75t_L g4985 ( 
.A(n_4304),
.Y(n_4985)
);

INVx2_ASAP7_75t_L g4986 ( 
.A(n_4304),
.Y(n_4986)
);

AOI22xp33_ASAP7_75t_L g4987 ( 
.A1(n_4520),
.A2(n_3994),
.B1(n_4027),
.B2(n_3697),
.Y(n_4987)
);

INVx4_ASAP7_75t_L g4988 ( 
.A(n_4484),
.Y(n_4988)
);

INVx1_ASAP7_75t_L g4989 ( 
.A(n_4306),
.Y(n_4989)
);

INVx1_ASAP7_75t_L g4990 ( 
.A(n_4306),
.Y(n_4990)
);

AOI21xp5_ASAP7_75t_SL g4991 ( 
.A1(n_4494),
.A2(n_4481),
.B(n_4396),
.Y(n_4991)
);

HB1xp67_ASAP7_75t_L g4992 ( 
.A(n_4573),
.Y(n_4992)
);

AO21x2_ASAP7_75t_L g4993 ( 
.A1(n_4571),
.A2(n_4029),
.B(n_4019),
.Y(n_4993)
);

BUFx3_ASAP7_75t_L g4994 ( 
.A(n_4484),
.Y(n_4994)
);

INVx1_ASAP7_75t_L g4995 ( 
.A(n_4311),
.Y(n_4995)
);

INVx3_ASAP7_75t_L g4996 ( 
.A(n_4613),
.Y(n_4996)
);

CKINVDCx5p33_ASAP7_75t_R g4997 ( 
.A(n_4411),
.Y(n_4997)
);

BUFx2_ASAP7_75t_R g4998 ( 
.A(n_4216),
.Y(n_4998)
);

OAI22xp5_ASAP7_75t_L g4999 ( 
.A1(n_4165),
.A2(n_4412),
.B1(n_4325),
.B2(n_4273),
.Y(n_4999)
);

INVx2_ASAP7_75t_L g5000 ( 
.A(n_4304),
.Y(n_5000)
);

NAND2xp5_ASAP7_75t_L g5001 ( 
.A(n_4628),
.B(n_4294),
.Y(n_5001)
);

INVx1_ASAP7_75t_L g5002 ( 
.A(n_4311),
.Y(n_5002)
);

INVx1_ASAP7_75t_L g5003 ( 
.A(n_4315),
.Y(n_5003)
);

INVx1_ASAP7_75t_L g5004 ( 
.A(n_4315),
.Y(n_5004)
);

INVx2_ASAP7_75t_L g5005 ( 
.A(n_4304),
.Y(n_5005)
);

INVx4_ASAP7_75t_SL g5006 ( 
.A(n_4484),
.Y(n_5006)
);

INVx2_ASAP7_75t_L g5007 ( 
.A(n_4304),
.Y(n_5007)
);

INVx2_ASAP7_75t_L g5008 ( 
.A(n_4304),
.Y(n_5008)
);

CKINVDCx20_ASAP7_75t_R g5009 ( 
.A(n_4411),
.Y(n_5009)
);

INVx1_ASAP7_75t_L g5010 ( 
.A(n_4317),
.Y(n_5010)
);

INVx1_ASAP7_75t_L g5011 ( 
.A(n_4317),
.Y(n_5011)
);

INVx6_ASAP7_75t_L g5012 ( 
.A(n_4161),
.Y(n_5012)
);

OAI21x1_ASAP7_75t_L g5013 ( 
.A1(n_4151),
.A2(n_3721),
.B(n_3714),
.Y(n_5013)
);

INVx1_ASAP7_75t_L g5014 ( 
.A(n_4321),
.Y(n_5014)
);

AOI22xp33_ASAP7_75t_L g5015 ( 
.A1(n_4479),
.A2(n_3994),
.B1(n_4027),
.B2(n_3697),
.Y(n_5015)
);

BUFx3_ASAP7_75t_L g5016 ( 
.A(n_4490),
.Y(n_5016)
);

INVx1_ASAP7_75t_L g5017 ( 
.A(n_4321),
.Y(n_5017)
);

INVx1_ASAP7_75t_L g5018 ( 
.A(n_4327),
.Y(n_5018)
);

AO21x2_ASAP7_75t_L g5019 ( 
.A1(n_4571),
.A2(n_4029),
.B(n_4019),
.Y(n_5019)
);

AOI22xp33_ASAP7_75t_SL g5020 ( 
.A1(n_4289),
.A2(n_3827),
.B1(n_3885),
.B2(n_3819),
.Y(n_5020)
);

AOI22xp5_ASAP7_75t_L g5021 ( 
.A1(n_4214),
.A2(n_3819),
.B1(n_3946),
.B2(n_3956),
.Y(n_5021)
);

INVx2_ASAP7_75t_SL g5022 ( 
.A(n_4500),
.Y(n_5022)
);

INVx2_ASAP7_75t_L g5023 ( 
.A(n_4351),
.Y(n_5023)
);

AND2x4_ASAP7_75t_L g5024 ( 
.A(n_4260),
.B(n_3680),
.Y(n_5024)
);

INVx1_ASAP7_75t_L g5025 ( 
.A(n_4327),
.Y(n_5025)
);

OR2x2_ASAP7_75t_L g5026 ( 
.A(n_4155),
.B(n_3956),
.Y(n_5026)
);

HB1xp67_ASAP7_75t_L g5027 ( 
.A(n_4578),
.Y(n_5027)
);

INVx2_ASAP7_75t_L g5028 ( 
.A(n_4351),
.Y(n_5028)
);

INVx1_ASAP7_75t_L g5029 ( 
.A(n_4328),
.Y(n_5029)
);

OAI21x1_ASAP7_75t_L g5030 ( 
.A1(n_4240),
.A2(n_3721),
.B(n_3714),
.Y(n_5030)
);

INVx2_ASAP7_75t_L g5031 ( 
.A(n_4351),
.Y(n_5031)
);

NAND2xp5_ASAP7_75t_L g5032 ( 
.A(n_4628),
.B(n_3895),
.Y(n_5032)
);

BUFx10_ASAP7_75t_L g5033 ( 
.A(n_4536),
.Y(n_5033)
);

INVx2_ASAP7_75t_L g5034 ( 
.A(n_4351),
.Y(n_5034)
);

AOI22xp33_ASAP7_75t_L g5035 ( 
.A1(n_4134),
.A2(n_4027),
.B1(n_3994),
.B2(n_3885),
.Y(n_5035)
);

AOI21x1_ASAP7_75t_L g5036 ( 
.A1(n_4190),
.A2(n_4116),
.B(n_4106),
.Y(n_5036)
);

BUFx6f_ASAP7_75t_L g5037 ( 
.A(n_4139),
.Y(n_5037)
);

NAND3xp33_ASAP7_75t_L g5038 ( 
.A(n_4134),
.B(n_3962),
.C(n_3992),
.Y(n_5038)
);

AOI22xp33_ASAP7_75t_L g5039 ( 
.A1(n_4324),
.A2(n_4027),
.B1(n_3994),
.B2(n_3885),
.Y(n_5039)
);

NAND2x1p5_ASAP7_75t_L g5040 ( 
.A(n_4395),
.B(n_3910),
.Y(n_5040)
);

INVx2_ASAP7_75t_L g5041 ( 
.A(n_4351),
.Y(n_5041)
);

BUFx2_ASAP7_75t_R g5042 ( 
.A(n_4216),
.Y(n_5042)
);

NAND2xp5_ASAP7_75t_L g5043 ( 
.A(n_4294),
.B(n_3896),
.Y(n_5043)
);

INVx4_ASAP7_75t_L g5044 ( 
.A(n_4490),
.Y(n_5044)
);

INVx1_ASAP7_75t_L g5045 ( 
.A(n_4328),
.Y(n_5045)
);

NAND2x1p5_ASAP7_75t_L g5046 ( 
.A(n_4460),
.B(n_3910),
.Y(n_5046)
);

OAI22xp33_ASAP7_75t_L g5047 ( 
.A1(n_4289),
.A2(n_3885),
.B1(n_3827),
.B2(n_3910),
.Y(n_5047)
);

INVx1_ASAP7_75t_L g5048 ( 
.A(n_4329),
.Y(n_5048)
);

INVx1_ASAP7_75t_SL g5049 ( 
.A(n_4209),
.Y(n_5049)
);

BUFx2_ASAP7_75t_L g5050 ( 
.A(n_4456),
.Y(n_5050)
);

INVx6_ASAP7_75t_L g5051 ( 
.A(n_4260),
.Y(n_5051)
);

INVx1_ASAP7_75t_L g5052 ( 
.A(n_4329),
.Y(n_5052)
);

INVx1_ASAP7_75t_L g5053 ( 
.A(n_4333),
.Y(n_5053)
);

INVx1_ASAP7_75t_L g5054 ( 
.A(n_4333),
.Y(n_5054)
);

INVx5_ASAP7_75t_L g5055 ( 
.A(n_4579),
.Y(n_5055)
);

INVx2_ASAP7_75t_L g5056 ( 
.A(n_4351),
.Y(n_5056)
);

INVx1_ASAP7_75t_L g5057 ( 
.A(n_4345),
.Y(n_5057)
);

AOI22xp33_ASAP7_75t_L g5058 ( 
.A1(n_4324),
.A2(n_3827),
.B1(n_3670),
.B2(n_3686),
.Y(n_5058)
);

OAI22xp33_ASAP7_75t_L g5059 ( 
.A1(n_4273),
.A2(n_3827),
.B1(n_3919),
.B2(n_4063),
.Y(n_5059)
);

BUFx2_ASAP7_75t_L g5060 ( 
.A(n_4504),
.Y(n_5060)
);

INVxp67_ASAP7_75t_L g5061 ( 
.A(n_4360),
.Y(n_5061)
);

AOI21x1_ASAP7_75t_L g5062 ( 
.A1(n_4190),
.A2(n_4391),
.B(n_4319),
.Y(n_5062)
);

CKINVDCx5p33_ASAP7_75t_R g5063 ( 
.A(n_4490),
.Y(n_5063)
);

OAI21x1_ASAP7_75t_L g5064 ( 
.A1(n_4240),
.A2(n_3769),
.B(n_3721),
.Y(n_5064)
);

INVx2_ASAP7_75t_L g5065 ( 
.A(n_4451),
.Y(n_5065)
);

INVx1_ASAP7_75t_L g5066 ( 
.A(n_4345),
.Y(n_5066)
);

HB1xp67_ASAP7_75t_L g5067 ( 
.A(n_4607),
.Y(n_5067)
);

NOR2xp33_ASAP7_75t_L g5068 ( 
.A(n_4192),
.B(n_3750),
.Y(n_5068)
);

AND2x2_ASAP7_75t_L g5069 ( 
.A(n_4208),
.B(n_4119),
.Y(n_5069)
);

AO21x2_ASAP7_75t_L g5070 ( 
.A1(n_4419),
.A2(n_4032),
.B(n_4029),
.Y(n_5070)
);

BUFx6f_ASAP7_75t_L g5071 ( 
.A(n_4287),
.Y(n_5071)
);

INVx2_ASAP7_75t_L g5072 ( 
.A(n_4451),
.Y(n_5072)
);

AO21x1_ASAP7_75t_SL g5073 ( 
.A1(n_4469),
.A2(n_3904),
.B(n_3896),
.Y(n_5073)
);

AO21x1_ASAP7_75t_L g5074 ( 
.A1(n_4330),
.A2(n_4009),
.B(n_3992),
.Y(n_5074)
);

INVx1_ASAP7_75t_L g5075 ( 
.A(n_4347),
.Y(n_5075)
);

AOI21x1_ASAP7_75t_L g5076 ( 
.A1(n_4319),
.A2(n_4116),
.B(n_4106),
.Y(n_5076)
);

INVx1_ASAP7_75t_L g5077 ( 
.A(n_4347),
.Y(n_5077)
);

AOI22xp33_ASAP7_75t_L g5078 ( 
.A1(n_4250),
.A2(n_3670),
.B1(n_3686),
.B2(n_3652),
.Y(n_5078)
);

AND2x2_ASAP7_75t_L g5079 ( 
.A(n_4208),
.B(n_4119),
.Y(n_5079)
);

INVx2_ASAP7_75t_L g5080 ( 
.A(n_4451),
.Y(n_5080)
);

BUFx3_ASAP7_75t_L g5081 ( 
.A(n_4216),
.Y(n_5081)
);

AND2x2_ASAP7_75t_L g5082 ( 
.A(n_4261),
.B(n_3913),
.Y(n_5082)
);

INVx1_ASAP7_75t_L g5083 ( 
.A(n_4348),
.Y(n_5083)
);

INVx4_ASAP7_75t_L g5084 ( 
.A(n_4277),
.Y(n_5084)
);

BUFx6f_ASAP7_75t_L g5085 ( 
.A(n_4287),
.Y(n_5085)
);

AOI21x1_ASAP7_75t_L g5086 ( 
.A1(n_4391),
.A2(n_3903),
.B(n_3897),
.Y(n_5086)
);

INVx1_ASAP7_75t_L g5087 ( 
.A(n_4348),
.Y(n_5087)
);

AOI22xp33_ASAP7_75t_L g5088 ( 
.A1(n_4250),
.A2(n_3670),
.B1(n_3686),
.B2(n_3652),
.Y(n_5088)
);

BUFx6f_ASAP7_75t_L g5089 ( 
.A(n_4287),
.Y(n_5089)
);

INVx5_ASAP7_75t_L g5090 ( 
.A(n_4579),
.Y(n_5090)
);

INVx2_ASAP7_75t_L g5091 ( 
.A(n_4451),
.Y(n_5091)
);

AOI22xp5_ASAP7_75t_SL g5092 ( 
.A1(n_4373),
.A2(n_3963),
.B1(n_3968),
.B2(n_3909),
.Y(n_5092)
);

INVx2_ASAP7_75t_L g5093 ( 
.A(n_4451),
.Y(n_5093)
);

HB1xp67_ASAP7_75t_L g5094 ( 
.A(n_4625),
.Y(n_5094)
);

INVx1_ASAP7_75t_L g5095 ( 
.A(n_4353),
.Y(n_5095)
);

INVx2_ASAP7_75t_L g5096 ( 
.A(n_4466),
.Y(n_5096)
);

INVx1_ASAP7_75t_SL g5097 ( 
.A(n_4209),
.Y(n_5097)
);

INVx2_ASAP7_75t_L g5098 ( 
.A(n_4466),
.Y(n_5098)
);

INVx2_ASAP7_75t_L g5099 ( 
.A(n_4466),
.Y(n_5099)
);

INVx1_ASAP7_75t_L g5100 ( 
.A(n_4353),
.Y(n_5100)
);

INVx1_ASAP7_75t_L g5101 ( 
.A(n_4355),
.Y(n_5101)
);

INVx3_ASAP7_75t_L g5102 ( 
.A(n_4491),
.Y(n_5102)
);

NAND2xp5_ASAP7_75t_L g5103 ( 
.A(n_4316),
.B(n_3904),
.Y(n_5103)
);

AOI22xp33_ASAP7_75t_L g5104 ( 
.A1(n_4298),
.A2(n_3670),
.B1(n_3686),
.B2(n_3652),
.Y(n_5104)
);

AOI22xp33_ASAP7_75t_SL g5105 ( 
.A1(n_4350),
.A2(n_4340),
.B1(n_4230),
.B2(n_4339),
.Y(n_5105)
);

BUFx2_ASAP7_75t_SL g5106 ( 
.A(n_4597),
.Y(n_5106)
);

AOI21x1_ASAP7_75t_L g5107 ( 
.A1(n_4583),
.A2(n_3903),
.B(n_3897),
.Y(n_5107)
);

CKINVDCx11_ASAP7_75t_R g5108 ( 
.A(n_4147),
.Y(n_5108)
);

INVx2_ASAP7_75t_SL g5109 ( 
.A(n_4504),
.Y(n_5109)
);

AOI21x1_ASAP7_75t_L g5110 ( 
.A1(n_4583),
.A2(n_3897),
.B(n_3980),
.Y(n_5110)
);

INVx2_ASAP7_75t_L g5111 ( 
.A(n_4466),
.Y(n_5111)
);

OA21x2_ASAP7_75t_L g5112 ( 
.A1(n_4246),
.A2(n_3972),
.B(n_4032),
.Y(n_5112)
);

BUFx6f_ASAP7_75t_L g5113 ( 
.A(n_4287),
.Y(n_5113)
);

INVx1_ASAP7_75t_SL g5114 ( 
.A(n_4253),
.Y(n_5114)
);

INVx2_ASAP7_75t_L g5115 ( 
.A(n_4466),
.Y(n_5115)
);

AOI22xp33_ASAP7_75t_L g5116 ( 
.A1(n_4268),
.A2(n_3670),
.B1(n_3686),
.B2(n_3652),
.Y(n_5116)
);

INVx1_ASAP7_75t_L g5117 ( 
.A(n_4355),
.Y(n_5117)
);

INVx1_ASAP7_75t_L g5118 ( 
.A(n_4357),
.Y(n_5118)
);

AOI22xp33_ASAP7_75t_L g5119 ( 
.A1(n_4326),
.A2(n_3818),
.B1(n_3652),
.B2(n_3893),
.Y(n_5119)
);

BUFx3_ASAP7_75t_L g5120 ( 
.A(n_4272),
.Y(n_5120)
);

AND2x4_ASAP7_75t_L g5121 ( 
.A(n_4260),
.B(n_3680),
.Y(n_5121)
);

BUFx3_ASAP7_75t_L g5122 ( 
.A(n_4272),
.Y(n_5122)
);

AOI21xp5_ASAP7_75t_SL g5123 ( 
.A1(n_4417),
.A2(n_3675),
.B(n_3766),
.Y(n_5123)
);

CKINVDCx11_ASAP7_75t_R g5124 ( 
.A(n_4147),
.Y(n_5124)
);

INVx2_ASAP7_75t_L g5125 ( 
.A(n_4594),
.Y(n_5125)
);

INVx4_ASAP7_75t_L g5126 ( 
.A(n_4277),
.Y(n_5126)
);

BUFx2_ASAP7_75t_L g5127 ( 
.A(n_4514),
.Y(n_5127)
);

CKINVDCx11_ASAP7_75t_R g5128 ( 
.A(n_4207),
.Y(n_5128)
);

INVx1_ASAP7_75t_L g5129 ( 
.A(n_4357),
.Y(n_5129)
);

AND2x4_ASAP7_75t_L g5130 ( 
.A(n_4260),
.B(n_3680),
.Y(n_5130)
);

CKINVDCx6p67_ASAP7_75t_R g5131 ( 
.A(n_4272),
.Y(n_5131)
);

AND2x2_ASAP7_75t_L g5132 ( 
.A(n_4261),
.B(n_4365),
.Y(n_5132)
);

AND2x2_ASAP7_75t_L g5133 ( 
.A(n_4365),
.B(n_3968),
.Y(n_5133)
);

BUFx3_ASAP7_75t_L g5134 ( 
.A(n_4342),
.Y(n_5134)
);

OAI22xp5_ASAP7_75t_L g5135 ( 
.A1(n_4339),
.A2(n_4230),
.B1(n_4142),
.B2(n_4162),
.Y(n_5135)
);

INVx4_ASAP7_75t_L g5136 ( 
.A(n_4277),
.Y(n_5136)
);

CKINVDCx20_ASAP7_75t_R g5137 ( 
.A(n_4367),
.Y(n_5137)
);

AND2x2_ASAP7_75t_L g5138 ( 
.A(n_4381),
.B(n_4387),
.Y(n_5138)
);

BUFx2_ASAP7_75t_SL g5139 ( 
.A(n_4597),
.Y(n_5139)
);

INVx1_ASAP7_75t_L g5140 ( 
.A(n_4359),
.Y(n_5140)
);

OAI21xp5_ASAP7_75t_L g5141 ( 
.A1(n_4199),
.A2(n_3957),
.B(n_3887),
.Y(n_5141)
);

AOI21x1_ASAP7_75t_L g5142 ( 
.A1(n_4143),
.A2(n_3986),
.B(n_3980),
.Y(n_5142)
);

AND2x2_ASAP7_75t_L g5143 ( 
.A(n_4381),
.B(n_3976),
.Y(n_5143)
);

INVx1_ASAP7_75t_L g5144 ( 
.A(n_4359),
.Y(n_5144)
);

INVx4_ASAP7_75t_L g5145 ( 
.A(n_4342),
.Y(n_5145)
);

INVx3_ASAP7_75t_L g5146 ( 
.A(n_4491),
.Y(n_5146)
);

INVxp67_ASAP7_75t_L g5147 ( 
.A(n_4310),
.Y(n_5147)
);

INVx1_ASAP7_75t_L g5148 ( 
.A(n_4361),
.Y(n_5148)
);

HB1xp67_ASAP7_75t_SL g5149 ( 
.A(n_4342),
.Y(n_5149)
);

NOR2xp33_ASAP7_75t_L g5150 ( 
.A(n_4206),
.B(n_3750),
.Y(n_5150)
);

BUFx6f_ASAP7_75t_SL g5151 ( 
.A(n_4392),
.Y(n_5151)
);

INVx2_ASAP7_75t_L g5152 ( 
.A(n_4594),
.Y(n_5152)
);

AOI21x1_ASAP7_75t_L g5153 ( 
.A1(n_4143),
.A2(n_4130),
.B(n_4570),
.Y(n_5153)
);

BUFx2_ASAP7_75t_R g5154 ( 
.A(n_4392),
.Y(n_5154)
);

INVx2_ASAP7_75t_L g5155 ( 
.A(n_4594),
.Y(n_5155)
);

AOI21x1_ASAP7_75t_L g5156 ( 
.A1(n_4130),
.A2(n_3986),
.B(n_3685),
.Y(n_5156)
);

BUFx2_ASAP7_75t_SL g5157 ( 
.A(n_4597),
.Y(n_5157)
);

HB1xp67_ASAP7_75t_L g5158 ( 
.A(n_4631),
.Y(n_5158)
);

INVx3_ASAP7_75t_L g5159 ( 
.A(n_4491),
.Y(n_5159)
);

HB1xp67_ASAP7_75t_L g5160 ( 
.A(n_4635),
.Y(n_5160)
);

INVx1_ASAP7_75t_L g5161 ( 
.A(n_4361),
.Y(n_5161)
);

INVx1_ASAP7_75t_L g5162 ( 
.A(n_4369),
.Y(n_5162)
);

INVx6_ASAP7_75t_L g5163 ( 
.A(n_4260),
.Y(n_5163)
);

BUFx3_ASAP7_75t_L g5164 ( 
.A(n_4392),
.Y(n_5164)
);

HB1xp67_ASAP7_75t_L g5165 ( 
.A(n_4657),
.Y(n_5165)
);

INVx1_ASAP7_75t_L g5166 ( 
.A(n_4369),
.Y(n_5166)
);

INVx2_ASAP7_75t_L g5167 ( 
.A(n_4594),
.Y(n_5167)
);

AND2x2_ASAP7_75t_L g5168 ( 
.A(n_4387),
.B(n_3976),
.Y(n_5168)
);

INVx1_ASAP7_75t_SL g5169 ( 
.A(n_4253),
.Y(n_5169)
);

INVx2_ASAP7_75t_L g5170 ( 
.A(n_4594),
.Y(n_5170)
);

INVx2_ASAP7_75t_L g5171 ( 
.A(n_4534),
.Y(n_5171)
);

OAI22xp5_ASAP7_75t_L g5172 ( 
.A1(n_4142),
.A2(n_4377),
.B1(n_4248),
.B2(n_4157),
.Y(n_5172)
);

INVx1_ASAP7_75t_L g5173 ( 
.A(n_4372),
.Y(n_5173)
);

HB1xp67_ASAP7_75t_L g5174 ( 
.A(n_4662),
.Y(n_5174)
);

BUFx2_ASAP7_75t_SL g5175 ( 
.A(n_4207),
.Y(n_5175)
);

OAI22xp33_ASAP7_75t_L g5176 ( 
.A1(n_4340),
.A2(n_3919),
.B1(n_4064),
.B2(n_4063),
.Y(n_5176)
);

INVx1_ASAP7_75t_L g5177 ( 
.A(n_4372),
.Y(n_5177)
);

INVx1_ASAP7_75t_L g5178 ( 
.A(n_4375),
.Y(n_5178)
);

INVx1_ASAP7_75t_L g5179 ( 
.A(n_4375),
.Y(n_5179)
);

INVx6_ASAP7_75t_L g5180 ( 
.A(n_4577),
.Y(n_5180)
);

BUFx2_ASAP7_75t_R g5181 ( 
.A(n_4415),
.Y(n_5181)
);

INVx2_ASAP7_75t_L g5182 ( 
.A(n_4534),
.Y(n_5182)
);

NOR2xp33_ASAP7_75t_L g5183 ( 
.A(n_4210),
.B(n_3798),
.Y(n_5183)
);

INVx2_ASAP7_75t_L g5184 ( 
.A(n_4534),
.Y(n_5184)
);

BUFx2_ASAP7_75t_R g5185 ( 
.A(n_4415),
.Y(n_5185)
);

INVx1_ASAP7_75t_L g5186 ( 
.A(n_4376),
.Y(n_5186)
);

AOI22xp33_ASAP7_75t_L g5187 ( 
.A1(n_4364),
.A2(n_3818),
.B1(n_3893),
.B2(n_3803),
.Y(n_5187)
);

INVx2_ASAP7_75t_L g5188 ( 
.A(n_4553),
.Y(n_5188)
);

NAND2xp5_ASAP7_75t_L g5189 ( 
.A(n_4316),
.B(n_3912),
.Y(n_5189)
);

AOI22xp33_ASAP7_75t_SL g5190 ( 
.A1(n_4350),
.A2(n_3807),
.B1(n_3834),
.B2(n_3988),
.Y(n_5190)
);

AND2x2_ASAP7_75t_L g5191 ( 
.A(n_4136),
.B(n_3976),
.Y(n_5191)
);

OAI22xp5_ASAP7_75t_L g5192 ( 
.A1(n_4377),
.A2(n_4011),
.B1(n_3983),
.B2(n_3889),
.Y(n_5192)
);

CKINVDCx5p33_ASAP7_75t_R g5193 ( 
.A(n_4415),
.Y(n_5193)
);

BUFx2_ASAP7_75t_SL g5194 ( 
.A(n_4429),
.Y(n_5194)
);

OAI22xp33_ASAP7_75t_R g5195 ( 
.A1(n_4213),
.A2(n_3977),
.B1(n_3866),
.B2(n_3954),
.Y(n_5195)
);

INVx1_ASAP7_75t_L g5196 ( 
.A(n_4376),
.Y(n_5196)
);

INVx1_ASAP7_75t_L g5197 ( 
.A(n_4379),
.Y(n_5197)
);

INVx2_ASAP7_75t_SL g5198 ( 
.A(n_4514),
.Y(n_5198)
);

INVx2_ASAP7_75t_SL g5199 ( 
.A(n_4522),
.Y(n_5199)
);

NOR2xp33_ASAP7_75t_L g5200 ( 
.A(n_4478),
.B(n_4499),
.Y(n_5200)
);

AND2x4_ASAP7_75t_L g5201 ( 
.A(n_4158),
.B(n_3726),
.Y(n_5201)
);

AOI22xp33_ASAP7_75t_L g5202 ( 
.A1(n_4352),
.A2(n_3818),
.B1(n_3893),
.B2(n_3803),
.Y(n_5202)
);

BUFx3_ASAP7_75t_L g5203 ( 
.A(n_4429),
.Y(n_5203)
);

BUFx6f_ASAP7_75t_L g5204 ( 
.A(n_4287),
.Y(n_5204)
);

CKINVDCx14_ASAP7_75t_R g5205 ( 
.A(n_4605),
.Y(n_5205)
);

INVx1_ASAP7_75t_L g5206 ( 
.A(n_4379),
.Y(n_5206)
);

INVx2_ASAP7_75t_L g5207 ( 
.A(n_4553),
.Y(n_5207)
);

NAND2x1p5_ASAP7_75t_L g5208 ( 
.A(n_4460),
.B(n_4063),
.Y(n_5208)
);

INVx2_ASAP7_75t_L g5209 ( 
.A(n_4553),
.Y(n_5209)
);

AOI22xp33_ASAP7_75t_L g5210 ( 
.A1(n_4356),
.A2(n_3818),
.B1(n_3893),
.B2(n_3803),
.Y(n_5210)
);

INVx1_ASAP7_75t_SL g5211 ( 
.A(n_4258),
.Y(n_5211)
);

INVx1_ASAP7_75t_L g5212 ( 
.A(n_4380),
.Y(n_5212)
);

AOI22xp33_ASAP7_75t_L g5213 ( 
.A1(n_4384),
.A2(n_3818),
.B1(n_3893),
.B2(n_3803),
.Y(n_5213)
);

INVx3_ASAP7_75t_L g5214 ( 
.A(n_4541),
.Y(n_5214)
);

INVx1_ASAP7_75t_L g5215 ( 
.A(n_4380),
.Y(n_5215)
);

INVx2_ASAP7_75t_L g5216 ( 
.A(n_4557),
.Y(n_5216)
);

BUFx3_ASAP7_75t_L g5217 ( 
.A(n_4429),
.Y(n_5217)
);

INVx2_ASAP7_75t_L g5218 ( 
.A(n_4557),
.Y(n_5218)
);

INVx1_ASAP7_75t_L g5219 ( 
.A(n_4398),
.Y(n_5219)
);

INVx1_ASAP7_75t_L g5220 ( 
.A(n_4398),
.Y(n_5220)
);

BUFx6f_ASAP7_75t_L g5221 ( 
.A(n_4287),
.Y(n_5221)
);

INVx1_ASAP7_75t_L g5222 ( 
.A(n_4408),
.Y(n_5222)
);

INVx2_ASAP7_75t_L g5223 ( 
.A(n_4557),
.Y(n_5223)
);

BUFx10_ASAP7_75t_L g5224 ( 
.A(n_4371),
.Y(n_5224)
);

BUFx6f_ASAP7_75t_L g5225 ( 
.A(n_4402),
.Y(n_5225)
);

INVx1_ASAP7_75t_L g5226 ( 
.A(n_4408),
.Y(n_5226)
);

INVx1_ASAP7_75t_L g5227 ( 
.A(n_4416),
.Y(n_5227)
);

BUFx10_ASAP7_75t_L g5228 ( 
.A(n_4371),
.Y(n_5228)
);

INVx11_ASAP7_75t_L g5229 ( 
.A(n_4443),
.Y(n_5229)
);

INVx1_ASAP7_75t_L g5230 ( 
.A(n_4416),
.Y(n_5230)
);

HB1xp67_ASAP7_75t_L g5231 ( 
.A(n_4439),
.Y(n_5231)
);

INVx2_ASAP7_75t_L g5232 ( 
.A(n_4560),
.Y(n_5232)
);

AOI22xp5_ASAP7_75t_L g5233 ( 
.A1(n_4403),
.A2(n_4010),
.B1(n_4023),
.B2(n_4009),
.Y(n_5233)
);

INVx1_ASAP7_75t_L g5234 ( 
.A(n_4447),
.Y(n_5234)
);

HB1xp67_ASAP7_75t_L g5235 ( 
.A(n_4472),
.Y(n_5235)
);

INVx1_ASAP7_75t_L g5236 ( 
.A(n_4447),
.Y(n_5236)
);

NAND2x1p5_ASAP7_75t_L g5237 ( 
.A(n_4614),
.B(n_4063),
.Y(n_5237)
);

AND2x4_ASAP7_75t_L g5238 ( 
.A(n_4158),
.B(n_4193),
.Y(n_5238)
);

BUFx12f_ASAP7_75t_L g5239 ( 
.A(n_4443),
.Y(n_5239)
);

AOI22xp33_ASAP7_75t_L g5240 ( 
.A1(n_4388),
.A2(n_4104),
.B1(n_4102),
.B2(n_4066),
.Y(n_5240)
);

AOI22xp33_ASAP7_75t_SL g5241 ( 
.A1(n_4305),
.A2(n_3807),
.B1(n_3834),
.B2(n_3988),
.Y(n_5241)
);

AOI22xp33_ASAP7_75t_SL g5242 ( 
.A1(n_4435),
.A2(n_3988),
.B1(n_3999),
.B2(n_3766),
.Y(n_5242)
);

NAND2xp5_ASAP7_75t_L g5243 ( 
.A(n_4527),
.B(n_3912),
.Y(n_5243)
);

AND2x2_ASAP7_75t_L g5244 ( 
.A(n_4136),
.B(n_3983),
.Y(n_5244)
);

AOI222xp33_ASAP7_75t_L g5245 ( 
.A1(n_4176),
.A2(n_4010),
.B1(n_4125),
.B2(n_4023),
.C1(n_4043),
.C2(n_4112),
.Y(n_5245)
);

BUFx2_ASAP7_75t_L g5246 ( 
.A(n_4522),
.Y(n_5246)
);

AOI21x1_ASAP7_75t_L g5247 ( 
.A1(n_4570),
.A2(n_4426),
.B(n_4555),
.Y(n_5247)
);

HB1xp67_ASAP7_75t_L g5248 ( 
.A(n_4155),
.Y(n_5248)
);

OAI22xp33_ASAP7_75t_L g5249 ( 
.A1(n_4435),
.A2(n_4064),
.B1(n_4063),
.B2(n_3967),
.Y(n_5249)
);

AOI22xp33_ASAP7_75t_L g5250 ( 
.A1(n_4471),
.A2(n_4104),
.B1(n_4102),
.B2(n_4066),
.Y(n_5250)
);

BUFx6f_ASAP7_75t_L g5251 ( 
.A(n_4402),
.Y(n_5251)
);

AO21x2_ASAP7_75t_L g5252 ( 
.A1(n_4419),
.A2(n_4067),
.B(n_4061),
.Y(n_5252)
);

INVx1_ASAP7_75t_L g5253 ( 
.A(n_4449),
.Y(n_5253)
);

AO21x2_ASAP7_75t_L g5254 ( 
.A1(n_4397),
.A2(n_4070),
.B(n_4067),
.Y(n_5254)
);

AOI22xp33_ASAP7_75t_L g5255 ( 
.A1(n_4471),
.A2(n_4066),
.B1(n_4085),
.B2(n_4069),
.Y(n_5255)
);

BUFx3_ASAP7_75t_L g5256 ( 
.A(n_4443),
.Y(n_5256)
);

HB1xp67_ASAP7_75t_L g5257 ( 
.A(n_4212),
.Y(n_5257)
);

INVx1_ASAP7_75t_SL g5258 ( 
.A(n_4258),
.Y(n_5258)
);

INVx2_ASAP7_75t_L g5259 ( 
.A(n_4560),
.Y(n_5259)
);

INVxp67_ASAP7_75t_SL g5260 ( 
.A(n_4404),
.Y(n_5260)
);

INVx2_ASAP7_75t_L g5261 ( 
.A(n_4560),
.Y(n_5261)
);

INVx2_ASAP7_75t_L g5262 ( 
.A(n_4564),
.Y(n_5262)
);

BUFx2_ASAP7_75t_SL g5263 ( 
.A(n_4507),
.Y(n_5263)
);

INVx1_ASAP7_75t_L g5264 ( 
.A(n_4449),
.Y(n_5264)
);

AOI22xp33_ASAP7_75t_L g5265 ( 
.A1(n_4410),
.A2(n_4069),
.B1(n_4091),
.B2(n_4085),
.Y(n_5265)
);

HB1xp67_ASAP7_75t_L g5266 ( 
.A(n_4295),
.Y(n_5266)
);

AOI22xp33_ASAP7_75t_L g5267 ( 
.A1(n_4410),
.A2(n_4069),
.B1(n_4091),
.B2(n_4085),
.Y(n_5267)
);

CKINVDCx20_ASAP7_75t_R g5268 ( 
.A(n_4517),
.Y(n_5268)
);

CKINVDCx11_ASAP7_75t_R g5269 ( 
.A(n_4259),
.Y(n_5269)
);

INVx1_ASAP7_75t_L g5270 ( 
.A(n_4450),
.Y(n_5270)
);

INVx1_ASAP7_75t_SL g5271 ( 
.A(n_4259),
.Y(n_5271)
);

AOI22xp33_ASAP7_75t_SL g5272 ( 
.A1(n_4305),
.A2(n_3999),
.B1(n_3766),
.B2(n_3842),
.Y(n_5272)
);

INVx2_ASAP7_75t_SL g5273 ( 
.A(n_4641),
.Y(n_5273)
);

BUFx12f_ASAP7_75t_L g5274 ( 
.A(n_4577),
.Y(n_5274)
);

AOI22xp33_ASAP7_75t_L g5275 ( 
.A1(n_4399),
.A2(n_4091),
.B1(n_4096),
.B2(n_4093),
.Y(n_5275)
);

AOI22xp33_ASAP7_75t_L g5276 ( 
.A1(n_4399),
.A2(n_4401),
.B1(n_4566),
.B2(n_4561),
.Y(n_5276)
);

INVx1_ASAP7_75t_L g5277 ( 
.A(n_4450),
.Y(n_5277)
);

INVx1_ASAP7_75t_L g5278 ( 
.A(n_4454),
.Y(n_5278)
);

CKINVDCx5p33_ASAP7_75t_R g5279 ( 
.A(n_4308),
.Y(n_5279)
);

INVx2_ASAP7_75t_L g5280 ( 
.A(n_4564),
.Y(n_5280)
);

INVx1_ASAP7_75t_L g5281 ( 
.A(n_4454),
.Y(n_5281)
);

INVx1_ASAP7_75t_L g5282 ( 
.A(n_4492),
.Y(n_5282)
);

AND2x2_ASAP7_75t_L g5283 ( 
.A(n_4159),
.B(n_3983),
.Y(n_5283)
);

INVx1_ASAP7_75t_L g5284 ( 
.A(n_4492),
.Y(n_5284)
);

NAND2xp5_ASAP7_75t_L g5285 ( 
.A(n_4527),
.B(n_3915),
.Y(n_5285)
);

BUFx5_ASAP7_75t_L g5286 ( 
.A(n_4579),
.Y(n_5286)
);

AOI22xp33_ASAP7_75t_L g5287 ( 
.A1(n_4399),
.A2(n_4093),
.B1(n_4097),
.B2(n_4096),
.Y(n_5287)
);

BUFx2_ASAP7_75t_R g5288 ( 
.A(n_4238),
.Y(n_5288)
);

INVx6_ASAP7_75t_L g5289 ( 
.A(n_4577),
.Y(n_5289)
);

INVx2_ASAP7_75t_L g5290 ( 
.A(n_4564),
.Y(n_5290)
);

AOI22xp33_ASAP7_75t_L g5291 ( 
.A1(n_4399),
.A2(n_4093),
.B1(n_4097),
.B2(n_4096),
.Y(n_5291)
);

CKINVDCx16_ASAP7_75t_R g5292 ( 
.A(n_4533),
.Y(n_5292)
);

AND2x2_ASAP7_75t_L g5293 ( 
.A(n_4159),
.B(n_4011),
.Y(n_5293)
);

AOI22xp33_ASAP7_75t_SL g5294 ( 
.A1(n_4374),
.A2(n_3999),
.B1(n_3766),
.B2(n_3842),
.Y(n_5294)
);

AOI22xp33_ASAP7_75t_L g5295 ( 
.A1(n_4399),
.A2(n_4401),
.B1(n_4566),
.B2(n_4561),
.Y(n_5295)
);

INVx1_ASAP7_75t_L g5296 ( 
.A(n_4493),
.Y(n_5296)
);

AND2x2_ASAP7_75t_L g5297 ( 
.A(n_4171),
.B(n_4011),
.Y(n_5297)
);

INVx1_ASAP7_75t_L g5298 ( 
.A(n_4493),
.Y(n_5298)
);

INVx2_ASAP7_75t_L g5299 ( 
.A(n_4568),
.Y(n_5299)
);

INVx3_ASAP7_75t_L g5300 ( 
.A(n_4541),
.Y(n_5300)
);

HB1xp67_ASAP7_75t_L g5301 ( 
.A(n_4358),
.Y(n_5301)
);

INVxp67_ASAP7_75t_SL g5302 ( 
.A(n_4404),
.Y(n_5302)
);

AND2x2_ASAP7_75t_L g5303 ( 
.A(n_4171),
.B(n_4120),
.Y(n_5303)
);

AOI22xp33_ASAP7_75t_L g5304 ( 
.A1(n_4399),
.A2(n_4122),
.B1(n_4124),
.B2(n_4097),
.Y(n_5304)
);

INVx1_ASAP7_75t_L g5305 ( 
.A(n_4496),
.Y(n_5305)
);

INVx1_ASAP7_75t_L g5306 ( 
.A(n_4496),
.Y(n_5306)
);

NAND2x1p5_ASAP7_75t_L g5307 ( 
.A(n_4614),
.B(n_4063),
.Y(n_5307)
);

OR2x6_ASAP7_75t_L g5308 ( 
.A(n_4160),
.B(n_4056),
.Y(n_5308)
);

INVx1_ASAP7_75t_L g5309 ( 
.A(n_4498),
.Y(n_5309)
);

AOI22xp33_ASAP7_75t_L g5310 ( 
.A1(n_4401),
.A2(n_4529),
.B1(n_4511),
.B2(n_4605),
.Y(n_5310)
);

OAI22xp33_ASAP7_75t_L g5311 ( 
.A1(n_4373),
.A2(n_4064),
.B1(n_4063),
.B2(n_3967),
.Y(n_5311)
);

NAND2x1p5_ASAP7_75t_L g5312 ( 
.A(n_4645),
.B(n_4064),
.Y(n_5312)
);

BUFx12f_ASAP7_75t_L g5313 ( 
.A(n_4577),
.Y(n_5313)
);

INVx2_ASAP7_75t_L g5314 ( 
.A(n_4568),
.Y(n_5314)
);

BUFx3_ASAP7_75t_L g5315 ( 
.A(n_4530),
.Y(n_5315)
);

AND2x2_ASAP7_75t_L g5316 ( 
.A(n_4179),
.B(n_4120),
.Y(n_5316)
);

AOI22xp33_ASAP7_75t_L g5317 ( 
.A1(n_4401),
.A2(n_4124),
.B1(n_4122),
.B2(n_3967),
.Y(n_5317)
);

INVx1_ASAP7_75t_L g5318 ( 
.A(n_4498),
.Y(n_5318)
);

INVx4_ASAP7_75t_L g5319 ( 
.A(n_4182),
.Y(n_5319)
);

INVx1_ASAP7_75t_L g5320 ( 
.A(n_4510),
.Y(n_5320)
);

HB1xp67_ASAP7_75t_L g5321 ( 
.A(n_4608),
.Y(n_5321)
);

BUFx2_ASAP7_75t_R g5322 ( 
.A(n_4238),
.Y(n_5322)
);

HB1xp67_ASAP7_75t_L g5323 ( 
.A(n_4580),
.Y(n_5323)
);

HB1xp67_ASAP7_75t_L g5324 ( 
.A(n_4580),
.Y(n_5324)
);

AO21x2_ASAP7_75t_L g5325 ( 
.A1(n_4397),
.A2(n_4126),
.B(n_4081),
.Y(n_5325)
);

INVx1_ASAP7_75t_L g5326 ( 
.A(n_4510),
.Y(n_5326)
);

INVx1_ASAP7_75t_L g5327 ( 
.A(n_4518),
.Y(n_5327)
);

OR2x2_ASAP7_75t_L g5328 ( 
.A(n_4363),
.B(n_4043),
.Y(n_5328)
);

AOI22xp33_ASAP7_75t_L g5329 ( 
.A1(n_4401),
.A2(n_4122),
.B1(n_4124),
.B2(n_3942),
.Y(n_5329)
);

AOI22xp5_ASAP7_75t_L g5330 ( 
.A1(n_4141),
.A2(n_4072),
.B1(n_4076),
.B2(n_4048),
.Y(n_5330)
);

INVx2_ASAP7_75t_L g5331 ( 
.A(n_4512),
.Y(n_5331)
);

OAI22xp5_ASAP7_75t_L g5332 ( 
.A1(n_4157),
.A2(n_3889),
.B1(n_3800),
.B2(n_3957),
.Y(n_5332)
);

BUFx2_ASAP7_75t_R g5333 ( 
.A(n_4420),
.Y(n_5333)
);

INVx1_ASAP7_75t_L g5334 ( 
.A(n_4518),
.Y(n_5334)
);

AOI21xp5_ASAP7_75t_L g5335 ( 
.A1(n_4150),
.A2(n_4051),
.B(n_3957),
.Y(n_5335)
);

INVx1_ASAP7_75t_L g5336 ( 
.A(n_4547),
.Y(n_5336)
);

INVx1_ASAP7_75t_L g5337 ( 
.A(n_4547),
.Y(n_5337)
);

AOI22xp33_ASAP7_75t_L g5338 ( 
.A1(n_4401),
.A2(n_3942),
.B1(n_3937),
.B2(n_3926),
.Y(n_5338)
);

INVx2_ASAP7_75t_L g5339 ( 
.A(n_4512),
.Y(n_5339)
);

INVx2_ASAP7_75t_L g5340 ( 
.A(n_4512),
.Y(n_5340)
);

AOI22xp33_ASAP7_75t_L g5341 ( 
.A1(n_4511),
.A2(n_4529),
.B1(n_4382),
.B2(n_4546),
.Y(n_5341)
);

BUFx12f_ASAP7_75t_L g5342 ( 
.A(n_4182),
.Y(n_5342)
);

INVx1_ASAP7_75t_L g5343 ( 
.A(n_4562),
.Y(n_5343)
);

INVx1_ASAP7_75t_L g5344 ( 
.A(n_4562),
.Y(n_5344)
);

AOI22xp33_ASAP7_75t_L g5345 ( 
.A1(n_4511),
.A2(n_3942),
.B1(n_3937),
.B2(n_3926),
.Y(n_5345)
);

AOI22xp33_ASAP7_75t_L g5346 ( 
.A1(n_4511),
.A2(n_3937),
.B1(n_3989),
.B2(n_3926),
.Y(n_5346)
);

INVx3_ASAP7_75t_SL g5347 ( 
.A(n_4371),
.Y(n_5347)
);

INVx2_ASAP7_75t_L g5348 ( 
.A(n_4512),
.Y(n_5348)
);

AOI22xp33_ASAP7_75t_SL g5349 ( 
.A1(n_4374),
.A2(n_3842),
.B1(n_4114),
.B2(n_4056),
.Y(n_5349)
);

INVx2_ASAP7_75t_L g5350 ( 
.A(n_4389),
.Y(n_5350)
);

INVx3_ASAP7_75t_L g5351 ( 
.A(n_4541),
.Y(n_5351)
);

AO21x1_ASAP7_75t_L g5352 ( 
.A1(n_4169),
.A2(n_4072),
.B(n_4048),
.Y(n_5352)
);

AOI22xp33_ASAP7_75t_SL g5353 ( 
.A1(n_4596),
.A2(n_3937),
.B1(n_3989),
.B2(n_3926),
.Y(n_5353)
);

CKINVDCx6p67_ASAP7_75t_R g5354 ( 
.A(n_4276),
.Y(n_5354)
);

INVx1_ASAP7_75t_L g5355 ( 
.A(n_4563),
.Y(n_5355)
);

INVx2_ASAP7_75t_L g5356 ( 
.A(n_4389),
.Y(n_5356)
);

INVx1_ASAP7_75t_L g5357 ( 
.A(n_4563),
.Y(n_5357)
);

BUFx2_ASAP7_75t_L g5358 ( 
.A(n_4641),
.Y(n_5358)
);

AO21x1_ASAP7_75t_L g5359 ( 
.A1(n_4169),
.A2(n_4086),
.B(n_4076),
.Y(n_5359)
);

AOI21xp33_ASAP7_75t_SL g5360 ( 
.A1(n_4281),
.A2(n_4468),
.B(n_4174),
.Y(n_5360)
);

AOI22xp33_ASAP7_75t_L g5361 ( 
.A1(n_4529),
.A2(n_3937),
.B1(n_3989),
.B2(n_3926),
.Y(n_5361)
);

INVx1_ASAP7_75t_SL g5362 ( 
.A(n_4276),
.Y(n_5362)
);

INVx2_ASAP7_75t_L g5363 ( 
.A(n_4389),
.Y(n_5363)
);

INVx2_ASAP7_75t_SL g5364 ( 
.A(n_4643),
.Y(n_5364)
);

INVx1_ASAP7_75t_L g5365 ( 
.A(n_4572),
.Y(n_5365)
);

INVx2_ASAP7_75t_L g5366 ( 
.A(n_4389),
.Y(n_5366)
);

INVx1_ASAP7_75t_L g5367 ( 
.A(n_4572),
.Y(n_5367)
);

AND2x2_ASAP7_75t_L g5368 ( 
.A(n_4679),
.B(n_4179),
.Y(n_5368)
);

AO21x1_ASAP7_75t_SL g5369 ( 
.A1(n_4791),
.A2(n_4349),
.B(n_4440),
.Y(n_5369)
);

INVx2_ASAP7_75t_L g5370 ( 
.A(n_5350),
.Y(n_5370)
);

HB1xp67_ASAP7_75t_L g5371 ( 
.A(n_4682),
.Y(n_5371)
);

INVx1_ASAP7_75t_L g5372 ( 
.A(n_4704),
.Y(n_5372)
);

INVx1_ASAP7_75t_L g5373 ( 
.A(n_4704),
.Y(n_5373)
);

NAND2xp5_ASAP7_75t_L g5374 ( 
.A(n_5074),
.B(n_4464),
.Y(n_5374)
);

INVx1_ASAP7_75t_L g5375 ( 
.A(n_4710),
.Y(n_5375)
);

AO21x2_ASAP7_75t_L g5376 ( 
.A1(n_4766),
.A2(n_4582),
.B(n_4341),
.Y(n_5376)
);

INVx1_ASAP7_75t_SL g5377 ( 
.A(n_4685),
.Y(n_5377)
);

INVx1_ASAP7_75t_L g5378 ( 
.A(n_4710),
.Y(n_5378)
);

NOR2xp33_ASAP7_75t_L g5379 ( 
.A(n_4773),
.B(n_4478),
.Y(n_5379)
);

INVx2_ASAP7_75t_L g5380 ( 
.A(n_5350),
.Y(n_5380)
);

INVx2_ASAP7_75t_SL g5381 ( 
.A(n_4675),
.Y(n_5381)
);

INVx2_ASAP7_75t_L g5382 ( 
.A(n_5350),
.Y(n_5382)
);

INVx1_ASAP7_75t_L g5383 ( 
.A(n_4719),
.Y(n_5383)
);

INVx1_ASAP7_75t_L g5384 ( 
.A(n_4719),
.Y(n_5384)
);

BUFx6f_ASAP7_75t_L g5385 ( 
.A(n_4713),
.Y(n_5385)
);

INVx2_ASAP7_75t_L g5386 ( 
.A(n_5356),
.Y(n_5386)
);

INVx5_ASAP7_75t_L g5387 ( 
.A(n_4675),
.Y(n_5387)
);

OR2x2_ASAP7_75t_L g5388 ( 
.A(n_5001),
.B(n_4195),
.Y(n_5388)
);

INVx2_ASAP7_75t_L g5389 ( 
.A(n_5356),
.Y(n_5389)
);

INVx4_ASAP7_75t_L g5390 ( 
.A(n_4680),
.Y(n_5390)
);

INVx1_ASAP7_75t_L g5391 ( 
.A(n_4727),
.Y(n_5391)
);

AND2x2_ASAP7_75t_L g5392 ( 
.A(n_4679),
.B(n_4612),
.Y(n_5392)
);

NAND2xp5_ASAP7_75t_L g5393 ( 
.A(n_5074),
.B(n_4464),
.Y(n_5393)
);

AND2x2_ASAP7_75t_L g5394 ( 
.A(n_4693),
.B(n_4612),
.Y(n_5394)
);

CKINVDCx5p33_ASAP7_75t_R g5395 ( 
.A(n_4670),
.Y(n_5395)
);

INVx1_ASAP7_75t_L g5396 ( 
.A(n_4727),
.Y(n_5396)
);

AND2x2_ASAP7_75t_L g5397 ( 
.A(n_4693),
.B(n_4630),
.Y(n_5397)
);

CKINVDCx5p33_ASAP7_75t_R g5398 ( 
.A(n_4747),
.Y(n_5398)
);

INVx2_ASAP7_75t_L g5399 ( 
.A(n_5356),
.Y(n_5399)
);

OR2x2_ASAP7_75t_L g5400 ( 
.A(n_5001),
.B(n_4195),
.Y(n_5400)
);

NOR2xp33_ASAP7_75t_L g5401 ( 
.A(n_4773),
.B(n_4732),
.Y(n_5401)
);

HB1xp67_ASAP7_75t_L g5402 ( 
.A(n_4695),
.Y(n_5402)
);

BUFx6f_ASAP7_75t_L g5403 ( 
.A(n_4732),
.Y(n_5403)
);

AND2x2_ASAP7_75t_L g5404 ( 
.A(n_4718),
.B(n_4630),
.Y(n_5404)
);

HB1xp67_ASAP7_75t_L g5405 ( 
.A(n_4709),
.Y(n_5405)
);

INVx2_ASAP7_75t_L g5406 ( 
.A(n_5363),
.Y(n_5406)
);

INVx2_ASAP7_75t_SL g5407 ( 
.A(n_4675),
.Y(n_5407)
);

BUFx2_ASAP7_75t_L g5408 ( 
.A(n_5315),
.Y(n_5408)
);

INVx2_ASAP7_75t_L g5409 ( 
.A(n_5363),
.Y(n_5409)
);

INVx2_ASAP7_75t_L g5410 ( 
.A(n_5363),
.Y(n_5410)
);

INVx1_ASAP7_75t_L g5411 ( 
.A(n_4730),
.Y(n_5411)
);

INVx3_ASAP7_75t_L g5412 ( 
.A(n_4715),
.Y(n_5412)
);

INVx2_ASAP7_75t_L g5413 ( 
.A(n_5366),
.Y(n_5413)
);

INVx2_ASAP7_75t_SL g5414 ( 
.A(n_4675),
.Y(n_5414)
);

AND2x2_ASAP7_75t_L g5415 ( 
.A(n_4718),
.B(n_4642),
.Y(n_5415)
);

AOI21xp5_ASAP7_75t_L g5416 ( 
.A1(n_4766),
.A2(n_5172),
.B(n_4991),
.Y(n_5416)
);

INVx1_ASAP7_75t_L g5417 ( 
.A(n_4730),
.Y(n_5417)
);

AOI21x1_ASAP7_75t_L g5418 ( 
.A1(n_5062),
.A2(n_4555),
.B(n_4426),
.Y(n_5418)
);

INVx1_ASAP7_75t_L g5419 ( 
.A(n_4739),
.Y(n_5419)
);

INVx2_ASAP7_75t_L g5420 ( 
.A(n_5366),
.Y(n_5420)
);

INVx1_ASAP7_75t_L g5421 ( 
.A(n_4739),
.Y(n_5421)
);

OA21x2_ASAP7_75t_L g5422 ( 
.A1(n_5260),
.A2(n_4600),
.B(n_4599),
.Y(n_5422)
);

INVx1_ASAP7_75t_L g5423 ( 
.A(n_4758),
.Y(n_5423)
);

INVx1_ASAP7_75t_L g5424 ( 
.A(n_4758),
.Y(n_5424)
);

OR2x2_ASAP7_75t_L g5425 ( 
.A(n_4792),
.B(n_4642),
.Y(n_5425)
);

AND2x2_ASAP7_75t_L g5426 ( 
.A(n_4683),
.B(n_4658),
.Y(n_5426)
);

INVx1_ASAP7_75t_L g5427 ( 
.A(n_4760),
.Y(n_5427)
);

INVx1_ASAP7_75t_L g5428 ( 
.A(n_4760),
.Y(n_5428)
);

BUFx3_ASAP7_75t_L g5429 ( 
.A(n_4735),
.Y(n_5429)
);

INVx2_ASAP7_75t_SL g5430 ( 
.A(n_4675),
.Y(n_5430)
);

AND2x2_ASAP7_75t_L g5431 ( 
.A(n_4683),
.B(n_4658),
.Y(n_5431)
);

INVx2_ASAP7_75t_SL g5432 ( 
.A(n_5229),
.Y(n_5432)
);

NOR2xp33_ASAP7_75t_SL g5433 ( 
.A(n_5288),
.B(n_4465),
.Y(n_5433)
);

INVx2_ASAP7_75t_SL g5434 ( 
.A(n_5229),
.Y(n_5434)
);

INVx2_ASAP7_75t_L g5435 ( 
.A(n_5366),
.Y(n_5435)
);

BUFx2_ASAP7_75t_L g5436 ( 
.A(n_5315),
.Y(n_5436)
);

OAI21x1_ASAP7_75t_L g5437 ( 
.A1(n_5247),
.A2(n_4600),
.B(n_4599),
.Y(n_5437)
);

INVx1_ASAP7_75t_L g5438 ( 
.A(n_4764),
.Y(n_5438)
);

INVx3_ASAP7_75t_L g5439 ( 
.A(n_4715),
.Y(n_5439)
);

BUFx3_ASAP7_75t_L g5440 ( 
.A(n_4735),
.Y(n_5440)
);

AND2x2_ASAP7_75t_L g5441 ( 
.A(n_4823),
.B(n_4837),
.Y(n_5441)
);

INVx1_ASAP7_75t_L g5442 ( 
.A(n_4764),
.Y(n_5442)
);

AOI21x1_ASAP7_75t_L g5443 ( 
.A1(n_5062),
.A2(n_4243),
.B(n_4432),
.Y(n_5443)
);

INVx1_ASAP7_75t_L g5444 ( 
.A(n_4767),
.Y(n_5444)
);

INVx1_ASAP7_75t_L g5445 ( 
.A(n_4767),
.Y(n_5445)
);

INVx1_ASAP7_75t_L g5446 ( 
.A(n_4775),
.Y(n_5446)
);

OA21x2_ASAP7_75t_L g5447 ( 
.A1(n_5302),
.A2(n_4954),
.B(n_4802),
.Y(n_5447)
);

INVx1_ASAP7_75t_L g5448 ( 
.A(n_4775),
.Y(n_5448)
);

OA21x2_ASAP7_75t_L g5449 ( 
.A1(n_4793),
.A2(n_4600),
.B(n_4599),
.Y(n_5449)
);

INVx1_ASAP7_75t_L g5450 ( 
.A(n_4783),
.Y(n_5450)
);

INVx1_ASAP7_75t_L g5451 ( 
.A(n_4783),
.Y(n_5451)
);

NOR2xp33_ASAP7_75t_L g5452 ( 
.A(n_4732),
.B(n_4499),
.Y(n_5452)
);

AND2x2_ASAP7_75t_L g5453 ( 
.A(n_4823),
.B(n_4418),
.Y(n_5453)
);

NOR2xp33_ASAP7_75t_L g5454 ( 
.A(n_4680),
.B(n_4621),
.Y(n_5454)
);

INVx1_ASAP7_75t_L g5455 ( 
.A(n_4786),
.Y(n_5455)
);

INVx1_ASAP7_75t_L g5456 ( 
.A(n_4786),
.Y(n_5456)
);

HB1xp67_ASAP7_75t_L g5457 ( 
.A(n_4731),
.Y(n_5457)
);

INVx2_ASAP7_75t_L g5458 ( 
.A(n_5096),
.Y(n_5458)
);

AO31x2_ASAP7_75t_L g5459 ( 
.A1(n_4700),
.A2(n_4624),
.A3(n_4595),
.B(n_4414),
.Y(n_5459)
);

AOI22xp33_ASAP7_75t_L g5460 ( 
.A1(n_4999),
.A2(n_5172),
.B1(n_4700),
.B2(n_5105),
.Y(n_5460)
);

INVx4_ASAP7_75t_SL g5461 ( 
.A(n_4752),
.Y(n_5461)
);

INVx2_ASAP7_75t_L g5462 ( 
.A(n_5096),
.Y(n_5462)
);

INVx2_ASAP7_75t_L g5463 ( 
.A(n_5096),
.Y(n_5463)
);

INVx1_ASAP7_75t_L g5464 ( 
.A(n_4799),
.Y(n_5464)
);

NAND2xp5_ASAP7_75t_L g5465 ( 
.A(n_5245),
.B(n_4241),
.Y(n_5465)
);

INVxp33_ASAP7_75t_L g5466 ( 
.A(n_4801),
.Y(n_5466)
);

INVx1_ASAP7_75t_L g5467 ( 
.A(n_4799),
.Y(n_5467)
);

BUFx6f_ASAP7_75t_L g5468 ( 
.A(n_4681),
.Y(n_5468)
);

INVx1_ASAP7_75t_L g5469 ( 
.A(n_4803),
.Y(n_5469)
);

INVx3_ASAP7_75t_L g5470 ( 
.A(n_4715),
.Y(n_5470)
);

BUFx3_ASAP7_75t_L g5471 ( 
.A(n_4735),
.Y(n_5471)
);

INVx1_ASAP7_75t_SL g5472 ( 
.A(n_5108),
.Y(n_5472)
);

NOR2xp33_ASAP7_75t_L g5473 ( 
.A(n_4680),
.B(n_4609),
.Y(n_5473)
);

AOI22xp33_ASAP7_75t_L g5474 ( 
.A1(n_4999),
.A2(n_4529),
.B1(n_4546),
.B2(n_4596),
.Y(n_5474)
);

INVx2_ASAP7_75t_L g5475 ( 
.A(n_5098),
.Y(n_5475)
);

INVx1_ASAP7_75t_L g5476 ( 
.A(n_4803),
.Y(n_5476)
);

INVx1_ASAP7_75t_L g5477 ( 
.A(n_4806),
.Y(n_5477)
);

INVx2_ASAP7_75t_L g5478 ( 
.A(n_5098),
.Y(n_5478)
);

HB1xp67_ASAP7_75t_L g5479 ( 
.A(n_4733),
.Y(n_5479)
);

AND2x2_ASAP7_75t_L g5480 ( 
.A(n_4837),
.B(n_4843),
.Y(n_5480)
);

BUFx3_ASAP7_75t_L g5481 ( 
.A(n_4735),
.Y(n_5481)
);

INVx2_ASAP7_75t_L g5482 ( 
.A(n_5098),
.Y(n_5482)
);

INVx2_ASAP7_75t_L g5483 ( 
.A(n_5099),
.Y(n_5483)
);

INVx1_ASAP7_75t_L g5484 ( 
.A(n_4806),
.Y(n_5484)
);

INVxp67_ASAP7_75t_L g5485 ( 
.A(n_5175),
.Y(n_5485)
);

INVx2_ASAP7_75t_L g5486 ( 
.A(n_5099),
.Y(n_5486)
);

HB1xp67_ASAP7_75t_L g5487 ( 
.A(n_4768),
.Y(n_5487)
);

OAI22xp33_ASAP7_75t_L g5488 ( 
.A1(n_4944),
.A2(n_4428),
.B1(n_4363),
.B2(n_4445),
.Y(n_5488)
);

INVx1_ASAP7_75t_SL g5489 ( 
.A(n_5124),
.Y(n_5489)
);

INVx2_ASAP7_75t_L g5490 ( 
.A(n_5099),
.Y(n_5490)
);

INVx1_ASAP7_75t_L g5491 ( 
.A(n_4811),
.Y(n_5491)
);

INVx1_ASAP7_75t_L g5492 ( 
.A(n_4811),
.Y(n_5492)
);

HB1xp67_ASAP7_75t_L g5493 ( 
.A(n_4943),
.Y(n_5493)
);

BUFx2_ASAP7_75t_L g5494 ( 
.A(n_5315),
.Y(n_5494)
);

INVx1_ASAP7_75t_L g5495 ( 
.A(n_4824),
.Y(n_5495)
);

NOR2xp33_ASAP7_75t_L g5496 ( 
.A(n_4753),
.B(n_4609),
.Y(n_5496)
);

BUFx2_ASAP7_75t_L g5497 ( 
.A(n_4853),
.Y(n_5497)
);

BUFx2_ASAP7_75t_SL g5498 ( 
.A(n_5137),
.Y(n_5498)
);

INVx2_ASAP7_75t_L g5499 ( 
.A(n_5111),
.Y(n_5499)
);

INVx1_ASAP7_75t_L g5500 ( 
.A(n_4824),
.Y(n_5500)
);

INVxp67_ASAP7_75t_L g5501 ( 
.A(n_5175),
.Y(n_5501)
);

INVx6_ASAP7_75t_L g5502 ( 
.A(n_4748),
.Y(n_5502)
);

HB1xp67_ASAP7_75t_L g5503 ( 
.A(n_4967),
.Y(n_5503)
);

OR2x2_ASAP7_75t_L g5504 ( 
.A(n_4792),
.B(n_4337),
.Y(n_5504)
);

HB1xp67_ASAP7_75t_L g5505 ( 
.A(n_4992),
.Y(n_5505)
);

AOI22xp33_ASAP7_75t_L g5506 ( 
.A1(n_5105),
.A2(n_4546),
.B1(n_4480),
.B2(n_4194),
.Y(n_5506)
);

AND2x2_ASAP7_75t_L g5507 ( 
.A(n_4843),
.B(n_4769),
.Y(n_5507)
);

AO21x1_ASAP7_75t_L g5508 ( 
.A1(n_5135),
.A2(n_4150),
.B(n_4194),
.Y(n_5508)
);

OR2x2_ASAP7_75t_L g5509 ( 
.A(n_4818),
.B(n_4888),
.Y(n_5509)
);

INVx1_ASAP7_75t_L g5510 ( 
.A(n_4829),
.Y(n_5510)
);

INVx1_ASAP7_75t_L g5511 ( 
.A(n_4829),
.Y(n_5511)
);

OAI21xp5_ASAP7_75t_L g5512 ( 
.A1(n_4861),
.A2(n_4156),
.B(n_4297),
.Y(n_5512)
);

OAI211xp5_ASAP7_75t_L g5513 ( 
.A1(n_4861),
.A2(n_5245),
.B(n_4991),
.C(n_5360),
.Y(n_5513)
);

INVx1_ASAP7_75t_L g5514 ( 
.A(n_4830),
.Y(n_5514)
);

INVx5_ASAP7_75t_SL g5515 ( 
.A(n_4805),
.Y(n_5515)
);

AO31x2_ASAP7_75t_L g5516 ( 
.A1(n_4927),
.A2(n_4551),
.A3(n_4217),
.B(n_4235),
.Y(n_5516)
);

INVx2_ASAP7_75t_SL g5517 ( 
.A(n_4681),
.Y(n_5517)
);

INVx1_ASAP7_75t_L g5518 ( 
.A(n_4830),
.Y(n_5518)
);

INVx1_ASAP7_75t_L g5519 ( 
.A(n_4835),
.Y(n_5519)
);

INVx2_ASAP7_75t_L g5520 ( 
.A(n_5111),
.Y(n_5520)
);

INVx3_ASAP7_75t_L g5521 ( 
.A(n_4715),
.Y(n_5521)
);

INVx1_ASAP7_75t_L g5522 ( 
.A(n_4835),
.Y(n_5522)
);

INVx1_ASAP7_75t_L g5523 ( 
.A(n_4840),
.Y(n_5523)
);

INVx2_ASAP7_75t_L g5524 ( 
.A(n_5111),
.Y(n_5524)
);

AND2x4_ASAP7_75t_L g5525 ( 
.A(n_4865),
.B(n_4507),
.Y(n_5525)
);

INVx1_ASAP7_75t_L g5526 ( 
.A(n_4840),
.Y(n_5526)
);

OAI21x1_ASAP7_75t_L g5527 ( 
.A1(n_5247),
.A2(n_4610),
.B(n_4603),
.Y(n_5527)
);

INVx2_ASAP7_75t_SL g5528 ( 
.A(n_4681),
.Y(n_5528)
);

OAI21x1_ASAP7_75t_L g5529 ( 
.A1(n_5156),
.A2(n_4610),
.B(n_4603),
.Y(n_5529)
);

INVx1_ASAP7_75t_L g5530 ( 
.A(n_4841),
.Y(n_5530)
);

INVx1_ASAP7_75t_L g5531 ( 
.A(n_4841),
.Y(n_5531)
);

OAI21x1_ASAP7_75t_L g5532 ( 
.A1(n_5156),
.A2(n_4610),
.B(n_4603),
.Y(n_5532)
);

INVx1_ASAP7_75t_L g5533 ( 
.A(n_4857),
.Y(n_5533)
);

OA21x2_ASAP7_75t_L g5534 ( 
.A1(n_4793),
.A2(n_4816),
.B(n_4802),
.Y(n_5534)
);

HB1xp67_ASAP7_75t_L g5535 ( 
.A(n_5027),
.Y(n_5535)
);

INVx1_ASAP7_75t_L g5536 ( 
.A(n_4857),
.Y(n_5536)
);

INVx1_ASAP7_75t_L g5537 ( 
.A(n_4866),
.Y(n_5537)
);

INVx2_ASAP7_75t_L g5538 ( 
.A(n_5115),
.Y(n_5538)
);

NAND2xp5_ASAP7_75t_L g5539 ( 
.A(n_5330),
.B(n_4241),
.Y(n_5539)
);

NAND2xp5_ASAP7_75t_L g5540 ( 
.A(n_5330),
.B(n_4436),
.Y(n_5540)
);

INVx2_ASAP7_75t_L g5541 ( 
.A(n_5115),
.Y(n_5541)
);

HB1xp67_ASAP7_75t_L g5542 ( 
.A(n_5067),
.Y(n_5542)
);

BUFx6f_ASAP7_75t_L g5543 ( 
.A(n_4753),
.Y(n_5543)
);

AOI22xp33_ASAP7_75t_L g5544 ( 
.A1(n_4784),
.A2(n_4546),
.B1(n_4480),
.B2(n_4428),
.Y(n_5544)
);

INVx1_ASAP7_75t_L g5545 ( 
.A(n_4866),
.Y(n_5545)
);

NAND2xp5_ASAP7_75t_L g5546 ( 
.A(n_5200),
.B(n_4436),
.Y(n_5546)
);

AOI21x1_ASAP7_75t_L g5547 ( 
.A1(n_5076),
.A2(n_4243),
.B(n_4432),
.Y(n_5547)
);

INVx1_ASAP7_75t_L g5548 ( 
.A(n_4870),
.Y(n_5548)
);

BUFx3_ASAP7_75t_L g5549 ( 
.A(n_4748),
.Y(n_5549)
);

INVx1_ASAP7_75t_L g5550 ( 
.A(n_4870),
.Y(n_5550)
);

BUFx6f_ASAP7_75t_L g5551 ( 
.A(n_4753),
.Y(n_5551)
);

BUFx10_ASAP7_75t_L g5552 ( 
.A(n_5151),
.Y(n_5552)
);

INVx1_ASAP7_75t_L g5553 ( 
.A(n_4875),
.Y(n_5553)
);

INVx2_ASAP7_75t_L g5554 ( 
.A(n_5115),
.Y(n_5554)
);

AND2x2_ASAP7_75t_L g5555 ( 
.A(n_4769),
.B(n_4418),
.Y(n_5555)
);

INVx2_ASAP7_75t_L g5556 ( 
.A(n_4674),
.Y(n_5556)
);

HB1xp67_ASAP7_75t_L g5557 ( 
.A(n_5094),
.Y(n_5557)
);

NAND2xp5_ASAP7_75t_L g5558 ( 
.A(n_4784),
.B(n_4184),
.Y(n_5558)
);

INVx1_ASAP7_75t_SL g5559 ( 
.A(n_5128),
.Y(n_5559)
);

NAND2xp33_ASAP7_75t_R g5560 ( 
.A(n_4746),
.B(n_4186),
.Y(n_5560)
);

INVx2_ASAP7_75t_L g5561 ( 
.A(n_4674),
.Y(n_5561)
);

INVx1_ASAP7_75t_L g5562 ( 
.A(n_4875),
.Y(n_5562)
);

HB1xp67_ASAP7_75t_L g5563 ( 
.A(n_5158),
.Y(n_5563)
);

AND2x4_ASAP7_75t_L g5564 ( 
.A(n_4865),
.B(n_4444),
.Y(n_5564)
);

INVx1_ASAP7_75t_L g5565 ( 
.A(n_4877),
.Y(n_5565)
);

HB1xp67_ASAP7_75t_L g5566 ( 
.A(n_5160),
.Y(n_5566)
);

INVx1_ASAP7_75t_L g5567 ( 
.A(n_4877),
.Y(n_5567)
);

BUFx6f_ASAP7_75t_L g5568 ( 
.A(n_4884),
.Y(n_5568)
);

INVx2_ASAP7_75t_L g5569 ( 
.A(n_4674),
.Y(n_5569)
);

INVx1_ASAP7_75t_L g5570 ( 
.A(n_4878),
.Y(n_5570)
);

INVx1_ASAP7_75t_L g5571 ( 
.A(n_4878),
.Y(n_5571)
);

INVx1_ASAP7_75t_L g5572 ( 
.A(n_4883),
.Y(n_5572)
);

INVx1_ASAP7_75t_L g5573 ( 
.A(n_4883),
.Y(n_5573)
);

OA21x2_ASAP7_75t_L g5574 ( 
.A1(n_4793),
.A2(n_4617),
.B(n_4615),
.Y(n_5574)
);

INVx1_ASAP7_75t_L g5575 ( 
.A(n_4900),
.Y(n_5575)
);

INVx1_ASAP7_75t_L g5576 ( 
.A(n_4900),
.Y(n_5576)
);

INVx1_ASAP7_75t_L g5577 ( 
.A(n_4903),
.Y(n_5577)
);

AOI21xp5_ASAP7_75t_L g5578 ( 
.A1(n_4899),
.A2(n_4312),
.B(n_4309),
.Y(n_5578)
);

INVxp67_ASAP7_75t_L g5579 ( 
.A(n_4746),
.Y(n_5579)
);

INVx1_ASAP7_75t_L g5580 ( 
.A(n_4903),
.Y(n_5580)
);

INVx1_ASAP7_75t_L g5581 ( 
.A(n_4905),
.Y(n_5581)
);

INVx2_ASAP7_75t_L g5582 ( 
.A(n_4678),
.Y(n_5582)
);

INVx2_ASAP7_75t_L g5583 ( 
.A(n_4678),
.Y(n_5583)
);

INVx2_ASAP7_75t_L g5584 ( 
.A(n_4678),
.Y(n_5584)
);

INVx1_ASAP7_75t_L g5585 ( 
.A(n_4905),
.Y(n_5585)
);

INVx2_ASAP7_75t_L g5586 ( 
.A(n_4687),
.Y(n_5586)
);

INVx2_ASAP7_75t_SL g5587 ( 
.A(n_5016),
.Y(n_5587)
);

NAND2x1p5_ASAP7_75t_L g5588 ( 
.A(n_5319),
.B(n_4645),
.Y(n_5588)
);

AND2x2_ASAP7_75t_L g5589 ( 
.A(n_4673),
.B(n_4433),
.Y(n_5589)
);

INVx1_ASAP7_75t_L g5590 ( 
.A(n_4908),
.Y(n_5590)
);

INVx3_ASAP7_75t_L g5591 ( 
.A(n_4715),
.Y(n_5591)
);

INVx2_ASAP7_75t_L g5592 ( 
.A(n_4687),
.Y(n_5592)
);

AO21x1_ASAP7_75t_L g5593 ( 
.A1(n_5135),
.A2(n_4156),
.B(n_4341),
.Y(n_5593)
);

INVx2_ASAP7_75t_L g5594 ( 
.A(n_4687),
.Y(n_5594)
);

INVx1_ASAP7_75t_L g5595 ( 
.A(n_4908),
.Y(n_5595)
);

INVx2_ASAP7_75t_L g5596 ( 
.A(n_4696),
.Y(n_5596)
);

INVx1_ASAP7_75t_L g5597 ( 
.A(n_4915),
.Y(n_5597)
);

INVx1_ASAP7_75t_L g5598 ( 
.A(n_4915),
.Y(n_5598)
);

INVx1_ASAP7_75t_L g5599 ( 
.A(n_4916),
.Y(n_5599)
);

INVx2_ASAP7_75t_L g5600 ( 
.A(n_4696),
.Y(n_5600)
);

AND2x4_ASAP7_75t_L g5601 ( 
.A(n_4865),
.B(n_4444),
.Y(n_5601)
);

HB1xp67_ASAP7_75t_L g5602 ( 
.A(n_5165),
.Y(n_5602)
);

BUFx3_ASAP7_75t_L g5603 ( 
.A(n_4748),
.Y(n_5603)
);

INVx3_ASAP7_75t_L g5604 ( 
.A(n_4715),
.Y(n_5604)
);

INVx1_ASAP7_75t_L g5605 ( 
.A(n_4916),
.Y(n_5605)
);

INVx1_ASAP7_75t_L g5606 ( 
.A(n_4919),
.Y(n_5606)
);

AOI22xp5_ASAP7_75t_L g5607 ( 
.A1(n_4738),
.A2(n_4517),
.B1(n_4445),
.B2(n_4438),
.Y(n_5607)
);

BUFx12f_ASAP7_75t_L g5608 ( 
.A(n_4748),
.Y(n_5608)
);

INVx3_ASAP7_75t_L g5609 ( 
.A(n_4865),
.Y(n_5609)
);

OAI21x1_ASAP7_75t_L g5610 ( 
.A1(n_5153),
.A2(n_4617),
.B(n_4615),
.Y(n_5610)
);

INVx1_ASAP7_75t_L g5611 ( 
.A(n_4919),
.Y(n_5611)
);

INVx1_ASAP7_75t_L g5612 ( 
.A(n_4930),
.Y(n_5612)
);

INVx1_ASAP7_75t_L g5613 ( 
.A(n_4930),
.Y(n_5613)
);

INVx2_ASAP7_75t_L g5614 ( 
.A(n_4696),
.Y(n_5614)
);

INVx1_ASAP7_75t_L g5615 ( 
.A(n_4933),
.Y(n_5615)
);

INVx2_ASAP7_75t_L g5616 ( 
.A(n_4698),
.Y(n_5616)
);

AND2x2_ASAP7_75t_L g5617 ( 
.A(n_4673),
.B(n_4433),
.Y(n_5617)
);

AND2x2_ASAP7_75t_L g5618 ( 
.A(n_4673),
.B(n_4441),
.Y(n_5618)
);

INVx2_ASAP7_75t_L g5619 ( 
.A(n_4698),
.Y(n_5619)
);

INVx2_ASAP7_75t_L g5620 ( 
.A(n_4698),
.Y(n_5620)
);

INVx3_ASAP7_75t_L g5621 ( 
.A(n_4937),
.Y(n_5621)
);

INVx2_ASAP7_75t_L g5622 ( 
.A(n_4723),
.Y(n_5622)
);

INVx1_ASAP7_75t_L g5623 ( 
.A(n_4933),
.Y(n_5623)
);

INVx2_ASAP7_75t_L g5624 ( 
.A(n_4723),
.Y(n_5624)
);

INVx2_ASAP7_75t_L g5625 ( 
.A(n_4723),
.Y(n_5625)
);

OA21x2_ASAP7_75t_L g5626 ( 
.A1(n_4802),
.A2(n_4828),
.B(n_4816),
.Y(n_5626)
);

OR2x6_ASAP7_75t_L g5627 ( 
.A(n_5123),
.B(n_4312),
.Y(n_5627)
);

HB1xp67_ASAP7_75t_L g5628 ( 
.A(n_5174),
.Y(n_5628)
);

OR2x6_ASAP7_75t_L g5629 ( 
.A(n_5123),
.B(n_4182),
.Y(n_5629)
);

INVx1_ASAP7_75t_L g5630 ( 
.A(n_4950),
.Y(n_5630)
);

INVx2_ASAP7_75t_L g5631 ( 
.A(n_4728),
.Y(n_5631)
);

INVx2_ASAP7_75t_L g5632 ( 
.A(n_4728),
.Y(n_5632)
);

INVxp33_ASAP7_75t_L g5633 ( 
.A(n_5269),
.Y(n_5633)
);

INVxp67_ASAP7_75t_SL g5634 ( 
.A(n_4927),
.Y(n_5634)
);

INVx1_ASAP7_75t_L g5635 ( 
.A(n_4950),
.Y(n_5635)
);

HB1xp67_ASAP7_75t_L g5636 ( 
.A(n_4825),
.Y(n_5636)
);

AOI211xp5_ASAP7_75t_L g5637 ( 
.A1(n_5352),
.A2(n_4440),
.B(n_4576),
.C(n_4293),
.Y(n_5637)
);

HB1xp67_ASAP7_75t_L g5638 ( 
.A(n_4867),
.Y(n_5638)
);

NAND2xp5_ASAP7_75t_L g5639 ( 
.A(n_5359),
.B(n_5352),
.Y(n_5639)
);

INVx1_ASAP7_75t_L g5640 ( 
.A(n_4951),
.Y(n_5640)
);

INVx1_ASAP7_75t_L g5641 ( 
.A(n_4951),
.Y(n_5641)
);

INVx1_ASAP7_75t_L g5642 ( 
.A(n_4955),
.Y(n_5642)
);

INVx3_ASAP7_75t_L g5643 ( 
.A(n_4937),
.Y(n_5643)
);

AOI22xp33_ASAP7_75t_L g5644 ( 
.A1(n_4690),
.A2(n_4480),
.B1(n_4281),
.B2(n_4228),
.Y(n_5644)
);

BUFx12f_ASAP7_75t_L g5645 ( 
.A(n_4796),
.Y(n_5645)
);

INVx1_ASAP7_75t_L g5646 ( 
.A(n_4955),
.Y(n_5646)
);

INVx1_ASAP7_75t_L g5647 ( 
.A(n_4956),
.Y(n_5647)
);

INVx2_ASAP7_75t_L g5648 ( 
.A(n_4728),
.Y(n_5648)
);

AND2x2_ASAP7_75t_L g5649 ( 
.A(n_4673),
.B(n_4708),
.Y(n_5649)
);

AOI21xp5_ASAP7_75t_L g5650 ( 
.A1(n_4936),
.A2(n_4405),
.B(n_4626),
.Y(n_5650)
);

INVxp33_ASAP7_75t_L g5651 ( 
.A(n_5183),
.Y(n_5651)
);

INVx2_ASAP7_75t_L g5652 ( 
.A(n_4734),
.Y(n_5652)
);

INVx1_ASAP7_75t_SL g5653 ( 
.A(n_4684),
.Y(n_5653)
);

INVx1_ASAP7_75t_L g5654 ( 
.A(n_4956),
.Y(n_5654)
);

OAI22xp33_ASAP7_75t_L g5655 ( 
.A1(n_4944),
.A2(n_4343),
.B1(n_4266),
.B2(n_4413),
.Y(n_5655)
);

INVx2_ASAP7_75t_L g5656 ( 
.A(n_4734),
.Y(n_5656)
);

INVx1_ASAP7_75t_L g5657 ( 
.A(n_4964),
.Y(n_5657)
);

INVx1_ASAP7_75t_L g5658 ( 
.A(n_4964),
.Y(n_5658)
);

INVx1_ASAP7_75t_L g5659 ( 
.A(n_4968),
.Y(n_5659)
);

BUFx2_ASAP7_75t_L g5660 ( 
.A(n_4765),
.Y(n_5660)
);

AND2x2_ASAP7_75t_L g5661 ( 
.A(n_4708),
.B(n_4441),
.Y(n_5661)
);

CKINVDCx20_ASAP7_75t_R g5662 ( 
.A(n_4697),
.Y(n_5662)
);

INVx1_ASAP7_75t_L g5663 ( 
.A(n_4968),
.Y(n_5663)
);

BUFx3_ASAP7_75t_L g5664 ( 
.A(n_4884),
.Y(n_5664)
);

INVx3_ASAP7_75t_L g5665 ( 
.A(n_4937),
.Y(n_5665)
);

INVx2_ASAP7_75t_L g5666 ( 
.A(n_4734),
.Y(n_5666)
);

INVx1_ASAP7_75t_L g5667 ( 
.A(n_4970),
.Y(n_5667)
);

INVx2_ASAP7_75t_L g5668 ( 
.A(n_4745),
.Y(n_5668)
);

AND2x4_ASAP7_75t_L g5669 ( 
.A(n_4852),
.B(n_4431),
.Y(n_5669)
);

AOI22xp5_ASAP7_75t_L g5670 ( 
.A1(n_4738),
.A2(n_5061),
.B1(n_5268),
.B2(n_5233),
.Y(n_5670)
);

INVx2_ASAP7_75t_SL g5671 ( 
.A(n_5016),
.Y(n_5671)
);

BUFx2_ASAP7_75t_L g5672 ( 
.A(n_4765),
.Y(n_5672)
);

AND2x4_ASAP7_75t_L g5673 ( 
.A(n_4852),
.B(n_4431),
.Y(n_5673)
);

AND2x4_ASAP7_75t_L g5674 ( 
.A(n_4852),
.B(n_4480),
.Y(n_5674)
);

INVx1_ASAP7_75t_L g5675 ( 
.A(n_4970),
.Y(n_5675)
);

INVx1_ASAP7_75t_L g5676 ( 
.A(n_4977),
.Y(n_5676)
);

AOI211xp5_ASAP7_75t_L g5677 ( 
.A1(n_5359),
.A2(n_4293),
.B(n_4245),
.C(n_4413),
.Y(n_5677)
);

INVx2_ASAP7_75t_SL g5678 ( 
.A(n_5016),
.Y(n_5678)
);

AND2x2_ASAP7_75t_L g5679 ( 
.A(n_4708),
.B(n_4170),
.Y(n_5679)
);

INVx1_ASAP7_75t_L g5680 ( 
.A(n_4977),
.Y(n_5680)
);

INVx2_ASAP7_75t_L g5681 ( 
.A(n_4745),
.Y(n_5681)
);

BUFx6f_ASAP7_75t_L g5682 ( 
.A(n_4884),
.Y(n_5682)
);

AND2x2_ASAP7_75t_L g5683 ( 
.A(n_4708),
.B(n_4170),
.Y(n_5683)
);

BUFx2_ASAP7_75t_L g5684 ( 
.A(n_4958),
.Y(n_5684)
);

INVx2_ASAP7_75t_L g5685 ( 
.A(n_4745),
.Y(n_5685)
);

BUFx2_ASAP7_75t_L g5686 ( 
.A(n_4958),
.Y(n_5686)
);

AOI21xp5_ASAP7_75t_L g5687 ( 
.A1(n_4936),
.A2(n_4406),
.B(n_4245),
.Y(n_5687)
);

INVx1_ASAP7_75t_L g5688 ( 
.A(n_4979),
.Y(n_5688)
);

AND2x2_ASAP7_75t_L g5689 ( 
.A(n_4722),
.B(n_4170),
.Y(n_5689)
);

AOI22xp33_ASAP7_75t_SL g5690 ( 
.A1(n_5205),
.A2(n_4180),
.B1(n_4205),
.B2(n_4225),
.Y(n_5690)
);

INVx2_ASAP7_75t_L g5691 ( 
.A(n_4754),
.Y(n_5691)
);

OAI21x1_ASAP7_75t_L g5692 ( 
.A1(n_5153),
.A2(n_4617),
.B(n_4615),
.Y(n_5692)
);

INVx1_ASAP7_75t_L g5693 ( 
.A(n_4979),
.Y(n_5693)
);

AO31x2_ASAP7_75t_L g5694 ( 
.A1(n_5331),
.A2(n_4218),
.A3(n_4235),
.B(n_4217),
.Y(n_5694)
);

NOR2x1_ASAP7_75t_SL g5695 ( 
.A(n_5073),
.B(n_4442),
.Y(n_5695)
);

BUFx3_ASAP7_75t_L g5696 ( 
.A(n_4891),
.Y(n_5696)
);

INVx1_ASAP7_75t_L g5697 ( 
.A(n_4980),
.Y(n_5697)
);

INVx1_ASAP7_75t_L g5698 ( 
.A(n_4980),
.Y(n_5698)
);

INVx4_ASAP7_75t_L g5699 ( 
.A(n_4891),
.Y(n_5699)
);

INVx1_ASAP7_75t_L g5700 ( 
.A(n_4984),
.Y(n_5700)
);

INVx1_ASAP7_75t_L g5701 ( 
.A(n_4984),
.Y(n_5701)
);

INVx1_ASAP7_75t_L g5702 ( 
.A(n_4989),
.Y(n_5702)
);

INVx2_ASAP7_75t_L g5703 ( 
.A(n_4754),
.Y(n_5703)
);

INVx2_ASAP7_75t_L g5704 ( 
.A(n_4754),
.Y(n_5704)
);

INVx2_ASAP7_75t_L g5705 ( 
.A(n_5065),
.Y(n_5705)
);

AOI21xp5_ASAP7_75t_L g5706 ( 
.A1(n_4910),
.A2(n_4406),
.B(n_4174),
.Y(n_5706)
);

INVx1_ASAP7_75t_L g5707 ( 
.A(n_4989),
.Y(n_5707)
);

AND2x4_ASAP7_75t_L g5708 ( 
.A(n_4852),
.B(n_4170),
.Y(n_5708)
);

INVx2_ASAP7_75t_L g5709 ( 
.A(n_5065),
.Y(n_5709)
);

BUFx3_ASAP7_75t_L g5710 ( 
.A(n_4891),
.Y(n_5710)
);

INVxp67_ASAP7_75t_L g5711 ( 
.A(n_5149),
.Y(n_5711)
);

INVx2_ASAP7_75t_SL g5712 ( 
.A(n_5033),
.Y(n_5712)
);

A2O1A1Ixp33_ASAP7_75t_L g5713 ( 
.A1(n_5038),
.A2(n_4343),
.B(n_4266),
.C(n_4619),
.Y(n_5713)
);

OR2x2_ASAP7_75t_L g5714 ( 
.A(n_4818),
.B(n_4337),
.Y(n_5714)
);

AND2x2_ASAP7_75t_L g5715 ( 
.A(n_4722),
.B(n_4173),
.Y(n_5715)
);

INVx3_ASAP7_75t_L g5716 ( 
.A(n_4937),
.Y(n_5716)
);

AOI21xp5_ASAP7_75t_L g5717 ( 
.A1(n_4910),
.A2(n_5032),
.B(n_5038),
.Y(n_5717)
);

INVx3_ASAP7_75t_L g5718 ( 
.A(n_4946),
.Y(n_5718)
);

BUFx2_ASAP7_75t_L g5719 ( 
.A(n_4958),
.Y(n_5719)
);

INVx2_ASAP7_75t_L g5720 ( 
.A(n_5065),
.Y(n_5720)
);

AOI21x1_ASAP7_75t_L g5721 ( 
.A1(n_5076),
.A2(n_4434),
.B(n_4643),
.Y(n_5721)
);

INVx2_ASAP7_75t_L g5722 ( 
.A(n_5072),
.Y(n_5722)
);

INVx1_ASAP7_75t_L g5723 ( 
.A(n_4990),
.Y(n_5723)
);

INVx3_ASAP7_75t_L g5724 ( 
.A(n_4946),
.Y(n_5724)
);

INVx1_ASAP7_75t_SL g5725 ( 
.A(n_4684),
.Y(n_5725)
);

AND2x2_ASAP7_75t_L g5726 ( 
.A(n_4722),
.B(n_4173),
.Y(n_5726)
);

NOR2xp33_ASAP7_75t_SL g5727 ( 
.A(n_5288),
.B(n_4528),
.Y(n_5727)
);

INVx1_ASAP7_75t_L g5728 ( 
.A(n_4990),
.Y(n_5728)
);

OAI21xp5_ASAP7_75t_L g5729 ( 
.A1(n_5021),
.A2(n_4601),
.B(n_4636),
.Y(n_5729)
);

INVx2_ASAP7_75t_L g5730 ( 
.A(n_5072),
.Y(n_5730)
);

INVx1_ASAP7_75t_L g5731 ( 
.A(n_4995),
.Y(n_5731)
);

INVx1_ASAP7_75t_L g5732 ( 
.A(n_4995),
.Y(n_5732)
);

AO21x2_ASAP7_75t_L g5733 ( 
.A1(n_5331),
.A2(n_4582),
.B(n_4423),
.Y(n_5733)
);

INVx2_ASAP7_75t_L g5734 ( 
.A(n_5072),
.Y(n_5734)
);

INVx2_ASAP7_75t_L g5735 ( 
.A(n_5080),
.Y(n_5735)
);

INVx1_ASAP7_75t_L g5736 ( 
.A(n_5002),
.Y(n_5736)
);

INVx1_ASAP7_75t_L g5737 ( 
.A(n_5002),
.Y(n_5737)
);

INVx1_ASAP7_75t_L g5738 ( 
.A(n_5003),
.Y(n_5738)
);

INVx2_ASAP7_75t_L g5739 ( 
.A(n_5080),
.Y(n_5739)
);

INVx2_ASAP7_75t_L g5740 ( 
.A(n_5080),
.Y(n_5740)
);

AND2x4_ASAP7_75t_L g5741 ( 
.A(n_4852),
.B(n_4173),
.Y(n_5741)
);

BUFx2_ASAP7_75t_SL g5742 ( 
.A(n_4938),
.Y(n_5742)
);

INVx2_ASAP7_75t_L g5743 ( 
.A(n_5091),
.Y(n_5743)
);

INVx2_ASAP7_75t_L g5744 ( 
.A(n_5091),
.Y(n_5744)
);

AND2x2_ASAP7_75t_L g5745 ( 
.A(n_4722),
.B(n_4173),
.Y(n_5745)
);

INVx1_ASAP7_75t_L g5746 ( 
.A(n_5003),
.Y(n_5746)
);

AND2x2_ASAP7_75t_L g5747 ( 
.A(n_4782),
.B(n_4231),
.Y(n_5747)
);

INVx1_ASAP7_75t_L g5748 ( 
.A(n_5004),
.Y(n_5748)
);

HB1xp67_ASAP7_75t_L g5749 ( 
.A(n_4886),
.Y(n_5749)
);

HB1xp67_ASAP7_75t_L g5750 ( 
.A(n_4890),
.Y(n_5750)
);

INVx2_ASAP7_75t_L g5751 ( 
.A(n_5091),
.Y(n_5751)
);

INVx1_ASAP7_75t_L g5752 ( 
.A(n_5004),
.Y(n_5752)
);

NAND2x1p5_ASAP7_75t_L g5753 ( 
.A(n_5319),
.B(n_4645),
.Y(n_5753)
);

INVx2_ASAP7_75t_L g5754 ( 
.A(n_5093),
.Y(n_5754)
);

NOR2xp33_ASAP7_75t_L g5755 ( 
.A(n_5147),
.B(n_4622),
.Y(n_5755)
);

INVx1_ASAP7_75t_L g5756 ( 
.A(n_5010),
.Y(n_5756)
);

INVx1_ASAP7_75t_L g5757 ( 
.A(n_5010),
.Y(n_5757)
);

INVx2_ASAP7_75t_SL g5758 ( 
.A(n_5033),
.Y(n_5758)
);

INVx1_ASAP7_75t_L g5759 ( 
.A(n_5011),
.Y(n_5759)
);

INVx1_ASAP7_75t_L g5760 ( 
.A(n_5011),
.Y(n_5760)
);

INVx1_ASAP7_75t_L g5761 ( 
.A(n_5014),
.Y(n_5761)
);

INVx2_ASAP7_75t_SL g5762 ( 
.A(n_5033),
.Y(n_5762)
);

NAND2xp5_ASAP7_75t_L g5763 ( 
.A(n_5233),
.B(n_4184),
.Y(n_5763)
);

OAI21x1_ASAP7_75t_L g5764 ( 
.A1(n_5142),
.A2(n_4627),
.B(n_4618),
.Y(n_5764)
);

INVx1_ASAP7_75t_L g5765 ( 
.A(n_5014),
.Y(n_5765)
);

INVx2_ASAP7_75t_L g5766 ( 
.A(n_5093),
.Y(n_5766)
);

INVx3_ASAP7_75t_L g5767 ( 
.A(n_4946),
.Y(n_5767)
);

INVx1_ASAP7_75t_L g5768 ( 
.A(n_5017),
.Y(n_5768)
);

INVx1_ASAP7_75t_L g5769 ( 
.A(n_5017),
.Y(n_5769)
);

INVx1_ASAP7_75t_L g5770 ( 
.A(n_5018),
.Y(n_5770)
);

INVx2_ASAP7_75t_L g5771 ( 
.A(n_5093),
.Y(n_5771)
);

INVx2_ASAP7_75t_SL g5772 ( 
.A(n_5033),
.Y(n_5772)
);

INVx1_ASAP7_75t_L g5773 ( 
.A(n_5018),
.Y(n_5773)
);

INVx1_ASAP7_75t_L g5774 ( 
.A(n_5025),
.Y(n_5774)
);

BUFx3_ASAP7_75t_L g5775 ( 
.A(n_4901),
.Y(n_5775)
);

OAI21x1_ASAP7_75t_L g5776 ( 
.A1(n_5142),
.A2(n_4627),
.B(n_4618),
.Y(n_5776)
);

INVx1_ASAP7_75t_L g5777 ( 
.A(n_5025),
.Y(n_5777)
);

INVx2_ASAP7_75t_L g5778 ( 
.A(n_4985),
.Y(n_5778)
);

OAI21xp5_ASAP7_75t_L g5779 ( 
.A1(n_5021),
.A2(n_4601),
.B(n_4636),
.Y(n_5779)
);

INVx2_ASAP7_75t_SL g5780 ( 
.A(n_4969),
.Y(n_5780)
);

INVx2_ASAP7_75t_L g5781 ( 
.A(n_4985),
.Y(n_5781)
);

INVx2_ASAP7_75t_SL g5782 ( 
.A(n_4969),
.Y(n_5782)
);

NOR2xp33_ASAP7_75t_L g5783 ( 
.A(n_4901),
.B(n_4622),
.Y(n_5783)
);

OAI21x1_ASAP7_75t_L g5784 ( 
.A1(n_4743),
.A2(n_4627),
.B(n_4618),
.Y(n_5784)
);

AND2x2_ASAP7_75t_L g5785 ( 
.A(n_4782),
.B(n_4231),
.Y(n_5785)
);

OAI21x1_ASAP7_75t_L g5786 ( 
.A1(n_4743),
.A2(n_4598),
.B(n_4462),
.Y(n_5786)
);

HB1xp67_ASAP7_75t_L g5787 ( 
.A(n_5231),
.Y(n_5787)
);

INVx1_ASAP7_75t_L g5788 ( 
.A(n_5029),
.Y(n_5788)
);

INVx3_ASAP7_75t_L g5789 ( 
.A(n_4946),
.Y(n_5789)
);

OAI22xp33_ASAP7_75t_SL g5790 ( 
.A1(n_4699),
.A2(n_4705),
.B1(n_4707),
.B2(n_4949),
.Y(n_5790)
);

INVx3_ASAP7_75t_L g5791 ( 
.A(n_5024),
.Y(n_5791)
);

HB1xp67_ASAP7_75t_L g5792 ( 
.A(n_5235),
.Y(n_5792)
);

HB1xp67_ASAP7_75t_L g5793 ( 
.A(n_5257),
.Y(n_5793)
);

INVx2_ASAP7_75t_L g5794 ( 
.A(n_4985),
.Y(n_5794)
);

INVx2_ASAP7_75t_L g5795 ( 
.A(n_4986),
.Y(n_5795)
);

INVx2_ASAP7_75t_L g5796 ( 
.A(n_4986),
.Y(n_5796)
);

AOI21x1_ASAP7_75t_L g5797 ( 
.A1(n_5086),
.A2(n_4434),
.B(n_4218),
.Y(n_5797)
);

OA21x2_ASAP7_75t_L g5798 ( 
.A1(n_4816),
.A2(n_4598),
.B(n_4200),
.Y(n_5798)
);

OR2x2_ASAP7_75t_L g5799 ( 
.A(n_4888),
.B(n_4362),
.Y(n_5799)
);

INVx1_ASAP7_75t_L g5800 ( 
.A(n_5029),
.Y(n_5800)
);

BUFx2_ASAP7_75t_SL g5801 ( 
.A(n_5009),
.Y(n_5801)
);

HB1xp67_ASAP7_75t_SL g5802 ( 
.A(n_4998),
.Y(n_5802)
);

AND2x2_ASAP7_75t_L g5803 ( 
.A(n_4790),
.B(n_4231),
.Y(n_5803)
);

NAND2xp5_ASAP7_75t_L g5804 ( 
.A(n_5032),
.B(n_4185),
.Y(n_5804)
);

INVx2_ASAP7_75t_L g5805 ( 
.A(n_4986),
.Y(n_5805)
);

BUFx2_ASAP7_75t_L g5806 ( 
.A(n_4812),
.Y(n_5806)
);

INVx1_ASAP7_75t_L g5807 ( 
.A(n_5045),
.Y(n_5807)
);

INVx3_ASAP7_75t_L g5808 ( 
.A(n_5024),
.Y(n_5808)
);

AO21x1_ASAP7_75t_SL g5809 ( 
.A1(n_5310),
.A2(n_4185),
.B(n_4229),
.Y(n_5809)
);

INVx3_ASAP7_75t_L g5810 ( 
.A(n_5024),
.Y(n_5810)
);

NAND2xp5_ASAP7_75t_L g5811 ( 
.A(n_4912),
.B(n_4229),
.Y(n_5811)
);

HB1xp67_ASAP7_75t_L g5812 ( 
.A(n_5266),
.Y(n_5812)
);

AND2x2_ASAP7_75t_L g5813 ( 
.A(n_4790),
.B(n_4231),
.Y(n_5813)
);

NAND2xp5_ASAP7_75t_L g5814 ( 
.A(n_4912),
.B(n_4362),
.Y(n_5814)
);

INVx1_ASAP7_75t_L g5815 ( 
.A(n_5045),
.Y(n_5815)
);

HB1xp67_ASAP7_75t_L g5816 ( 
.A(n_5301),
.Y(n_5816)
);

BUFx2_ASAP7_75t_L g5817 ( 
.A(n_4812),
.Y(n_5817)
);

INVx3_ASAP7_75t_L g5818 ( 
.A(n_5024),
.Y(n_5818)
);

INVx2_ASAP7_75t_L g5819 ( 
.A(n_5000),
.Y(n_5819)
);

HB1xp67_ASAP7_75t_L g5820 ( 
.A(n_5321),
.Y(n_5820)
);

INVx2_ASAP7_75t_L g5821 ( 
.A(n_5000),
.Y(n_5821)
);

INVx2_ASAP7_75t_L g5822 ( 
.A(n_5000),
.Y(n_5822)
);

OAI21x1_ASAP7_75t_L g5823 ( 
.A1(n_4779),
.A2(n_4598),
.B(n_4462),
.Y(n_5823)
);

INVx3_ASAP7_75t_L g5824 ( 
.A(n_5121),
.Y(n_5824)
);

INVx1_ASAP7_75t_L g5825 ( 
.A(n_5048),
.Y(n_5825)
);

INVx1_ASAP7_75t_L g5826 ( 
.A(n_5048),
.Y(n_5826)
);

INVx1_ASAP7_75t_L g5827 ( 
.A(n_5052),
.Y(n_5827)
);

INVx1_ASAP7_75t_L g5828 ( 
.A(n_5052),
.Y(n_5828)
);

OR2x6_ASAP7_75t_L g5829 ( 
.A(n_4969),
.B(n_4160),
.Y(n_5829)
);

INVx2_ASAP7_75t_L g5830 ( 
.A(n_5005),
.Y(n_5830)
);

AND2x2_ASAP7_75t_L g5831 ( 
.A(n_4699),
.B(n_4705),
.Y(n_5831)
);

OAI21xp5_ASAP7_75t_L g5832 ( 
.A1(n_5360),
.A2(n_4638),
.B(n_4659),
.Y(n_5832)
);

INVx1_ASAP7_75t_L g5833 ( 
.A(n_5053),
.Y(n_5833)
);

OA21x2_ASAP7_75t_L g5834 ( 
.A1(n_4828),
.A2(n_4200),
.B(n_4197),
.Y(n_5834)
);

INVx1_ASAP7_75t_L g5835 ( 
.A(n_5053),
.Y(n_5835)
);

NAND2x1p5_ASAP7_75t_L g5836 ( 
.A(n_5319),
.B(n_4647),
.Y(n_5836)
);

INVx2_ASAP7_75t_L g5837 ( 
.A(n_5005),
.Y(n_5837)
);

AND2x4_ASAP7_75t_L g5838 ( 
.A(n_4852),
.B(n_4275),
.Y(n_5838)
);

OR2x6_ASAP7_75t_L g5839 ( 
.A(n_4969),
.B(n_4160),
.Y(n_5839)
);

HB1xp67_ASAP7_75t_L g5840 ( 
.A(n_4772),
.Y(n_5840)
);

BUFx3_ASAP7_75t_L g5841 ( 
.A(n_4901),
.Y(n_5841)
);

AOI22xp5_ASAP7_75t_L g5842 ( 
.A1(n_4949),
.A2(n_5141),
.B1(n_4844),
.B2(n_4690),
.Y(n_5842)
);

INVx1_ASAP7_75t_L g5843 ( 
.A(n_5054),
.Y(n_5843)
);

INVx1_ASAP7_75t_L g5844 ( 
.A(n_5054),
.Y(n_5844)
);

INVx1_ASAP7_75t_L g5845 ( 
.A(n_5057),
.Y(n_5845)
);

INVx1_ASAP7_75t_L g5846 ( 
.A(n_5057),
.Y(n_5846)
);

AND2x2_ASAP7_75t_L g5847 ( 
.A(n_4707),
.B(n_4275),
.Y(n_5847)
);

NAND2xp5_ASAP7_75t_L g5848 ( 
.A(n_4921),
.B(n_4370),
.Y(n_5848)
);

NAND2xp5_ASAP7_75t_L g5849 ( 
.A(n_4921),
.B(n_4370),
.Y(n_5849)
);

AOI22xp5_ASAP7_75t_L g5850 ( 
.A1(n_5141),
.A2(n_4477),
.B1(n_4344),
.B2(n_4225),
.Y(n_5850)
);

INVx1_ASAP7_75t_L g5851 ( 
.A(n_5066),
.Y(n_5851)
);

INVx1_ASAP7_75t_L g5852 ( 
.A(n_5066),
.Y(n_5852)
);

AND2x2_ASAP7_75t_L g5853 ( 
.A(n_4785),
.B(n_4275),
.Y(n_5853)
);

INVx1_ASAP7_75t_L g5854 ( 
.A(n_5075),
.Y(n_5854)
);

AND2x4_ASAP7_75t_L g5855 ( 
.A(n_4852),
.B(n_4275),
.Y(n_5855)
);

INVx1_ASAP7_75t_L g5856 ( 
.A(n_5075),
.Y(n_5856)
);

AND2x2_ASAP7_75t_L g5857 ( 
.A(n_4785),
.B(n_4322),
.Y(n_5857)
);

INVxp67_ASAP7_75t_L g5858 ( 
.A(n_5149),
.Y(n_5858)
);

AO21x2_ASAP7_75t_L g5859 ( 
.A1(n_5331),
.A2(n_4423),
.B(n_4448),
.Y(n_5859)
);

INVx2_ASAP7_75t_L g5860 ( 
.A(n_5005),
.Y(n_5860)
);

BUFx2_ASAP7_75t_L g5861 ( 
.A(n_5121),
.Y(n_5861)
);

AOI22xp33_ASAP7_75t_SL g5862 ( 
.A1(n_4690),
.A2(n_4180),
.B1(n_4205),
.B2(n_4225),
.Y(n_5862)
);

INVx2_ASAP7_75t_L g5863 ( 
.A(n_5007),
.Y(n_5863)
);

INVx1_ASAP7_75t_L g5864 ( 
.A(n_5077),
.Y(n_5864)
);

AND2x2_ASAP7_75t_L g5865 ( 
.A(n_4800),
.B(n_4322),
.Y(n_5865)
);

INVx1_ASAP7_75t_L g5866 ( 
.A(n_5077),
.Y(n_5866)
);

HB1xp67_ASAP7_75t_L g5867 ( 
.A(n_4772),
.Y(n_5867)
);

AO21x2_ASAP7_75t_L g5868 ( 
.A1(n_5339),
.A2(n_4448),
.B(n_4424),
.Y(n_5868)
);

OAI21x1_ASAP7_75t_L g5869 ( 
.A1(n_4779),
.A2(n_4462),
.B(n_4459),
.Y(n_5869)
);

INVx1_ASAP7_75t_L g5870 ( 
.A(n_5083),
.Y(n_5870)
);

INVx1_ASAP7_75t_L g5871 ( 
.A(n_5083),
.Y(n_5871)
);

INVx1_ASAP7_75t_L g5872 ( 
.A(n_5087),
.Y(n_5872)
);

INVx1_ASAP7_75t_L g5873 ( 
.A(n_5087),
.Y(n_5873)
);

INVx2_ASAP7_75t_L g5874 ( 
.A(n_5007),
.Y(n_5874)
);

INVx1_ASAP7_75t_L g5875 ( 
.A(n_5095),
.Y(n_5875)
);

INVx1_ASAP7_75t_L g5876 ( 
.A(n_5095),
.Y(n_5876)
);

BUFx3_ASAP7_75t_L g5877 ( 
.A(n_4750),
.Y(n_5877)
);

BUFx2_ASAP7_75t_L g5878 ( 
.A(n_5121),
.Y(n_5878)
);

BUFx4f_ASAP7_75t_SL g5879 ( 
.A(n_4750),
.Y(n_5879)
);

OAI21x1_ASAP7_75t_L g5880 ( 
.A1(n_5110),
.A2(n_4474),
.B(n_4459),
.Y(n_5880)
);

HB1xp67_ASAP7_75t_L g5881 ( 
.A(n_4778),
.Y(n_5881)
);

OAI21x1_ASAP7_75t_L g5882 ( 
.A1(n_5110),
.A2(n_4474),
.B(n_4459),
.Y(n_5882)
);

INVx2_ASAP7_75t_L g5883 ( 
.A(n_5007),
.Y(n_5883)
);

BUFx3_ASAP7_75t_L g5884 ( 
.A(n_4750),
.Y(n_5884)
);

INVx1_ASAP7_75t_L g5885 ( 
.A(n_5100),
.Y(n_5885)
);

INVx1_ASAP7_75t_L g5886 ( 
.A(n_5100),
.Y(n_5886)
);

INVx1_ASAP7_75t_L g5887 ( 
.A(n_5101),
.Y(n_5887)
);

INVx1_ASAP7_75t_L g5888 ( 
.A(n_5101),
.Y(n_5888)
);

INVx2_ASAP7_75t_L g5889 ( 
.A(n_5008),
.Y(n_5889)
);

INVx2_ASAP7_75t_L g5890 ( 
.A(n_5008),
.Y(n_5890)
);

BUFx2_ASAP7_75t_L g5891 ( 
.A(n_5121),
.Y(n_5891)
);

INVx1_ASAP7_75t_L g5892 ( 
.A(n_5117),
.Y(n_5892)
);

INVx1_ASAP7_75t_L g5893 ( 
.A(n_5117),
.Y(n_5893)
);

INVx1_ASAP7_75t_L g5894 ( 
.A(n_5118),
.Y(n_5894)
);

AND2x4_ASAP7_75t_L g5895 ( 
.A(n_5055),
.B(n_4323),
.Y(n_5895)
);

INVx2_ASAP7_75t_L g5896 ( 
.A(n_5008),
.Y(n_5896)
);

HB1xp67_ASAP7_75t_L g5897 ( 
.A(n_4778),
.Y(n_5897)
);

OAI22xp33_ASAP7_75t_SL g5898 ( 
.A1(n_4672),
.A2(n_4565),
.B1(n_4590),
.B2(n_4589),
.Y(n_5898)
);

INVx1_ASAP7_75t_L g5899 ( 
.A(n_5118),
.Y(n_5899)
);

INVx2_ASAP7_75t_L g5900 ( 
.A(n_5023),
.Y(n_5900)
);

INVx2_ASAP7_75t_L g5901 ( 
.A(n_5023),
.Y(n_5901)
);

INVx2_ASAP7_75t_L g5902 ( 
.A(n_5023),
.Y(n_5902)
);

AO21x2_ASAP7_75t_L g5903 ( 
.A1(n_5339),
.A2(n_4424),
.B(n_4237),
.Y(n_5903)
);

AOI22xp33_ASAP7_75t_L g5904 ( 
.A1(n_4690),
.A2(n_4228),
.B1(n_4579),
.B2(n_4314),
.Y(n_5904)
);

NOR2xp33_ASAP7_75t_L g5905 ( 
.A(n_4805),
.B(n_4895),
.Y(n_5905)
);

INVx2_ASAP7_75t_L g5906 ( 
.A(n_5028),
.Y(n_5906)
);

INVx1_ASAP7_75t_L g5907 ( 
.A(n_5129),
.Y(n_5907)
);

INVx2_ASAP7_75t_L g5908 ( 
.A(n_5028),
.Y(n_5908)
);

OAI21xp5_ASAP7_75t_L g5909 ( 
.A1(n_4844),
.A2(n_4638),
.B(n_4659),
.Y(n_5909)
);

INVx2_ASAP7_75t_L g5910 ( 
.A(n_5028),
.Y(n_5910)
);

INVx2_ASAP7_75t_L g5911 ( 
.A(n_5031),
.Y(n_5911)
);

AND2x4_ASAP7_75t_L g5912 ( 
.A(n_5055),
.B(n_4323),
.Y(n_5912)
);

INVx3_ASAP7_75t_L g5913 ( 
.A(n_5130),
.Y(n_5913)
);

INVx1_ASAP7_75t_L g5914 ( 
.A(n_5129),
.Y(n_5914)
);

INVx1_ASAP7_75t_L g5915 ( 
.A(n_5140),
.Y(n_5915)
);

INVx1_ASAP7_75t_L g5916 ( 
.A(n_5140),
.Y(n_5916)
);

AND2x2_ASAP7_75t_L g5917 ( 
.A(n_4800),
.B(n_4322),
.Y(n_5917)
);

INVx2_ASAP7_75t_L g5918 ( 
.A(n_5031),
.Y(n_5918)
);

AOI21xp5_ASAP7_75t_L g5919 ( 
.A1(n_5195),
.A2(n_4648),
.B(n_4640),
.Y(n_5919)
);

INVx2_ASAP7_75t_SL g5920 ( 
.A(n_4969),
.Y(n_5920)
);

INVx3_ASAP7_75t_L g5921 ( 
.A(n_5130),
.Y(n_5921)
);

HB1xp67_ASAP7_75t_L g5922 ( 
.A(n_4872),
.Y(n_5922)
);

AND2x2_ASAP7_75t_L g5923 ( 
.A(n_4804),
.B(n_4873),
.Y(n_5923)
);

INVx2_ASAP7_75t_L g5924 ( 
.A(n_5031),
.Y(n_5924)
);

INVx1_ASAP7_75t_L g5925 ( 
.A(n_5144),
.Y(n_5925)
);

INVx1_ASAP7_75t_L g5926 ( 
.A(n_5144),
.Y(n_5926)
);

AOI21xp33_ASAP7_75t_L g5927 ( 
.A1(n_4671),
.A2(n_4344),
.B(n_4521),
.Y(n_5927)
);

INVx2_ASAP7_75t_L g5928 ( 
.A(n_5034),
.Y(n_5928)
);

INVx2_ASAP7_75t_L g5929 ( 
.A(n_5034),
.Y(n_5929)
);

INVx1_ASAP7_75t_L g5930 ( 
.A(n_5148),
.Y(n_5930)
);

INVxp67_ASAP7_75t_L g5931 ( 
.A(n_4998),
.Y(n_5931)
);

AND2x2_ASAP7_75t_L g5932 ( 
.A(n_4804),
.B(n_4322),
.Y(n_5932)
);

OAI22xp33_ASAP7_75t_L g5933 ( 
.A1(n_4959),
.A2(n_4371),
.B1(n_4181),
.B2(n_4168),
.Y(n_5933)
);

OAI21x1_ASAP7_75t_L g5934 ( 
.A1(n_4789),
.A2(n_4476),
.B(n_4474),
.Y(n_5934)
);

INVx1_ASAP7_75t_L g5935 ( 
.A(n_5148),
.Y(n_5935)
);

INVx4_ASAP7_75t_L g5936 ( 
.A(n_4794),
.Y(n_5936)
);

INVx2_ASAP7_75t_L g5937 ( 
.A(n_5034),
.Y(n_5937)
);

NAND2xp5_ASAP7_75t_L g5938 ( 
.A(n_4941),
.B(n_4407),
.Y(n_5938)
);

OAI21x1_ASAP7_75t_L g5939 ( 
.A1(n_4789),
.A2(n_4476),
.B(n_4400),
.Y(n_5939)
);

INVx2_ASAP7_75t_SL g5940 ( 
.A(n_5012),
.Y(n_5940)
);

NAND2xp5_ASAP7_75t_L g5941 ( 
.A(n_4941),
.B(n_4945),
.Y(n_5941)
);

INVx1_ASAP7_75t_L g5942 ( 
.A(n_5161),
.Y(n_5942)
);

INVxp67_ASAP7_75t_SL g5943 ( 
.A(n_4672),
.Y(n_5943)
);

BUFx3_ASAP7_75t_L g5944 ( 
.A(n_5239),
.Y(n_5944)
);

OAI21x1_ASAP7_75t_L g5945 ( 
.A1(n_4952),
.A2(n_4476),
.B(n_4400),
.Y(n_5945)
);

INVx2_ASAP7_75t_L g5946 ( 
.A(n_5041),
.Y(n_5946)
);

BUFx3_ASAP7_75t_L g5947 ( 
.A(n_5239),
.Y(n_5947)
);

INVx1_ASAP7_75t_L g5948 ( 
.A(n_5161),
.Y(n_5948)
);

INVx2_ASAP7_75t_L g5949 ( 
.A(n_5041),
.Y(n_5949)
);

INVx1_ASAP7_75t_L g5950 ( 
.A(n_5162),
.Y(n_5950)
);

INVx2_ASAP7_75t_L g5951 ( 
.A(n_5041),
.Y(n_5951)
);

HB1xp67_ASAP7_75t_L g5952 ( 
.A(n_4872),
.Y(n_5952)
);

INVx1_ASAP7_75t_L g5953 ( 
.A(n_5162),
.Y(n_5953)
);

INVx1_ASAP7_75t_L g5954 ( 
.A(n_5166),
.Y(n_5954)
);

AND2x2_ASAP7_75t_L g5955 ( 
.A(n_4873),
.B(n_4323),
.Y(n_5955)
);

INVx2_ASAP7_75t_L g5956 ( 
.A(n_5056),
.Y(n_5956)
);

INVx1_ASAP7_75t_L g5957 ( 
.A(n_5166),
.Y(n_5957)
);

OAI21x1_ASAP7_75t_L g5958 ( 
.A1(n_4952),
.A2(n_4400),
.B(n_4409),
.Y(n_5958)
);

INVx1_ASAP7_75t_L g5959 ( 
.A(n_5173),
.Y(n_5959)
);

OR2x2_ASAP7_75t_L g5960 ( 
.A(n_4909),
.B(n_4407),
.Y(n_5960)
);

INVx1_ASAP7_75t_L g5961 ( 
.A(n_5173),
.Y(n_5961)
);

INVx1_ASAP7_75t_L g5962 ( 
.A(n_5177),
.Y(n_5962)
);

BUFx3_ASAP7_75t_L g5963 ( 
.A(n_5239),
.Y(n_5963)
);

INVx6_ASAP7_75t_L g5964 ( 
.A(n_4781),
.Y(n_5964)
);

INVx1_ASAP7_75t_L g5965 ( 
.A(n_5177),
.Y(n_5965)
);

INVx2_ASAP7_75t_L g5966 ( 
.A(n_5056),
.Y(n_5966)
);

BUFx3_ASAP7_75t_L g5967 ( 
.A(n_4923),
.Y(n_5967)
);

INVx1_ASAP7_75t_L g5968 ( 
.A(n_5178),
.Y(n_5968)
);

INVx1_ASAP7_75t_L g5969 ( 
.A(n_5178),
.Y(n_5969)
);

INVx1_ASAP7_75t_L g5970 ( 
.A(n_5179),
.Y(n_5970)
);

INVx3_ASAP7_75t_L g5971 ( 
.A(n_5130),
.Y(n_5971)
);

INVx1_ASAP7_75t_L g5972 ( 
.A(n_5179),
.Y(n_5972)
);

AND2x2_ASAP7_75t_L g5973 ( 
.A(n_4897),
.B(n_4323),
.Y(n_5973)
);

OR2x2_ASAP7_75t_L g5974 ( 
.A(n_4909),
.B(n_4667),
.Y(n_5974)
);

BUFx6f_ASAP7_75t_L g5975 ( 
.A(n_4794),
.Y(n_5975)
);

INVx2_ASAP7_75t_SL g5976 ( 
.A(n_5012),
.Y(n_5976)
);

INVx1_ASAP7_75t_L g5977 ( 
.A(n_5186),
.Y(n_5977)
);

OR2x2_ASAP7_75t_L g5978 ( 
.A(n_5243),
.B(n_4667),
.Y(n_5978)
);

INVx1_ASAP7_75t_L g5979 ( 
.A(n_5186),
.Y(n_5979)
);

AND2x2_ASAP7_75t_L g5980 ( 
.A(n_4897),
.B(n_4331),
.Y(n_5980)
);

OAI21xp5_ASAP7_75t_L g5981 ( 
.A1(n_4959),
.A2(n_4390),
.B(n_4521),
.Y(n_5981)
);

INVx1_ASAP7_75t_L g5982 ( 
.A(n_5196),
.Y(n_5982)
);

AOI21x1_ASAP7_75t_L g5983 ( 
.A1(n_5086),
.A2(n_4218),
.B(n_4217),
.Y(n_5983)
);

INVx4_ASAP7_75t_L g5984 ( 
.A(n_4794),
.Y(n_5984)
);

HB1xp67_ASAP7_75t_L g5985 ( 
.A(n_4947),
.Y(n_5985)
);

INVx1_ASAP7_75t_L g5986 ( 
.A(n_5196),
.Y(n_5986)
);

INVx1_ASAP7_75t_L g5987 ( 
.A(n_5197),
.Y(n_5987)
);

INVx1_ASAP7_75t_L g5988 ( 
.A(n_5197),
.Y(n_5988)
);

NAND2xp5_ASAP7_75t_SL g5989 ( 
.A(n_4932),
.B(n_5292),
.Y(n_5989)
);

INVxp33_ASAP7_75t_L g5990 ( 
.A(n_5068),
.Y(n_5990)
);

INVx3_ASAP7_75t_L g5991 ( 
.A(n_5130),
.Y(n_5991)
);

INVx2_ASAP7_75t_SL g5992 ( 
.A(n_5012),
.Y(n_5992)
);

INVx1_ASAP7_75t_L g5993 ( 
.A(n_5206),
.Y(n_5993)
);

CKINVDCx5p33_ASAP7_75t_R g5994 ( 
.A(n_4706),
.Y(n_5994)
);

BUFx12f_ASAP7_75t_L g5995 ( 
.A(n_4848),
.Y(n_5995)
);

AOI22xp33_ASAP7_75t_L g5996 ( 
.A1(n_4725),
.A2(n_4228),
.B1(n_4579),
.B2(n_4314),
.Y(n_5996)
);

INVx1_ASAP7_75t_L g5997 ( 
.A(n_5206),
.Y(n_5997)
);

BUFx2_ASAP7_75t_L g5998 ( 
.A(n_5006),
.Y(n_5998)
);

OA21x2_ASAP7_75t_L g5999 ( 
.A1(n_4828),
.A2(n_4200),
.B(n_4197),
.Y(n_5999)
);

AND2x2_ASAP7_75t_L g6000 ( 
.A(n_4911),
.B(n_4331),
.Y(n_6000)
);

HB1xp67_ASAP7_75t_L g6001 ( 
.A(n_4947),
.Y(n_6001)
);

AO21x2_ASAP7_75t_L g6002 ( 
.A1(n_5339),
.A2(n_4237),
.B(n_4233),
.Y(n_6002)
);

AND2x4_ASAP7_75t_L g6003 ( 
.A(n_5055),
.B(n_5090),
.Y(n_6003)
);

BUFx3_ASAP7_75t_L g6004 ( 
.A(n_4997),
.Y(n_6004)
);

OAI22xp5_ASAP7_75t_SL g6005 ( 
.A1(n_4932),
.A2(n_3866),
.B1(n_3954),
.B2(n_3886),
.Y(n_6005)
);

HB1xp67_ASAP7_75t_L g6006 ( 
.A(n_5248),
.Y(n_6006)
);

INVx1_ASAP7_75t_L g6007 ( 
.A(n_5212),
.Y(n_6007)
);

INVx1_ASAP7_75t_L g6008 ( 
.A(n_5212),
.Y(n_6008)
);

INVx1_ASAP7_75t_L g6009 ( 
.A(n_5215),
.Y(n_6009)
);

INVx1_ASAP7_75t_L g6010 ( 
.A(n_5215),
.Y(n_6010)
);

INVx1_ASAP7_75t_L g6011 ( 
.A(n_5219),
.Y(n_6011)
);

INVx2_ASAP7_75t_SL g6012 ( 
.A(n_5012),
.Y(n_6012)
);

INVx1_ASAP7_75t_SL g6013 ( 
.A(n_5042),
.Y(n_6013)
);

AO21x2_ASAP7_75t_L g6014 ( 
.A1(n_5340),
.A2(n_4237),
.B(n_4233),
.Y(n_6014)
);

AND2x2_ASAP7_75t_L g6015 ( 
.A(n_5426),
.B(n_4973),
.Y(n_6015)
);

INVx3_ASAP7_75t_L g6016 ( 
.A(n_5418),
.Y(n_6016)
);

INVx1_ASAP7_75t_L g6017 ( 
.A(n_5384),
.Y(n_6017)
);

AO21x2_ASAP7_75t_L g6018 ( 
.A1(n_5634),
.A2(n_5152),
.B(n_5125),
.Y(n_6018)
);

INVx1_ASAP7_75t_L g6019 ( 
.A(n_5384),
.Y(n_6019)
);

INVx1_ASAP7_75t_L g6020 ( 
.A(n_5417),
.Y(n_6020)
);

AND2x2_ASAP7_75t_L g6021 ( 
.A(n_5426),
.B(n_5431),
.Y(n_6021)
);

AND2x2_ASAP7_75t_L g6022 ( 
.A(n_5431),
.B(n_4973),
.Y(n_6022)
);

INVx2_ASAP7_75t_L g6023 ( 
.A(n_5516),
.Y(n_6023)
);

INVx2_ASAP7_75t_SL g6024 ( 
.A(n_5502),
.Y(n_6024)
);

INVx1_ASAP7_75t_L g6025 ( 
.A(n_5417),
.Y(n_6025)
);

HB1xp67_ASAP7_75t_L g6026 ( 
.A(n_5840),
.Y(n_6026)
);

AND2x2_ASAP7_75t_L g6027 ( 
.A(n_5998),
.B(n_5050),
.Y(n_6027)
);

INVx3_ASAP7_75t_L g6028 ( 
.A(n_5418),
.Y(n_6028)
);

AND2x2_ASAP7_75t_L g6029 ( 
.A(n_5998),
.B(n_5923),
.Y(n_6029)
);

INVx1_ASAP7_75t_L g6030 ( 
.A(n_5419),
.Y(n_6030)
);

INVx1_ASAP7_75t_L g6031 ( 
.A(n_5419),
.Y(n_6031)
);

OR2x2_ASAP7_75t_L g6032 ( 
.A(n_5558),
.B(n_4787),
.Y(n_6032)
);

INVx1_ASAP7_75t_L g6033 ( 
.A(n_5438),
.Y(n_6033)
);

INVx1_ASAP7_75t_L g6034 ( 
.A(n_5372),
.Y(n_6034)
);

INVx2_ASAP7_75t_L g6035 ( 
.A(n_5516),
.Y(n_6035)
);

INVx1_ASAP7_75t_L g6036 ( 
.A(n_5372),
.Y(n_6036)
);

INVxp67_ASAP7_75t_L g6037 ( 
.A(n_5802),
.Y(n_6037)
);

AND2x2_ASAP7_75t_L g6038 ( 
.A(n_5923),
.B(n_5050),
.Y(n_6038)
);

INVx2_ASAP7_75t_L g6039 ( 
.A(n_5516),
.Y(n_6039)
);

INVx1_ASAP7_75t_L g6040 ( 
.A(n_5373),
.Y(n_6040)
);

INVx2_ASAP7_75t_L g6041 ( 
.A(n_5516),
.Y(n_6041)
);

AOI21xp5_ASAP7_75t_L g6042 ( 
.A1(n_5416),
.A2(n_5195),
.B(n_4787),
.Y(n_6042)
);

OR2x2_ASAP7_75t_L g6043 ( 
.A(n_5388),
.B(n_5243),
.Y(n_6043)
);

BUFx2_ASAP7_75t_L g6044 ( 
.A(n_5403),
.Y(n_6044)
);

AND2x2_ASAP7_75t_L g6045 ( 
.A(n_5441),
.B(n_5292),
.Y(n_6045)
);

OAI21x1_ASAP7_75t_L g6046 ( 
.A1(n_5721),
.A2(n_5036),
.B(n_5102),
.Y(n_6046)
);

BUFx2_ASAP7_75t_L g6047 ( 
.A(n_5403),
.Y(n_6047)
);

INVx2_ASAP7_75t_L g6048 ( 
.A(n_5516),
.Y(n_6048)
);

INVx2_ASAP7_75t_L g6049 ( 
.A(n_5376),
.Y(n_6049)
);

INVx1_ASAP7_75t_L g6050 ( 
.A(n_5448),
.Y(n_6050)
);

OR2x2_ASAP7_75t_L g6051 ( 
.A(n_5388),
.B(n_5285),
.Y(n_6051)
);

OR2x2_ASAP7_75t_L g6052 ( 
.A(n_5400),
.B(n_5285),
.Y(n_6052)
);

HB1xp67_ASAP7_75t_L g6053 ( 
.A(n_5867),
.Y(n_6053)
);

AND2x2_ASAP7_75t_L g6054 ( 
.A(n_5441),
.B(n_4720),
.Y(n_6054)
);

INVx1_ASAP7_75t_L g6055 ( 
.A(n_5411),
.Y(n_6055)
);

INVx1_ASAP7_75t_L g6056 ( 
.A(n_5411),
.Y(n_6056)
);

INVx1_ASAP7_75t_L g6057 ( 
.A(n_5424),
.Y(n_6057)
);

BUFx6f_ASAP7_75t_L g6058 ( 
.A(n_5385),
.Y(n_6058)
);

INVx2_ASAP7_75t_L g6059 ( 
.A(n_5376),
.Y(n_6059)
);

OR2x6_ASAP7_75t_L g6060 ( 
.A(n_5627),
.B(n_5012),
.Y(n_6060)
);

INVx1_ASAP7_75t_L g6061 ( 
.A(n_5424),
.Y(n_6061)
);

HB1xp67_ASAP7_75t_L g6062 ( 
.A(n_5881),
.Y(n_6062)
);

AND2x2_ASAP7_75t_L g6063 ( 
.A(n_5480),
.B(n_4720),
.Y(n_6063)
);

HB1xp67_ASAP7_75t_L g6064 ( 
.A(n_5897),
.Y(n_6064)
);

INVx3_ASAP7_75t_L g6065 ( 
.A(n_5564),
.Y(n_6065)
);

INVx1_ASAP7_75t_L g6066 ( 
.A(n_5444),
.Y(n_6066)
);

NAND2xp5_ASAP7_75t_L g6067 ( 
.A(n_5374),
.B(n_4945),
.Y(n_6067)
);

AO31x2_ASAP7_75t_L g6068 ( 
.A1(n_5593),
.A2(n_5348),
.A3(n_5340),
.B(n_4716),
.Y(n_6068)
);

OR2x2_ASAP7_75t_L g6069 ( 
.A(n_5400),
.B(n_5043),
.Y(n_6069)
);

INVx1_ASAP7_75t_L g6070 ( 
.A(n_5378),
.Y(n_6070)
);

AND2x2_ASAP7_75t_L g6071 ( 
.A(n_5480),
.B(n_4720),
.Y(n_6071)
);

INVx1_ASAP7_75t_L g6072 ( 
.A(n_5378),
.Y(n_6072)
);

AND2x2_ASAP7_75t_L g6073 ( 
.A(n_5507),
.B(n_4720),
.Y(n_6073)
);

INVx1_ASAP7_75t_L g6074 ( 
.A(n_5373),
.Y(n_6074)
);

INVx2_ASAP7_75t_SL g6075 ( 
.A(n_5502),
.Y(n_6075)
);

INVx2_ASAP7_75t_L g6076 ( 
.A(n_5376),
.Y(n_6076)
);

INVx1_ASAP7_75t_L g6077 ( 
.A(n_5375),
.Y(n_6077)
);

OR2x2_ASAP7_75t_L g6078 ( 
.A(n_5763),
.B(n_5043),
.Y(n_6078)
);

AND2x2_ASAP7_75t_L g6079 ( 
.A(n_5507),
.B(n_4724),
.Y(n_6079)
);

INVx2_ASAP7_75t_L g6080 ( 
.A(n_5447),
.Y(n_6080)
);

AO21x2_ASAP7_75t_L g6081 ( 
.A1(n_5639),
.A2(n_5152),
.B(n_5125),
.Y(n_6081)
);

HB1xp67_ASAP7_75t_L g6082 ( 
.A(n_5922),
.Y(n_6082)
);

OAI21x1_ASAP7_75t_L g6083 ( 
.A1(n_5721),
.A2(n_5036),
.B(n_5102),
.Y(n_6083)
);

OA21x2_ASAP7_75t_L g6084 ( 
.A1(n_5512),
.A2(n_5152),
.B(n_5125),
.Y(n_6084)
);

INVx1_ASAP7_75t_L g6085 ( 
.A(n_5391),
.Y(n_6085)
);

INVxp67_ASAP7_75t_SL g6086 ( 
.A(n_5593),
.Y(n_6086)
);

INVx2_ASAP7_75t_L g6087 ( 
.A(n_5447),
.Y(n_6087)
);

OA21x2_ASAP7_75t_L g6088 ( 
.A1(n_5460),
.A2(n_5167),
.B(n_5155),
.Y(n_6088)
);

AND2x2_ASAP7_75t_L g6089 ( 
.A(n_5589),
.B(n_4724),
.Y(n_6089)
);

AOI22xp33_ASAP7_75t_L g6090 ( 
.A1(n_5508),
.A2(n_5369),
.B1(n_5540),
.B2(n_5488),
.Y(n_6090)
);

INVx2_ASAP7_75t_L g6091 ( 
.A(n_5447),
.Y(n_6091)
);

INVx1_ASAP7_75t_L g6092 ( 
.A(n_5391),
.Y(n_6092)
);

OA21x2_ASAP7_75t_L g6093 ( 
.A1(n_5393),
.A2(n_5513),
.B(n_5717),
.Y(n_6093)
);

INVx2_ASAP7_75t_L g6094 ( 
.A(n_5447),
.Y(n_6094)
);

HB1xp67_ASAP7_75t_L g6095 ( 
.A(n_5952),
.Y(n_6095)
);

BUFx3_ASAP7_75t_L g6096 ( 
.A(n_5645),
.Y(n_6096)
);

AO21x2_ASAP7_75t_L g6097 ( 
.A1(n_5842),
.A2(n_5167),
.B(n_5155),
.Y(n_6097)
);

AO31x2_ASAP7_75t_L g6098 ( 
.A1(n_5508),
.A2(n_5348),
.A3(n_5340),
.B(n_4716),
.Y(n_6098)
);

OR2x2_ASAP7_75t_L g6099 ( 
.A(n_5804),
.B(n_5103),
.Y(n_6099)
);

INVx1_ASAP7_75t_L g6100 ( 
.A(n_5423),
.Y(n_6100)
);

OR2x6_ASAP7_75t_L g6101 ( 
.A(n_5627),
.B(n_5051),
.Y(n_6101)
);

OA21x2_ASAP7_75t_L g6102 ( 
.A1(n_5934),
.A2(n_5167),
.B(n_5155),
.Y(n_6102)
);

INVx2_ASAP7_75t_L g6103 ( 
.A(n_5983),
.Y(n_6103)
);

AND2x2_ASAP7_75t_L g6104 ( 
.A(n_5589),
.B(n_4724),
.Y(n_6104)
);

INVx2_ASAP7_75t_L g6105 ( 
.A(n_5983),
.Y(n_6105)
);

INVx2_ASAP7_75t_L g6106 ( 
.A(n_5412),
.Y(n_6106)
);

OAI21x1_ASAP7_75t_L g6107 ( 
.A1(n_5797),
.A2(n_5146),
.B(n_5102),
.Y(n_6107)
);

AND2x2_ASAP7_75t_L g6108 ( 
.A(n_5617),
.B(n_4724),
.Y(n_6108)
);

INVx1_ASAP7_75t_L g6109 ( 
.A(n_5423),
.Y(n_6109)
);

INVx2_ASAP7_75t_L g6110 ( 
.A(n_5412),
.Y(n_6110)
);

INVx1_ASAP7_75t_L g6111 ( 
.A(n_5444),
.Y(n_6111)
);

INVxp67_ASAP7_75t_SL g6112 ( 
.A(n_5677),
.Y(n_6112)
);

INVx2_ASAP7_75t_L g6113 ( 
.A(n_5412),
.Y(n_6113)
);

INVx1_ASAP7_75t_L g6114 ( 
.A(n_5427),
.Y(n_6114)
);

AOI21xp5_ASAP7_75t_SL g6115 ( 
.A1(n_5627),
.A2(n_4404),
.B(n_5151),
.Y(n_6115)
);

AO21x2_ASAP7_75t_L g6116 ( 
.A1(n_5842),
.A2(n_5927),
.B(n_5443),
.Y(n_6116)
);

INVx1_ASAP7_75t_L g6117 ( 
.A(n_5427),
.Y(n_6117)
);

AND2x2_ASAP7_75t_L g6118 ( 
.A(n_5617),
.B(n_4777),
.Y(n_6118)
);

INVx1_ASAP7_75t_L g6119 ( 
.A(n_5428),
.Y(n_6119)
);

OAI22xp5_ASAP7_75t_L g6120 ( 
.A1(n_5607),
.A2(n_5333),
.B1(n_5265),
.B2(n_5267),
.Y(n_6120)
);

INVx2_ASAP7_75t_L g6121 ( 
.A(n_5439),
.Y(n_6121)
);

NOR2xp33_ASAP7_75t_L g6122 ( 
.A(n_5385),
.B(n_5042),
.Y(n_6122)
);

OR2x2_ASAP7_75t_L g6123 ( 
.A(n_5941),
.B(n_5103),
.Y(n_6123)
);

BUFx3_ASAP7_75t_L g6124 ( 
.A(n_5645),
.Y(n_6124)
);

OR2x6_ASAP7_75t_L g6125 ( 
.A(n_5627),
.B(n_5051),
.Y(n_6125)
);

INVx1_ASAP7_75t_L g6126 ( 
.A(n_5428),
.Y(n_6126)
);

BUFx2_ASAP7_75t_L g6127 ( 
.A(n_5403),
.Y(n_6127)
);

INVx2_ASAP7_75t_L g6128 ( 
.A(n_5439),
.Y(n_6128)
);

BUFx2_ASAP7_75t_L g6129 ( 
.A(n_5403),
.Y(n_6129)
);

INVx1_ASAP7_75t_L g6130 ( 
.A(n_5438),
.Y(n_6130)
);

INVx2_ASAP7_75t_L g6131 ( 
.A(n_5439),
.Y(n_6131)
);

OR2x2_ASAP7_75t_L g6132 ( 
.A(n_5811),
.B(n_5189),
.Y(n_6132)
);

INVx1_ASAP7_75t_L g6133 ( 
.A(n_5451),
.Y(n_6133)
);

INVx2_ASAP7_75t_L g6134 ( 
.A(n_5470),
.Y(n_6134)
);

BUFx2_ASAP7_75t_L g6135 ( 
.A(n_5403),
.Y(n_6135)
);

NAND2x1_ASAP7_75t_L g6136 ( 
.A(n_5564),
.B(n_5051),
.Y(n_6136)
);

BUFx6f_ASAP7_75t_L g6137 ( 
.A(n_5385),
.Y(n_6137)
);

INVx1_ASAP7_75t_L g6138 ( 
.A(n_5442),
.Y(n_6138)
);

INVx2_ASAP7_75t_L g6139 ( 
.A(n_5470),
.Y(n_6139)
);

INVx1_ASAP7_75t_L g6140 ( 
.A(n_5442),
.Y(n_6140)
);

INVx2_ASAP7_75t_L g6141 ( 
.A(n_5470),
.Y(n_6141)
);

OR2x2_ASAP7_75t_L g6142 ( 
.A(n_5539),
.B(n_5425),
.Y(n_6142)
);

INVx2_ASAP7_75t_L g6143 ( 
.A(n_5521),
.Y(n_6143)
);

INVx2_ASAP7_75t_L g6144 ( 
.A(n_5521),
.Y(n_6144)
);

INVx2_ASAP7_75t_L g6145 ( 
.A(n_5521),
.Y(n_6145)
);

AO21x2_ASAP7_75t_L g6146 ( 
.A1(n_5443),
.A2(n_5170),
.B(n_4832),
.Y(n_6146)
);

AOI22xp33_ASAP7_75t_L g6147 ( 
.A1(n_5369),
.A2(n_4725),
.B1(n_4876),
.B2(n_4688),
.Y(n_6147)
);

AO21x2_ASAP7_75t_L g6148 ( 
.A1(n_5729),
.A2(n_5170),
.B(n_4832),
.Y(n_6148)
);

INVx2_ASAP7_75t_L g6149 ( 
.A(n_5591),
.Y(n_6149)
);

AND2x2_ASAP7_75t_L g6150 ( 
.A(n_5618),
.B(n_4777),
.Y(n_6150)
);

INVx3_ASAP7_75t_L g6151 ( 
.A(n_5564),
.Y(n_6151)
);

HB1xp67_ASAP7_75t_L g6152 ( 
.A(n_5985),
.Y(n_6152)
);

BUFx2_ASAP7_75t_L g6153 ( 
.A(n_5608),
.Y(n_6153)
);

NOR2xp33_ASAP7_75t_L g6154 ( 
.A(n_5385),
.B(n_5154),
.Y(n_6154)
);

OAI222xp33_ASAP7_75t_L g6155 ( 
.A1(n_5670),
.A2(n_4688),
.B1(n_5190),
.B2(n_4981),
.C1(n_5353),
.C2(n_5295),
.Y(n_6155)
);

INVx1_ASAP7_75t_L g6156 ( 
.A(n_5446),
.Y(n_6156)
);

INVx1_ASAP7_75t_L g6157 ( 
.A(n_5446),
.Y(n_6157)
);

INVx1_ASAP7_75t_L g6158 ( 
.A(n_5448),
.Y(n_6158)
);

INVxp67_ASAP7_75t_L g6159 ( 
.A(n_5498),
.Y(n_6159)
);

NAND2xp5_ASAP7_75t_L g6160 ( 
.A(n_5546),
.B(n_4821),
.Y(n_6160)
);

INVx1_ASAP7_75t_SL g6161 ( 
.A(n_5498),
.Y(n_6161)
);

INVx3_ASAP7_75t_L g6162 ( 
.A(n_5564),
.Y(n_6162)
);

INVx2_ASAP7_75t_L g6163 ( 
.A(n_5591),
.Y(n_6163)
);

INVx3_ASAP7_75t_L g6164 ( 
.A(n_5601),
.Y(n_6164)
);

AND2x4_ASAP7_75t_L g6165 ( 
.A(n_5387),
.B(n_5006),
.Y(n_6165)
);

INVx1_ASAP7_75t_L g6166 ( 
.A(n_5484),
.Y(n_6166)
);

INVx4_ASAP7_75t_SL g6167 ( 
.A(n_5502),
.Y(n_6167)
);

NAND2xp5_ASAP7_75t_L g6168 ( 
.A(n_5687),
.B(n_4821),
.Y(n_6168)
);

INVx1_ASAP7_75t_L g6169 ( 
.A(n_5484),
.Y(n_6169)
);

INVx1_ASAP7_75t_L g6170 ( 
.A(n_5533),
.Y(n_6170)
);

INVx2_ASAP7_75t_L g6171 ( 
.A(n_5591),
.Y(n_6171)
);

INVx2_ASAP7_75t_L g6172 ( 
.A(n_5604),
.Y(n_6172)
);

INVx2_ASAP7_75t_L g6173 ( 
.A(n_5604),
.Y(n_6173)
);

INVx2_ASAP7_75t_L g6174 ( 
.A(n_5604),
.Y(n_6174)
);

INVx1_ASAP7_75t_L g6175 ( 
.A(n_5533),
.Y(n_6175)
);

INVx2_ASAP7_75t_L g6176 ( 
.A(n_5797),
.Y(n_6176)
);

BUFx3_ASAP7_75t_L g6177 ( 
.A(n_5385),
.Y(n_6177)
);

INVx2_ASAP7_75t_L g6178 ( 
.A(n_6002),
.Y(n_6178)
);

INVx2_ASAP7_75t_L g6179 ( 
.A(n_6002),
.Y(n_6179)
);

AND2x2_ASAP7_75t_L g6180 ( 
.A(n_5618),
.B(n_4777),
.Y(n_6180)
);

INVx1_ASAP7_75t_SL g6181 ( 
.A(n_5472),
.Y(n_6181)
);

INVx1_ASAP7_75t_L g6182 ( 
.A(n_5450),
.Y(n_6182)
);

OA21x2_ASAP7_75t_L g6183 ( 
.A1(n_5934),
.A2(n_5532),
.B(n_5529),
.Y(n_6183)
);

INVx2_ASAP7_75t_L g6184 ( 
.A(n_6002),
.Y(n_6184)
);

INVx2_ASAP7_75t_L g6185 ( 
.A(n_6014),
.Y(n_6185)
);

INVx2_ASAP7_75t_L g6186 ( 
.A(n_6014),
.Y(n_6186)
);

AND2x2_ASAP7_75t_L g6187 ( 
.A(n_5661),
.B(n_4777),
.Y(n_6187)
);

INVx1_ASAP7_75t_SL g6188 ( 
.A(n_5489),
.Y(n_6188)
);

INVx2_ASAP7_75t_L g6189 ( 
.A(n_6014),
.Y(n_6189)
);

INVx2_ASAP7_75t_L g6190 ( 
.A(n_5556),
.Y(n_6190)
);

INVx2_ASAP7_75t_L g6191 ( 
.A(n_5556),
.Y(n_6191)
);

INVxp67_ASAP7_75t_L g6192 ( 
.A(n_5497),
.Y(n_6192)
);

INVx1_ASAP7_75t_L g6193 ( 
.A(n_5375),
.Y(n_6193)
);

INVx2_ASAP7_75t_L g6194 ( 
.A(n_5561),
.Y(n_6194)
);

OA21x2_ASAP7_75t_L g6195 ( 
.A1(n_5529),
.A2(n_5170),
.B(n_4832),
.Y(n_6195)
);

INVx1_ASAP7_75t_L g6196 ( 
.A(n_5383),
.Y(n_6196)
);

OR2x6_ASAP7_75t_L g6197 ( 
.A(n_5627),
.B(n_5051),
.Y(n_6197)
);

INVx2_ASAP7_75t_L g6198 ( 
.A(n_5561),
.Y(n_6198)
);

INVx1_ASAP7_75t_L g6199 ( 
.A(n_5383),
.Y(n_6199)
);

INVx1_ASAP7_75t_L g6200 ( 
.A(n_5396),
.Y(n_6200)
);

INVx1_ASAP7_75t_L g6201 ( 
.A(n_5396),
.Y(n_6201)
);

AND2x2_ASAP7_75t_L g6202 ( 
.A(n_5661),
.B(n_4911),
.Y(n_6202)
);

AO21x2_ASAP7_75t_L g6203 ( 
.A1(n_5779),
.A2(n_4677),
.B(n_4676),
.Y(n_6203)
);

INVx1_ASAP7_75t_L g6204 ( 
.A(n_5421),
.Y(n_6204)
);

AND2x2_ASAP7_75t_L g6205 ( 
.A(n_5392),
.B(n_4966),
.Y(n_6205)
);

INVx1_ASAP7_75t_L g6206 ( 
.A(n_5421),
.Y(n_6206)
);

INVx2_ASAP7_75t_L g6207 ( 
.A(n_5569),
.Y(n_6207)
);

INVx4_ASAP7_75t_L g6208 ( 
.A(n_5608),
.Y(n_6208)
);

HB1xp67_ASAP7_75t_L g6209 ( 
.A(n_6001),
.Y(n_6209)
);

INVx1_ASAP7_75t_L g6210 ( 
.A(n_5445),
.Y(n_6210)
);

OA21x2_ASAP7_75t_L g6211 ( 
.A1(n_5532),
.A2(n_5348),
.B(n_4763),
.Y(n_6211)
);

OAI21xp5_ASAP7_75t_L g6212 ( 
.A1(n_5578),
.A2(n_5241),
.B(n_5190),
.Y(n_6212)
);

AND2x2_ASAP7_75t_L g6213 ( 
.A(n_5392),
.B(n_4966),
.Y(n_6213)
);

AND2x2_ASAP7_75t_L g6214 ( 
.A(n_5394),
.B(n_5082),
.Y(n_6214)
);

INVx2_ASAP7_75t_L g6215 ( 
.A(n_5569),
.Y(n_6215)
);

INVx1_ASAP7_75t_L g6216 ( 
.A(n_5445),
.Y(n_6216)
);

AND2x4_ASAP7_75t_L g6217 ( 
.A(n_5387),
.B(n_5006),
.Y(n_6217)
);

AND2x2_ASAP7_75t_L g6218 ( 
.A(n_5394),
.B(n_5082),
.Y(n_6218)
);

INVx3_ASAP7_75t_L g6219 ( 
.A(n_5601),
.Y(n_6219)
);

INVx2_ASAP7_75t_L g6220 ( 
.A(n_5582),
.Y(n_6220)
);

AND2x2_ASAP7_75t_L g6221 ( 
.A(n_5397),
.B(n_4795),
.Y(n_6221)
);

OAI22xp5_ASAP7_75t_L g6222 ( 
.A1(n_5607),
.A2(n_5333),
.B1(n_5349),
.B2(n_5241),
.Y(n_6222)
);

INVx2_ASAP7_75t_L g6223 ( 
.A(n_5582),
.Y(n_6223)
);

OR2x6_ASAP7_75t_L g6224 ( 
.A(n_5829),
.B(n_5051),
.Y(n_6224)
);

INVx2_ASAP7_75t_L g6225 ( 
.A(n_5583),
.Y(n_6225)
);

INVx11_ASAP7_75t_L g6226 ( 
.A(n_5995),
.Y(n_6226)
);

BUFx6f_ASAP7_75t_L g6227 ( 
.A(n_5543),
.Y(n_6227)
);

OR2x2_ASAP7_75t_L g6228 ( 
.A(n_5425),
.B(n_5189),
.Y(n_6228)
);

HB1xp67_ASAP7_75t_L g6229 ( 
.A(n_5636),
.Y(n_6229)
);

AND2x4_ASAP7_75t_L g6230 ( 
.A(n_5387),
.B(n_5006),
.Y(n_6230)
);

INVx2_ASAP7_75t_L g6231 ( 
.A(n_5583),
.Y(n_6231)
);

INVx1_ASAP7_75t_L g6232 ( 
.A(n_5450),
.Y(n_6232)
);

HB1xp67_ASAP7_75t_L g6233 ( 
.A(n_5638),
.Y(n_6233)
);

INVx2_ASAP7_75t_L g6234 ( 
.A(n_5584),
.Y(n_6234)
);

AND2x2_ASAP7_75t_L g6235 ( 
.A(n_5397),
.B(n_4795),
.Y(n_6235)
);

AOI21x1_ASAP7_75t_L g6236 ( 
.A1(n_5684),
.A2(n_5107),
.B(n_5060),
.Y(n_6236)
);

OA222x2_ASAP7_75t_L g6237 ( 
.A1(n_5629),
.A2(n_4839),
.B1(n_4976),
.B2(n_4664),
.C1(n_5308),
.C2(n_4371),
.Y(n_6237)
);

INVx2_ASAP7_75t_L g6238 ( 
.A(n_5584),
.Y(n_6238)
);

INVx1_ASAP7_75t_L g6239 ( 
.A(n_5469),
.Y(n_6239)
);

AND2x2_ASAP7_75t_L g6240 ( 
.A(n_5404),
.B(n_4795),
.Y(n_6240)
);

AND2x2_ASAP7_75t_L g6241 ( 
.A(n_5404),
.B(n_5415),
.Y(n_6241)
);

AND2x2_ASAP7_75t_L g6242 ( 
.A(n_5415),
.B(n_4795),
.Y(n_6242)
);

INVx2_ASAP7_75t_L g6243 ( 
.A(n_5586),
.Y(n_6243)
);

HB1xp67_ASAP7_75t_L g6244 ( 
.A(n_5749),
.Y(n_6244)
);

OA21x2_ASAP7_75t_L g6245 ( 
.A1(n_5610),
.A2(n_4763),
.B(n_4759),
.Y(n_6245)
);

OR2x6_ASAP7_75t_L g6246 ( 
.A(n_5829),
.B(n_5163),
.Y(n_6246)
);

INVx2_ASAP7_75t_SL g6247 ( 
.A(n_5502),
.Y(n_6247)
);

HB1xp67_ASAP7_75t_L g6248 ( 
.A(n_5750),
.Y(n_6248)
);

INVx1_ASAP7_75t_L g6249 ( 
.A(n_5536),
.Y(n_6249)
);

INVx2_ASAP7_75t_L g6250 ( 
.A(n_5586),
.Y(n_6250)
);

INVxp67_ASAP7_75t_L g6251 ( 
.A(n_5497),
.Y(n_6251)
);

INVx1_ASAP7_75t_L g6252 ( 
.A(n_5526),
.Y(n_6252)
);

INVx2_ASAP7_75t_L g6253 ( 
.A(n_5592),
.Y(n_6253)
);

AND2x4_ASAP7_75t_L g6254 ( 
.A(n_5387),
.B(n_5006),
.Y(n_6254)
);

BUFx3_ASAP7_75t_L g6255 ( 
.A(n_5995),
.Y(n_6255)
);

AND2x2_ASAP7_75t_L g6256 ( 
.A(n_5649),
.B(n_4814),
.Y(n_6256)
);

OR2x2_ASAP7_75t_L g6257 ( 
.A(n_5814),
.B(n_4929),
.Y(n_6257)
);

AND2x2_ASAP7_75t_L g6258 ( 
.A(n_5649),
.B(n_4814),
.Y(n_6258)
);

AOI21xp33_ASAP7_75t_L g6259 ( 
.A1(n_5465),
.A2(n_5637),
.B(n_5943),
.Y(n_6259)
);

NAND2xp5_ASAP7_75t_L g6260 ( 
.A(n_5755),
.B(n_5049),
.Y(n_6260)
);

BUFx2_ASAP7_75t_L g6261 ( 
.A(n_5931),
.Y(n_6261)
);

INVx1_ASAP7_75t_L g6262 ( 
.A(n_5518),
.Y(n_6262)
);

AND2x2_ASAP7_75t_L g6263 ( 
.A(n_5601),
.B(n_4814),
.Y(n_6263)
);

INVx3_ASAP7_75t_L g6264 ( 
.A(n_5601),
.Y(n_6264)
);

AOI21xp5_ASAP7_75t_SL g6265 ( 
.A1(n_5650),
.A2(n_4404),
.B(n_5151),
.Y(n_6265)
);

BUFx3_ASAP7_75t_L g6266 ( 
.A(n_5395),
.Y(n_6266)
);

INVx1_ASAP7_75t_L g6267 ( 
.A(n_5518),
.Y(n_6267)
);

INVx2_ASAP7_75t_L g6268 ( 
.A(n_5592),
.Y(n_6268)
);

OR2x2_ASAP7_75t_L g6269 ( 
.A(n_5848),
.B(n_4929),
.Y(n_6269)
);

INVx2_ASAP7_75t_L g6270 ( 
.A(n_5594),
.Y(n_6270)
);

INVx1_ASAP7_75t_L g6271 ( 
.A(n_5451),
.Y(n_6271)
);

OR2x2_ASAP7_75t_L g6272 ( 
.A(n_5849),
.B(n_5026),
.Y(n_6272)
);

INVx1_ASAP7_75t_L g6273 ( 
.A(n_5455),
.Y(n_6273)
);

INVx1_ASAP7_75t_L g6274 ( 
.A(n_5455),
.Y(n_6274)
);

OR2x2_ASAP7_75t_L g6275 ( 
.A(n_5938),
.B(n_5026),
.Y(n_6275)
);

INVx1_ASAP7_75t_L g6276 ( 
.A(n_5456),
.Y(n_6276)
);

HB1xp67_ASAP7_75t_L g6277 ( 
.A(n_5371),
.Y(n_6277)
);

INVx2_ASAP7_75t_L g6278 ( 
.A(n_5594),
.Y(n_6278)
);

INVx1_ASAP7_75t_L g6279 ( 
.A(n_5456),
.Y(n_6279)
);

INVx2_ASAP7_75t_L g6280 ( 
.A(n_5596),
.Y(n_6280)
);

HB1xp67_ASAP7_75t_L g6281 ( 
.A(n_5402),
.Y(n_6281)
);

OR2x6_ASAP7_75t_L g6282 ( 
.A(n_5829),
.B(n_5163),
.Y(n_6282)
);

AND2x4_ASAP7_75t_L g6283 ( 
.A(n_5387),
.B(n_5092),
.Y(n_6283)
);

INVx2_ASAP7_75t_L g6284 ( 
.A(n_5596),
.Y(n_6284)
);

INVx1_ASAP7_75t_L g6285 ( 
.A(n_5464),
.Y(n_6285)
);

INVx2_ASAP7_75t_L g6286 ( 
.A(n_5600),
.Y(n_6286)
);

OR2x2_ASAP7_75t_L g6287 ( 
.A(n_5504),
.B(n_4863),
.Y(n_6287)
);

INVx1_ASAP7_75t_L g6288 ( 
.A(n_5464),
.Y(n_6288)
);

INVx2_ASAP7_75t_L g6289 ( 
.A(n_5600),
.Y(n_6289)
);

NOR2xp33_ASAP7_75t_L g6290 ( 
.A(n_5466),
.B(n_5154),
.Y(n_6290)
);

AO21x2_ASAP7_75t_L g6291 ( 
.A1(n_5547),
.A2(n_4677),
.B(n_4676),
.Y(n_6291)
);

INVx2_ASAP7_75t_L g6292 ( 
.A(n_5614),
.Y(n_6292)
);

BUFx3_ASAP7_75t_L g6293 ( 
.A(n_5395),
.Y(n_6293)
);

AND2x2_ASAP7_75t_L g6294 ( 
.A(n_5525),
.B(n_4814),
.Y(n_6294)
);

INVx1_ASAP7_75t_L g6295 ( 
.A(n_5467),
.Y(n_6295)
);

AND2x2_ASAP7_75t_L g6296 ( 
.A(n_5525),
.B(n_5453),
.Y(n_6296)
);

INVx1_ASAP7_75t_L g6297 ( 
.A(n_5467),
.Y(n_6297)
);

INVx1_ASAP7_75t_L g6298 ( 
.A(n_5469),
.Y(n_6298)
);

OR2x2_ASAP7_75t_L g6299 ( 
.A(n_5504),
.B(n_4863),
.Y(n_6299)
);

OR2x6_ASAP7_75t_L g6300 ( 
.A(n_5829),
.B(n_5163),
.Y(n_6300)
);

INVx1_ASAP7_75t_L g6301 ( 
.A(n_5476),
.Y(n_6301)
);

AO21x2_ASAP7_75t_L g6302 ( 
.A1(n_5547),
.A2(n_4692),
.B(n_4686),
.Y(n_6302)
);

INVx2_ASAP7_75t_L g6303 ( 
.A(n_5614),
.Y(n_6303)
);

AND2x2_ASAP7_75t_L g6304 ( 
.A(n_5525),
.B(n_5453),
.Y(n_6304)
);

NOR2xp33_ASAP7_75t_L g6305 ( 
.A(n_5633),
.B(n_5181),
.Y(n_6305)
);

AO21x2_ASAP7_75t_L g6306 ( 
.A1(n_5859),
.A2(n_4692),
.B(n_4686),
.Y(n_6306)
);

HB1xp67_ASAP7_75t_L g6307 ( 
.A(n_5405),
.Y(n_6307)
);

INVx2_ASAP7_75t_L g6308 ( 
.A(n_5616),
.Y(n_6308)
);

HB1xp67_ASAP7_75t_L g6309 ( 
.A(n_5457),
.Y(n_6309)
);

AND2x2_ASAP7_75t_L g6310 ( 
.A(n_5525),
.B(n_5555),
.Y(n_6310)
);

AND2x2_ASAP7_75t_L g6311 ( 
.A(n_5555),
.B(n_4902),
.Y(n_6311)
);

INVx2_ASAP7_75t_L g6312 ( 
.A(n_5616),
.Y(n_6312)
);

HB1xp67_ASAP7_75t_L g6313 ( 
.A(n_5479),
.Y(n_6313)
);

INVx1_ASAP7_75t_L g6314 ( 
.A(n_5476),
.Y(n_6314)
);

INVx2_ASAP7_75t_L g6315 ( 
.A(n_5619),
.Y(n_6315)
);

NOR2xp33_ASAP7_75t_L g6316 ( 
.A(n_6013),
.B(n_5181),
.Y(n_6316)
);

BUFx2_ASAP7_75t_L g6317 ( 
.A(n_5660),
.Y(n_6317)
);

NAND2xp5_ASAP7_75t_L g6318 ( 
.A(n_5793),
.B(n_5049),
.Y(n_6318)
);

NAND2xp5_ASAP7_75t_L g6319 ( 
.A(n_5812),
.B(n_5097),
.Y(n_6319)
);

AO21x2_ASAP7_75t_L g6320 ( 
.A1(n_5859),
.A2(n_4701),
.B(n_4694),
.Y(n_6320)
);

OR2x2_ASAP7_75t_L g6321 ( 
.A(n_5714),
.B(n_5328),
.Y(n_6321)
);

INVx1_ASAP7_75t_L g6322 ( 
.A(n_5477),
.Y(n_6322)
);

INVx1_ASAP7_75t_L g6323 ( 
.A(n_5477),
.Y(n_6323)
);

BUFx3_ASAP7_75t_L g6324 ( 
.A(n_5662),
.Y(n_6324)
);

INVx1_ASAP7_75t_L g6325 ( 
.A(n_5491),
.Y(n_6325)
);

INVx1_ASAP7_75t_L g6326 ( 
.A(n_5491),
.Y(n_6326)
);

BUFx2_ASAP7_75t_L g6327 ( 
.A(n_5660),
.Y(n_6327)
);

OR2x2_ASAP7_75t_L g6328 ( 
.A(n_5714),
.B(n_5328),
.Y(n_6328)
);

INVx2_ASAP7_75t_L g6329 ( 
.A(n_5619),
.Y(n_6329)
);

AO21x2_ASAP7_75t_L g6330 ( 
.A1(n_5859),
.A2(n_4701),
.B(n_4694),
.Y(n_6330)
);

INVx4_ASAP7_75t_L g6331 ( 
.A(n_5543),
.Y(n_6331)
);

BUFx3_ASAP7_75t_L g6332 ( 
.A(n_5398),
.Y(n_6332)
);

INVx1_ASAP7_75t_L g6333 ( 
.A(n_5492),
.Y(n_6333)
);

INVx1_ASAP7_75t_L g6334 ( 
.A(n_5492),
.Y(n_6334)
);

AO21x2_ASAP7_75t_L g6335 ( 
.A1(n_5909),
.A2(n_4716),
.B(n_4714),
.Y(n_6335)
);

AO21x2_ASAP7_75t_L g6336 ( 
.A1(n_5733),
.A2(n_5868),
.B(n_5903),
.Y(n_6336)
);

AOI21xp33_ASAP7_75t_L g6337 ( 
.A1(n_5832),
.A2(n_4671),
.B(n_4876),
.Y(n_6337)
);

AND2x2_ASAP7_75t_L g6338 ( 
.A(n_5861),
.B(n_4902),
.Y(n_6338)
);

INVx1_ASAP7_75t_L g6339 ( 
.A(n_5495),
.Y(n_6339)
);

INVx3_ASAP7_75t_L g6340 ( 
.A(n_5708),
.Y(n_6340)
);

INVx1_ASAP7_75t_L g6341 ( 
.A(n_5495),
.Y(n_6341)
);

BUFx2_ASAP7_75t_L g6342 ( 
.A(n_5672),
.Y(n_6342)
);

INVx1_ASAP7_75t_SL g6343 ( 
.A(n_5559),
.Y(n_6343)
);

INVx1_ASAP7_75t_L g6344 ( 
.A(n_5500),
.Y(n_6344)
);

AND2x2_ASAP7_75t_L g6345 ( 
.A(n_5861),
.B(n_4902),
.Y(n_6345)
);

INVxp67_ASAP7_75t_L g6346 ( 
.A(n_5379),
.Y(n_6346)
);

INVx2_ASAP7_75t_SL g6347 ( 
.A(n_5429),
.Y(n_6347)
);

HB1xp67_ASAP7_75t_L g6348 ( 
.A(n_5487),
.Y(n_6348)
);

BUFx3_ASAP7_75t_L g6349 ( 
.A(n_5398),
.Y(n_6349)
);

INVx2_ASAP7_75t_L g6350 ( 
.A(n_5620),
.Y(n_6350)
);

AO21x2_ASAP7_75t_L g6351 ( 
.A1(n_5733),
.A2(n_4717),
.B(n_4714),
.Y(n_6351)
);

INVx1_ASAP7_75t_L g6352 ( 
.A(n_5500),
.Y(n_6352)
);

INVx1_ASAP7_75t_L g6353 ( 
.A(n_5510),
.Y(n_6353)
);

BUFx6f_ASAP7_75t_L g6354 ( 
.A(n_5543),
.Y(n_6354)
);

OR2x6_ASAP7_75t_L g6355 ( 
.A(n_5829),
.B(n_5163),
.Y(n_6355)
);

AND2x2_ASAP7_75t_L g6356 ( 
.A(n_5878),
.B(n_4902),
.Y(n_6356)
);

INVx1_ASAP7_75t_L g6357 ( 
.A(n_5510),
.Y(n_6357)
);

AO21x2_ASAP7_75t_L g6358 ( 
.A1(n_5733),
.A2(n_4717),
.B(n_4714),
.Y(n_6358)
);

OR2x6_ASAP7_75t_L g6359 ( 
.A(n_5839),
.B(n_5163),
.Y(n_6359)
);

INVx2_ASAP7_75t_L g6360 ( 
.A(n_5620),
.Y(n_6360)
);

INVx1_ASAP7_75t_L g6361 ( 
.A(n_5511),
.Y(n_6361)
);

INVx2_ASAP7_75t_L g6362 ( 
.A(n_5370),
.Y(n_6362)
);

AND2x4_ASAP7_75t_L g6363 ( 
.A(n_5387),
.B(n_5092),
.Y(n_6363)
);

INVx1_ASAP7_75t_SL g6364 ( 
.A(n_5377),
.Y(n_6364)
);

HB1xp67_ASAP7_75t_L g6365 ( 
.A(n_5493),
.Y(n_6365)
);

HB1xp67_ASAP7_75t_L g6366 ( 
.A(n_5503),
.Y(n_6366)
);

AND2x2_ASAP7_75t_L g6367 ( 
.A(n_5878),
.B(n_5069),
.Y(n_6367)
);

INVx3_ASAP7_75t_L g6368 ( 
.A(n_5708),
.Y(n_6368)
);

AOI22xp5_ASAP7_75t_L g6369 ( 
.A1(n_5670),
.A2(n_5655),
.B1(n_5690),
.B2(n_5474),
.Y(n_6369)
);

AO21x2_ASAP7_75t_L g6370 ( 
.A1(n_5868),
.A2(n_4721),
.B(n_4717),
.Y(n_6370)
);

INVx3_ASAP7_75t_L g6371 ( 
.A(n_5708),
.Y(n_6371)
);

BUFx2_ASAP7_75t_L g6372 ( 
.A(n_5672),
.Y(n_6372)
);

AND2x2_ASAP7_75t_L g6373 ( 
.A(n_5891),
.B(n_5609),
.Y(n_6373)
);

INVx2_ASAP7_75t_L g6374 ( 
.A(n_5370),
.Y(n_6374)
);

AO21x2_ASAP7_75t_L g6375 ( 
.A1(n_5868),
.A2(n_4721),
.B(n_4842),
.Y(n_6375)
);

OAI321xp33_ASAP7_75t_L g6376 ( 
.A1(n_5850),
.A2(n_5276),
.A3(n_4987),
.B1(n_4691),
.B2(n_4935),
.C(n_4712),
.Y(n_6376)
);

INVx1_ASAP7_75t_L g6377 ( 
.A(n_5511),
.Y(n_6377)
);

OAI21x1_ASAP7_75t_L g6378 ( 
.A1(n_5437),
.A2(n_5146),
.B(n_5102),
.Y(n_6378)
);

INVx2_ASAP7_75t_SL g6379 ( 
.A(n_5429),
.Y(n_6379)
);

BUFx2_ASAP7_75t_L g6380 ( 
.A(n_5390),
.Y(n_6380)
);

OAI21xp5_ASAP7_75t_L g6381 ( 
.A1(n_5713),
.A2(n_4935),
.B(n_4960),
.Y(n_6381)
);

AO21x2_ASAP7_75t_L g6382 ( 
.A1(n_5903),
.A2(n_4721),
.B(n_4842),
.Y(n_6382)
);

OAI21x1_ASAP7_75t_L g6383 ( 
.A1(n_5437),
.A2(n_5159),
.B(n_5146),
.Y(n_6383)
);

INVx2_ASAP7_75t_L g6384 ( 
.A(n_5380),
.Y(n_6384)
);

INVx2_ASAP7_75t_L g6385 ( 
.A(n_5380),
.Y(n_6385)
);

BUFx2_ASAP7_75t_L g6386 ( 
.A(n_5390),
.Y(n_6386)
);

BUFx2_ASAP7_75t_L g6387 ( 
.A(n_5390),
.Y(n_6387)
);

INVx2_ASAP7_75t_L g6388 ( 
.A(n_5382),
.Y(n_6388)
);

INVx2_ASAP7_75t_L g6389 ( 
.A(n_5382),
.Y(n_6389)
);

AND2x2_ASAP7_75t_L g6390 ( 
.A(n_5891),
.B(n_5069),
.Y(n_6390)
);

INVx2_ASAP7_75t_L g6391 ( 
.A(n_5386),
.Y(n_6391)
);

INVx2_ASAP7_75t_SL g6392 ( 
.A(n_5440),
.Y(n_6392)
);

OR2x6_ASAP7_75t_L g6393 ( 
.A(n_5839),
.B(n_5194),
.Y(n_6393)
);

NAND2xp5_ASAP7_75t_L g6394 ( 
.A(n_5816),
.B(n_5097),
.Y(n_6394)
);

OA21x2_ASAP7_75t_L g6395 ( 
.A1(n_5610),
.A2(n_4763),
.B(n_4759),
.Y(n_6395)
);

INVx2_ASAP7_75t_L g6396 ( 
.A(n_5386),
.Y(n_6396)
);

AND2x2_ASAP7_75t_L g6397 ( 
.A(n_5609),
.B(n_5079),
.Y(n_6397)
);

AND2x2_ASAP7_75t_L g6398 ( 
.A(n_5609),
.B(n_5079),
.Y(n_6398)
);

INVx2_ASAP7_75t_L g6399 ( 
.A(n_5389),
.Y(n_6399)
);

NOR2xp33_ASAP7_75t_L g6400 ( 
.A(n_5699),
.B(n_5185),
.Y(n_6400)
);

INVx1_ASAP7_75t_L g6401 ( 
.A(n_5514),
.Y(n_6401)
);

NOR2xp33_ASAP7_75t_L g6402 ( 
.A(n_5699),
.B(n_5185),
.Y(n_6402)
);

AND2x2_ASAP7_75t_L g6403 ( 
.A(n_5695),
.B(n_5132),
.Y(n_6403)
);

BUFx2_ASAP7_75t_L g6404 ( 
.A(n_5390),
.Y(n_6404)
);

HB1xp67_ASAP7_75t_L g6405 ( 
.A(n_5505),
.Y(n_6405)
);

INVx1_ASAP7_75t_L g6406 ( 
.A(n_5514),
.Y(n_6406)
);

INVx3_ASAP7_75t_L g6407 ( 
.A(n_5708),
.Y(n_6407)
);

OR2x6_ASAP7_75t_L g6408 ( 
.A(n_5839),
.B(n_5194),
.Y(n_6408)
);

INVx1_ASAP7_75t_L g6409 ( 
.A(n_5519),
.Y(n_6409)
);

INVx1_ASAP7_75t_L g6410 ( 
.A(n_5519),
.Y(n_6410)
);

INVx1_ASAP7_75t_L g6411 ( 
.A(n_5522),
.Y(n_6411)
);

NOR2xp33_ASAP7_75t_L g6412 ( 
.A(n_5699),
.B(n_5063),
.Y(n_6412)
);

OR2x2_ASAP7_75t_L g6413 ( 
.A(n_5799),
.B(n_5323),
.Y(n_6413)
);

AND2x2_ASAP7_75t_L g6414 ( 
.A(n_5695),
.B(n_5132),
.Y(n_6414)
);

HB1xp67_ASAP7_75t_L g6415 ( 
.A(n_5535),
.Y(n_6415)
);

INVx2_ASAP7_75t_L g6416 ( 
.A(n_5389),
.Y(n_6416)
);

INVx2_ASAP7_75t_L g6417 ( 
.A(n_5399),
.Y(n_6417)
);

AO21x2_ASAP7_75t_L g6418 ( 
.A1(n_5903),
.A2(n_4850),
.B(n_4842),
.Y(n_6418)
);

AND2x2_ASAP7_75t_L g6419 ( 
.A(n_5780),
.B(n_5782),
.Y(n_6419)
);

OR2x6_ASAP7_75t_L g6420 ( 
.A(n_5839),
.B(n_6003),
.Y(n_6420)
);

NOR2xp33_ASAP7_75t_SL g6421 ( 
.A(n_5401),
.B(n_5322),
.Y(n_6421)
);

NAND2xp5_ASAP7_75t_L g6422 ( 
.A(n_5820),
.B(n_5114),
.Y(n_6422)
);

INVx2_ASAP7_75t_L g6423 ( 
.A(n_5399),
.Y(n_6423)
);

OR2x2_ASAP7_75t_L g6424 ( 
.A(n_5799),
.B(n_5324),
.Y(n_6424)
);

OAI211xp5_ASAP7_75t_L g6425 ( 
.A1(n_5706),
.A2(n_5850),
.B(n_5981),
.C(n_5501),
.Y(n_6425)
);

BUFx3_ASAP7_75t_L g6426 ( 
.A(n_5543),
.Y(n_6426)
);

OR2x2_ASAP7_75t_L g6427 ( 
.A(n_5960),
.B(n_4455),
.Y(n_6427)
);

AND2x2_ASAP7_75t_L g6428 ( 
.A(n_5780),
.B(n_5138),
.Y(n_6428)
);

OR2x2_ASAP7_75t_L g6429 ( 
.A(n_5960),
.B(n_4455),
.Y(n_6429)
);

HB1xp67_ASAP7_75t_L g6430 ( 
.A(n_5542),
.Y(n_6430)
);

INVx1_ASAP7_75t_L g6431 ( 
.A(n_5522),
.Y(n_6431)
);

AO21x2_ASAP7_75t_L g6432 ( 
.A1(n_5958),
.A2(n_4851),
.B(n_4850),
.Y(n_6432)
);

INVx2_ASAP7_75t_L g6433 ( 
.A(n_5406),
.Y(n_6433)
);

AND2x2_ASAP7_75t_L g6434 ( 
.A(n_5782),
.B(n_5138),
.Y(n_6434)
);

INVx2_ASAP7_75t_L g6435 ( 
.A(n_5406),
.Y(n_6435)
);

INVx2_ASAP7_75t_L g6436 ( 
.A(n_5409),
.Y(n_6436)
);

INVx1_ASAP7_75t_L g6437 ( 
.A(n_5523),
.Y(n_6437)
);

AND2x2_ASAP7_75t_L g6438 ( 
.A(n_5920),
.B(n_5201),
.Y(n_6438)
);

OAI21x1_ASAP7_75t_L g6439 ( 
.A1(n_5527),
.A2(n_5159),
.B(n_5146),
.Y(n_6439)
);

INVx3_ASAP7_75t_L g6440 ( 
.A(n_5741),
.Y(n_6440)
);

AND2x4_ASAP7_75t_L g6441 ( 
.A(n_5920),
.B(n_5238),
.Y(n_6441)
);

AND2x2_ASAP7_75t_L g6442 ( 
.A(n_5940),
.B(n_5201),
.Y(n_6442)
);

INVx1_ASAP7_75t_L g6443 ( 
.A(n_5523),
.Y(n_6443)
);

AND2x2_ASAP7_75t_L g6444 ( 
.A(n_5940),
.B(n_5201),
.Y(n_6444)
);

INVx1_ASAP7_75t_L g6445 ( 
.A(n_5526),
.Y(n_6445)
);

AO21x2_ASAP7_75t_L g6446 ( 
.A1(n_5958),
.A2(n_4851),
.B(n_4850),
.Y(n_6446)
);

INVx1_ASAP7_75t_L g6447 ( 
.A(n_5530),
.Y(n_6447)
);

INVx1_ASAP7_75t_L g6448 ( 
.A(n_5530),
.Y(n_6448)
);

AO21x2_ASAP7_75t_L g6449 ( 
.A1(n_5939),
.A2(n_4858),
.B(n_4851),
.Y(n_6449)
);

BUFx2_ASAP7_75t_L g6450 ( 
.A(n_5440),
.Y(n_6450)
);

AND2x2_ASAP7_75t_L g6451 ( 
.A(n_5976),
.B(n_5201),
.Y(n_6451)
);

NAND2xp5_ASAP7_75t_L g6452 ( 
.A(n_5452),
.B(n_5114),
.Y(n_6452)
);

INVx1_ASAP7_75t_L g6453 ( 
.A(n_5531),
.Y(n_6453)
);

NAND2xp5_ASAP7_75t_L g6454 ( 
.A(n_5557),
.B(n_5169),
.Y(n_6454)
);

AOI221xp5_ASAP7_75t_L g6455 ( 
.A1(n_5790),
.A2(n_4876),
.B1(n_4871),
.B2(n_4845),
.C(n_5240),
.Y(n_6455)
);

HB1xp67_ASAP7_75t_L g6456 ( 
.A(n_5563),
.Y(n_6456)
);

INVx1_ASAP7_75t_L g6457 ( 
.A(n_5531),
.Y(n_6457)
);

INVx2_ASAP7_75t_L g6458 ( 
.A(n_5409),
.Y(n_6458)
);

INVx1_ASAP7_75t_L g6459 ( 
.A(n_5536),
.Y(n_6459)
);

OA21x2_ASAP7_75t_L g6460 ( 
.A1(n_5692),
.A2(n_4776),
.B(n_4759),
.Y(n_6460)
);

AND2x2_ASAP7_75t_L g6461 ( 
.A(n_5976),
.B(n_5354),
.Y(n_6461)
);

INVx1_ASAP7_75t_L g6462 ( 
.A(n_5537),
.Y(n_6462)
);

INVx1_ASAP7_75t_L g6463 ( 
.A(n_5537),
.Y(n_6463)
);

AOI21x1_ASAP7_75t_L g6464 ( 
.A1(n_5684),
.A2(n_5107),
.B(n_5060),
.Y(n_6464)
);

AO21x2_ASAP7_75t_L g6465 ( 
.A1(n_5939),
.A2(n_4880),
.B(n_4858),
.Y(n_6465)
);

NAND3xp33_ASAP7_75t_L g6466 ( 
.A(n_5862),
.B(n_4344),
.C(n_5294),
.Y(n_6466)
);

AO21x2_ASAP7_75t_L g6467 ( 
.A1(n_5945),
.A2(n_5413),
.B(n_5410),
.Y(n_6467)
);

INVx2_ASAP7_75t_L g6468 ( 
.A(n_5410),
.Y(n_6468)
);

OAI21x1_ASAP7_75t_L g6469 ( 
.A1(n_5527),
.A2(n_5214),
.B(n_5159),
.Y(n_6469)
);

INVx2_ASAP7_75t_L g6470 ( 
.A(n_5413),
.Y(n_6470)
);

INVx1_ASAP7_75t_L g6471 ( 
.A(n_5545),
.Y(n_6471)
);

INVx1_ASAP7_75t_L g6472 ( 
.A(n_5545),
.Y(n_6472)
);

BUFx2_ASAP7_75t_L g6473 ( 
.A(n_5471),
.Y(n_6473)
);

OR2x2_ASAP7_75t_L g6474 ( 
.A(n_5509),
.B(n_5169),
.Y(n_6474)
);

HB1xp67_ASAP7_75t_L g6475 ( 
.A(n_5566),
.Y(n_6475)
);

INVx3_ASAP7_75t_L g6476 ( 
.A(n_5741),
.Y(n_6476)
);

OR2x6_ASAP7_75t_L g6477 ( 
.A(n_5839),
.B(n_4839),
.Y(n_6477)
);

AOI221xp5_ASAP7_75t_L g6478 ( 
.A1(n_5790),
.A2(n_4876),
.B1(n_4871),
.B2(n_4845),
.C(n_4858),
.Y(n_6478)
);

NAND2xp5_ASAP7_75t_L g6479 ( 
.A(n_5602),
.B(n_5211),
.Y(n_6479)
);

AND2x2_ASAP7_75t_L g6480 ( 
.A(n_5992),
.B(n_5354),
.Y(n_6480)
);

BUFx2_ASAP7_75t_L g6481 ( 
.A(n_5471),
.Y(n_6481)
);

INVx1_ASAP7_75t_L g6482 ( 
.A(n_5548),
.Y(n_6482)
);

INVx1_ASAP7_75t_L g6483 ( 
.A(n_5548),
.Y(n_6483)
);

INVx2_ASAP7_75t_L g6484 ( 
.A(n_5420),
.Y(n_6484)
);

BUFx3_ASAP7_75t_L g6485 ( 
.A(n_5543),
.Y(n_6485)
);

BUFx3_ASAP7_75t_L g6486 ( 
.A(n_5551),
.Y(n_6486)
);

NAND2xp5_ASAP7_75t_L g6487 ( 
.A(n_5628),
.B(n_5211),
.Y(n_6487)
);

INVx1_ASAP7_75t_L g6488 ( 
.A(n_5550),
.Y(n_6488)
);

AO21x2_ASAP7_75t_L g6489 ( 
.A1(n_5945),
.A2(n_4881),
.B(n_4880),
.Y(n_6489)
);

INVx2_ASAP7_75t_SL g6490 ( 
.A(n_5481),
.Y(n_6490)
);

INVxp67_ASAP7_75t_L g6491 ( 
.A(n_5742),
.Y(n_6491)
);

INVx2_ASAP7_75t_L g6492 ( 
.A(n_5420),
.Y(n_6492)
);

OA21x2_ASAP7_75t_L g6493 ( 
.A1(n_5692),
.A2(n_4788),
.B(n_4776),
.Y(n_6493)
);

INVx1_ASAP7_75t_L g6494 ( 
.A(n_5550),
.Y(n_6494)
);

NOR2xp33_ASAP7_75t_L g6495 ( 
.A(n_5879),
.B(n_5279),
.Y(n_6495)
);

INVxp67_ASAP7_75t_SL g6496 ( 
.A(n_5485),
.Y(n_6496)
);

INVx1_ASAP7_75t_L g6497 ( 
.A(n_5553),
.Y(n_6497)
);

CKINVDCx20_ASAP7_75t_R g6498 ( 
.A(n_5994),
.Y(n_6498)
);

INVx1_ASAP7_75t_L g6499 ( 
.A(n_5553),
.Y(n_6499)
);

INVx1_ASAP7_75t_L g6500 ( 
.A(n_5562),
.Y(n_6500)
);

NAND2xp5_ASAP7_75t_L g6501 ( 
.A(n_5787),
.B(n_5258),
.Y(n_6501)
);

NOR2xp33_ASAP7_75t_L g6502 ( 
.A(n_5653),
.B(n_5193),
.Y(n_6502)
);

HB1xp67_ASAP7_75t_L g6503 ( 
.A(n_5792),
.Y(n_6503)
);

BUFx2_ASAP7_75t_L g6504 ( 
.A(n_5481),
.Y(n_6504)
);

INVx1_ASAP7_75t_L g6505 ( 
.A(n_5562),
.Y(n_6505)
);

AO21x2_ASAP7_75t_L g6506 ( 
.A1(n_5435),
.A2(n_4881),
.B(n_4880),
.Y(n_6506)
);

INVx2_ASAP7_75t_L g6507 ( 
.A(n_5435),
.Y(n_6507)
);

AOI21xp5_ASAP7_75t_L g6508 ( 
.A1(n_5433),
.A2(n_4794),
.B(n_4960),
.Y(n_6508)
);

AO21x1_ASAP7_75t_SL g6509 ( 
.A1(n_6006),
.A2(n_5255),
.B(n_5322),
.Y(n_6509)
);

INVx1_ASAP7_75t_L g6510 ( 
.A(n_5565),
.Y(n_6510)
);

INVx2_ASAP7_75t_SL g6511 ( 
.A(n_5549),
.Y(n_6511)
);

INVx1_ASAP7_75t_L g6512 ( 
.A(n_5565),
.Y(n_6512)
);

INVx1_ASAP7_75t_L g6513 ( 
.A(n_5567),
.Y(n_6513)
);

INVx2_ASAP7_75t_L g6514 ( 
.A(n_5705),
.Y(n_6514)
);

INVx1_ASAP7_75t_L g6515 ( 
.A(n_5567),
.Y(n_6515)
);

INVx3_ASAP7_75t_L g6516 ( 
.A(n_5741),
.Y(n_6516)
);

INVx1_ASAP7_75t_L g6517 ( 
.A(n_5570),
.Y(n_6517)
);

OR2x6_ASAP7_75t_L g6518 ( 
.A(n_6003),
.B(n_4839),
.Y(n_6518)
);

AND2x2_ASAP7_75t_L g6519 ( 
.A(n_5992),
.B(n_5354),
.Y(n_6519)
);

INVx2_ASAP7_75t_L g6520 ( 
.A(n_5705),
.Y(n_6520)
);

INVx1_ASAP7_75t_L g6521 ( 
.A(n_5570),
.Y(n_6521)
);

INVx2_ASAP7_75t_L g6522 ( 
.A(n_5709),
.Y(n_6522)
);

INVx2_ASAP7_75t_L g6523 ( 
.A(n_5709),
.Y(n_6523)
);

INVx2_ASAP7_75t_L g6524 ( 
.A(n_5720),
.Y(n_6524)
);

NAND2xp5_ASAP7_75t_L g6525 ( 
.A(n_5473),
.B(n_5579),
.Y(n_6525)
);

INVx1_ASAP7_75t_L g6526 ( 
.A(n_5571),
.Y(n_6526)
);

BUFx8_ASAP7_75t_L g6527 ( 
.A(n_5551),
.Y(n_6527)
);

NAND2xp5_ASAP7_75t_L g6528 ( 
.A(n_5509),
.B(n_5258),
.Y(n_6528)
);

AND2x2_ASAP7_75t_L g6529 ( 
.A(n_6012),
.B(n_5238),
.Y(n_6529)
);

HB1xp67_ASAP7_75t_L g6530 ( 
.A(n_5806),
.Y(n_6530)
);

BUFx3_ASAP7_75t_L g6531 ( 
.A(n_5551),
.Y(n_6531)
);

NAND2xp5_ASAP7_75t_L g6532 ( 
.A(n_5806),
.B(n_5271),
.Y(n_6532)
);

INVx1_ASAP7_75t_L g6533 ( 
.A(n_5571),
.Y(n_6533)
);

INVx1_ASAP7_75t_L g6534 ( 
.A(n_5572),
.Y(n_6534)
);

BUFx5_ASAP7_75t_L g6535 ( 
.A(n_5552),
.Y(n_6535)
);

OA21x2_ASAP7_75t_L g6536 ( 
.A1(n_5880),
.A2(n_4788),
.B(n_4776),
.Y(n_6536)
);

INVx1_ASAP7_75t_L g6537 ( 
.A(n_5572),
.Y(n_6537)
);

OR2x2_ASAP7_75t_L g6538 ( 
.A(n_5974),
.B(n_5271),
.Y(n_6538)
);

INVx1_ASAP7_75t_L g6539 ( 
.A(n_5573),
.Y(n_6539)
);

INVx2_ASAP7_75t_L g6540 ( 
.A(n_5720),
.Y(n_6540)
);

INVx2_ASAP7_75t_L g6541 ( 
.A(n_5722),
.Y(n_6541)
);

AO21x2_ASAP7_75t_L g6542 ( 
.A1(n_5722),
.A2(n_4893),
.B(n_4881),
.Y(n_6542)
);

INVx3_ASAP7_75t_L g6543 ( 
.A(n_5741),
.Y(n_6543)
);

INVx1_ASAP7_75t_L g6544 ( 
.A(n_5573),
.Y(n_6544)
);

AND2x4_ASAP7_75t_L g6545 ( 
.A(n_6012),
.B(n_5238),
.Y(n_6545)
);

AOI22xp33_ASAP7_75t_L g6546 ( 
.A1(n_5831),
.A2(n_4845),
.B1(n_4871),
.B2(n_4770),
.Y(n_6546)
);

INVx1_ASAP7_75t_L g6547 ( 
.A(n_6011),
.Y(n_6547)
);

INVx1_ASAP7_75t_L g6548 ( 
.A(n_6011),
.Y(n_6548)
);

BUFx4f_ASAP7_75t_SL g6549 ( 
.A(n_5725),
.Y(n_6549)
);

BUFx3_ASAP7_75t_L g6550 ( 
.A(n_5551),
.Y(n_6550)
);

INVx2_ASAP7_75t_L g6551 ( 
.A(n_5730),
.Y(n_6551)
);

INVx1_ASAP7_75t_L g6552 ( 
.A(n_6010),
.Y(n_6552)
);

OR2x2_ASAP7_75t_L g6553 ( 
.A(n_5974),
.B(n_5362),
.Y(n_6553)
);

OR2x2_ASAP7_75t_L g6554 ( 
.A(n_5978),
.B(n_5362),
.Y(n_6554)
);

AO21x2_ASAP7_75t_L g6555 ( 
.A1(n_5730),
.A2(n_4898),
.B(n_4893),
.Y(n_6555)
);

AND2x2_ASAP7_75t_L g6556 ( 
.A(n_5381),
.B(n_5238),
.Y(n_6556)
);

INVx3_ASAP7_75t_L g6557 ( 
.A(n_6283),
.Y(n_6557)
);

INVx2_ASAP7_75t_SL g6558 ( 
.A(n_6058),
.Y(n_6558)
);

INVx2_ASAP7_75t_L g6559 ( 
.A(n_6336),
.Y(n_6559)
);

HB1xp67_ASAP7_75t_L g6560 ( 
.A(n_6086),
.Y(n_6560)
);

INVx2_ASAP7_75t_L g6561 ( 
.A(n_6336),
.Y(n_6561)
);

INVx1_ASAP7_75t_L g6562 ( 
.A(n_6026),
.Y(n_6562)
);

NAND2xp5_ASAP7_75t_L g6563 ( 
.A(n_6112),
.B(n_5817),
.Y(n_6563)
);

INVx1_ASAP7_75t_L g6564 ( 
.A(n_6053),
.Y(n_6564)
);

INVx2_ASAP7_75t_L g6565 ( 
.A(n_6336),
.Y(n_6565)
);

AND2x4_ASAP7_75t_L g6566 ( 
.A(n_6045),
.B(n_6003),
.Y(n_6566)
);

AND2x2_ASAP7_75t_L g6567 ( 
.A(n_6241),
.B(n_5686),
.Y(n_6567)
);

NAND2xp5_ASAP7_75t_L g6568 ( 
.A(n_6093),
.B(n_5817),
.Y(n_6568)
);

NAND2xp5_ASAP7_75t_L g6569 ( 
.A(n_6093),
.B(n_6142),
.Y(n_6569)
);

AND2x4_ASAP7_75t_SL g6570 ( 
.A(n_6058),
.B(n_6137),
.Y(n_6570)
);

HB1xp67_ASAP7_75t_L g6571 ( 
.A(n_6261),
.Y(n_6571)
);

AND2x4_ASAP7_75t_L g6572 ( 
.A(n_6045),
.B(n_6003),
.Y(n_6572)
);

AND2x2_ASAP7_75t_L g6573 ( 
.A(n_6241),
.B(n_5686),
.Y(n_6573)
);

BUFx2_ASAP7_75t_L g6574 ( 
.A(n_6261),
.Y(n_6574)
);

INVx2_ASAP7_75t_L g6575 ( 
.A(n_6018),
.Y(n_6575)
);

INVxp67_ASAP7_75t_L g6576 ( 
.A(n_6450),
.Y(n_6576)
);

INVx1_ASAP7_75t_L g6577 ( 
.A(n_6062),
.Y(n_6577)
);

BUFx3_ASAP7_75t_L g6578 ( 
.A(n_6498),
.Y(n_6578)
);

INVx1_ASAP7_75t_L g6579 ( 
.A(n_6064),
.Y(n_6579)
);

AND2x2_ASAP7_75t_L g6580 ( 
.A(n_6021),
.B(n_5719),
.Y(n_6580)
);

AND2x2_ASAP7_75t_L g6581 ( 
.A(n_6021),
.B(n_5719),
.Y(n_6581)
);

BUFx3_ASAP7_75t_L g6582 ( 
.A(n_6498),
.Y(n_6582)
);

INVx1_ASAP7_75t_L g6583 ( 
.A(n_6082),
.Y(n_6583)
);

NAND2xp5_ASAP7_75t_L g6584 ( 
.A(n_6093),
.B(n_6142),
.Y(n_6584)
);

AND2x4_ASAP7_75t_L g6585 ( 
.A(n_6221),
.B(n_5408),
.Y(n_6585)
);

HB1xp67_ASAP7_75t_L g6586 ( 
.A(n_6192),
.Y(n_6586)
);

AOI22xp33_ASAP7_75t_L g6587 ( 
.A1(n_6090),
.A2(n_4845),
.B1(n_4871),
.B2(n_5254),
.Y(n_6587)
);

AND2x2_ASAP7_75t_L g6588 ( 
.A(n_6205),
.B(n_5711),
.Y(n_6588)
);

INVx1_ASAP7_75t_L g6589 ( 
.A(n_6095),
.Y(n_6589)
);

AND2x2_ASAP7_75t_L g6590 ( 
.A(n_6205),
.B(n_5858),
.Y(n_6590)
);

AND2x2_ASAP7_75t_L g6591 ( 
.A(n_6213),
.B(n_5381),
.Y(n_6591)
);

INVx2_ASAP7_75t_L g6592 ( 
.A(n_6018),
.Y(n_6592)
);

INVx1_ASAP7_75t_L g6593 ( 
.A(n_6152),
.Y(n_6593)
);

BUFx2_ASAP7_75t_L g6594 ( 
.A(n_6177),
.Y(n_6594)
);

NAND2x1_ASAP7_75t_L g6595 ( 
.A(n_6265),
.B(n_5621),
.Y(n_6595)
);

INVx1_ASAP7_75t_L g6596 ( 
.A(n_6209),
.Y(n_6596)
);

OR2x2_ASAP7_75t_SL g6597 ( 
.A(n_6058),
.B(n_6137),
.Y(n_6597)
);

OR2x2_ASAP7_75t_L g6598 ( 
.A(n_6160),
.B(n_5978),
.Y(n_6598)
);

OAI21x1_ASAP7_75t_L g6599 ( 
.A1(n_6265),
.A2(n_5989),
.B(n_5643),
.Y(n_6599)
);

AND2x2_ASAP7_75t_L g6600 ( 
.A(n_6213),
.B(n_5407),
.Y(n_6600)
);

OR2x2_ASAP7_75t_L g6601 ( 
.A(n_6228),
.B(n_5831),
.Y(n_6601)
);

NAND2x1p5_ASAP7_75t_SL g6602 ( 
.A(n_6347),
.B(n_5517),
.Y(n_6602)
);

INVx1_ASAP7_75t_L g6603 ( 
.A(n_6034),
.Y(n_6603)
);

INVxp67_ASAP7_75t_SL g6604 ( 
.A(n_6080),
.Y(n_6604)
);

BUFx12f_ASAP7_75t_L g6605 ( 
.A(n_6208),
.Y(n_6605)
);

AND2x4_ASAP7_75t_SL g6606 ( 
.A(n_6058),
.B(n_5551),
.Y(n_6606)
);

AND2x2_ASAP7_75t_L g6607 ( 
.A(n_6221),
.B(n_5407),
.Y(n_6607)
);

INVx1_ASAP7_75t_L g6608 ( 
.A(n_6034),
.Y(n_6608)
);

INVx2_ASAP7_75t_L g6609 ( 
.A(n_6018),
.Y(n_6609)
);

AND2x2_ASAP7_75t_L g6610 ( 
.A(n_6235),
.B(n_5414),
.Y(n_6610)
);

HB1xp67_ASAP7_75t_L g6611 ( 
.A(n_6251),
.Y(n_6611)
);

INVx2_ASAP7_75t_L g6612 ( 
.A(n_6023),
.Y(n_6612)
);

INVx2_ASAP7_75t_L g6613 ( 
.A(n_6023),
.Y(n_6613)
);

AND2x2_ASAP7_75t_L g6614 ( 
.A(n_6235),
.B(n_5414),
.Y(n_6614)
);

HB1xp67_ASAP7_75t_L g6615 ( 
.A(n_6530),
.Y(n_6615)
);

NAND2xp5_ASAP7_75t_L g6616 ( 
.A(n_6067),
.B(n_5517),
.Y(n_6616)
);

INVx2_ASAP7_75t_L g6617 ( 
.A(n_6035),
.Y(n_6617)
);

HB1xp67_ASAP7_75t_L g6618 ( 
.A(n_6229),
.Y(n_6618)
);

INVx1_ASAP7_75t_L g6619 ( 
.A(n_6036),
.Y(n_6619)
);

NAND2xp5_ASAP7_75t_L g6620 ( 
.A(n_6042),
.B(n_5528),
.Y(n_6620)
);

INVx2_ASAP7_75t_L g6621 ( 
.A(n_6035),
.Y(n_6621)
);

NAND2xp5_ASAP7_75t_L g6622 ( 
.A(n_6259),
.B(n_5528),
.Y(n_6622)
);

INVx2_ASAP7_75t_L g6623 ( 
.A(n_6039),
.Y(n_6623)
);

NAND2xp5_ASAP7_75t_L g6624 ( 
.A(n_6233),
.B(n_5408),
.Y(n_6624)
);

BUFx6f_ASAP7_75t_L g6625 ( 
.A(n_6096),
.Y(n_6625)
);

BUFx3_ASAP7_75t_L g6626 ( 
.A(n_6266),
.Y(n_6626)
);

AND2x2_ASAP7_75t_L g6627 ( 
.A(n_6240),
.B(n_5430),
.Y(n_6627)
);

BUFx3_ASAP7_75t_L g6628 ( 
.A(n_6266),
.Y(n_6628)
);

INVx2_ASAP7_75t_L g6629 ( 
.A(n_6039),
.Y(n_6629)
);

OR2x2_ASAP7_75t_L g6630 ( 
.A(n_6228),
.B(n_5430),
.Y(n_6630)
);

NAND2xp5_ASAP7_75t_L g6631 ( 
.A(n_6244),
.B(n_5436),
.Y(n_6631)
);

INVx2_ASAP7_75t_L g6632 ( 
.A(n_6041),
.Y(n_6632)
);

INVx1_ASAP7_75t_L g6633 ( 
.A(n_6036),
.Y(n_6633)
);

NAND2xp5_ASAP7_75t_L g6634 ( 
.A(n_6248),
.B(n_5436),
.Y(n_6634)
);

AND2x2_ASAP7_75t_L g6635 ( 
.A(n_6240),
.B(n_5944),
.Y(n_6635)
);

AND2x2_ASAP7_75t_L g6636 ( 
.A(n_6242),
.B(n_5944),
.Y(n_6636)
);

INVx1_ASAP7_75t_L g6637 ( 
.A(n_6040),
.Y(n_6637)
);

INVx1_ASAP7_75t_L g6638 ( 
.A(n_6040),
.Y(n_6638)
);

INVx2_ASAP7_75t_SL g6639 ( 
.A(n_6058),
.Y(n_6639)
);

INVx1_ASAP7_75t_L g6640 ( 
.A(n_6074),
.Y(n_6640)
);

AND2x2_ASAP7_75t_L g6641 ( 
.A(n_6242),
.B(n_5947),
.Y(n_6641)
);

INVx3_ASAP7_75t_L g6642 ( 
.A(n_6283),
.Y(n_6642)
);

INVx2_ASAP7_75t_L g6643 ( 
.A(n_6041),
.Y(n_6643)
);

INVx1_ASAP7_75t_L g6644 ( 
.A(n_6074),
.Y(n_6644)
);

INVx1_ASAP7_75t_L g6645 ( 
.A(n_6077),
.Y(n_6645)
);

AND2x2_ASAP7_75t_L g6646 ( 
.A(n_6214),
.B(n_5947),
.Y(n_6646)
);

INVx3_ASAP7_75t_L g6647 ( 
.A(n_6283),
.Y(n_6647)
);

NAND2xp5_ASAP7_75t_L g6648 ( 
.A(n_6277),
.B(n_5494),
.Y(n_6648)
);

INVx2_ASAP7_75t_L g6649 ( 
.A(n_6048),
.Y(n_6649)
);

NAND2xp5_ASAP7_75t_L g6650 ( 
.A(n_6281),
.B(n_5494),
.Y(n_6650)
);

INVx3_ASAP7_75t_L g6651 ( 
.A(n_6363),
.Y(n_6651)
);

AND2x4_ASAP7_75t_L g6652 ( 
.A(n_6165),
.B(n_5877),
.Y(n_6652)
);

AND2x2_ASAP7_75t_L g6653 ( 
.A(n_6214),
.B(n_5963),
.Y(n_6653)
);

AND2x4_ASAP7_75t_L g6654 ( 
.A(n_6165),
.B(n_6217),
.Y(n_6654)
);

AND2x6_ASAP7_75t_L g6655 ( 
.A(n_6137),
.B(n_5515),
.Y(n_6655)
);

HB1xp67_ASAP7_75t_L g6656 ( 
.A(n_6307),
.Y(n_6656)
);

AND2x2_ASAP7_75t_L g6657 ( 
.A(n_6218),
.B(n_5963),
.Y(n_6657)
);

HB1xp67_ASAP7_75t_L g6658 ( 
.A(n_6309),
.Y(n_6658)
);

NAND2xp5_ASAP7_75t_L g6659 ( 
.A(n_6313),
.B(n_5468),
.Y(n_6659)
);

AND2x2_ASAP7_75t_L g6660 ( 
.A(n_6218),
.B(n_5587),
.Y(n_6660)
);

INVxp67_ASAP7_75t_SL g6661 ( 
.A(n_6080),
.Y(n_6661)
);

INVx1_ASAP7_75t_L g6662 ( 
.A(n_6077),
.Y(n_6662)
);

INVx2_ASAP7_75t_L g6663 ( 
.A(n_6048),
.Y(n_6663)
);

AND2x2_ASAP7_75t_L g6664 ( 
.A(n_6029),
.B(n_5587),
.Y(n_6664)
);

INVx1_ASAP7_75t_L g6665 ( 
.A(n_6193),
.Y(n_6665)
);

AND2x2_ASAP7_75t_L g6666 ( 
.A(n_6029),
.B(n_5671),
.Y(n_6666)
);

OR2x2_ASAP7_75t_L g6667 ( 
.A(n_6078),
.B(n_6474),
.Y(n_6667)
);

OAI22xp33_ASAP7_75t_L g6668 ( 
.A1(n_6369),
.A2(n_6168),
.B1(n_6222),
.B2(n_6212),
.Y(n_6668)
);

BUFx3_ASAP7_75t_L g6669 ( 
.A(n_6293),
.Y(n_6669)
);

INVx11_ASAP7_75t_L g6670 ( 
.A(n_6527),
.Y(n_6670)
);

INVx2_ASAP7_75t_L g6671 ( 
.A(n_6148),
.Y(n_6671)
);

INVx1_ASAP7_75t_L g6672 ( 
.A(n_6193),
.Y(n_6672)
);

INVx2_ASAP7_75t_L g6673 ( 
.A(n_6148),
.Y(n_6673)
);

INVx1_ASAP7_75t_L g6674 ( 
.A(n_6196),
.Y(n_6674)
);

INVx2_ASAP7_75t_SL g6675 ( 
.A(n_6137),
.Y(n_6675)
);

INVx1_ASAP7_75t_L g6676 ( 
.A(n_6196),
.Y(n_6676)
);

BUFx3_ASAP7_75t_L g6677 ( 
.A(n_6293),
.Y(n_6677)
);

INVx2_ASAP7_75t_L g6678 ( 
.A(n_6148),
.Y(n_6678)
);

HB1xp67_ASAP7_75t_L g6679 ( 
.A(n_6348),
.Y(n_6679)
);

INVx1_ASAP7_75t_L g6680 ( 
.A(n_6199),
.Y(n_6680)
);

AND2x4_ASAP7_75t_L g6681 ( 
.A(n_6165),
.B(n_5877),
.Y(n_6681)
);

OAI22xp33_ASAP7_75t_L g6682 ( 
.A1(n_6120),
.A2(n_5727),
.B1(n_5629),
.B2(n_5990),
.Y(n_6682)
);

INVx1_ASAP7_75t_L g6683 ( 
.A(n_6199),
.Y(n_6683)
);

INVx1_ASAP7_75t_L g6684 ( 
.A(n_6200),
.Y(n_6684)
);

NOR2xp33_ASAP7_75t_L g6685 ( 
.A(n_6037),
.B(n_5568),
.Y(n_6685)
);

INVx1_ASAP7_75t_L g6686 ( 
.A(n_6200),
.Y(n_6686)
);

AND2x4_ASAP7_75t_L g6687 ( 
.A(n_6217),
.B(n_5884),
.Y(n_6687)
);

OR2x2_ASAP7_75t_L g6688 ( 
.A(n_6078),
.B(n_4632),
.Y(n_6688)
);

INVx2_ASAP7_75t_L g6689 ( 
.A(n_6087),
.Y(n_6689)
);

BUFx3_ASAP7_75t_L g6690 ( 
.A(n_6324),
.Y(n_6690)
);

INVx2_ASAP7_75t_L g6691 ( 
.A(n_6087),
.Y(n_6691)
);

AND2x2_ASAP7_75t_L g6692 ( 
.A(n_6428),
.B(n_5671),
.Y(n_6692)
);

AND2x2_ASAP7_75t_L g6693 ( 
.A(n_6428),
.B(n_5678),
.Y(n_6693)
);

INVx1_ASAP7_75t_L g6694 ( 
.A(n_6201),
.Y(n_6694)
);

INVx1_ASAP7_75t_L g6695 ( 
.A(n_6201),
.Y(n_6695)
);

NAND2xp5_ASAP7_75t_L g6696 ( 
.A(n_6365),
.B(n_5468),
.Y(n_6696)
);

OA21x2_ASAP7_75t_L g6697 ( 
.A1(n_6337),
.A2(n_5882),
.B(n_5880),
.Y(n_6697)
);

HB1xp67_ASAP7_75t_L g6698 ( 
.A(n_6366),
.Y(n_6698)
);

AND2x4_ASAP7_75t_L g6699 ( 
.A(n_6217),
.B(n_5884),
.Y(n_6699)
);

INVx1_ASAP7_75t_L g6700 ( 
.A(n_6204),
.Y(n_6700)
);

INVx1_ASAP7_75t_L g6701 ( 
.A(n_6204),
.Y(n_6701)
);

OR2x2_ASAP7_75t_L g6702 ( 
.A(n_6474),
.B(n_4632),
.Y(n_6702)
);

INVx2_ASAP7_75t_SL g6703 ( 
.A(n_6137),
.Y(n_6703)
);

INVx2_ASAP7_75t_L g6704 ( 
.A(n_6091),
.Y(n_6704)
);

INVx2_ASAP7_75t_L g6705 ( 
.A(n_6091),
.Y(n_6705)
);

INVx2_ASAP7_75t_L g6706 ( 
.A(n_6094),
.Y(n_6706)
);

HB1xp67_ASAP7_75t_L g6707 ( 
.A(n_6405),
.Y(n_6707)
);

AND2x2_ASAP7_75t_L g6708 ( 
.A(n_6434),
.B(n_5678),
.Y(n_6708)
);

AND2x2_ASAP7_75t_L g6709 ( 
.A(n_6434),
.B(n_5468),
.Y(n_6709)
);

OR2x2_ASAP7_75t_L g6710 ( 
.A(n_6538),
.B(n_4649),
.Y(n_6710)
);

AND2x2_ASAP7_75t_L g6711 ( 
.A(n_6230),
.B(n_6254),
.Y(n_6711)
);

INVx1_ASAP7_75t_L g6712 ( 
.A(n_6206),
.Y(n_6712)
);

AND2x4_ASAP7_75t_L g6713 ( 
.A(n_6230),
.B(n_5984),
.Y(n_6713)
);

INVxp67_ASAP7_75t_SL g6714 ( 
.A(n_6094),
.Y(n_6714)
);

INVx2_ASAP7_75t_SL g6715 ( 
.A(n_6177),
.Y(n_6715)
);

AND2x2_ASAP7_75t_L g6716 ( 
.A(n_6230),
.B(n_5468),
.Y(n_6716)
);

INVx2_ASAP7_75t_L g6717 ( 
.A(n_6068),
.Y(n_6717)
);

HB1xp67_ASAP7_75t_L g6718 ( 
.A(n_6415),
.Y(n_6718)
);

AOI22xp33_ASAP7_75t_L g6719 ( 
.A1(n_6116),
.A2(n_5325),
.B1(n_5254),
.B2(n_5809),
.Y(n_6719)
);

AND2x2_ASAP7_75t_L g6720 ( 
.A(n_6254),
.B(n_5468),
.Y(n_6720)
);

OR2x2_ASAP7_75t_L g6721 ( 
.A(n_6538),
.B(n_4649),
.Y(n_6721)
);

INVx2_ASAP7_75t_L g6722 ( 
.A(n_6068),
.Y(n_6722)
);

INVx1_ASAP7_75t_L g6723 ( 
.A(n_6206),
.Y(n_6723)
);

AND2x2_ASAP7_75t_L g6724 ( 
.A(n_6254),
.B(n_5454),
.Y(n_6724)
);

AND2x2_ASAP7_75t_L g6725 ( 
.A(n_6015),
.B(n_5461),
.Y(n_6725)
);

INVx2_ASAP7_75t_SL g6726 ( 
.A(n_6549),
.Y(n_6726)
);

AND2x2_ASAP7_75t_L g6727 ( 
.A(n_6015),
.B(n_5461),
.Y(n_6727)
);

NAND2xp5_ASAP7_75t_L g6728 ( 
.A(n_6430),
.B(n_5496),
.Y(n_6728)
);

INVx3_ASAP7_75t_L g6729 ( 
.A(n_6363),
.Y(n_6729)
);

INVx2_ASAP7_75t_L g6730 ( 
.A(n_6068),
.Y(n_6730)
);

NAND2xp5_ASAP7_75t_L g6731 ( 
.A(n_6456),
.B(n_5783),
.Y(n_6731)
);

INVx1_ASAP7_75t_L g6732 ( 
.A(n_6210),
.Y(n_6732)
);

INVx1_ASAP7_75t_SL g6733 ( 
.A(n_6324),
.Y(n_6733)
);

INVx2_ASAP7_75t_L g6734 ( 
.A(n_6068),
.Y(n_6734)
);

INVx2_ASAP7_75t_L g6735 ( 
.A(n_6068),
.Y(n_6735)
);

AOI22xp33_ASAP7_75t_L g6736 ( 
.A1(n_6116),
.A2(n_5325),
.B1(n_5254),
.B2(n_5809),
.Y(n_6736)
);

AND2x2_ASAP7_75t_L g6737 ( 
.A(n_6022),
.B(n_5461),
.Y(n_6737)
);

AND2x2_ASAP7_75t_L g6738 ( 
.A(n_6022),
.B(n_5461),
.Y(n_6738)
);

AND2x4_ASAP7_75t_SL g6739 ( 
.A(n_6208),
.B(n_5568),
.Y(n_6739)
);

NOR2xp33_ASAP7_75t_L g6740 ( 
.A(n_6161),
.B(n_5568),
.Y(n_6740)
);

NAND2xp5_ASAP7_75t_L g6741 ( 
.A(n_6475),
.B(n_5506),
.Y(n_6741)
);

INVx1_ASAP7_75t_L g6742 ( 
.A(n_6210),
.Y(n_6742)
);

AND2x2_ASAP7_75t_L g6743 ( 
.A(n_6556),
.B(n_6024),
.Y(n_6743)
);

INVx2_ASAP7_75t_L g6744 ( 
.A(n_6146),
.Y(n_6744)
);

INVx1_ASAP7_75t_L g6745 ( 
.A(n_6216),
.Y(n_6745)
);

HB1xp67_ASAP7_75t_L g6746 ( 
.A(n_6503),
.Y(n_6746)
);

AND2x2_ASAP7_75t_L g6747 ( 
.A(n_6556),
.B(n_5712),
.Y(n_6747)
);

BUFx3_ASAP7_75t_L g6748 ( 
.A(n_6332),
.Y(n_6748)
);

INVx1_ASAP7_75t_L g6749 ( 
.A(n_6216),
.Y(n_6749)
);

AND2x2_ASAP7_75t_L g6750 ( 
.A(n_6024),
.B(n_5712),
.Y(n_6750)
);

INVx3_ASAP7_75t_L g6751 ( 
.A(n_6363),
.Y(n_6751)
);

AOI221xp5_ASAP7_75t_L g6752 ( 
.A1(n_6455),
.A2(n_5898),
.B1(n_5544),
.B2(n_5734),
.C(n_5739),
.Y(n_6752)
);

AND2x2_ASAP7_75t_L g6753 ( 
.A(n_6075),
.B(n_5758),
.Y(n_6753)
);

NAND3xp33_ASAP7_75t_L g6754 ( 
.A(n_6425),
.B(n_5644),
.C(n_5984),
.Y(n_6754)
);

INVx2_ASAP7_75t_L g6755 ( 
.A(n_6146),
.Y(n_6755)
);

INVx2_ASAP7_75t_L g6756 ( 
.A(n_6146),
.Y(n_6756)
);

AOI22xp5_ASAP7_75t_L g6757 ( 
.A1(n_6116),
.A2(n_5904),
.B1(n_5325),
.B2(n_5254),
.Y(n_6757)
);

AND2x2_ASAP7_75t_L g6758 ( 
.A(n_6075),
.B(n_5758),
.Y(n_6758)
);

AND2x2_ASAP7_75t_L g6759 ( 
.A(n_6247),
.B(n_5762),
.Y(n_6759)
);

INVx1_ASAP7_75t_L g6760 ( 
.A(n_6232),
.Y(n_6760)
);

AND2x2_ASAP7_75t_L g6761 ( 
.A(n_6247),
.B(n_5762),
.Y(n_6761)
);

OR2x2_ASAP7_75t_L g6762 ( 
.A(n_6553),
.B(n_4665),
.Y(n_6762)
);

INVx2_ASAP7_75t_L g6763 ( 
.A(n_6098),
.Y(n_6763)
);

NAND2xp5_ASAP7_75t_L g6764 ( 
.A(n_6317),
.B(n_5459),
.Y(n_6764)
);

NAND2xp5_ASAP7_75t_L g6765 ( 
.A(n_6317),
.B(n_5459),
.Y(n_6765)
);

INVx1_ASAP7_75t_L g6766 ( 
.A(n_6232),
.Y(n_6766)
);

OR2x6_ASAP7_75t_L g6767 ( 
.A(n_6115),
.B(n_5568),
.Y(n_6767)
);

INVx1_ASAP7_75t_L g6768 ( 
.A(n_6325),
.Y(n_6768)
);

AND2x2_ASAP7_75t_L g6769 ( 
.A(n_6529),
.B(n_5772),
.Y(n_6769)
);

AND2x2_ASAP7_75t_L g6770 ( 
.A(n_6529),
.B(n_5772),
.Y(n_6770)
);

AND2x2_ASAP7_75t_L g6771 ( 
.A(n_6461),
.B(n_5549),
.Y(n_6771)
);

INVx2_ASAP7_75t_L g6772 ( 
.A(n_6098),
.Y(n_6772)
);

BUFx6f_ASAP7_75t_L g6773 ( 
.A(n_6096),
.Y(n_6773)
);

OR2x2_ASAP7_75t_L g6774 ( 
.A(n_6553),
.B(n_4665),
.Y(n_6774)
);

INVx2_ASAP7_75t_L g6775 ( 
.A(n_6098),
.Y(n_6775)
);

INVx2_ASAP7_75t_L g6776 ( 
.A(n_6098),
.Y(n_6776)
);

HB1xp67_ASAP7_75t_L g6777 ( 
.A(n_6327),
.Y(n_6777)
);

AND2x2_ASAP7_75t_L g6778 ( 
.A(n_6461),
.B(n_5603),
.Y(n_6778)
);

AND2x4_ASAP7_75t_L g6779 ( 
.A(n_6167),
.B(n_5984),
.Y(n_6779)
);

BUFx6f_ASAP7_75t_L g6780 ( 
.A(n_6124),
.Y(n_6780)
);

AND2x2_ASAP7_75t_L g6781 ( 
.A(n_6480),
.B(n_5603),
.Y(n_6781)
);

AND2x2_ASAP7_75t_L g6782 ( 
.A(n_6480),
.B(n_5432),
.Y(n_6782)
);

AND2x2_ASAP7_75t_SL g6783 ( 
.A(n_6421),
.B(n_5984),
.Y(n_6783)
);

AND2x4_ASAP7_75t_L g6784 ( 
.A(n_6167),
.B(n_5936),
.Y(n_6784)
);

INVx1_ASAP7_75t_SL g6785 ( 
.A(n_6332),
.Y(n_6785)
);

AO31x2_ASAP7_75t_L g6786 ( 
.A1(n_6049),
.A2(n_5735),
.A3(n_5739),
.B(n_5734),
.Y(n_6786)
);

INVxp67_ASAP7_75t_SL g6787 ( 
.A(n_6016),
.Y(n_6787)
);

AOI22xp33_ASAP7_75t_L g6788 ( 
.A1(n_6088),
.A2(n_5325),
.B1(n_5070),
.B2(n_5252),
.Y(n_6788)
);

INVx2_ASAP7_75t_L g6789 ( 
.A(n_6098),
.Y(n_6789)
);

INVx1_ASAP7_75t_L g6790 ( 
.A(n_6325),
.Y(n_6790)
);

INVx3_ASAP7_75t_L g6791 ( 
.A(n_6349),
.Y(n_6791)
);

AOI22xp33_ASAP7_75t_SL g6792 ( 
.A1(n_6088),
.A2(n_5898),
.B1(n_4404),
.B2(n_4736),
.Y(n_6792)
);

AND2x4_ASAP7_75t_L g6793 ( 
.A(n_6167),
.B(n_6327),
.Y(n_6793)
);

INVx4_ASAP7_75t_L g6794 ( 
.A(n_6226),
.Y(n_6794)
);

INVx2_ASAP7_75t_L g6795 ( 
.A(n_6291),
.Y(n_6795)
);

INVx2_ASAP7_75t_L g6796 ( 
.A(n_6291),
.Y(n_6796)
);

INVx3_ASAP7_75t_L g6797 ( 
.A(n_6349),
.Y(n_6797)
);

INVx2_ASAP7_75t_L g6798 ( 
.A(n_6291),
.Y(n_6798)
);

INVx1_ASAP7_75t_L g6799 ( 
.A(n_6431),
.Y(n_6799)
);

AND2x2_ASAP7_75t_L g6800 ( 
.A(n_6519),
.B(n_5432),
.Y(n_6800)
);

HB1xp67_ASAP7_75t_L g6801 ( 
.A(n_6342),
.Y(n_6801)
);

INVx1_ASAP7_75t_L g6802 ( 
.A(n_6431),
.Y(n_6802)
);

INVx1_ASAP7_75t_L g6803 ( 
.A(n_6437),
.Y(n_6803)
);

INVx2_ASAP7_75t_L g6804 ( 
.A(n_6302),
.Y(n_6804)
);

BUFx2_ASAP7_75t_L g6805 ( 
.A(n_6159),
.Y(n_6805)
);

INVx1_ASAP7_75t_L g6806 ( 
.A(n_6437),
.Y(n_6806)
);

AND2x4_ASAP7_75t_SL g6807 ( 
.A(n_6208),
.B(n_5568),
.Y(n_6807)
);

AND2x2_ASAP7_75t_L g6808 ( 
.A(n_6519),
.B(n_5434),
.Y(n_6808)
);

INVx5_ASAP7_75t_SL g6809 ( 
.A(n_6226),
.Y(n_6809)
);

AND2x4_ASAP7_75t_L g6810 ( 
.A(n_6167),
.B(n_5936),
.Y(n_6810)
);

AND2x2_ASAP7_75t_L g6811 ( 
.A(n_6509),
.B(n_5434),
.Y(n_6811)
);

INVx2_ASAP7_75t_L g6812 ( 
.A(n_6302),
.Y(n_6812)
);

AND2x2_ASAP7_75t_L g6813 ( 
.A(n_6509),
.B(n_5742),
.Y(n_6813)
);

AND2x2_ASAP7_75t_L g6814 ( 
.A(n_6296),
.B(n_5801),
.Y(n_6814)
);

INVx2_ASAP7_75t_L g6815 ( 
.A(n_6302),
.Y(n_6815)
);

INVx1_ASAP7_75t_L g6816 ( 
.A(n_6443),
.Y(n_6816)
);

INVx1_ASAP7_75t_L g6817 ( 
.A(n_6443),
.Y(n_6817)
);

INVx2_ASAP7_75t_SL g6818 ( 
.A(n_6527),
.Y(n_6818)
);

HB1xp67_ASAP7_75t_L g6819 ( 
.A(n_6342),
.Y(n_6819)
);

INVxp67_ASAP7_75t_L g6820 ( 
.A(n_6450),
.Y(n_6820)
);

OR2x2_ASAP7_75t_L g6821 ( 
.A(n_6554),
.B(n_4668),
.Y(n_6821)
);

OR2x2_ASAP7_75t_L g6822 ( 
.A(n_6554),
.B(n_4668),
.Y(n_6822)
);

INVx1_ASAP7_75t_L g6823 ( 
.A(n_6445),
.Y(n_6823)
);

INVx2_ASAP7_75t_L g6824 ( 
.A(n_6084),
.Y(n_6824)
);

INVx1_ASAP7_75t_L g6825 ( 
.A(n_6445),
.Y(n_6825)
);

INVx2_ASAP7_75t_L g6826 ( 
.A(n_6084),
.Y(n_6826)
);

NAND2xp5_ASAP7_75t_L g6827 ( 
.A(n_6372),
.B(n_5459),
.Y(n_6827)
);

HB1xp67_ASAP7_75t_L g6828 ( 
.A(n_6372),
.Y(n_6828)
);

INVx1_ASAP7_75t_L g6829 ( 
.A(n_6447),
.Y(n_6829)
);

AND2x2_ASAP7_75t_L g6830 ( 
.A(n_6296),
.B(n_5801),
.Y(n_6830)
);

AND2x2_ASAP7_75t_L g6831 ( 
.A(n_6304),
.B(n_5552),
.Y(n_6831)
);

INVx1_ASAP7_75t_L g6832 ( 
.A(n_6447),
.Y(n_6832)
);

INVx1_ASAP7_75t_L g6833 ( 
.A(n_6448),
.Y(n_6833)
);

INVx3_ASAP7_75t_L g6834 ( 
.A(n_6136),
.Y(n_6834)
);

INVx1_ASAP7_75t_L g6835 ( 
.A(n_6448),
.Y(n_6835)
);

INVx1_ASAP7_75t_L g6836 ( 
.A(n_6453),
.Y(n_6836)
);

AND2x2_ASAP7_75t_L g6837 ( 
.A(n_6304),
.B(n_5552),
.Y(n_6837)
);

NAND2xp5_ASAP7_75t_L g6838 ( 
.A(n_6496),
.B(n_5459),
.Y(n_6838)
);

NAND3xp33_ASAP7_75t_L g6839 ( 
.A(n_6466),
.B(n_5936),
.C(n_4344),
.Y(n_6839)
);

INVx3_ASAP7_75t_L g6840 ( 
.A(n_6136),
.Y(n_6840)
);

OR2x2_ASAP7_75t_L g6841 ( 
.A(n_6257),
.B(n_4669),
.Y(n_6841)
);

INVx3_ASAP7_75t_L g6842 ( 
.A(n_6441),
.Y(n_6842)
);

INVx2_ASAP7_75t_L g6843 ( 
.A(n_6084),
.Y(n_6843)
);

INVx1_ASAP7_75t_L g6844 ( 
.A(n_6453),
.Y(n_6844)
);

INVx1_ASAP7_75t_L g6845 ( 
.A(n_6457),
.Y(n_6845)
);

AND2x2_ASAP7_75t_L g6846 ( 
.A(n_6310),
.B(n_5552),
.Y(n_6846)
);

AND2x2_ASAP7_75t_L g6847 ( 
.A(n_6310),
.B(n_5145),
.Y(n_6847)
);

NOR2x1p5_ASAP7_75t_L g6848 ( 
.A(n_6255),
.B(n_5664),
.Y(n_6848)
);

OAI22xp5_ASAP7_75t_L g6849 ( 
.A1(n_6381),
.A2(n_5996),
.B1(n_5349),
.B2(n_5919),
.Y(n_6849)
);

BUFx12f_ASAP7_75t_L g6850 ( 
.A(n_6153),
.Y(n_6850)
);

INVxp67_ASAP7_75t_SL g6851 ( 
.A(n_6016),
.Y(n_6851)
);

INVx1_ASAP7_75t_L g6852 ( 
.A(n_6457),
.Y(n_6852)
);

INVx2_ASAP7_75t_L g6853 ( 
.A(n_6097),
.Y(n_6853)
);

NAND2xp5_ASAP7_75t_L g6854 ( 
.A(n_6032),
.B(n_5459),
.Y(n_6854)
);

CKINVDCx20_ASAP7_75t_R g6855 ( 
.A(n_6124),
.Y(n_6855)
);

OR2x2_ASAP7_75t_L g6856 ( 
.A(n_6257),
.B(n_4669),
.Y(n_6856)
);

INVx3_ASAP7_75t_L g6857 ( 
.A(n_6441),
.Y(n_6857)
);

NAND2xp5_ASAP7_75t_L g6858 ( 
.A(n_6032),
.B(n_6099),
.Y(n_6858)
);

INVx3_ASAP7_75t_L g6859 ( 
.A(n_6441),
.Y(n_6859)
);

HB1xp67_ASAP7_75t_L g6860 ( 
.A(n_6176),
.Y(n_6860)
);

AND2x2_ASAP7_75t_L g6861 ( 
.A(n_6545),
.B(n_6367),
.Y(n_6861)
);

AND2x2_ASAP7_75t_L g6862 ( 
.A(n_6545),
.B(n_5145),
.Y(n_6862)
);

INVx2_ASAP7_75t_L g6863 ( 
.A(n_6097),
.Y(n_6863)
);

NAND2xp5_ASAP7_75t_L g6864 ( 
.A(n_6099),
.B(n_5368),
.Y(n_6864)
);

INVx3_ASAP7_75t_L g6865 ( 
.A(n_6545),
.Y(n_6865)
);

INVx2_ASAP7_75t_L g6866 ( 
.A(n_6097),
.Y(n_6866)
);

AND2x2_ASAP7_75t_L g6867 ( 
.A(n_6367),
.B(n_5145),
.Y(n_6867)
);

NAND2xp5_ASAP7_75t_L g6868 ( 
.A(n_6069),
.B(n_5368),
.Y(n_6868)
);

INVx2_ASAP7_75t_L g6869 ( 
.A(n_6467),
.Y(n_6869)
);

BUFx2_ASAP7_75t_L g6870 ( 
.A(n_6527),
.Y(n_6870)
);

INVx1_ASAP7_75t_L g6871 ( 
.A(n_6459),
.Y(n_6871)
);

BUFx3_ASAP7_75t_L g6872 ( 
.A(n_6255),
.Y(n_6872)
);

INVx1_ASAP7_75t_SL g6873 ( 
.A(n_6364),
.Y(n_6873)
);

AND2x2_ASAP7_75t_L g6874 ( 
.A(n_6390),
.B(n_5145),
.Y(n_6874)
);

INVx3_ASAP7_75t_L g6875 ( 
.A(n_6227),
.Y(n_6875)
);

AND2x4_ASAP7_75t_L g6876 ( 
.A(n_6060),
.B(n_5621),
.Y(n_6876)
);

NAND2xp5_ASAP7_75t_L g6877 ( 
.A(n_6069),
.B(n_5997),
.Y(n_6877)
);

AND2x2_ASAP7_75t_L g6878 ( 
.A(n_6390),
.B(n_5131),
.Y(n_6878)
);

HB1xp67_ASAP7_75t_L g6879 ( 
.A(n_6176),
.Y(n_6879)
);

OR2x2_ASAP7_75t_L g6880 ( 
.A(n_6269),
.B(n_5997),
.Y(n_6880)
);

INVx2_ASAP7_75t_L g6881 ( 
.A(n_6467),
.Y(n_6881)
);

INVx3_ASAP7_75t_L g6882 ( 
.A(n_6183),
.Y(n_6882)
);

AND2x2_ASAP7_75t_L g6883 ( 
.A(n_6473),
.B(n_5131),
.Y(n_6883)
);

OAI22xp5_ASAP7_75t_L g6884 ( 
.A1(n_6147),
.A2(n_5294),
.B1(n_4737),
.B2(n_5651),
.Y(n_6884)
);

AND2x2_ASAP7_75t_L g6885 ( 
.A(n_6473),
.B(n_5131),
.Y(n_6885)
);

AND2x2_ASAP7_75t_L g6886 ( 
.A(n_6481),
.B(n_5682),
.Y(n_6886)
);

INVx1_ASAP7_75t_L g6887 ( 
.A(n_6459),
.Y(n_6887)
);

OAI22xp33_ASAP7_75t_L g6888 ( 
.A1(n_6376),
.A2(n_5629),
.B1(n_5192),
.B2(n_4737),
.Y(n_6888)
);

AND2x2_ASAP7_75t_L g6889 ( 
.A(n_6481),
.B(n_5682),
.Y(n_6889)
);

AND2x2_ASAP7_75t_L g6890 ( 
.A(n_6504),
.B(n_5682),
.Y(n_6890)
);

INVx1_ASAP7_75t_L g6891 ( 
.A(n_6462),
.Y(n_6891)
);

INVx1_ASAP7_75t_L g6892 ( 
.A(n_6462),
.Y(n_6892)
);

AND2x2_ASAP7_75t_L g6893 ( 
.A(n_6504),
.B(n_5682),
.Y(n_6893)
);

INVx1_ASAP7_75t_L g6894 ( 
.A(n_6017),
.Y(n_6894)
);

BUFx3_ASAP7_75t_L g6895 ( 
.A(n_6153),
.Y(n_6895)
);

INVx2_ASAP7_75t_L g6896 ( 
.A(n_6467),
.Y(n_6896)
);

AND2x4_ASAP7_75t_L g6897 ( 
.A(n_6060),
.B(n_5621),
.Y(n_6897)
);

INVx2_ASAP7_75t_L g6898 ( 
.A(n_6306),
.Y(n_6898)
);

INVx2_ASAP7_75t_L g6899 ( 
.A(n_6306),
.Y(n_6899)
);

INVx2_ASAP7_75t_L g6900 ( 
.A(n_6306),
.Y(n_6900)
);

INVx1_ASAP7_75t_L g6901 ( 
.A(n_6019),
.Y(n_6901)
);

NAND2xp5_ASAP7_75t_L g6902 ( 
.A(n_6260),
.B(n_6007),
.Y(n_6902)
);

INVx3_ASAP7_75t_L g6903 ( 
.A(n_6183),
.Y(n_6903)
);

OAI33xp33_ASAP7_75t_L g6904 ( 
.A1(n_6346),
.A2(n_5933),
.A3(n_6005),
.B1(n_5743),
.B2(n_5735),
.B3(n_5751),
.Y(n_6904)
);

AND2x2_ASAP7_75t_L g6905 ( 
.A(n_6256),
.B(n_5682),
.Y(n_6905)
);

INVx1_ASAP7_75t_L g6906 ( 
.A(n_6020),
.Y(n_6906)
);

NOR2xp67_ASAP7_75t_L g6907 ( 
.A(n_6491),
.B(n_5718),
.Y(n_6907)
);

AOI221xp5_ASAP7_75t_L g6908 ( 
.A1(n_6478),
.A2(n_5744),
.B1(n_5751),
.B2(n_5743),
.C(n_5740),
.Y(n_6908)
);

NAND2xp5_ASAP7_75t_L g6909 ( 
.A(n_6043),
.B(n_5982),
.Y(n_6909)
);

INVx1_ASAP7_75t_L g6910 ( 
.A(n_6025),
.Y(n_6910)
);

INVx2_ASAP7_75t_L g6911 ( 
.A(n_6320),
.Y(n_6911)
);

INVx2_ASAP7_75t_L g6912 ( 
.A(n_6320),
.Y(n_6912)
);

INVx3_ASAP7_75t_L g6913 ( 
.A(n_6183),
.Y(n_6913)
);

INVx2_ASAP7_75t_L g6914 ( 
.A(n_6320),
.Y(n_6914)
);

INVx2_ASAP7_75t_L g6915 ( 
.A(n_6330),
.Y(n_6915)
);

AND2x2_ASAP7_75t_L g6916 ( 
.A(n_6256),
.B(n_5967),
.Y(n_6916)
);

INVx3_ASAP7_75t_L g6917 ( 
.A(n_6236),
.Y(n_6917)
);

BUFx6f_ASAP7_75t_L g6918 ( 
.A(n_6227),
.Y(n_6918)
);

HB1xp67_ASAP7_75t_L g6919 ( 
.A(n_6318),
.Y(n_6919)
);

NAND2xp5_ASAP7_75t_L g6920 ( 
.A(n_6043),
.B(n_5982),
.Y(n_6920)
);

INVxp67_ASAP7_75t_L g6921 ( 
.A(n_6316),
.Y(n_6921)
);

INVx1_ASAP7_75t_L g6922 ( 
.A(n_6030),
.Y(n_6922)
);

OR2x2_ASAP7_75t_L g6923 ( 
.A(n_6269),
.B(n_5986),
.Y(n_6923)
);

AND2x2_ASAP7_75t_L g6924 ( 
.A(n_6258),
.B(n_5967),
.Y(n_6924)
);

INVx1_ASAP7_75t_L g6925 ( 
.A(n_6031),
.Y(n_6925)
);

BUFx3_ASAP7_75t_L g6926 ( 
.A(n_6122),
.Y(n_6926)
);

INVx2_ASAP7_75t_L g6927 ( 
.A(n_6330),
.Y(n_6927)
);

OA21x2_ASAP7_75t_L g6928 ( 
.A1(n_6049),
.A2(n_5882),
.B(n_5869),
.Y(n_6928)
);

BUFx2_ASAP7_75t_L g6929 ( 
.A(n_6426),
.Y(n_6929)
);

AND2x2_ASAP7_75t_L g6930 ( 
.A(n_6258),
.B(n_6004),
.Y(n_6930)
);

AND2x4_ASAP7_75t_L g6931 ( 
.A(n_6060),
.B(n_5643),
.Y(n_6931)
);

INVx1_ASAP7_75t_SL g6932 ( 
.A(n_6181),
.Y(n_6932)
);

AND2x2_ASAP7_75t_SL g6933 ( 
.A(n_6088),
.B(n_5084),
.Y(n_6933)
);

NOR2x1_ASAP7_75t_SL g6934 ( 
.A(n_6060),
.B(n_5106),
.Y(n_6934)
);

INVx2_ASAP7_75t_L g6935 ( 
.A(n_6330),
.Y(n_6935)
);

OR2x2_ASAP7_75t_L g6936 ( 
.A(n_6272),
.B(n_5988),
.Y(n_6936)
);

BUFx2_ASAP7_75t_L g6937 ( 
.A(n_6426),
.Y(n_6937)
);

INVx1_ASAP7_75t_SL g6938 ( 
.A(n_6188),
.Y(n_6938)
);

INVx1_ASAP7_75t_L g6939 ( 
.A(n_6033),
.Y(n_6939)
);

BUFx3_ASAP7_75t_L g6940 ( 
.A(n_6154),
.Y(n_6940)
);

INVx2_ASAP7_75t_L g6941 ( 
.A(n_6203),
.Y(n_6941)
);

NAND2xp5_ASAP7_75t_L g6942 ( 
.A(n_6051),
.B(n_5988),
.Y(n_6942)
);

INVx2_ASAP7_75t_SL g6943 ( 
.A(n_6343),
.Y(n_6943)
);

AND2x2_ASAP7_75t_L g6944 ( 
.A(n_6202),
.B(n_6004),
.Y(n_6944)
);

AND2x2_ASAP7_75t_L g6945 ( 
.A(n_6202),
.B(n_4755),
.Y(n_6945)
);

INVx1_ASAP7_75t_L g6946 ( 
.A(n_6050),
.Y(n_6946)
);

INVx2_ASAP7_75t_SL g6947 ( 
.A(n_6227),
.Y(n_6947)
);

AND2x2_ASAP7_75t_L g6948 ( 
.A(n_6311),
.B(n_4755),
.Y(n_6948)
);

BUFx2_ASAP7_75t_SL g6949 ( 
.A(n_6227),
.Y(n_6949)
);

OR2x2_ASAP7_75t_L g6950 ( 
.A(n_6272),
.B(n_5993),
.Y(n_6950)
);

INVx1_ASAP7_75t_L g6951 ( 
.A(n_6055),
.Y(n_6951)
);

OR2x2_ASAP7_75t_L g6952 ( 
.A(n_6275),
.B(n_5993),
.Y(n_6952)
);

NOR2xp33_ASAP7_75t_L g6953 ( 
.A(n_6305),
.B(n_5664),
.Y(n_6953)
);

AND2x2_ASAP7_75t_L g6954 ( 
.A(n_6311),
.B(n_4755),
.Y(n_6954)
);

AND2x2_ASAP7_75t_L g6955 ( 
.A(n_6347),
.B(n_4761),
.Y(n_6955)
);

OR2x2_ASAP7_75t_L g6956 ( 
.A(n_6275),
.B(n_6007),
.Y(n_6956)
);

INVx2_ASAP7_75t_SL g6957 ( 
.A(n_6227),
.Y(n_6957)
);

AO31x2_ASAP7_75t_L g6958 ( 
.A1(n_6059),
.A2(n_5744),
.A3(n_5754),
.B(n_5740),
.Y(n_6958)
);

BUFx2_ASAP7_75t_L g6959 ( 
.A(n_6485),
.Y(n_6959)
);

INVx1_ASAP7_75t_L g6960 ( 
.A(n_6056),
.Y(n_6960)
);

INVx2_ASAP7_75t_L g6961 ( 
.A(n_6203),
.Y(n_6961)
);

INVx1_ASAP7_75t_L g6962 ( 
.A(n_6057),
.Y(n_6962)
);

BUFx2_ASAP7_75t_L g6963 ( 
.A(n_6485),
.Y(n_6963)
);

INVx1_ASAP7_75t_L g6964 ( 
.A(n_6061),
.Y(n_6964)
);

AND2x2_ASAP7_75t_L g6965 ( 
.A(n_6379),
.B(n_4761),
.Y(n_6965)
);

INVx1_ASAP7_75t_L g6966 ( 
.A(n_6066),
.Y(n_6966)
);

INVx1_ASAP7_75t_L g6967 ( 
.A(n_6070),
.Y(n_6967)
);

INVx1_ASAP7_75t_L g6968 ( 
.A(n_6072),
.Y(n_6968)
);

AND2x2_ASAP7_75t_L g6969 ( 
.A(n_6379),
.B(n_4761),
.Y(n_6969)
);

INVx1_ASAP7_75t_L g6970 ( 
.A(n_6085),
.Y(n_6970)
);

AND2x4_ASAP7_75t_L g6971 ( 
.A(n_6101),
.B(n_5643),
.Y(n_6971)
);

NAND2xp5_ASAP7_75t_L g6972 ( 
.A(n_6051),
.B(n_6009),
.Y(n_6972)
);

INVx2_ASAP7_75t_L g6973 ( 
.A(n_6203),
.Y(n_6973)
);

AND2x2_ASAP7_75t_L g6974 ( 
.A(n_6392),
.B(n_4798),
.Y(n_6974)
);

INVx1_ASAP7_75t_L g6975 ( 
.A(n_6092),
.Y(n_6975)
);

AND2x2_ASAP7_75t_L g6976 ( 
.A(n_6392),
.B(n_4798),
.Y(n_6976)
);

NAND4xp25_ASAP7_75t_L g6977 ( 
.A(n_6400),
.B(n_5560),
.C(n_5905),
.D(n_5710),
.Y(n_6977)
);

INVx4_ASAP7_75t_L g6978 ( 
.A(n_6354),
.Y(n_6978)
);

INVx2_ASAP7_75t_L g6979 ( 
.A(n_6351),
.Y(n_6979)
);

NAND2xp5_ASAP7_75t_L g6980 ( 
.A(n_6052),
.B(n_5575),
.Y(n_6980)
);

AND2x2_ASAP7_75t_L g6981 ( 
.A(n_6490),
.B(n_4798),
.Y(n_6981)
);

INVxp67_ASAP7_75t_L g6982 ( 
.A(n_6490),
.Y(n_6982)
);

AND2x2_ASAP7_75t_L g6983 ( 
.A(n_6511),
.B(n_5665),
.Y(n_6983)
);

INVx2_ASAP7_75t_L g6984 ( 
.A(n_6351),
.Y(n_6984)
);

INVx2_ASAP7_75t_L g6985 ( 
.A(n_6351),
.Y(n_6985)
);

AND2x2_ASAP7_75t_L g6986 ( 
.A(n_6511),
.B(n_5665),
.Y(n_6986)
);

INVx1_ASAP7_75t_L g6987 ( 
.A(n_6100),
.Y(n_6987)
);

HB1xp67_ASAP7_75t_L g6988 ( 
.A(n_6319),
.Y(n_6988)
);

NAND2xp5_ASAP7_75t_L g6989 ( 
.A(n_6052),
.B(n_5977),
.Y(n_6989)
);

AOI22xp33_ASAP7_75t_SL g6990 ( 
.A1(n_6335),
.A2(n_4736),
.B1(n_4689),
.B2(n_4180),
.Y(n_6990)
);

AND2x4_ASAP7_75t_L g6991 ( 
.A(n_6101),
.B(n_5665),
.Y(n_6991)
);

INVxp67_ASAP7_75t_SL g6992 ( 
.A(n_6016),
.Y(n_6992)
);

OR2x2_ASAP7_75t_L g6993 ( 
.A(n_6528),
.B(n_5977),
.Y(n_6993)
);

AND2x2_ASAP7_75t_L g6994 ( 
.A(n_6038),
.B(n_5716),
.Y(n_6994)
);

BUFx3_ASAP7_75t_L g6995 ( 
.A(n_6402),
.Y(n_6995)
);

AND2x4_ASAP7_75t_L g6996 ( 
.A(n_6101),
.B(n_5716),
.Y(n_6996)
);

HB1xp67_ASAP7_75t_L g6997 ( 
.A(n_6394),
.Y(n_6997)
);

NAND2xp5_ASAP7_75t_L g6998 ( 
.A(n_6422),
.B(n_5979),
.Y(n_6998)
);

OR2x2_ASAP7_75t_L g6999 ( 
.A(n_6287),
.B(n_6299),
.Y(n_6999)
);

INVx1_ASAP7_75t_L g7000 ( 
.A(n_6109),
.Y(n_7000)
);

INVx1_ASAP7_75t_L g7001 ( 
.A(n_6111),
.Y(n_7001)
);

INVx1_ASAP7_75t_L g7002 ( 
.A(n_6114),
.Y(n_7002)
);

AND2x2_ASAP7_75t_L g7003 ( 
.A(n_6038),
.B(n_6438),
.Y(n_7003)
);

NOR2x1_ASAP7_75t_L g7004 ( 
.A(n_6331),
.B(n_5696),
.Y(n_7004)
);

INVx2_ASAP7_75t_L g7005 ( 
.A(n_6358),
.Y(n_7005)
);

INVxp67_ASAP7_75t_L g7006 ( 
.A(n_6380),
.Y(n_7006)
);

OA21x2_ASAP7_75t_L g7007 ( 
.A1(n_6059),
.A2(n_5869),
.B(n_5776),
.Y(n_7007)
);

INVx2_ASAP7_75t_L g7008 ( 
.A(n_6358),
.Y(n_7008)
);

OAI211xp5_ASAP7_75t_L g7009 ( 
.A1(n_6115),
.A2(n_5126),
.B(n_5136),
.C(n_5084),
.Y(n_7009)
);

BUFx2_ASAP7_75t_L g7010 ( 
.A(n_6486),
.Y(n_7010)
);

AOI22xp33_ASAP7_75t_L g7011 ( 
.A1(n_6668),
.A2(n_6335),
.B1(n_6076),
.B2(n_6081),
.Y(n_7011)
);

AND2x2_ASAP7_75t_L g7012 ( 
.A(n_6813),
.B(n_6419),
.Y(n_7012)
);

INVx2_ASAP7_75t_SL g7013 ( 
.A(n_6690),
.Y(n_7013)
);

INVx1_ASAP7_75t_L g7014 ( 
.A(n_6586),
.Y(n_7014)
);

BUFx2_ASAP7_75t_L g7015 ( 
.A(n_6690),
.Y(n_7015)
);

AND2x2_ASAP7_75t_L g7016 ( 
.A(n_6783),
.B(n_6943),
.Y(n_7016)
);

AND2x2_ASAP7_75t_L g7017 ( 
.A(n_6574),
.B(n_6419),
.Y(n_7017)
);

HB1xp67_ASAP7_75t_L g7018 ( 
.A(n_6560),
.Y(n_7018)
);

AND2x4_ASAP7_75t_L g7019 ( 
.A(n_6814),
.B(n_6486),
.Y(n_7019)
);

INVx2_ASAP7_75t_SL g7020 ( 
.A(n_6670),
.Y(n_7020)
);

INVx2_ASAP7_75t_L g7021 ( 
.A(n_6853),
.Y(n_7021)
);

INVx1_ASAP7_75t_L g7022 ( 
.A(n_6586),
.Y(n_7022)
);

AND2x2_ASAP7_75t_L g7023 ( 
.A(n_6783),
.B(n_6290),
.Y(n_7023)
);

INVx1_ASAP7_75t_L g7024 ( 
.A(n_6611),
.Y(n_7024)
);

NAND2xp5_ASAP7_75t_L g7025 ( 
.A(n_6571),
.B(n_6454),
.Y(n_7025)
);

NOR2x1_ASAP7_75t_SL g7026 ( 
.A(n_6767),
.B(n_6101),
.Y(n_7026)
);

INVx2_ASAP7_75t_L g7027 ( 
.A(n_6853),
.Y(n_7027)
);

INVx1_ASAP7_75t_L g7028 ( 
.A(n_6611),
.Y(n_7028)
);

AND2x4_ASAP7_75t_L g7029 ( 
.A(n_6830),
.B(n_6531),
.Y(n_7029)
);

AND2x2_ASAP7_75t_L g7030 ( 
.A(n_6725),
.B(n_6550),
.Y(n_7030)
);

INVx1_ASAP7_75t_L g7031 ( 
.A(n_6618),
.Y(n_7031)
);

INVx2_ASAP7_75t_L g7032 ( 
.A(n_6863),
.Y(n_7032)
);

AND2x2_ASAP7_75t_L g7033 ( 
.A(n_6943),
.B(n_6531),
.Y(n_7033)
);

AND2x2_ASAP7_75t_L g7034 ( 
.A(n_6727),
.B(n_6550),
.Y(n_7034)
);

INVx2_ASAP7_75t_L g7035 ( 
.A(n_6863),
.Y(n_7035)
);

AOI22xp33_ASAP7_75t_L g7036 ( 
.A1(n_6668),
.A2(n_6335),
.B1(n_6076),
.B2(n_6081),
.Y(n_7036)
);

AOI22xp33_ASAP7_75t_L g7037 ( 
.A1(n_6560),
.A2(n_6081),
.B1(n_6546),
.B2(n_6105),
.Y(n_7037)
);

HB1xp67_ASAP7_75t_L g7038 ( 
.A(n_6571),
.Y(n_7038)
);

AND2x2_ASAP7_75t_L g7039 ( 
.A(n_6737),
.B(n_6354),
.Y(n_7039)
);

INVx2_ASAP7_75t_L g7040 ( 
.A(n_6866),
.Y(n_7040)
);

AND2x2_ASAP7_75t_L g7041 ( 
.A(n_6738),
.B(n_6354),
.Y(n_7041)
);

BUFx3_ASAP7_75t_L g7042 ( 
.A(n_6578),
.Y(n_7042)
);

INVx2_ASAP7_75t_SL g7043 ( 
.A(n_6726),
.Y(n_7043)
);

INVx1_ASAP7_75t_L g7044 ( 
.A(n_6618),
.Y(n_7044)
);

NAND2xp5_ASAP7_75t_L g7045 ( 
.A(n_6873),
.B(n_6479),
.Y(n_7045)
);

OR2x2_ASAP7_75t_L g7046 ( 
.A(n_6999),
.B(n_6287),
.Y(n_7046)
);

AO21x2_ASAP7_75t_L g7047 ( 
.A1(n_6569),
.A2(n_6464),
.B(n_6236),
.Y(n_7047)
);

INVx1_ASAP7_75t_SL g7048 ( 
.A(n_6578),
.Y(n_7048)
);

INVx2_ASAP7_75t_L g7049 ( 
.A(n_6866),
.Y(n_7049)
);

OR2x2_ASAP7_75t_L g7050 ( 
.A(n_6667),
.B(n_6299),
.Y(n_7050)
);

HB1xp67_ASAP7_75t_L g7051 ( 
.A(n_6882),
.Y(n_7051)
);

AND2x2_ASAP7_75t_L g7052 ( 
.A(n_6567),
.B(n_6354),
.Y(n_7052)
);

BUFx2_ASAP7_75t_SL g7053 ( 
.A(n_6855),
.Y(n_7053)
);

BUFx2_ASAP7_75t_L g7054 ( 
.A(n_6850),
.Y(n_7054)
);

INVx1_ASAP7_75t_L g7055 ( 
.A(n_6656),
.Y(n_7055)
);

INVx1_ASAP7_75t_L g7056 ( 
.A(n_6656),
.Y(n_7056)
);

NOR2xp67_ASAP7_75t_L g7057 ( 
.A(n_6726),
.B(n_6508),
.Y(n_7057)
);

AND2x2_ASAP7_75t_L g7058 ( 
.A(n_6932),
.B(n_5515),
.Y(n_7058)
);

INVx2_ASAP7_75t_L g7059 ( 
.A(n_6717),
.Y(n_7059)
);

INVx2_ASAP7_75t_L g7060 ( 
.A(n_6717),
.Y(n_7060)
);

BUFx6f_ASAP7_75t_L g7061 ( 
.A(n_6605),
.Y(n_7061)
);

INVx2_ASAP7_75t_L g7062 ( 
.A(n_6722),
.Y(n_7062)
);

INVx2_ASAP7_75t_L g7063 ( 
.A(n_6722),
.Y(n_7063)
);

BUFx2_ASAP7_75t_L g7064 ( 
.A(n_6850),
.Y(n_7064)
);

INVx2_ASAP7_75t_L g7065 ( 
.A(n_6730),
.Y(n_7065)
);

INVx2_ASAP7_75t_L g7066 ( 
.A(n_6730),
.Y(n_7066)
);

INVx1_ASAP7_75t_L g7067 ( 
.A(n_6658),
.Y(n_7067)
);

INVx2_ASAP7_75t_L g7068 ( 
.A(n_6734),
.Y(n_7068)
);

BUFx2_ASAP7_75t_L g7069 ( 
.A(n_6582),
.Y(n_7069)
);

INVx2_ASAP7_75t_L g7070 ( 
.A(n_6734),
.Y(n_7070)
);

INVx2_ASAP7_75t_L g7071 ( 
.A(n_6735),
.Y(n_7071)
);

AND2x2_ASAP7_75t_L g7072 ( 
.A(n_6573),
.B(n_6354),
.Y(n_7072)
);

HB1xp67_ASAP7_75t_L g7073 ( 
.A(n_6882),
.Y(n_7073)
);

AND2x2_ASAP7_75t_L g7074 ( 
.A(n_6861),
.B(n_6331),
.Y(n_7074)
);

HB1xp67_ASAP7_75t_L g7075 ( 
.A(n_6882),
.Y(n_7075)
);

AND2x2_ASAP7_75t_L g7076 ( 
.A(n_6944),
.B(n_6331),
.Y(n_7076)
);

BUFx2_ASAP7_75t_L g7077 ( 
.A(n_6582),
.Y(n_7077)
);

INVx1_ASAP7_75t_L g7078 ( 
.A(n_6658),
.Y(n_7078)
);

AND2x4_ASAP7_75t_L g7079 ( 
.A(n_6793),
.B(n_6380),
.Y(n_7079)
);

AND2x2_ASAP7_75t_L g7080 ( 
.A(n_6916),
.B(n_6044),
.Y(n_7080)
);

AND2x2_ASAP7_75t_L g7081 ( 
.A(n_6938),
.B(n_5515),
.Y(n_7081)
);

INVx1_ASAP7_75t_L g7082 ( 
.A(n_6679),
.Y(n_7082)
);

INVx1_ASAP7_75t_L g7083 ( 
.A(n_6679),
.Y(n_7083)
);

CKINVDCx20_ASAP7_75t_R g7084 ( 
.A(n_6855),
.Y(n_7084)
);

INVx1_ASAP7_75t_L g7085 ( 
.A(n_6698),
.Y(n_7085)
);

INVx1_ASAP7_75t_L g7086 ( 
.A(n_6698),
.Y(n_7086)
);

BUFx3_ASAP7_75t_L g7087 ( 
.A(n_6605),
.Y(n_7087)
);

NAND2xp5_ASAP7_75t_L g7088 ( 
.A(n_6584),
.B(n_6487),
.Y(n_7088)
);

AND2x2_ASAP7_75t_L g7089 ( 
.A(n_6924),
.B(n_5515),
.Y(n_7089)
);

AND2x4_ASAP7_75t_SL g7090 ( 
.A(n_6930),
.B(n_6502),
.Y(n_7090)
);

HB1xp67_ASAP7_75t_L g7091 ( 
.A(n_6903),
.Y(n_7091)
);

INVx1_ASAP7_75t_L g7092 ( 
.A(n_6707),
.Y(n_7092)
);

INVx1_ASAP7_75t_L g7093 ( 
.A(n_6707),
.Y(n_7093)
);

INVx1_ASAP7_75t_L g7094 ( 
.A(n_6718),
.Y(n_7094)
);

BUFx3_ASAP7_75t_L g7095 ( 
.A(n_6626),
.Y(n_7095)
);

AND2x2_ASAP7_75t_L g7096 ( 
.A(n_7003),
.B(n_5696),
.Y(n_7096)
);

AND2x2_ASAP7_75t_L g7097 ( 
.A(n_6646),
.B(n_5710),
.Y(n_7097)
);

INVx1_ASAP7_75t_L g7098 ( 
.A(n_6718),
.Y(n_7098)
);

BUFx3_ASAP7_75t_L g7099 ( 
.A(n_6626),
.Y(n_7099)
);

NAND2xp5_ASAP7_75t_L g7100 ( 
.A(n_6733),
.B(n_6027),
.Y(n_7100)
);

INVx2_ASAP7_75t_L g7101 ( 
.A(n_6735),
.Y(n_7101)
);

INVx1_ASAP7_75t_L g7102 ( 
.A(n_6746),
.Y(n_7102)
);

AND2x2_ASAP7_75t_L g7103 ( 
.A(n_6653),
.B(n_5775),
.Y(n_7103)
);

INVx1_ASAP7_75t_L g7104 ( 
.A(n_6746),
.Y(n_7104)
);

INVx3_ASAP7_75t_L g7105 ( 
.A(n_6595),
.Y(n_7105)
);

AND2x2_ASAP7_75t_L g7106 ( 
.A(n_6570),
.B(n_6044),
.Y(n_7106)
);

BUFx2_ASAP7_75t_L g7107 ( 
.A(n_6628),
.Y(n_7107)
);

INVx2_ASAP7_75t_L g7108 ( 
.A(n_6763),
.Y(n_7108)
);

INVx1_ASAP7_75t_L g7109 ( 
.A(n_6615),
.Y(n_7109)
);

INVx1_ASAP7_75t_L g7110 ( 
.A(n_6615),
.Y(n_7110)
);

HB1xp67_ASAP7_75t_L g7111 ( 
.A(n_6903),
.Y(n_7111)
);

HB1xp67_ASAP7_75t_L g7112 ( 
.A(n_6903),
.Y(n_7112)
);

INVx1_ASAP7_75t_L g7113 ( 
.A(n_6777),
.Y(n_7113)
);

OR2x2_ASAP7_75t_L g7114 ( 
.A(n_6601),
.B(n_6413),
.Y(n_7114)
);

HB1xp67_ASAP7_75t_L g7115 ( 
.A(n_6913),
.Y(n_7115)
);

OR2x2_ASAP7_75t_L g7116 ( 
.A(n_6598),
.B(n_6858),
.Y(n_7116)
);

INVx1_ASAP7_75t_L g7117 ( 
.A(n_6777),
.Y(n_7117)
);

AND2x4_ASAP7_75t_L g7118 ( 
.A(n_6793),
.B(n_6386),
.Y(n_7118)
);

INVx2_ASAP7_75t_L g7119 ( 
.A(n_6763),
.Y(n_7119)
);

OR2x2_ASAP7_75t_L g7120 ( 
.A(n_6841),
.B(n_6413),
.Y(n_7120)
);

INVxp67_ASAP7_75t_L g7121 ( 
.A(n_6685),
.Y(n_7121)
);

AND2x2_ASAP7_75t_L g7122 ( 
.A(n_6570),
.B(n_6657),
.Y(n_7122)
);

INVx1_ASAP7_75t_L g7123 ( 
.A(n_6801),
.Y(n_7123)
);

AND2x2_ASAP7_75t_L g7124 ( 
.A(n_6995),
.B(n_5775),
.Y(n_7124)
);

INVx1_ASAP7_75t_L g7125 ( 
.A(n_6801),
.Y(n_7125)
);

INVx2_ASAP7_75t_L g7126 ( 
.A(n_6772),
.Y(n_7126)
);

INVx1_ASAP7_75t_L g7127 ( 
.A(n_6819),
.Y(n_7127)
);

INVx2_ASAP7_75t_L g7128 ( 
.A(n_6772),
.Y(n_7128)
);

INVx2_ASAP7_75t_L g7129 ( 
.A(n_6775),
.Y(n_7129)
);

NOR2xp33_ASAP7_75t_L g7130 ( 
.A(n_6794),
.B(n_5841),
.Y(n_7130)
);

INVx1_ASAP7_75t_L g7131 ( 
.A(n_6819),
.Y(n_7131)
);

NAND2xp5_ASAP7_75t_L g7132 ( 
.A(n_6576),
.B(n_6027),
.Y(n_7132)
);

AND2x2_ASAP7_75t_L g7133 ( 
.A(n_6995),
.B(n_5841),
.Y(n_7133)
);

AND2x2_ASAP7_75t_L g7134 ( 
.A(n_6711),
.B(n_6412),
.Y(n_7134)
);

INVx2_ASAP7_75t_L g7135 ( 
.A(n_6775),
.Y(n_7135)
);

AND2x2_ASAP7_75t_L g7136 ( 
.A(n_6580),
.B(n_6438),
.Y(n_7136)
);

AND2x2_ASAP7_75t_L g7137 ( 
.A(n_6581),
.B(n_6442),
.Y(n_7137)
);

INVx2_ASAP7_75t_L g7138 ( 
.A(n_6776),
.Y(n_7138)
);

INVx2_ASAP7_75t_L g7139 ( 
.A(n_6776),
.Y(n_7139)
);

INVx2_ASAP7_75t_L g7140 ( 
.A(n_6789),
.Y(n_7140)
);

INVx1_ASAP7_75t_L g7141 ( 
.A(n_6828),
.Y(n_7141)
);

INVx2_ASAP7_75t_L g7142 ( 
.A(n_6789),
.Y(n_7142)
);

AO21x2_ASAP7_75t_L g7143 ( 
.A1(n_6568),
.A2(n_6464),
.B(n_6105),
.Y(n_7143)
);

OR2x2_ASAP7_75t_L g7144 ( 
.A(n_6856),
.B(n_6424),
.Y(n_7144)
);

BUFx3_ASAP7_75t_L g7145 ( 
.A(n_6628),
.Y(n_7145)
);

AND2x2_ASAP7_75t_L g7146 ( 
.A(n_6771),
.B(n_6778),
.Y(n_7146)
);

HB1xp67_ASAP7_75t_L g7147 ( 
.A(n_6913),
.Y(n_7147)
);

AND2x2_ASAP7_75t_L g7148 ( 
.A(n_6781),
.B(n_6442),
.Y(n_7148)
);

AND2x2_ASAP7_75t_L g7149 ( 
.A(n_6591),
.B(n_6444),
.Y(n_7149)
);

HB1xp67_ASAP7_75t_L g7150 ( 
.A(n_6913),
.Y(n_7150)
);

INVx2_ASAP7_75t_L g7151 ( 
.A(n_6575),
.Y(n_7151)
);

AND2x2_ASAP7_75t_L g7152 ( 
.A(n_6600),
.B(n_6444),
.Y(n_7152)
);

INVx2_ASAP7_75t_L g7153 ( 
.A(n_6575),
.Y(n_7153)
);

INVx2_ASAP7_75t_L g7154 ( 
.A(n_6592),
.Y(n_7154)
);

AND2x2_ASAP7_75t_L g7155 ( 
.A(n_6660),
.B(n_6451),
.Y(n_7155)
);

INVx2_ASAP7_75t_L g7156 ( 
.A(n_6592),
.Y(n_7156)
);

INVx2_ASAP7_75t_L g7157 ( 
.A(n_6609),
.Y(n_7157)
);

AND2x4_ASAP7_75t_L g7158 ( 
.A(n_6793),
.B(n_6386),
.Y(n_7158)
);

INVx1_ASAP7_75t_L g7159 ( 
.A(n_6828),
.Y(n_7159)
);

INVx2_ASAP7_75t_L g7160 ( 
.A(n_6609),
.Y(n_7160)
);

HB1xp67_ASAP7_75t_L g7161 ( 
.A(n_6576),
.Y(n_7161)
);

AND2x2_ASAP7_75t_L g7162 ( 
.A(n_6566),
.B(n_6047),
.Y(n_7162)
);

AOI22xp33_ASAP7_75t_L g7163 ( 
.A1(n_6839),
.A2(n_6103),
.B1(n_6028),
.B2(n_4344),
.Y(n_7163)
);

AO21x2_ASAP7_75t_L g7164 ( 
.A1(n_6838),
.A2(n_6103),
.B(n_6155),
.Y(n_7164)
);

INVx2_ASAP7_75t_SL g7165 ( 
.A(n_6848),
.Y(n_7165)
);

NAND2xp5_ASAP7_75t_L g7166 ( 
.A(n_6820),
.B(n_6452),
.Y(n_7166)
);

OR2x2_ASAP7_75t_L g7167 ( 
.A(n_6688),
.B(n_6424),
.Y(n_7167)
);

INVx5_ASAP7_75t_L g7168 ( 
.A(n_6809),
.Y(n_7168)
);

INVx1_ASAP7_75t_L g7169 ( 
.A(n_6860),
.Y(n_7169)
);

INVx2_ASAP7_75t_L g7170 ( 
.A(n_6824),
.Y(n_7170)
);

BUFx6f_ASAP7_75t_L g7171 ( 
.A(n_6625),
.Y(n_7171)
);

INVx2_ASAP7_75t_L g7172 ( 
.A(n_6824),
.Y(n_7172)
);

INVx2_ASAP7_75t_L g7173 ( 
.A(n_6826),
.Y(n_7173)
);

AND2x2_ASAP7_75t_L g7174 ( 
.A(n_6566),
.B(n_6047),
.Y(n_7174)
);

HB1xp67_ASAP7_75t_L g7175 ( 
.A(n_6820),
.Y(n_7175)
);

INVx1_ASAP7_75t_L g7176 ( 
.A(n_6860),
.Y(n_7176)
);

INVx1_ASAP7_75t_L g7177 ( 
.A(n_6879),
.Y(n_7177)
);

NOR2xp33_ASAP7_75t_SL g7178 ( 
.A(n_6785),
.B(n_6495),
.Y(n_7178)
);

OR2x2_ASAP7_75t_L g7179 ( 
.A(n_6710),
.B(n_6132),
.Y(n_7179)
);

INVx1_ASAP7_75t_L g7180 ( 
.A(n_6879),
.Y(n_7180)
);

INVx1_ASAP7_75t_L g7181 ( 
.A(n_6603),
.Y(n_7181)
);

INVx4_ASAP7_75t_L g7182 ( 
.A(n_6794),
.Y(n_7182)
);

AND2x4_ASAP7_75t_SL g7183 ( 
.A(n_6811),
.B(n_5044),
.Y(n_7183)
);

AO21x2_ASAP7_75t_L g7184 ( 
.A1(n_6764),
.A2(n_6179),
.B(n_6178),
.Y(n_7184)
);

AND2x2_ASAP7_75t_L g7185 ( 
.A(n_6566),
.B(n_6127),
.Y(n_7185)
);

AND2x2_ASAP7_75t_L g7186 ( 
.A(n_6572),
.B(n_6127),
.Y(n_7186)
);

AND2x2_ASAP7_75t_L g7187 ( 
.A(n_6572),
.B(n_6129),
.Y(n_7187)
);

NAND2xp5_ASAP7_75t_L g7188 ( 
.A(n_6919),
.B(n_6501),
.Y(n_7188)
);

AND2x2_ASAP7_75t_L g7189 ( 
.A(n_6572),
.B(n_6129),
.Y(n_7189)
);

INVx1_ASAP7_75t_L g7190 ( 
.A(n_6608),
.Y(n_7190)
);

INVx1_ASAP7_75t_L g7191 ( 
.A(n_6619),
.Y(n_7191)
);

AND2x2_ASAP7_75t_L g7192 ( 
.A(n_6635),
.B(n_6135),
.Y(n_7192)
);

AND2x2_ASAP7_75t_L g7193 ( 
.A(n_6636),
.B(n_6135),
.Y(n_7193)
);

OR2x2_ASAP7_75t_L g7194 ( 
.A(n_6721),
.B(n_6132),
.Y(n_7194)
);

BUFx6f_ASAP7_75t_L g7195 ( 
.A(n_6625),
.Y(n_7195)
);

OR2x2_ASAP7_75t_L g7196 ( 
.A(n_6762),
.B(n_6774),
.Y(n_7196)
);

INVx1_ASAP7_75t_SL g7197 ( 
.A(n_6669),
.Y(n_7197)
);

INVx1_ASAP7_75t_L g7198 ( 
.A(n_6633),
.Y(n_7198)
);

INVx2_ASAP7_75t_L g7199 ( 
.A(n_6826),
.Y(n_7199)
);

INVx1_ASAP7_75t_L g7200 ( 
.A(n_6637),
.Y(n_7200)
);

NAND2xp5_ASAP7_75t_L g7201 ( 
.A(n_6919),
.B(n_6525),
.Y(n_7201)
);

NAND2xp5_ASAP7_75t_L g7202 ( 
.A(n_6988),
.B(n_6123),
.Y(n_7202)
);

AND2x4_ASAP7_75t_L g7203 ( 
.A(n_6654),
.B(n_6387),
.Y(n_7203)
);

AND2x2_ASAP7_75t_L g7204 ( 
.A(n_6641),
.B(n_6403),
.Y(n_7204)
);

INVx2_ASAP7_75t_L g7205 ( 
.A(n_6843),
.Y(n_7205)
);

NAND2xp5_ASAP7_75t_L g7206 ( 
.A(n_6988),
.B(n_6997),
.Y(n_7206)
);

INVx2_ASAP7_75t_L g7207 ( 
.A(n_6843),
.Y(n_7207)
);

AND2x2_ASAP7_75t_L g7208 ( 
.A(n_6654),
.B(n_6403),
.Y(n_7208)
);

AND2x4_ASAP7_75t_L g7209 ( 
.A(n_6654),
.B(n_6387),
.Y(n_7209)
);

AOI22xp33_ASAP7_75t_L g7210 ( 
.A1(n_6904),
.A2(n_6028),
.B1(n_6191),
.B2(n_6190),
.Y(n_7210)
);

INVx3_ASAP7_75t_L g7211 ( 
.A(n_6767),
.Y(n_7211)
);

BUFx2_ASAP7_75t_L g7212 ( 
.A(n_6669),
.Y(n_7212)
);

INVx2_ASAP7_75t_L g7213 ( 
.A(n_6744),
.Y(n_7213)
);

HB1xp67_ASAP7_75t_L g7214 ( 
.A(n_6765),
.Y(n_7214)
);

NAND2xp5_ASAP7_75t_L g7215 ( 
.A(n_6997),
.B(n_6123),
.Y(n_7215)
);

INVx1_ASAP7_75t_L g7216 ( 
.A(n_6638),
.Y(n_7216)
);

AND2x2_ASAP7_75t_L g7217 ( 
.A(n_6905),
.B(n_6451),
.Y(n_7217)
);

NAND2xp5_ASAP7_75t_L g7218 ( 
.A(n_6588),
.B(n_6404),
.Y(n_7218)
);

AND2x2_ASAP7_75t_L g7219 ( 
.A(n_6921),
.B(n_6791),
.Y(n_7219)
);

AND2x2_ASAP7_75t_L g7220 ( 
.A(n_6921),
.B(n_6338),
.Y(n_7220)
);

INVx1_ASAP7_75t_L g7221 ( 
.A(n_6640),
.Y(n_7221)
);

BUFx3_ASAP7_75t_L g7222 ( 
.A(n_6677),
.Y(n_7222)
);

AND2x2_ASAP7_75t_L g7223 ( 
.A(n_6791),
.B(n_6338),
.Y(n_7223)
);

HB1xp67_ASAP7_75t_L g7224 ( 
.A(n_6827),
.Y(n_7224)
);

INVx2_ASAP7_75t_L g7225 ( 
.A(n_6744),
.Y(n_7225)
);

AND2x2_ASAP7_75t_L g7226 ( 
.A(n_6797),
.B(n_6345),
.Y(n_7226)
);

NAND2xp5_ASAP7_75t_L g7227 ( 
.A(n_6590),
.B(n_6404),
.Y(n_7227)
);

AND2x2_ASAP7_75t_L g7228 ( 
.A(n_6797),
.B(n_6345),
.Y(n_7228)
);

HB1xp67_ASAP7_75t_L g7229 ( 
.A(n_6805),
.Y(n_7229)
);

AND2x2_ASAP7_75t_L g7230 ( 
.A(n_6607),
.B(n_6356),
.Y(n_7230)
);

INVx1_ASAP7_75t_L g7231 ( 
.A(n_6644),
.Y(n_7231)
);

AND2x2_ASAP7_75t_L g7232 ( 
.A(n_6610),
.B(n_6356),
.Y(n_7232)
);

INVx2_ASAP7_75t_L g7233 ( 
.A(n_6755),
.Y(n_7233)
);

INVxp67_ASAP7_75t_L g7234 ( 
.A(n_6685),
.Y(n_7234)
);

INVx2_ASAP7_75t_L g7235 ( 
.A(n_6755),
.Y(n_7235)
);

AND2x2_ASAP7_75t_L g7236 ( 
.A(n_6614),
.B(n_6294),
.Y(n_7236)
);

OR2x2_ASAP7_75t_L g7237 ( 
.A(n_6821),
.B(n_6427),
.Y(n_7237)
);

INVx2_ASAP7_75t_L g7238 ( 
.A(n_6756),
.Y(n_7238)
);

AOI221xp5_ASAP7_75t_L g7239 ( 
.A1(n_6904),
.A2(n_6028),
.B1(n_5771),
.B2(n_5766),
.C(n_5754),
.Y(n_7239)
);

AND2x4_ASAP7_75t_L g7240 ( 
.A(n_6652),
.B(n_6125),
.Y(n_7240)
);

OR2x2_ASAP7_75t_L g7241 ( 
.A(n_6822),
.B(n_6427),
.Y(n_7241)
);

NAND2xp5_ASAP7_75t_L g7242 ( 
.A(n_6594),
.B(n_6532),
.Y(n_7242)
);

INVx2_ASAP7_75t_L g7243 ( 
.A(n_6756),
.Y(n_7243)
);

NAND2xp5_ASAP7_75t_L g7244 ( 
.A(n_6715),
.B(n_6321),
.Y(n_7244)
);

INVx1_ASAP7_75t_L g7245 ( 
.A(n_6645),
.Y(n_7245)
);

INVx1_ASAP7_75t_L g7246 ( 
.A(n_6662),
.Y(n_7246)
);

INVx2_ASAP7_75t_L g7247 ( 
.A(n_6795),
.Y(n_7247)
);

OR2x2_ASAP7_75t_L g7248 ( 
.A(n_6702),
.B(n_6429),
.Y(n_7248)
);

AND2x2_ASAP7_75t_L g7249 ( 
.A(n_6627),
.B(n_6294),
.Y(n_7249)
);

AND2x2_ASAP7_75t_L g7250 ( 
.A(n_6585),
.B(n_6397),
.Y(n_7250)
);

AND2x2_ASAP7_75t_L g7251 ( 
.A(n_6585),
.B(n_6397),
.Y(n_7251)
);

INVx1_ASAP7_75t_L g7252 ( 
.A(n_6665),
.Y(n_7252)
);

NAND2xp5_ASAP7_75t_L g7253 ( 
.A(n_6715),
.B(n_6982),
.Y(n_7253)
);

AND2x2_ASAP7_75t_L g7254 ( 
.A(n_6945),
.B(n_6414),
.Y(n_7254)
);

AND2x2_ASAP7_75t_L g7255 ( 
.A(n_6585),
.B(n_6398),
.Y(n_7255)
);

AND2x2_ASAP7_75t_L g7256 ( 
.A(n_6709),
.B(n_6398),
.Y(n_7256)
);

INVx1_ASAP7_75t_L g7257 ( 
.A(n_6672),
.Y(n_7257)
);

INVx1_ASAP7_75t_L g7258 ( 
.A(n_6674),
.Y(n_7258)
);

INVx3_ASAP7_75t_L g7259 ( 
.A(n_6767),
.Y(n_7259)
);

INVx2_ASAP7_75t_L g7260 ( 
.A(n_6795),
.Y(n_7260)
);

INVx1_ASAP7_75t_L g7261 ( 
.A(n_6676),
.Y(n_7261)
);

HB1xp67_ASAP7_75t_L g7262 ( 
.A(n_7006),
.Y(n_7262)
);

INVx1_ASAP7_75t_SL g7263 ( 
.A(n_6677),
.Y(n_7263)
);

AND2x2_ASAP7_75t_L g7264 ( 
.A(n_6878),
.B(n_6263),
.Y(n_7264)
);

AND2x2_ASAP7_75t_L g7265 ( 
.A(n_6886),
.B(n_6263),
.Y(n_7265)
);

NAND2x1p5_ASAP7_75t_L g7266 ( 
.A(n_6779),
.B(n_5044),
.Y(n_7266)
);

OR2x2_ASAP7_75t_L g7267 ( 
.A(n_6562),
.B(n_6429),
.Y(n_7267)
);

BUFx2_ASAP7_75t_L g7268 ( 
.A(n_6748),
.Y(n_7268)
);

AND2x2_ASAP7_75t_L g7269 ( 
.A(n_6889),
.B(n_6414),
.Y(n_7269)
);

INVx1_ASAP7_75t_L g7270 ( 
.A(n_6680),
.Y(n_7270)
);

AND2x2_ASAP7_75t_L g7271 ( 
.A(n_6890),
.B(n_6893),
.Y(n_7271)
);

INVx3_ASAP7_75t_L g7272 ( 
.A(n_6599),
.Y(n_7272)
);

AND2x2_ASAP7_75t_L g7273 ( 
.A(n_6664),
.B(n_6373),
.Y(n_7273)
);

NAND2xp5_ASAP7_75t_L g7274 ( 
.A(n_6982),
.B(n_6321),
.Y(n_7274)
);

AND2x2_ASAP7_75t_L g7275 ( 
.A(n_6666),
.B(n_6373),
.Y(n_7275)
);

AOI22xp33_ASAP7_75t_L g7276 ( 
.A1(n_6888),
.A2(n_6191),
.B1(n_6194),
.B2(n_6190),
.Y(n_7276)
);

INVx1_ASAP7_75t_L g7277 ( 
.A(n_6683),
.Y(n_7277)
);

NOR3xp33_ASAP7_75t_L g7278 ( 
.A(n_6563),
.B(n_6083),
.C(n_6046),
.Y(n_7278)
);

INVx2_ASAP7_75t_L g7279 ( 
.A(n_6796),
.Y(n_7279)
);

INVx2_ASAP7_75t_L g7280 ( 
.A(n_6796),
.Y(n_7280)
);

INVx1_ASAP7_75t_L g7281 ( 
.A(n_6684),
.Y(n_7281)
);

AND2x2_ASAP7_75t_L g7282 ( 
.A(n_6724),
.B(n_6065),
.Y(n_7282)
);

BUFx2_ASAP7_75t_L g7283 ( 
.A(n_6748),
.Y(n_7283)
);

INVx2_ASAP7_75t_L g7284 ( 
.A(n_6798),
.Y(n_7284)
);

BUFx2_ASAP7_75t_L g7285 ( 
.A(n_6926),
.Y(n_7285)
);

INVx1_ASAP7_75t_L g7286 ( 
.A(n_6686),
.Y(n_7286)
);

INVx2_ASAP7_75t_SL g7287 ( 
.A(n_6606),
.Y(n_7287)
);

AND2x2_ASAP7_75t_L g7288 ( 
.A(n_6926),
.B(n_6065),
.Y(n_7288)
);

OR2x2_ASAP7_75t_L g7289 ( 
.A(n_6564),
.B(n_6328),
.Y(n_7289)
);

INVx2_ASAP7_75t_L g7290 ( 
.A(n_6798),
.Y(n_7290)
);

INVx1_ASAP7_75t_L g7291 ( 
.A(n_6694),
.Y(n_7291)
);

INVx2_ASAP7_75t_L g7292 ( 
.A(n_6804),
.Y(n_7292)
);

INVx2_ASAP7_75t_L g7293 ( 
.A(n_6804),
.Y(n_7293)
);

AND2x2_ASAP7_75t_L g7294 ( 
.A(n_6940),
.B(n_6065),
.Y(n_7294)
);

BUFx2_ASAP7_75t_L g7295 ( 
.A(n_6940),
.Y(n_7295)
);

NAND2xp5_ASAP7_75t_L g7296 ( 
.A(n_7010),
.B(n_6328),
.Y(n_7296)
);

INVx1_ASAP7_75t_L g7297 ( 
.A(n_6695),
.Y(n_7297)
);

INVxp67_ASAP7_75t_SL g7298 ( 
.A(n_6917),
.Y(n_7298)
);

OR2x2_ASAP7_75t_L g7299 ( 
.A(n_6577),
.B(n_6117),
.Y(n_7299)
);

INVx2_ASAP7_75t_SL g7300 ( 
.A(n_6606),
.Y(n_7300)
);

AND2x2_ASAP7_75t_L g7301 ( 
.A(n_6934),
.B(n_6716),
.Y(n_7301)
);

INVx2_ASAP7_75t_L g7302 ( 
.A(n_6812),
.Y(n_7302)
);

INVx1_ASAP7_75t_L g7303 ( 
.A(n_6700),
.Y(n_7303)
);

AND2x2_ASAP7_75t_L g7304 ( 
.A(n_6720),
.B(n_6151),
.Y(n_7304)
);

INVx2_ASAP7_75t_L g7305 ( 
.A(n_6812),
.Y(n_7305)
);

AND2x2_ASAP7_75t_L g7306 ( 
.A(n_6948),
.B(n_6151),
.Y(n_7306)
);

INVx1_ASAP7_75t_L g7307 ( 
.A(n_6701),
.Y(n_7307)
);

INVx2_ASAP7_75t_L g7308 ( 
.A(n_6815),
.Y(n_7308)
);

AND2x4_ASAP7_75t_L g7309 ( 
.A(n_6652),
.B(n_6125),
.Y(n_7309)
);

INVx2_ASAP7_75t_L g7310 ( 
.A(n_6815),
.Y(n_7310)
);

INVx3_ASAP7_75t_L g7311 ( 
.A(n_6599),
.Y(n_7311)
);

AND2x2_ASAP7_75t_L g7312 ( 
.A(n_6954),
.B(n_6151),
.Y(n_7312)
);

NAND2xp5_ASAP7_75t_L g7313 ( 
.A(n_6929),
.B(n_6119),
.Y(n_7313)
);

OR2x2_ASAP7_75t_L g7314 ( 
.A(n_6579),
.B(n_6126),
.Y(n_7314)
);

INVx1_ASAP7_75t_L g7315 ( 
.A(n_6712),
.Y(n_7315)
);

INVx3_ASAP7_75t_L g7316 ( 
.A(n_6917),
.Y(n_7316)
);

INVx2_ASAP7_75t_SL g7317 ( 
.A(n_6739),
.Y(n_7317)
);

INVx3_ASAP7_75t_SL g7318 ( 
.A(n_6794),
.Y(n_7318)
);

AOI22xp33_ASAP7_75t_L g7319 ( 
.A1(n_6888),
.A2(n_6854),
.B1(n_6792),
.B2(n_6587),
.Y(n_7319)
);

INVxp67_ASAP7_75t_SL g7320 ( 
.A(n_6917),
.Y(n_7320)
);

INVx1_ASAP7_75t_L g7321 ( 
.A(n_6723),
.Y(n_7321)
);

INVx2_ASAP7_75t_L g7322 ( 
.A(n_6671),
.Y(n_7322)
);

AND2x2_ASAP7_75t_L g7323 ( 
.A(n_6831),
.B(n_6162),
.Y(n_7323)
);

NAND2xp5_ASAP7_75t_L g7324 ( 
.A(n_6937),
.B(n_6130),
.Y(n_7324)
);

AND2x2_ASAP7_75t_L g7325 ( 
.A(n_6652),
.B(n_6162),
.Y(n_7325)
);

AND2x2_ASAP7_75t_L g7326 ( 
.A(n_6681),
.B(n_6162),
.Y(n_7326)
);

AND2x2_ASAP7_75t_L g7327 ( 
.A(n_6681),
.B(n_6164),
.Y(n_7327)
);

HB1xp67_ASAP7_75t_L g7328 ( 
.A(n_7006),
.Y(n_7328)
);

AND2x2_ASAP7_75t_L g7329 ( 
.A(n_6681),
.B(n_6164),
.Y(n_7329)
);

AND2x2_ASAP7_75t_L g7330 ( 
.A(n_6687),
.B(n_6164),
.Y(n_7330)
);

INVxp67_ASAP7_75t_SL g7331 ( 
.A(n_6787),
.Y(n_7331)
);

NAND2xp5_ASAP7_75t_L g7332 ( 
.A(n_6959),
.B(n_6133),
.Y(n_7332)
);

INVx1_ASAP7_75t_L g7333 ( 
.A(n_6732),
.Y(n_7333)
);

BUFx6f_ASAP7_75t_L g7334 ( 
.A(n_6625),
.Y(n_7334)
);

AND2x2_ASAP7_75t_L g7335 ( 
.A(n_6687),
.B(n_6219),
.Y(n_7335)
);

AND2x2_ASAP7_75t_L g7336 ( 
.A(n_6687),
.B(n_6219),
.Y(n_7336)
);

INVx2_ASAP7_75t_L g7337 ( 
.A(n_6671),
.Y(n_7337)
);

AND2x2_ASAP7_75t_L g7338 ( 
.A(n_6699),
.B(n_6219),
.Y(n_7338)
);

INVx1_ASAP7_75t_L g7339 ( 
.A(n_6742),
.Y(n_7339)
);

NAND2xp5_ASAP7_75t_L g7340 ( 
.A(n_6963),
.B(n_6138),
.Y(n_7340)
);

AND2x2_ASAP7_75t_L g7341 ( 
.A(n_6837),
.B(n_6264),
.Y(n_7341)
);

INVx2_ASAP7_75t_L g7342 ( 
.A(n_6673),
.Y(n_7342)
);

AND2x2_ASAP7_75t_L g7343 ( 
.A(n_6846),
.B(n_6264),
.Y(n_7343)
);

INVx2_ASAP7_75t_L g7344 ( 
.A(n_6673),
.Y(n_7344)
);

INVx1_ASAP7_75t_L g7345 ( 
.A(n_6745),
.Y(n_7345)
);

INVx2_ASAP7_75t_L g7346 ( 
.A(n_6678),
.Y(n_7346)
);

OR2x2_ASAP7_75t_L g7347 ( 
.A(n_6583),
.B(n_6589),
.Y(n_7347)
);

OR2x2_ASAP7_75t_L g7348 ( 
.A(n_6593),
.B(n_6140),
.Y(n_7348)
);

AND2x2_ASAP7_75t_L g7349 ( 
.A(n_6883),
.B(n_6885),
.Y(n_7349)
);

INVx2_ASAP7_75t_L g7350 ( 
.A(n_6678),
.Y(n_7350)
);

NAND2xp5_ASAP7_75t_L g7351 ( 
.A(n_6596),
.B(n_6156),
.Y(n_7351)
);

AND2x4_ASAP7_75t_L g7352 ( 
.A(n_6699),
.B(n_6125),
.Y(n_7352)
);

INVxp67_ASAP7_75t_SL g7353 ( 
.A(n_6787),
.Y(n_7353)
);

AND2x4_ASAP7_75t_L g7354 ( 
.A(n_6699),
.B(n_6895),
.Y(n_7354)
);

INVx2_ASAP7_75t_L g7355 ( 
.A(n_6786),
.Y(n_7355)
);

NOR2xp67_ASAP7_75t_L g7356 ( 
.A(n_6834),
.B(n_6264),
.Y(n_7356)
);

INVx5_ASAP7_75t_L g7357 ( 
.A(n_6809),
.Y(n_7357)
);

INVx1_ASAP7_75t_L g7358 ( 
.A(n_6749),
.Y(n_7358)
);

OR2x2_ASAP7_75t_L g7359 ( 
.A(n_6902),
.B(n_6157),
.Y(n_7359)
);

AND2x2_ASAP7_75t_L g7360 ( 
.A(n_6743),
.B(n_6782),
.Y(n_7360)
);

BUFx6f_ASAP7_75t_L g7361 ( 
.A(n_6625),
.Y(n_7361)
);

OR2x2_ASAP7_75t_L g7362 ( 
.A(n_6993),
.B(n_6158),
.Y(n_7362)
);

AND2x2_ASAP7_75t_L g7363 ( 
.A(n_6800),
.B(n_6054),
.Y(n_7363)
);

AND2x2_ASAP7_75t_L g7364 ( 
.A(n_6808),
.B(n_6054),
.Y(n_7364)
);

NAND2xp5_ASAP7_75t_L g7365 ( 
.A(n_6895),
.B(n_6166),
.Y(n_7365)
);

AND2x2_ASAP7_75t_L g7366 ( 
.A(n_6955),
.B(n_6063),
.Y(n_7366)
);

INVx1_ASAP7_75t_L g7367 ( 
.A(n_6760),
.Y(n_7367)
);

AND2x2_ASAP7_75t_L g7368 ( 
.A(n_6965),
.B(n_6063),
.Y(n_7368)
);

AND2x2_ASAP7_75t_L g7369 ( 
.A(n_6969),
.B(n_6071),
.Y(n_7369)
);

NAND2xp5_ASAP7_75t_L g7370 ( 
.A(n_6630),
.B(n_6169),
.Y(n_7370)
);

INVx4_ASAP7_75t_L g7371 ( 
.A(n_6773),
.Y(n_7371)
);

AND2x2_ASAP7_75t_L g7372 ( 
.A(n_6974),
.B(n_6071),
.Y(n_7372)
);

CKINVDCx6p67_ASAP7_75t_R g7373 ( 
.A(n_6872),
.Y(n_7373)
);

INVx1_ASAP7_75t_L g7374 ( 
.A(n_6766),
.Y(n_7374)
);

INVx2_ASAP7_75t_L g7375 ( 
.A(n_6786),
.Y(n_7375)
);

INVx2_ASAP7_75t_L g7376 ( 
.A(n_6786),
.Y(n_7376)
);

INVx1_ASAP7_75t_L g7377 ( 
.A(n_6768),
.Y(n_7377)
);

NOR2xp33_ASAP7_75t_L g7378 ( 
.A(n_6809),
.B(n_5994),
.Y(n_7378)
);

NAND2xp5_ASAP7_75t_L g7379 ( 
.A(n_6616),
.B(n_6170),
.Y(n_7379)
);

INVx2_ASAP7_75t_L g7380 ( 
.A(n_6786),
.Y(n_7380)
);

AND2x4_ASAP7_75t_L g7381 ( 
.A(n_6557),
.B(n_6125),
.Y(n_7381)
);

AND2x2_ASAP7_75t_L g7382 ( 
.A(n_6976),
.B(n_6073),
.Y(n_7382)
);

NOR2xp33_ASAP7_75t_L g7383 ( 
.A(n_6773),
.B(n_4864),
.Y(n_7383)
);

INVx1_ASAP7_75t_L g7384 ( 
.A(n_6790),
.Y(n_7384)
);

INVx1_ASAP7_75t_L g7385 ( 
.A(n_6799),
.Y(n_7385)
);

INVx2_ASAP7_75t_L g7386 ( 
.A(n_6958),
.Y(n_7386)
);

HB1xp67_ASAP7_75t_L g7387 ( 
.A(n_6624),
.Y(n_7387)
);

AND2x2_ASAP7_75t_L g7388 ( 
.A(n_6981),
.B(n_6073),
.Y(n_7388)
);

INVx1_ASAP7_75t_L g7389 ( 
.A(n_6802),
.Y(n_7389)
);

INVx2_ASAP7_75t_L g7390 ( 
.A(n_6958),
.Y(n_7390)
);

AND2x2_ASAP7_75t_L g7391 ( 
.A(n_6692),
.B(n_6079),
.Y(n_7391)
);

AND2x2_ASAP7_75t_L g7392 ( 
.A(n_6693),
.B(n_6079),
.Y(n_7392)
);

INVx1_ASAP7_75t_L g7393 ( 
.A(n_6803),
.Y(n_7393)
);

AND2x2_ASAP7_75t_L g7394 ( 
.A(n_6708),
.B(n_6089),
.Y(n_7394)
);

AND2x2_ASAP7_75t_L g7395 ( 
.A(n_6870),
.B(n_6089),
.Y(n_7395)
);

INVx1_ASAP7_75t_L g7396 ( 
.A(n_6806),
.Y(n_7396)
);

HB1xp67_ASAP7_75t_L g7397 ( 
.A(n_6631),
.Y(n_7397)
);

AND2x2_ASAP7_75t_L g7398 ( 
.A(n_6953),
.B(n_6104),
.Y(n_7398)
);

INVx2_ASAP7_75t_L g7399 ( 
.A(n_6958),
.Y(n_7399)
);

INVxp67_ASAP7_75t_SL g7400 ( 
.A(n_6851),
.Y(n_7400)
);

INVx1_ASAP7_75t_L g7401 ( 
.A(n_6816),
.Y(n_7401)
);

NAND2xp5_ASAP7_75t_L g7402 ( 
.A(n_6620),
.B(n_6175),
.Y(n_7402)
);

OR2x2_ASAP7_75t_L g7403 ( 
.A(n_6864),
.B(n_6182),
.Y(n_7403)
);

AND2x2_ASAP7_75t_L g7404 ( 
.A(n_6953),
.B(n_6104),
.Y(n_7404)
);

AND2x2_ASAP7_75t_L g7405 ( 
.A(n_6818),
.B(n_6747),
.Y(n_7405)
);

AND2x2_ASAP7_75t_L g7406 ( 
.A(n_6818),
.B(n_6108),
.Y(n_7406)
);

AND2x2_ASAP7_75t_L g7407 ( 
.A(n_6769),
.B(n_6108),
.Y(n_7407)
);

OR2x2_ASAP7_75t_L g7408 ( 
.A(n_6868),
.B(n_6998),
.Y(n_7408)
);

INVx1_ASAP7_75t_L g7409 ( 
.A(n_6817),
.Y(n_7409)
);

INVx2_ASAP7_75t_L g7410 ( 
.A(n_6958),
.Y(n_7410)
);

INVx1_ASAP7_75t_L g7411 ( 
.A(n_6823),
.Y(n_7411)
);

AND2x2_ASAP7_75t_L g7412 ( 
.A(n_6770),
.B(n_6118),
.Y(n_7412)
);

INVx2_ASAP7_75t_SL g7413 ( 
.A(n_6739),
.Y(n_7413)
);

OR2x2_ASAP7_75t_L g7414 ( 
.A(n_6880),
.B(n_6239),
.Y(n_7414)
);

INVx2_ASAP7_75t_L g7415 ( 
.A(n_6941),
.Y(n_7415)
);

INVx3_ASAP7_75t_L g7416 ( 
.A(n_6933),
.Y(n_7416)
);

AND2x2_ASAP7_75t_L g7417 ( 
.A(n_6779),
.B(n_6340),
.Y(n_7417)
);

INVx2_ASAP7_75t_L g7418 ( 
.A(n_6941),
.Y(n_7418)
);

INVx2_ASAP7_75t_L g7419 ( 
.A(n_6961),
.Y(n_7419)
);

AND2x2_ASAP7_75t_L g7420 ( 
.A(n_6779),
.B(n_6784),
.Y(n_7420)
);

INVx1_ASAP7_75t_L g7421 ( 
.A(n_6825),
.Y(n_7421)
);

OR2x2_ASAP7_75t_L g7422 ( 
.A(n_6923),
.B(n_6249),
.Y(n_7422)
);

INVx2_ASAP7_75t_L g7423 ( 
.A(n_6961),
.Y(n_7423)
);

NAND2x1p5_ASAP7_75t_L g7424 ( 
.A(n_6784),
.B(n_6810),
.Y(n_7424)
);

AND2x2_ASAP7_75t_L g7425 ( 
.A(n_6784),
.B(n_6340),
.Y(n_7425)
);

INVx1_ASAP7_75t_L g7426 ( 
.A(n_6829),
.Y(n_7426)
);

NAND2xp5_ASAP7_75t_L g7427 ( 
.A(n_6634),
.B(n_6252),
.Y(n_7427)
);

INVx2_ASAP7_75t_L g7428 ( 
.A(n_6973),
.Y(n_7428)
);

AND2x2_ASAP7_75t_L g7429 ( 
.A(n_6810),
.B(n_6340),
.Y(n_7429)
);

INVx1_ASAP7_75t_L g7430 ( 
.A(n_6832),
.Y(n_7430)
);

INVx1_ASAP7_75t_L g7431 ( 
.A(n_6833),
.Y(n_7431)
);

INVxp67_ASAP7_75t_L g7432 ( 
.A(n_6872),
.Y(n_7432)
);

INVx1_ASAP7_75t_L g7433 ( 
.A(n_6835),
.Y(n_7433)
);

INVx1_ASAP7_75t_L g7434 ( 
.A(n_6836),
.Y(n_7434)
);

NAND2xp5_ASAP7_75t_L g7435 ( 
.A(n_6648),
.B(n_6262),
.Y(n_7435)
);

INVx3_ASAP7_75t_L g7436 ( 
.A(n_6933),
.Y(n_7436)
);

HB1xp67_ASAP7_75t_L g7437 ( 
.A(n_6650),
.Y(n_7437)
);

INVx3_ASAP7_75t_L g7438 ( 
.A(n_7007),
.Y(n_7438)
);

BUFx3_ASAP7_75t_L g7439 ( 
.A(n_6773),
.Y(n_7439)
);

BUFx3_ASAP7_75t_L g7440 ( 
.A(n_6773),
.Y(n_7440)
);

NOR2xp33_ASAP7_75t_L g7441 ( 
.A(n_6780),
.B(n_6807),
.Y(n_7441)
);

INVx1_ASAP7_75t_L g7442 ( 
.A(n_6844),
.Y(n_7442)
);

INVx3_ASAP7_75t_L g7443 ( 
.A(n_7007),
.Y(n_7443)
);

INVx2_ASAP7_75t_L g7444 ( 
.A(n_6973),
.Y(n_7444)
);

INVx2_ASAP7_75t_L g7445 ( 
.A(n_6898),
.Y(n_7445)
);

INVx1_ASAP7_75t_L g7446 ( 
.A(n_6845),
.Y(n_7446)
);

BUFx3_ASAP7_75t_L g7447 ( 
.A(n_6780),
.Y(n_7447)
);

NAND4xp25_ASAP7_75t_L g7448 ( 
.A(n_7011),
.B(n_6740),
.C(n_6754),
.D(n_6977),
.Y(n_7448)
);

INVxp67_ASAP7_75t_SL g7449 ( 
.A(n_7084),
.Y(n_7449)
);

BUFx6f_ASAP7_75t_L g7450 ( 
.A(n_7061),
.Y(n_7450)
);

INVx2_ASAP7_75t_L g7451 ( 
.A(n_7084),
.Y(n_7451)
);

INVx2_ASAP7_75t_SL g7452 ( 
.A(n_7168),
.Y(n_7452)
);

INVx1_ASAP7_75t_L g7453 ( 
.A(n_7018),
.Y(n_7453)
);

INVx4_ASAP7_75t_SL g7454 ( 
.A(n_7318),
.Y(n_7454)
);

INVx1_ASAP7_75t_L g7455 ( 
.A(n_7018),
.Y(n_7455)
);

OA21x2_ASAP7_75t_L g7456 ( 
.A1(n_7011),
.A2(n_6992),
.B(n_6851),
.Y(n_7456)
);

OAI21x1_ASAP7_75t_L g7457 ( 
.A1(n_7105),
.A2(n_6840),
.B(n_6834),
.Y(n_7457)
);

INVx1_ASAP7_75t_L g7458 ( 
.A(n_7331),
.Y(n_7458)
);

NAND2xp5_ASAP7_75t_L g7459 ( 
.A(n_7069),
.B(n_6780),
.Y(n_7459)
);

AND2x4_ASAP7_75t_L g7460 ( 
.A(n_7013),
.B(n_6807),
.Y(n_7460)
);

INVx1_ASAP7_75t_SL g7461 ( 
.A(n_7053),
.Y(n_7461)
);

BUFx6f_ASAP7_75t_L g7462 ( 
.A(n_7061),
.Y(n_7462)
);

HB1xp67_ASAP7_75t_L g7463 ( 
.A(n_7042),
.Y(n_7463)
);

AO21x2_ASAP7_75t_L g7464 ( 
.A1(n_7331),
.A2(n_6602),
.B(n_6992),
.Y(n_7464)
);

INVx1_ASAP7_75t_L g7465 ( 
.A(n_7353),
.Y(n_7465)
);

INVxp67_ASAP7_75t_L g7466 ( 
.A(n_7178),
.Y(n_7466)
);

NAND2xp5_ASAP7_75t_L g7467 ( 
.A(n_7077),
.B(n_7048),
.Y(n_7467)
);

AO21x2_ASAP7_75t_L g7468 ( 
.A1(n_7353),
.A2(n_6602),
.B(n_6682),
.Y(n_7468)
);

AND2x6_ASAP7_75t_L g7469 ( 
.A(n_7061),
.B(n_6780),
.Y(n_7469)
);

OR2x2_ASAP7_75t_L g7470 ( 
.A(n_7046),
.B(n_6936),
.Y(n_7470)
);

NOR2xp33_ASAP7_75t_L g7471 ( 
.A(n_7168),
.B(n_6740),
.Y(n_7471)
);

INVx2_ASAP7_75t_SL g7472 ( 
.A(n_7168),
.Y(n_7472)
);

INVx4_ASAP7_75t_L g7473 ( 
.A(n_7168),
.Y(n_7473)
);

HB1xp67_ASAP7_75t_L g7474 ( 
.A(n_7042),
.Y(n_7474)
);

AND2x2_ASAP7_75t_L g7475 ( 
.A(n_7146),
.B(n_6810),
.Y(n_7475)
);

INVx2_ASAP7_75t_L g7476 ( 
.A(n_7285),
.Y(n_7476)
);

INVx2_ASAP7_75t_L g7477 ( 
.A(n_7295),
.Y(n_7477)
);

INVx1_ASAP7_75t_L g7478 ( 
.A(n_7400),
.Y(n_7478)
);

AND2x2_ASAP7_75t_L g7479 ( 
.A(n_7015),
.B(n_6750),
.Y(n_7479)
);

INVx3_ASAP7_75t_L g7480 ( 
.A(n_7171),
.Y(n_7480)
);

NAND2xp5_ASAP7_75t_L g7481 ( 
.A(n_7229),
.B(n_7013),
.Y(n_7481)
);

INVx2_ASAP7_75t_SL g7482 ( 
.A(n_7357),
.Y(n_7482)
);

OAI21xp33_ASAP7_75t_SL g7483 ( 
.A1(n_7319),
.A2(n_6907),
.B(n_6840),
.Y(n_7483)
);

OAI21x1_ASAP7_75t_L g7484 ( 
.A1(n_7105),
.A2(n_6557),
.B(n_6642),
.Y(n_7484)
);

BUFx3_ASAP7_75t_L g7485 ( 
.A(n_7357),
.Y(n_7485)
);

NAND2xp5_ASAP7_75t_L g7486 ( 
.A(n_7229),
.B(n_7220),
.Y(n_7486)
);

INVx5_ASAP7_75t_L g7487 ( 
.A(n_7061),
.Y(n_7487)
);

AND2x2_ASAP7_75t_L g7488 ( 
.A(n_7016),
.B(n_6753),
.Y(n_7488)
);

A2O1A1Ixp33_ASAP7_75t_L g7489 ( 
.A1(n_7319),
.A2(n_6752),
.B(n_6792),
.C(n_6757),
.Y(n_7489)
);

BUFx2_ASAP7_75t_L g7490 ( 
.A(n_7095),
.Y(n_7490)
);

BUFx3_ASAP7_75t_L g7491 ( 
.A(n_7357),
.Y(n_7491)
);

AND2x2_ASAP7_75t_L g7492 ( 
.A(n_7360),
.B(n_6758),
.Y(n_7492)
);

AND2x2_ASAP7_75t_L g7493 ( 
.A(n_7124),
.B(n_6759),
.Y(n_7493)
);

OAI21x1_ASAP7_75t_L g7494 ( 
.A1(n_7105),
.A2(n_7311),
.B(n_7272),
.Y(n_7494)
);

INVx1_ASAP7_75t_L g7495 ( 
.A(n_7051),
.Y(n_7495)
);

INVx4_ASAP7_75t_SL g7496 ( 
.A(n_7318),
.Y(n_7496)
);

AND2x4_ASAP7_75t_L g7497 ( 
.A(n_7095),
.B(n_7004),
.Y(n_7497)
);

INVx1_ASAP7_75t_L g7498 ( 
.A(n_7051),
.Y(n_7498)
);

BUFx2_ASAP7_75t_L g7499 ( 
.A(n_7099),
.Y(n_7499)
);

AND2x2_ASAP7_75t_L g7500 ( 
.A(n_7133),
.B(n_6761),
.Y(n_7500)
);

INVx2_ASAP7_75t_L g7501 ( 
.A(n_7171),
.Y(n_7501)
);

INVx2_ASAP7_75t_SL g7502 ( 
.A(n_7357),
.Y(n_7502)
);

INVx1_ASAP7_75t_L g7503 ( 
.A(n_7073),
.Y(n_7503)
);

INVx1_ASAP7_75t_L g7504 ( 
.A(n_7073),
.Y(n_7504)
);

OAI21xp5_ASAP7_75t_L g7505 ( 
.A1(n_7036),
.A2(n_6884),
.B(n_6682),
.Y(n_7505)
);

INVx3_ASAP7_75t_L g7506 ( 
.A(n_7171),
.Y(n_7506)
);

HB1xp67_ASAP7_75t_L g7507 ( 
.A(n_7107),
.Y(n_7507)
);

INVx4_ASAP7_75t_L g7508 ( 
.A(n_7087),
.Y(n_7508)
);

BUFx3_ASAP7_75t_L g7509 ( 
.A(n_7099),
.Y(n_7509)
);

OAI211xp5_ASAP7_75t_L g7510 ( 
.A1(n_7036),
.A2(n_6622),
.B(n_6741),
.C(n_7009),
.Y(n_7510)
);

NAND4xp25_ASAP7_75t_L g7511 ( 
.A(n_7054),
.B(n_6728),
.C(n_6731),
.D(n_6557),
.Y(n_7511)
);

INVx1_ASAP7_75t_L g7512 ( 
.A(n_7075),
.Y(n_7512)
);

INVx2_ASAP7_75t_L g7513 ( 
.A(n_7171),
.Y(n_7513)
);

OR2x6_ASAP7_75t_L g7514 ( 
.A(n_7064),
.B(n_6197),
.Y(n_7514)
);

INVx1_ASAP7_75t_L g7515 ( 
.A(n_7075),
.Y(n_7515)
);

INVx2_ASAP7_75t_L g7516 ( 
.A(n_7195),
.Y(n_7516)
);

NAND2xp5_ASAP7_75t_L g7517 ( 
.A(n_7017),
.B(n_6950),
.Y(n_7517)
);

INVx1_ASAP7_75t_L g7518 ( 
.A(n_7091),
.Y(n_7518)
);

AOI21xp33_ASAP7_75t_L g7519 ( 
.A1(n_7164),
.A2(n_6661),
.B(n_6604),
.Y(n_7519)
);

HB1xp67_ASAP7_75t_L g7520 ( 
.A(n_7212),
.Y(n_7520)
);

BUFx3_ASAP7_75t_L g7521 ( 
.A(n_7145),
.Y(n_7521)
);

AND2x2_ASAP7_75t_L g7522 ( 
.A(n_7398),
.B(n_6713),
.Y(n_7522)
);

BUFx3_ASAP7_75t_L g7523 ( 
.A(n_7145),
.Y(n_7523)
);

NOR4xp75_ASAP7_75t_L g7524 ( 
.A(n_7043),
.B(n_6696),
.C(n_6659),
.D(n_6647),
.Y(n_7524)
);

INVx2_ASAP7_75t_L g7525 ( 
.A(n_7195),
.Y(n_7525)
);

OR2x2_ASAP7_75t_L g7526 ( 
.A(n_7050),
.B(n_6952),
.Y(n_7526)
);

INVx2_ASAP7_75t_L g7527 ( 
.A(n_7195),
.Y(n_7527)
);

OAI21xp33_ASAP7_75t_L g7528 ( 
.A1(n_7276),
.A2(n_6849),
.B(n_6983),
.Y(n_7528)
);

NAND4xp25_ASAP7_75t_L g7529 ( 
.A(n_7130),
.B(n_6713),
.C(n_6978),
.D(n_6647),
.Y(n_7529)
);

NAND2xp5_ASAP7_75t_L g7530 ( 
.A(n_7017),
.B(n_6956),
.Y(n_7530)
);

BUFx8_ASAP7_75t_L g7531 ( 
.A(n_7087),
.Y(n_7531)
);

INVxp67_ASAP7_75t_SL g7532 ( 
.A(n_7383),
.Y(n_7532)
);

INVx4_ASAP7_75t_SL g7533 ( 
.A(n_7195),
.Y(n_7533)
);

AND2x4_ASAP7_75t_L g7534 ( 
.A(n_7222),
.B(n_6642),
.Y(n_7534)
);

BUFx8_ASAP7_75t_L g7535 ( 
.A(n_7020),
.Y(n_7535)
);

NAND2xp5_ASAP7_75t_L g7536 ( 
.A(n_7268),
.B(n_6894),
.Y(n_7536)
);

BUFx3_ASAP7_75t_L g7537 ( 
.A(n_7222),
.Y(n_7537)
);

NAND2xp5_ASAP7_75t_L g7538 ( 
.A(n_7283),
.B(n_6901),
.Y(n_7538)
);

INVx1_ASAP7_75t_L g7539 ( 
.A(n_7400),
.Y(n_7539)
);

OAI21xp5_ASAP7_75t_L g7540 ( 
.A1(n_7276),
.A2(n_6587),
.B(n_6719),
.Y(n_7540)
);

NAND2xp5_ASAP7_75t_L g7541 ( 
.A(n_7219),
.B(n_6906),
.Y(n_7541)
);

INVx1_ASAP7_75t_L g7542 ( 
.A(n_7091),
.Y(n_7542)
);

OAI21xp5_ASAP7_75t_L g7543 ( 
.A1(n_7037),
.A2(n_6736),
.B(n_6719),
.Y(n_7543)
);

NAND2x1p5_ASAP7_75t_SL g7544 ( 
.A(n_7043),
.B(n_6558),
.Y(n_7544)
);

AND2x2_ASAP7_75t_L g7545 ( 
.A(n_7404),
.B(n_6713),
.Y(n_7545)
);

A2O1A1Ixp33_ASAP7_75t_L g7546 ( 
.A1(n_7037),
.A2(n_6736),
.B(n_6908),
.C(n_6990),
.Y(n_7546)
);

INVx1_ASAP7_75t_L g7547 ( 
.A(n_7111),
.Y(n_7547)
);

AND2x4_ASAP7_75t_SL g7548 ( 
.A(n_7058),
.B(n_5150),
.Y(n_7548)
);

HB1xp67_ASAP7_75t_L g7549 ( 
.A(n_7432),
.Y(n_7549)
);

INVx1_ASAP7_75t_L g7550 ( 
.A(n_7111),
.Y(n_7550)
);

INVx2_ASAP7_75t_L g7551 ( 
.A(n_7334),
.Y(n_7551)
);

INVx1_ASAP7_75t_L g7552 ( 
.A(n_7112),
.Y(n_7552)
);

BUFx3_ASAP7_75t_L g7553 ( 
.A(n_7373),
.Y(n_7553)
);

INVx1_ASAP7_75t_L g7554 ( 
.A(n_7112),
.Y(n_7554)
);

NOR2xp33_ASAP7_75t_L g7555 ( 
.A(n_7373),
.B(n_6651),
.Y(n_7555)
);

NAND2xp5_ASAP7_75t_L g7556 ( 
.A(n_7197),
.B(n_6910),
.Y(n_7556)
);

NAND2xp5_ASAP7_75t_L g7557 ( 
.A(n_7263),
.B(n_6922),
.Y(n_7557)
);

NAND2xp33_ASAP7_75t_L g7558 ( 
.A(n_7334),
.B(n_6655),
.Y(n_7558)
);

INVxp67_ASAP7_75t_SL g7559 ( 
.A(n_7383),
.Y(n_7559)
);

NAND2xp5_ASAP7_75t_L g7560 ( 
.A(n_7387),
.B(n_6925),
.Y(n_7560)
);

OA21x2_ASAP7_75t_L g7561 ( 
.A1(n_7298),
.A2(n_6899),
.B(n_6898),
.Y(n_7561)
);

O2A1O1Ixp33_ASAP7_75t_L g7562 ( 
.A1(n_7206),
.A2(n_6661),
.B(n_6714),
.C(n_6604),
.Y(n_7562)
);

INVx5_ASAP7_75t_L g7563 ( 
.A(n_7334),
.Y(n_7563)
);

HB1xp67_ASAP7_75t_L g7564 ( 
.A(n_7100),
.Y(n_7564)
);

OA21x2_ASAP7_75t_L g7565 ( 
.A1(n_7298),
.A2(n_6900),
.B(n_6899),
.Y(n_7565)
);

AND2x4_ASAP7_75t_L g7566 ( 
.A(n_7354),
.B(n_6651),
.Y(n_7566)
);

OAI21x1_ASAP7_75t_L g7567 ( 
.A1(n_7272),
.A2(n_6751),
.B(n_6729),
.Y(n_7567)
);

INVx1_ASAP7_75t_L g7568 ( 
.A(n_7115),
.Y(n_7568)
);

INVx2_ASAP7_75t_L g7569 ( 
.A(n_7334),
.Y(n_7569)
);

BUFx2_ASAP7_75t_L g7570 ( 
.A(n_7354),
.Y(n_7570)
);

OR2x2_ASAP7_75t_L g7571 ( 
.A(n_7114),
.B(n_6877),
.Y(n_7571)
);

BUFx6f_ASAP7_75t_L g7572 ( 
.A(n_7361),
.Y(n_7572)
);

NAND2x1p5_ASAP7_75t_SL g7573 ( 
.A(n_7020),
.B(n_6558),
.Y(n_7573)
);

INVx2_ASAP7_75t_SL g7574 ( 
.A(n_7090),
.Y(n_7574)
);

BUFx2_ASAP7_75t_L g7575 ( 
.A(n_7354),
.Y(n_7575)
);

NAND2xp33_ASAP7_75t_SL g7576 ( 
.A(n_7012),
.B(n_6005),
.Y(n_7576)
);

INVx1_ASAP7_75t_L g7577 ( 
.A(n_7115),
.Y(n_7577)
);

INVx4_ASAP7_75t_SL g7578 ( 
.A(n_7361),
.Y(n_7578)
);

INVx1_ASAP7_75t_L g7579 ( 
.A(n_7147),
.Y(n_7579)
);

INVx1_ASAP7_75t_L g7580 ( 
.A(n_7147),
.Y(n_7580)
);

AND2x2_ASAP7_75t_L g7581 ( 
.A(n_7090),
.B(n_6986),
.Y(n_7581)
);

BUFx2_ASAP7_75t_L g7582 ( 
.A(n_7439),
.Y(n_7582)
);

NOR2xp33_ASAP7_75t_L g7583 ( 
.A(n_7378),
.B(n_6729),
.Y(n_7583)
);

INVx1_ASAP7_75t_SL g7584 ( 
.A(n_7023),
.Y(n_7584)
);

BUFx2_ASAP7_75t_L g7585 ( 
.A(n_7439),
.Y(n_7585)
);

OA21x2_ASAP7_75t_L g7586 ( 
.A1(n_7320),
.A2(n_6911),
.B(n_6900),
.Y(n_7586)
);

INVx1_ASAP7_75t_L g7587 ( 
.A(n_7150),
.Y(n_7587)
);

INVx1_ASAP7_75t_L g7588 ( 
.A(n_7150),
.Y(n_7588)
);

OAI21x1_ASAP7_75t_L g7589 ( 
.A1(n_7272),
.A2(n_6751),
.B(n_6842),
.Y(n_7589)
);

BUFx2_ASAP7_75t_L g7590 ( 
.A(n_7440),
.Y(n_7590)
);

INVx3_ASAP7_75t_L g7591 ( 
.A(n_7361),
.Y(n_7591)
);

BUFx2_ASAP7_75t_SL g7592 ( 
.A(n_7440),
.Y(n_7592)
);

NAND4xp25_ASAP7_75t_L g7593 ( 
.A(n_7130),
.B(n_6978),
.C(n_6857),
.D(n_6859),
.Y(n_7593)
);

INVx2_ASAP7_75t_L g7594 ( 
.A(n_7361),
.Y(n_7594)
);

AND2x2_ASAP7_75t_L g7595 ( 
.A(n_7012),
.B(n_6842),
.Y(n_7595)
);

AND2x4_ASAP7_75t_L g7596 ( 
.A(n_7447),
.B(n_6857),
.Y(n_7596)
);

INVx4_ASAP7_75t_L g7597 ( 
.A(n_7182),
.Y(n_7597)
);

INVx1_ASAP7_75t_L g7598 ( 
.A(n_7038),
.Y(n_7598)
);

BUFx2_ASAP7_75t_L g7599 ( 
.A(n_7447),
.Y(n_7599)
);

OAI21x1_ASAP7_75t_L g7600 ( 
.A1(n_7311),
.A2(n_7210),
.B(n_7045),
.Y(n_7600)
);

INVx1_ASAP7_75t_L g7601 ( 
.A(n_7038),
.Y(n_7601)
);

AOI21xp5_ASAP7_75t_L g7602 ( 
.A1(n_7164),
.A2(n_6714),
.B(n_6697),
.Y(n_7602)
);

INVx2_ASAP7_75t_L g7603 ( 
.A(n_7371),
.Y(n_7603)
);

AND2x2_ASAP7_75t_L g7604 ( 
.A(n_7030),
.B(n_6859),
.Y(n_7604)
);

INVx1_ASAP7_75t_L g7605 ( 
.A(n_7161),
.Y(n_7605)
);

CKINVDCx5p33_ASAP7_75t_R g7606 ( 
.A(n_7378),
.Y(n_7606)
);

INVx1_ASAP7_75t_L g7607 ( 
.A(n_7161),
.Y(n_7607)
);

AOI211x1_ASAP7_75t_SL g7608 ( 
.A1(n_7132),
.A2(n_6691),
.B(n_6704),
.C(n_6689),
.Y(n_7608)
);

INVx1_ASAP7_75t_L g7609 ( 
.A(n_7175),
.Y(n_7609)
);

NOR2xp33_ASAP7_75t_L g7610 ( 
.A(n_7371),
.B(n_6978),
.Y(n_7610)
);

INVx2_ASAP7_75t_L g7611 ( 
.A(n_7371),
.Y(n_7611)
);

INVx4_ASAP7_75t_SL g7612 ( 
.A(n_7081),
.Y(n_7612)
);

INVx2_ASAP7_75t_L g7613 ( 
.A(n_7162),
.Y(n_7613)
);

NAND2xp5_ASAP7_75t_L g7614 ( 
.A(n_7387),
.B(n_7397),
.Y(n_7614)
);

AOI21xp5_ASAP7_75t_L g7615 ( 
.A1(n_7057),
.A2(n_6697),
.B(n_6990),
.Y(n_7615)
);

INVx1_ASAP7_75t_L g7616 ( 
.A(n_7175),
.Y(n_7616)
);

INVx1_ASAP7_75t_L g7617 ( 
.A(n_7262),
.Y(n_7617)
);

AND2x2_ASAP7_75t_L g7618 ( 
.A(n_7030),
.B(n_6865),
.Y(n_7618)
);

INVx1_ASAP7_75t_L g7619 ( 
.A(n_7262),
.Y(n_7619)
);

HB1xp67_ASAP7_75t_L g7620 ( 
.A(n_7328),
.Y(n_7620)
);

INVx1_ASAP7_75t_L g7621 ( 
.A(n_7328),
.Y(n_7621)
);

INVx2_ASAP7_75t_L g7622 ( 
.A(n_7162),
.Y(n_7622)
);

OAI21x1_ASAP7_75t_L g7623 ( 
.A1(n_7311),
.A2(n_6865),
.B(n_6875),
.Y(n_7623)
);

INVx2_ASAP7_75t_L g7624 ( 
.A(n_7174),
.Y(n_7624)
);

INVx2_ASAP7_75t_L g7625 ( 
.A(n_7174),
.Y(n_7625)
);

AND2x2_ASAP7_75t_L g7626 ( 
.A(n_7034),
.B(n_6847),
.Y(n_7626)
);

INVx2_ASAP7_75t_L g7627 ( 
.A(n_7185),
.Y(n_7627)
);

INVx1_ASAP7_75t_L g7628 ( 
.A(n_7170),
.Y(n_7628)
);

AND2x4_ASAP7_75t_L g7629 ( 
.A(n_7089),
.B(n_6876),
.Y(n_7629)
);

AND2x4_ASAP7_75t_L g7630 ( 
.A(n_7420),
.B(n_6876),
.Y(n_7630)
);

OAI21xp33_ASAP7_75t_L g7631 ( 
.A1(n_7163),
.A2(n_6994),
.B(n_6920),
.Y(n_7631)
);

BUFx3_ASAP7_75t_L g7632 ( 
.A(n_7033),
.Y(n_7632)
);

INVx1_ASAP7_75t_L g7633 ( 
.A(n_7170),
.Y(n_7633)
);

INVx1_ASAP7_75t_L g7634 ( 
.A(n_7172),
.Y(n_7634)
);

INVx1_ASAP7_75t_L g7635 ( 
.A(n_7172),
.Y(n_7635)
);

INVx2_ASAP7_75t_L g7636 ( 
.A(n_7185),
.Y(n_7636)
);

AND2x2_ASAP7_75t_L g7637 ( 
.A(n_7034),
.B(n_6862),
.Y(n_7637)
);

AND2x2_ASAP7_75t_L g7638 ( 
.A(n_7122),
.B(n_6867),
.Y(n_7638)
);

OAI21x1_ASAP7_75t_L g7639 ( 
.A1(n_7210),
.A2(n_6875),
.B(n_6691),
.Y(n_7639)
);

INVx1_ASAP7_75t_L g7640 ( 
.A(n_7173),
.Y(n_7640)
);

AO21x2_ASAP7_75t_L g7641 ( 
.A1(n_7320),
.A2(n_6565),
.B(n_6561),
.Y(n_7641)
);

INVx1_ASAP7_75t_L g7642 ( 
.A(n_7173),
.Y(n_7642)
);

OR2x6_ASAP7_75t_L g7643 ( 
.A(n_7165),
.B(n_6197),
.Y(n_7643)
);

AO21x2_ASAP7_75t_L g7644 ( 
.A1(n_7278),
.A2(n_6565),
.B(n_6561),
.Y(n_7644)
);

INVx2_ASAP7_75t_SL g7645 ( 
.A(n_7183),
.Y(n_7645)
);

INVx1_ASAP7_75t_L g7646 ( 
.A(n_7199),
.Y(n_7646)
);

INVx2_ASAP7_75t_L g7647 ( 
.A(n_7186),
.Y(n_7647)
);

INVx1_ASAP7_75t_L g7648 ( 
.A(n_7199),
.Y(n_7648)
);

A2O1A1Ixp33_ASAP7_75t_L g7649 ( 
.A1(n_7278),
.A2(n_6788),
.B(n_6704),
.C(n_6705),
.Y(n_7649)
);

INVx1_ASAP7_75t_L g7650 ( 
.A(n_7205),
.Y(n_7650)
);

OAI21x1_ASAP7_75t_L g7651 ( 
.A1(n_7416),
.A2(n_6705),
.B(n_6689),
.Y(n_7651)
);

INVx4_ASAP7_75t_L g7652 ( 
.A(n_7182),
.Y(n_7652)
);

INVx1_ASAP7_75t_L g7653 ( 
.A(n_7205),
.Y(n_7653)
);

INVxp67_ASAP7_75t_L g7654 ( 
.A(n_7441),
.Y(n_7654)
);

NOR2x1p5_ASAP7_75t_L g7655 ( 
.A(n_7218),
.B(n_5044),
.Y(n_7655)
);

AO21x2_ASAP7_75t_L g7656 ( 
.A1(n_7014),
.A2(n_6559),
.B(n_6911),
.Y(n_7656)
);

OR2x2_ASAP7_75t_L g7657 ( 
.A(n_7116),
.B(n_6909),
.Y(n_7657)
);

INVx5_ASAP7_75t_L g7658 ( 
.A(n_7182),
.Y(n_7658)
);

INVx3_ASAP7_75t_L g7659 ( 
.A(n_7240),
.Y(n_7659)
);

A2O1A1Ixp33_ASAP7_75t_L g7660 ( 
.A1(n_7163),
.A2(n_6788),
.B(n_6706),
.C(n_6083),
.Y(n_7660)
);

INVx2_ASAP7_75t_L g7661 ( 
.A(n_7186),
.Y(n_7661)
);

NAND2xp5_ASAP7_75t_L g7662 ( 
.A(n_7397),
.B(n_6939),
.Y(n_7662)
);

HB1xp67_ASAP7_75t_L g7663 ( 
.A(n_7121),
.Y(n_7663)
);

AOI21xp5_ASAP7_75t_L g7664 ( 
.A1(n_7201),
.A2(n_7047),
.B(n_7402),
.Y(n_7664)
);

AND2x4_ASAP7_75t_SL g7665 ( 
.A(n_7097),
.B(n_7103),
.Y(n_7665)
);

NOR2x1_ASAP7_75t_L g7666 ( 
.A(n_7441),
.B(n_6949),
.Y(n_7666)
);

A2O1A1Ixp33_ASAP7_75t_L g7667 ( 
.A1(n_7239),
.A2(n_6706),
.B(n_6046),
.C(n_6869),
.Y(n_7667)
);

INVxp67_ASAP7_75t_SL g7668 ( 
.A(n_7424),
.Y(n_7668)
);

HB1xp67_ASAP7_75t_L g7669 ( 
.A(n_7234),
.Y(n_7669)
);

INVx2_ASAP7_75t_L g7670 ( 
.A(n_7187),
.Y(n_7670)
);

INVx2_ASAP7_75t_L g7671 ( 
.A(n_7187),
.Y(n_7671)
);

INVx1_ASAP7_75t_L g7672 ( 
.A(n_7207),
.Y(n_7672)
);

INVx1_ASAP7_75t_L g7673 ( 
.A(n_7207),
.Y(n_7673)
);

OA21x2_ASAP7_75t_L g7674 ( 
.A1(n_7169),
.A2(n_6914),
.B(n_6912),
.Y(n_7674)
);

AOI21xp5_ASAP7_75t_L g7675 ( 
.A1(n_7047),
.A2(n_6697),
.B(n_6197),
.Y(n_7675)
);

INVx1_ASAP7_75t_L g7676 ( 
.A(n_7151),
.Y(n_7676)
);

AND2x4_ASAP7_75t_SL g7677 ( 
.A(n_7096),
.B(n_5044),
.Y(n_7677)
);

OR2x2_ASAP7_75t_L g7678 ( 
.A(n_7120),
.B(n_6942),
.Y(n_7678)
);

AND2x2_ASAP7_75t_L g7679 ( 
.A(n_7122),
.B(n_6874),
.Y(n_7679)
);

AND2x2_ASAP7_75t_L g7680 ( 
.A(n_7052),
.B(n_6639),
.Y(n_7680)
);

A2O1A1Ixp33_ASAP7_75t_L g7681 ( 
.A1(n_7438),
.A2(n_6869),
.B(n_6896),
.C(n_6881),
.Y(n_7681)
);

INVx4_ASAP7_75t_R g7682 ( 
.A(n_7165),
.Y(n_7682)
);

INVx2_ASAP7_75t_L g7683 ( 
.A(n_7189),
.Y(n_7683)
);

INVxp67_ASAP7_75t_L g7684 ( 
.A(n_7039),
.Y(n_7684)
);

INVx1_ASAP7_75t_L g7685 ( 
.A(n_7151),
.Y(n_7685)
);

INVxp67_ASAP7_75t_SL g7686 ( 
.A(n_7424),
.Y(n_7686)
);

AO21x2_ASAP7_75t_L g7687 ( 
.A1(n_7022),
.A2(n_6559),
.B(n_6912),
.Y(n_7687)
);

AO21x2_ASAP7_75t_L g7688 ( 
.A1(n_7024),
.A2(n_6915),
.B(n_6914),
.Y(n_7688)
);

INVx4_ASAP7_75t_L g7689 ( 
.A(n_7079),
.Y(n_7689)
);

NAND2xp5_ASAP7_75t_L g7690 ( 
.A(n_7437),
.B(n_6946),
.Y(n_7690)
);

INVxp67_ASAP7_75t_SL g7691 ( 
.A(n_7288),
.Y(n_7691)
);

BUFx2_ASAP7_75t_L g7692 ( 
.A(n_7019),
.Y(n_7692)
);

NAND2xp5_ASAP7_75t_L g7693 ( 
.A(n_7437),
.B(n_7296),
.Y(n_7693)
);

INVx2_ASAP7_75t_L g7694 ( 
.A(n_7189),
.Y(n_7694)
);

INVx1_ASAP7_75t_L g7695 ( 
.A(n_7153),
.Y(n_7695)
);

INVx1_ASAP7_75t_L g7696 ( 
.A(n_7153),
.Y(n_7696)
);

INVx2_ASAP7_75t_L g7697 ( 
.A(n_7381),
.Y(n_7697)
);

AOI22xp5_ASAP7_75t_L g7698 ( 
.A1(n_7438),
.A2(n_6881),
.B1(n_6896),
.B2(n_6197),
.Y(n_7698)
);

INVx1_ASAP7_75t_L g7699 ( 
.A(n_7154),
.Y(n_7699)
);

INVx1_ASAP7_75t_L g7700 ( 
.A(n_7154),
.Y(n_7700)
);

AND2x2_ASAP7_75t_L g7701 ( 
.A(n_7052),
.B(n_6639),
.Y(n_7701)
);

OAI21x1_ASAP7_75t_L g7702 ( 
.A1(n_7416),
.A2(n_6927),
.B(n_6915),
.Y(n_7702)
);

NAND2xp5_ASAP7_75t_L g7703 ( 
.A(n_7028),
.B(n_6951),
.Y(n_7703)
);

OR2x2_ASAP7_75t_L g7704 ( 
.A(n_7144),
.B(n_6972),
.Y(n_7704)
);

BUFx3_ASAP7_75t_L g7705 ( 
.A(n_7420),
.Y(n_7705)
);

INVx3_ASAP7_75t_L g7706 ( 
.A(n_7240),
.Y(n_7706)
);

BUFx6f_ASAP7_75t_L g7707 ( 
.A(n_7211),
.Y(n_7707)
);

INVx2_ASAP7_75t_L g7708 ( 
.A(n_7381),
.Y(n_7708)
);

INVx2_ASAP7_75t_L g7709 ( 
.A(n_7381),
.Y(n_7709)
);

INVx2_ASAP7_75t_L g7710 ( 
.A(n_7080),
.Y(n_7710)
);

NAND2xp5_ASAP7_75t_L g7711 ( 
.A(n_7244),
.B(n_6960),
.Y(n_7711)
);

AOI21xp33_ASAP7_75t_L g7712 ( 
.A1(n_7088),
.A2(n_6918),
.B(n_6703),
.Y(n_7712)
);

AO21x2_ASAP7_75t_L g7713 ( 
.A1(n_7176),
.A2(n_7180),
.B(n_7177),
.Y(n_7713)
);

INVx1_ASAP7_75t_L g7714 ( 
.A(n_7113),
.Y(n_7714)
);

AOI21xp33_ASAP7_75t_L g7715 ( 
.A1(n_7214),
.A2(n_6918),
.B(n_6703),
.Y(n_7715)
);

A2O1A1Ixp33_ASAP7_75t_L g7716 ( 
.A1(n_7438),
.A2(n_6107),
.B(n_6935),
.C(n_6927),
.Y(n_7716)
);

AOI21xp5_ASAP7_75t_L g7717 ( 
.A1(n_7202),
.A2(n_6675),
.B(n_6947),
.Y(n_7717)
);

INVxp67_ASAP7_75t_SL g7718 ( 
.A(n_7294),
.Y(n_7718)
);

INVx1_ASAP7_75t_L g7719 ( 
.A(n_7117),
.Y(n_7719)
);

HB1xp67_ASAP7_75t_L g7720 ( 
.A(n_7253),
.Y(n_7720)
);

NAND2xp5_ASAP7_75t_SL g7721 ( 
.A(n_7019),
.B(n_7029),
.Y(n_7721)
);

OAI31xp33_ASAP7_75t_SL g7722 ( 
.A1(n_7240),
.A2(n_6876),
.A3(n_6931),
.B(n_6897),
.Y(n_7722)
);

INVx2_ASAP7_75t_L g7723 ( 
.A(n_7080),
.Y(n_7723)
);

NAND2xp5_ASAP7_75t_L g7724 ( 
.A(n_7215),
.B(n_6962),
.Y(n_7724)
);

OR2x2_ASAP7_75t_L g7725 ( 
.A(n_7196),
.B(n_6980),
.Y(n_7725)
);

AOI21xp33_ASAP7_75t_L g7726 ( 
.A1(n_7214),
.A2(n_6918),
.B(n_6675),
.Y(n_7726)
);

NAND2xp5_ASAP7_75t_SL g7727 ( 
.A(n_7019),
.B(n_6991),
.Y(n_7727)
);

NAND2xp5_ASAP7_75t_SL g7728 ( 
.A(n_7029),
.B(n_6991),
.Y(n_7728)
);

INVx2_ASAP7_75t_L g7729 ( 
.A(n_7192),
.Y(n_7729)
);

NAND3xp33_ASAP7_75t_L g7730 ( 
.A(n_7031),
.B(n_6918),
.C(n_6947),
.Y(n_7730)
);

INVx2_ASAP7_75t_L g7731 ( 
.A(n_7192),
.Y(n_7731)
);

AOI21xp5_ASAP7_75t_L g7732 ( 
.A1(n_7188),
.A2(n_6957),
.B(n_6989),
.Y(n_7732)
);

AOI21xp5_ASAP7_75t_SL g7733 ( 
.A1(n_7026),
.A2(n_6957),
.B(n_6931),
.Y(n_7733)
);

INVx2_ASAP7_75t_L g7734 ( 
.A(n_7193),
.Y(n_7734)
);

AND2x2_ASAP7_75t_L g7735 ( 
.A(n_7072),
.B(n_6655),
.Y(n_7735)
);

INVx2_ASAP7_75t_L g7736 ( 
.A(n_7193),
.Y(n_7736)
);

AND2x2_ASAP7_75t_L g7737 ( 
.A(n_7072),
.B(n_6655),
.Y(n_7737)
);

INVx3_ASAP7_75t_L g7738 ( 
.A(n_7309),
.Y(n_7738)
);

OA21x2_ASAP7_75t_L g7739 ( 
.A1(n_7355),
.A2(n_6935),
.B(n_6979),
.Y(n_7739)
);

INVx2_ASAP7_75t_L g7740 ( 
.A(n_7211),
.Y(n_7740)
);

NAND2xp5_ASAP7_75t_SL g7741 ( 
.A(n_7029),
.B(n_6897),
.Y(n_7741)
);

INVx1_ASAP7_75t_L g7742 ( 
.A(n_7123),
.Y(n_7742)
);

INVx1_ASAP7_75t_L g7743 ( 
.A(n_7125),
.Y(n_7743)
);

INVx1_ASAP7_75t_L g7744 ( 
.A(n_7127),
.Y(n_7744)
);

OR2x2_ASAP7_75t_L g7745 ( 
.A(n_7167),
.B(n_6964),
.Y(n_7745)
);

NAND2xp5_ASAP7_75t_L g7746 ( 
.A(n_7274),
.B(n_6966),
.Y(n_7746)
);

AOI21xp33_ASAP7_75t_L g7747 ( 
.A1(n_7224),
.A2(n_6613),
.B(n_6612),
.Y(n_7747)
);

INVx2_ASAP7_75t_L g7748 ( 
.A(n_7211),
.Y(n_7748)
);

INVx1_ASAP7_75t_L g7749 ( 
.A(n_7131),
.Y(n_7749)
);

INVx1_ASAP7_75t_L g7750 ( 
.A(n_7141),
.Y(n_7750)
);

INVx1_ASAP7_75t_L g7751 ( 
.A(n_7159),
.Y(n_7751)
);

INVx1_ASAP7_75t_L g7752 ( 
.A(n_7156),
.Y(n_7752)
);

INVx1_ASAP7_75t_L g7753 ( 
.A(n_7156),
.Y(n_7753)
);

OA21x2_ASAP7_75t_L g7754 ( 
.A1(n_7355),
.A2(n_6984),
.B(n_6979),
.Y(n_7754)
);

INVx2_ASAP7_75t_L g7755 ( 
.A(n_7259),
.Y(n_7755)
);

INVx2_ASAP7_75t_L g7756 ( 
.A(n_7259),
.Y(n_7756)
);

INVx1_ASAP7_75t_L g7757 ( 
.A(n_7157),
.Y(n_7757)
);

OR2x2_ASAP7_75t_L g7758 ( 
.A(n_7179),
.B(n_6967),
.Y(n_7758)
);

OR2x2_ASAP7_75t_L g7759 ( 
.A(n_7194),
.B(n_6968),
.Y(n_7759)
);

NAND4xp25_ASAP7_75t_L g7760 ( 
.A(n_7227),
.B(n_7025),
.C(n_7166),
.D(n_7242),
.Y(n_7760)
);

INVx1_ASAP7_75t_L g7761 ( 
.A(n_7157),
.Y(n_7761)
);

INVx2_ASAP7_75t_L g7762 ( 
.A(n_7259),
.Y(n_7762)
);

OAI211xp5_ASAP7_75t_L g7763 ( 
.A1(n_7416),
.A2(n_6371),
.B(n_6407),
.C(n_6368),
.Y(n_7763)
);

AOI21x1_ASAP7_75t_L g7764 ( 
.A1(n_7044),
.A2(n_6931),
.B(n_6897),
.Y(n_7764)
);

OA21x2_ASAP7_75t_L g7765 ( 
.A1(n_7375),
.A2(n_7380),
.B(n_7376),
.Y(n_7765)
);

INVx2_ASAP7_75t_L g7766 ( 
.A(n_7148),
.Y(n_7766)
);

AND2x2_ASAP7_75t_L g7767 ( 
.A(n_7039),
.B(n_6655),
.Y(n_7767)
);

INVx1_ASAP7_75t_L g7768 ( 
.A(n_7160),
.Y(n_7768)
);

INVxp67_ASAP7_75t_SL g7769 ( 
.A(n_7436),
.Y(n_7769)
);

AOI22xp5_ASAP7_75t_L g7770 ( 
.A1(n_7443),
.A2(n_6420),
.B1(n_6408),
.B2(n_6393),
.Y(n_7770)
);

INVx1_ASAP7_75t_L g7771 ( 
.A(n_7160),
.Y(n_7771)
);

INVx1_ASAP7_75t_L g7772 ( 
.A(n_7109),
.Y(n_7772)
);

INVx2_ASAP7_75t_L g7773 ( 
.A(n_7203),
.Y(n_7773)
);

INVx1_ASAP7_75t_L g7774 ( 
.A(n_7110),
.Y(n_7774)
);

AOI21xp5_ASAP7_75t_L g7775 ( 
.A1(n_7143),
.A2(n_6991),
.B(n_6971),
.Y(n_7775)
);

AOI21xp33_ASAP7_75t_L g7776 ( 
.A1(n_7224),
.A2(n_6613),
.B(n_6612),
.Y(n_7776)
);

INVx4_ASAP7_75t_SL g7777 ( 
.A(n_7317),
.Y(n_7777)
);

INVx1_ASAP7_75t_L g7778 ( 
.A(n_7055),
.Y(n_7778)
);

INVx1_ASAP7_75t_SL g7779 ( 
.A(n_7041),
.Y(n_7779)
);

HB1xp67_ASAP7_75t_L g7780 ( 
.A(n_7223),
.Y(n_7780)
);

BUFx3_ASAP7_75t_L g7781 ( 
.A(n_7405),
.Y(n_7781)
);

NAND4xp25_ASAP7_75t_L g7782 ( 
.A(n_7271),
.B(n_6871),
.C(n_6887),
.D(n_6852),
.Y(n_7782)
);

NAND2xp5_ASAP7_75t_SL g7783 ( 
.A(n_7309),
.B(n_6971),
.Y(n_7783)
);

NAND2xp5_ASAP7_75t_SL g7784 ( 
.A(n_7309),
.B(n_6971),
.Y(n_7784)
);

OA21x2_ASAP7_75t_L g7785 ( 
.A1(n_7375),
.A2(n_6985),
.B(n_6984),
.Y(n_7785)
);

OR2x2_ASAP7_75t_L g7786 ( 
.A(n_7289),
.B(n_6970),
.Y(n_7786)
);

INVx1_ASAP7_75t_SL g7787 ( 
.A(n_7041),
.Y(n_7787)
);

O2A1O1Ixp33_ASAP7_75t_L g7788 ( 
.A1(n_7056),
.A2(n_7005),
.B(n_7008),
.C(n_6985),
.Y(n_7788)
);

NOR2xp33_ASAP7_75t_L g7789 ( 
.A(n_7317),
.B(n_6655),
.Y(n_7789)
);

INVx2_ASAP7_75t_L g7790 ( 
.A(n_7203),
.Y(n_7790)
);

BUFx3_ASAP7_75t_L g7791 ( 
.A(n_7203),
.Y(n_7791)
);

AND2x4_ASAP7_75t_L g7792 ( 
.A(n_7209),
.B(n_6996),
.Y(n_7792)
);

OAI21x1_ASAP7_75t_L g7793 ( 
.A1(n_7436),
.A2(n_7316),
.B(n_7443),
.Y(n_7793)
);

NOR3xp33_ASAP7_75t_L g7794 ( 
.A(n_7316),
.B(n_7005),
.C(n_7008),
.Y(n_7794)
);

INVx1_ASAP7_75t_L g7795 ( 
.A(n_7067),
.Y(n_7795)
);

AOI21x1_ASAP7_75t_L g7796 ( 
.A1(n_7078),
.A2(n_6996),
.B(n_6892),
.Y(n_7796)
);

OA21x2_ASAP7_75t_L g7797 ( 
.A1(n_7376),
.A2(n_6179),
.B(n_6178),
.Y(n_7797)
);

INVx2_ASAP7_75t_L g7798 ( 
.A(n_7209),
.Y(n_7798)
);

INVx1_ASAP7_75t_L g7799 ( 
.A(n_7082),
.Y(n_7799)
);

AO22x2_ASAP7_75t_L g7800 ( 
.A1(n_7083),
.A2(n_6621),
.B1(n_6623),
.B2(n_6617),
.Y(n_7800)
);

INVx1_ASAP7_75t_L g7801 ( 
.A(n_7085),
.Y(n_7801)
);

INVx2_ASAP7_75t_SL g7802 ( 
.A(n_7183),
.Y(n_7802)
);

NOR2xp67_ASAP7_75t_L g7803 ( 
.A(n_7413),
.B(n_6996),
.Y(n_7803)
);

A2O1A1Ixp33_ASAP7_75t_L g7804 ( 
.A1(n_7443),
.A2(n_6107),
.B(n_5771),
.C(n_5766),
.Y(n_7804)
);

AND2x2_ASAP7_75t_L g7805 ( 
.A(n_7363),
.B(n_6118),
.Y(n_7805)
);

INVx2_ASAP7_75t_L g7806 ( 
.A(n_7209),
.Y(n_7806)
);

INVx4_ASAP7_75t_SL g7807 ( 
.A(n_7413),
.Y(n_7807)
);

OAI21x1_ASAP7_75t_L g7808 ( 
.A1(n_7436),
.A2(n_6371),
.B(n_6368),
.Y(n_7808)
);

INVx2_ASAP7_75t_SL g7809 ( 
.A(n_7352),
.Y(n_7809)
);

OR2x6_ASAP7_75t_L g7810 ( 
.A(n_7134),
.B(n_6393),
.Y(n_7810)
);

OR2x2_ASAP7_75t_L g7811 ( 
.A(n_7237),
.B(n_6975),
.Y(n_7811)
);

AND2x2_ASAP7_75t_L g7812 ( 
.A(n_7364),
.B(n_7204),
.Y(n_7812)
);

OR2x2_ASAP7_75t_L g7813 ( 
.A(n_7241),
.B(n_7248),
.Y(n_7813)
);

HB1xp67_ASAP7_75t_L g7814 ( 
.A(n_7226),
.Y(n_7814)
);

AO21x2_ASAP7_75t_L g7815 ( 
.A1(n_7086),
.A2(n_6891),
.B(n_6987),
.Y(n_7815)
);

HB1xp67_ASAP7_75t_L g7816 ( 
.A(n_7228),
.Y(n_7816)
);

NAND2xp5_ASAP7_75t_L g7817 ( 
.A(n_7273),
.B(n_7000),
.Y(n_7817)
);

INVx1_ASAP7_75t_L g7818 ( 
.A(n_7092),
.Y(n_7818)
);

INVx2_ASAP7_75t_L g7819 ( 
.A(n_7250),
.Y(n_7819)
);

AND2x2_ASAP7_75t_L g7820 ( 
.A(n_7204),
.B(n_6150),
.Y(n_7820)
);

INVx2_ASAP7_75t_L g7821 ( 
.A(n_7251),
.Y(n_7821)
);

INVx1_ASAP7_75t_L g7822 ( 
.A(n_7449),
.Y(n_7822)
);

OR2x2_ASAP7_75t_L g7823 ( 
.A(n_7813),
.B(n_7347),
.Y(n_7823)
);

NAND2xp5_ASAP7_75t_SL g7824 ( 
.A(n_7466),
.B(n_7460),
.Y(n_7824)
);

AND2x2_ASAP7_75t_L g7825 ( 
.A(n_7451),
.B(n_7208),
.Y(n_7825)
);

AND2x2_ASAP7_75t_L g7826 ( 
.A(n_7812),
.B(n_7208),
.Y(n_7826)
);

OAI211xp5_ASAP7_75t_SL g7827 ( 
.A1(n_7608),
.A2(n_7094),
.B(n_7098),
.C(n_7093),
.Y(n_7827)
);

AOI21xp5_ASAP7_75t_L g7828 ( 
.A1(n_7602),
.A2(n_7143),
.B(n_7287),
.Y(n_7828)
);

INVx1_ASAP7_75t_L g7829 ( 
.A(n_7542),
.Y(n_7829)
);

NOR3xp33_ASAP7_75t_L g7830 ( 
.A(n_7519),
.B(n_7316),
.C(n_7300),
.Y(n_7830)
);

NOR2xp33_ASAP7_75t_L g7831 ( 
.A(n_7461),
.B(n_7079),
.Y(n_7831)
);

NOR3xp33_ASAP7_75t_L g7832 ( 
.A(n_7483),
.B(n_7300),
.C(n_7287),
.Y(n_7832)
);

AOI211x1_ASAP7_75t_L g7833 ( 
.A1(n_7505),
.A2(n_7104),
.B(n_7102),
.C(n_7365),
.Y(n_7833)
);

NAND3xp33_ASAP7_75t_SL g7834 ( 
.A(n_7489),
.B(n_7266),
.C(n_7076),
.Y(n_7834)
);

NAND2xp5_ASAP7_75t_L g7835 ( 
.A(n_7463),
.B(n_7275),
.Y(n_7835)
);

INVx2_ASAP7_75t_SL g7836 ( 
.A(n_7535),
.Y(n_7836)
);

NOR3xp33_ASAP7_75t_L g7837 ( 
.A(n_7510),
.B(n_7225),
.C(n_7213),
.Y(n_7837)
);

NOR2xp33_ASAP7_75t_L g7838 ( 
.A(n_7508),
.B(n_7079),
.Y(n_7838)
);

AND2x2_ASAP7_75t_L g7839 ( 
.A(n_7665),
.B(n_7076),
.Y(n_7839)
);

NOR2xp33_ASAP7_75t_L g7840 ( 
.A(n_7508),
.B(n_7118),
.Y(n_7840)
);

AO21x2_ASAP7_75t_L g7841 ( 
.A1(n_7458),
.A2(n_7260),
.B(n_7247),
.Y(n_7841)
);

NAND2xp5_ASAP7_75t_L g7842 ( 
.A(n_7474),
.B(n_7395),
.Y(n_7842)
);

NAND2xp5_ASAP7_75t_L g7843 ( 
.A(n_7490),
.B(n_7408),
.Y(n_7843)
);

OAI211xp5_ASAP7_75t_L g7844 ( 
.A1(n_7448),
.A2(n_7301),
.B(n_7356),
.C(n_7425),
.Y(n_7844)
);

NAND4xp75_ASAP7_75t_L g7845 ( 
.A(n_7456),
.B(n_7301),
.C(n_7326),
.D(n_7325),
.Y(n_7845)
);

INVx2_ASAP7_75t_L g7846 ( 
.A(n_7572),
.Y(n_7846)
);

AND2x2_ASAP7_75t_L g7847 ( 
.A(n_7475),
.B(n_7612),
.Y(n_7847)
);

INVx2_ASAP7_75t_L g7848 ( 
.A(n_7572),
.Y(n_7848)
);

AND2x2_ASAP7_75t_L g7849 ( 
.A(n_7612),
.B(n_7074),
.Y(n_7849)
);

INVx2_ASAP7_75t_L g7850 ( 
.A(n_7572),
.Y(n_7850)
);

NAND3xp33_ASAP7_75t_L g7851 ( 
.A(n_7546),
.B(n_7158),
.C(n_7118),
.Y(n_7851)
);

NOR3xp33_ASAP7_75t_L g7852 ( 
.A(n_7543),
.B(n_7225),
.C(n_7213),
.Y(n_7852)
);

NAND4xp75_ASAP7_75t_L g7853 ( 
.A(n_7456),
.B(n_7326),
.C(n_7327),
.D(n_7325),
.Y(n_7853)
);

INVx2_ASAP7_75t_L g7854 ( 
.A(n_7764),
.Y(n_7854)
);

AND2x2_ASAP7_75t_L g7855 ( 
.A(n_7604),
.B(n_7074),
.Y(n_7855)
);

AND2x2_ASAP7_75t_L g7856 ( 
.A(n_7618),
.B(n_7136),
.Y(n_7856)
);

NAND2xp5_ASAP7_75t_L g7857 ( 
.A(n_7499),
.B(n_7137),
.Y(n_7857)
);

AND2x2_ASAP7_75t_L g7858 ( 
.A(n_7692),
.B(n_7255),
.Y(n_7858)
);

AND2x4_ASAP7_75t_L g7859 ( 
.A(n_7777),
.B(n_7118),
.Y(n_7859)
);

NAND3xp33_ASAP7_75t_L g7860 ( 
.A(n_7667),
.B(n_7158),
.C(n_7313),
.Y(n_7860)
);

NAND2xp5_ASAP7_75t_L g7861 ( 
.A(n_7584),
.B(n_7158),
.Y(n_7861)
);

NAND4xp75_ASAP7_75t_L g7862 ( 
.A(n_7540),
.B(n_7329),
.C(n_7330),
.D(n_7327),
.Y(n_7862)
);

AOI211xp5_ASAP7_75t_L g7863 ( 
.A1(n_7664),
.A2(n_7615),
.B(n_7562),
.C(n_7600),
.Y(n_7863)
);

NAND2xp5_ASAP7_75t_L g7864 ( 
.A(n_7507),
.B(n_7230),
.Y(n_7864)
);

NAND3xp33_ASAP7_75t_L g7865 ( 
.A(n_7649),
.B(n_7332),
.C(n_7324),
.Y(n_7865)
);

NAND3xp33_ASAP7_75t_L g7866 ( 
.A(n_7660),
.B(n_7340),
.C(n_7106),
.Y(n_7866)
);

NOR2x1_ASAP7_75t_SL g7867 ( 
.A(n_7464),
.B(n_7425),
.Y(n_7867)
);

NAND4xp75_ASAP7_75t_L g7868 ( 
.A(n_7675),
.B(n_7583),
.C(n_7666),
.D(n_7803),
.Y(n_7868)
);

AND2x2_ASAP7_75t_L g7869 ( 
.A(n_7781),
.B(n_7264),
.Y(n_7869)
);

OR2x2_ASAP7_75t_L g7870 ( 
.A(n_7470),
.B(n_7267),
.Y(n_7870)
);

HB1xp67_ASAP7_75t_L g7871 ( 
.A(n_7713),
.Y(n_7871)
);

NAND2xp5_ASAP7_75t_L g7872 ( 
.A(n_7520),
.B(n_7232),
.Y(n_7872)
);

NAND2xp5_ASAP7_75t_L g7873 ( 
.A(n_7779),
.B(n_7406),
.Y(n_7873)
);

INVx2_ASAP7_75t_L g7874 ( 
.A(n_7533),
.Y(n_7874)
);

AOI221xp5_ASAP7_75t_L g7875 ( 
.A1(n_7528),
.A2(n_7238),
.B1(n_7243),
.B2(n_7235),
.C(n_7233),
.Y(n_7875)
);

INVx1_ASAP7_75t_L g7876 ( 
.A(n_7542),
.Y(n_7876)
);

NOR3xp33_ASAP7_75t_L g7877 ( 
.A(n_7473),
.B(n_7748),
.C(n_7740),
.Y(n_7877)
);

NAND4xp75_ASAP7_75t_L g7878 ( 
.A(n_7471),
.B(n_7330),
.C(n_7335),
.D(n_7329),
.Y(n_7878)
);

AND2x2_ASAP7_75t_L g7879 ( 
.A(n_7479),
.B(n_7282),
.Y(n_7879)
);

AO21x2_ASAP7_75t_L g7880 ( 
.A1(n_7458),
.A2(n_7293),
.B(n_7279),
.Y(n_7880)
);

INVx1_ASAP7_75t_L g7881 ( 
.A(n_7547),
.Y(n_7881)
);

NAND2xp5_ASAP7_75t_L g7882 ( 
.A(n_7787),
.B(n_7403),
.Y(n_7882)
);

NAND3xp33_ASAP7_75t_L g7883 ( 
.A(n_7620),
.B(n_7106),
.C(n_7351),
.Y(n_7883)
);

NAND3xp33_ASAP7_75t_L g7884 ( 
.A(n_7614),
.B(n_7430),
.C(n_7426),
.Y(n_7884)
);

NAND3xp33_ASAP7_75t_L g7885 ( 
.A(n_7730),
.B(n_7433),
.C(n_7431),
.Y(n_7885)
);

AND2x2_ASAP7_75t_L g7886 ( 
.A(n_7492),
.B(n_7265),
.Y(n_7886)
);

AND2x2_ASAP7_75t_L g7887 ( 
.A(n_7522),
.B(n_7335),
.Y(n_7887)
);

AND2x2_ASAP7_75t_L g7888 ( 
.A(n_7545),
.B(n_7336),
.Y(n_7888)
);

AND2x2_ASAP7_75t_L g7889 ( 
.A(n_7570),
.B(n_7336),
.Y(n_7889)
);

INVx2_ASAP7_75t_L g7890 ( 
.A(n_7533),
.Y(n_7890)
);

NOR3xp33_ASAP7_75t_L g7891 ( 
.A(n_7473),
.B(n_7235),
.C(n_7233),
.Y(n_7891)
);

AOI22xp5_ASAP7_75t_L g7892 ( 
.A1(n_7468),
.A2(n_7021),
.B1(n_7032),
.B2(n_7027),
.Y(n_7892)
);

NAND3xp33_ASAP7_75t_L g7893 ( 
.A(n_7575),
.B(n_7446),
.C(n_7442),
.Y(n_7893)
);

AND2x2_ASAP7_75t_L g7894 ( 
.A(n_7626),
.B(n_7338),
.Y(n_7894)
);

HB1xp67_ASAP7_75t_L g7895 ( 
.A(n_7815),
.Y(n_7895)
);

AND2x2_ASAP7_75t_L g7896 ( 
.A(n_7581),
.B(n_7595),
.Y(n_7896)
);

AND2x2_ASAP7_75t_L g7897 ( 
.A(n_7553),
.B(n_7338),
.Y(n_7897)
);

NAND3xp33_ASAP7_75t_L g7898 ( 
.A(n_7707),
.B(n_7190),
.C(n_7181),
.Y(n_7898)
);

NAND2xp5_ASAP7_75t_L g7899 ( 
.A(n_7691),
.B(n_7718),
.Y(n_7899)
);

AOI22xp5_ASAP7_75t_L g7900 ( 
.A1(n_7639),
.A2(n_7021),
.B1(n_7032),
.B2(n_7027),
.Y(n_7900)
);

NAND2xp5_ASAP7_75t_L g7901 ( 
.A(n_7582),
.B(n_7370),
.Y(n_7901)
);

NAND3xp33_ASAP7_75t_L g7902 ( 
.A(n_7707),
.B(n_7434),
.C(n_7421),
.Y(n_7902)
);

NOR3xp33_ASAP7_75t_L g7903 ( 
.A(n_7755),
.B(n_7243),
.C(n_7238),
.Y(n_7903)
);

NAND2xp5_ASAP7_75t_L g7904 ( 
.A(n_7585),
.B(n_7391),
.Y(n_7904)
);

NOR3xp33_ASAP7_75t_SL g7905 ( 
.A(n_7606),
.B(n_7435),
.C(n_7427),
.Y(n_7905)
);

OAI211xp5_ASAP7_75t_L g7906 ( 
.A1(n_7796),
.A2(n_7429),
.B(n_7417),
.C(n_7304),
.Y(n_7906)
);

NOR3xp33_ASAP7_75t_L g7907 ( 
.A(n_7756),
.B(n_7762),
.C(n_7506),
.Y(n_7907)
);

AOI221xp5_ASAP7_75t_L g7908 ( 
.A1(n_7800),
.A2(n_7279),
.B1(n_7280),
.B2(n_7260),
.C(n_7247),
.Y(n_7908)
);

OAI211xp5_ASAP7_75t_SL g7909 ( 
.A1(n_7558),
.A2(n_7379),
.B(n_7198),
.C(n_7200),
.Y(n_7909)
);

INVx1_ASAP7_75t_L g7910 ( 
.A(n_7547),
.Y(n_7910)
);

AOI211xp5_ASAP7_75t_L g7911 ( 
.A1(n_7733),
.A2(n_7191),
.B(n_7221),
.C(n_7216),
.Y(n_7911)
);

OR2x2_ASAP7_75t_L g7912 ( 
.A(n_7526),
.B(n_7362),
.Y(n_7912)
);

AOI22xp5_ASAP7_75t_L g7913 ( 
.A1(n_7800),
.A2(n_7035),
.B1(n_7049),
.B2(n_7040),
.Y(n_7913)
);

BUFx2_ASAP7_75t_L g7914 ( 
.A(n_7469),
.Y(n_7914)
);

AND2x2_ASAP7_75t_L g7915 ( 
.A(n_7493),
.B(n_7236),
.Y(n_7915)
);

AND2x2_ASAP7_75t_L g7916 ( 
.A(n_7500),
.B(n_7705),
.Y(n_7916)
);

AOI22xp33_ASAP7_75t_L g7917 ( 
.A1(n_7644),
.A2(n_7386),
.B1(n_7390),
.B2(n_7380),
.Y(n_7917)
);

AND2x2_ASAP7_75t_L g7918 ( 
.A(n_7509),
.B(n_7249),
.Y(n_7918)
);

NAND2xp5_ASAP7_75t_L g7919 ( 
.A(n_7590),
.B(n_7392),
.Y(n_7919)
);

NAND3xp33_ASAP7_75t_L g7920 ( 
.A(n_7465),
.B(n_7245),
.C(n_7231),
.Y(n_7920)
);

INVxp67_ASAP7_75t_SL g7921 ( 
.A(n_7535),
.Y(n_7921)
);

NAND2xp5_ASAP7_75t_L g7922 ( 
.A(n_7599),
.B(n_7155),
.Y(n_7922)
);

OAI211xp5_ASAP7_75t_SL g7923 ( 
.A1(n_7654),
.A2(n_7252),
.B(n_7257),
.C(n_7246),
.Y(n_7923)
);

AND2x2_ASAP7_75t_L g7924 ( 
.A(n_7521),
.B(n_7349),
.Y(n_7924)
);

NAND3xp33_ASAP7_75t_L g7925 ( 
.A(n_7465),
.B(n_7261),
.C(n_7258),
.Y(n_7925)
);

NOR2x1_ASAP7_75t_L g7926 ( 
.A(n_7523),
.B(n_7352),
.Y(n_7926)
);

AND2x2_ASAP7_75t_L g7927 ( 
.A(n_7537),
.B(n_7149),
.Y(n_7927)
);

NAND3xp33_ASAP7_75t_SL g7928 ( 
.A(n_7524),
.B(n_7266),
.C(n_7429),
.Y(n_7928)
);

AND2x2_ASAP7_75t_L g7929 ( 
.A(n_7632),
.B(n_7152),
.Y(n_7929)
);

NAND2xp5_ASAP7_75t_L g7930 ( 
.A(n_7780),
.B(n_7394),
.Y(n_7930)
);

OR2x2_ASAP7_75t_L g7931 ( 
.A(n_7486),
.B(n_7359),
.Y(n_7931)
);

NAND2xp5_ASAP7_75t_L g7932 ( 
.A(n_7814),
.B(n_7414),
.Y(n_7932)
);

OR2x2_ASAP7_75t_L g7933 ( 
.A(n_7467),
.B(n_7422),
.Y(n_7933)
);

AND2x2_ASAP7_75t_L g7934 ( 
.A(n_7816),
.B(n_7217),
.Y(n_7934)
);

AND2x2_ASAP7_75t_L g7935 ( 
.A(n_7637),
.B(n_7269),
.Y(n_7935)
);

NOR2xp33_ASAP7_75t_L g7936 ( 
.A(n_7450),
.B(n_7352),
.Y(n_7936)
);

NAND2xp5_ASAP7_75t_L g7937 ( 
.A(n_7766),
.B(n_7710),
.Y(n_7937)
);

XNOR2x1_ASAP7_75t_L g7938 ( 
.A(n_7697),
.B(n_7035),
.Y(n_7938)
);

NAND3xp33_ASAP7_75t_L g7939 ( 
.A(n_7707),
.B(n_7277),
.C(n_7270),
.Y(n_7939)
);

NOR2x1_ASAP7_75t_L g7940 ( 
.A(n_7485),
.B(n_7417),
.Y(n_7940)
);

NOR2xp33_ASAP7_75t_L g7941 ( 
.A(n_7450),
.B(n_7323),
.Y(n_7941)
);

INVx1_ASAP7_75t_SL g7942 ( 
.A(n_7576),
.Y(n_7942)
);

AOI22xp33_ASAP7_75t_L g7943 ( 
.A1(n_7635),
.A2(n_7390),
.B1(n_7399),
.B2(n_7386),
.Y(n_7943)
);

AND2x2_ASAP7_75t_L g7944 ( 
.A(n_7630),
.B(n_7366),
.Y(n_7944)
);

NOR3xp33_ASAP7_75t_L g7945 ( 
.A(n_7480),
.B(n_7284),
.C(n_7280),
.Y(n_7945)
);

AND2x2_ASAP7_75t_L g7946 ( 
.A(n_7630),
.B(n_7368),
.Y(n_7946)
);

OR2x2_ASAP7_75t_L g7947 ( 
.A(n_7693),
.B(n_7299),
.Y(n_7947)
);

INVx2_ASAP7_75t_L g7948 ( 
.A(n_7578),
.Y(n_7948)
);

INVx1_ASAP7_75t_L g7949 ( 
.A(n_7550),
.Y(n_7949)
);

OAI211xp5_ASAP7_75t_L g7950 ( 
.A1(n_7668),
.A2(n_7304),
.B(n_7281),
.C(n_7291),
.Y(n_7950)
);

NAND3xp33_ASAP7_75t_L g7951 ( 
.A(n_7549),
.B(n_7297),
.C(n_7286),
.Y(n_7951)
);

INVx1_ASAP7_75t_L g7952 ( 
.A(n_7550),
.Y(n_7952)
);

INVx1_ASAP7_75t_L g7953 ( 
.A(n_7552),
.Y(n_7953)
);

NAND3xp33_ASAP7_75t_L g7954 ( 
.A(n_7459),
.B(n_7307),
.C(n_7303),
.Y(n_7954)
);

INVx1_ASAP7_75t_L g7955 ( 
.A(n_7552),
.Y(n_7955)
);

AOI22xp33_ASAP7_75t_L g7956 ( 
.A1(n_7635),
.A2(n_7410),
.B1(n_7399),
.B2(n_7415),
.Y(n_7956)
);

NAND4xp75_ASAP7_75t_L g7957 ( 
.A(n_7555),
.B(n_7060),
.C(n_7062),
.D(n_7059),
.Y(n_7957)
);

OAI211xp5_ASAP7_75t_L g7958 ( 
.A1(n_7686),
.A2(n_7321),
.B(n_7333),
.C(n_7315),
.Y(n_7958)
);

AND2x2_ASAP7_75t_L g7959 ( 
.A(n_7638),
.B(n_7369),
.Y(n_7959)
);

NOR2x1_ASAP7_75t_L g7960 ( 
.A(n_7491),
.B(n_7339),
.Y(n_7960)
);

NAND4xp75_ASAP7_75t_L g7961 ( 
.A(n_7775),
.B(n_7809),
.C(n_7717),
.D(n_7726),
.Y(n_7961)
);

NAND2xp5_ASAP7_75t_L g7962 ( 
.A(n_7723),
.B(n_7407),
.Y(n_7962)
);

NOR2xp33_ASAP7_75t_L g7963 ( 
.A(n_7450),
.B(n_7341),
.Y(n_7963)
);

INVxp67_ASAP7_75t_L g7964 ( 
.A(n_7531),
.Y(n_7964)
);

INVx1_ASAP7_75t_L g7965 ( 
.A(n_7554),
.Y(n_7965)
);

NAND3xp33_ASAP7_75t_L g7966 ( 
.A(n_7478),
.B(n_7358),
.C(n_7345),
.Y(n_7966)
);

AND2x2_ASAP7_75t_L g7967 ( 
.A(n_7679),
.B(n_7729),
.Y(n_7967)
);

AND2x2_ASAP7_75t_L g7968 ( 
.A(n_7731),
.B(n_7372),
.Y(n_7968)
);

NAND3xp33_ASAP7_75t_L g7969 ( 
.A(n_7478),
.B(n_7374),
.C(n_7367),
.Y(n_7969)
);

NOR3xp33_ASAP7_75t_L g7970 ( 
.A(n_7480),
.B(n_7290),
.C(n_7284),
.Y(n_7970)
);

AND2x2_ASAP7_75t_L g7971 ( 
.A(n_7734),
.B(n_7382),
.Y(n_7971)
);

NOR3xp33_ASAP7_75t_L g7972 ( 
.A(n_7506),
.B(n_7292),
.C(n_7290),
.Y(n_7972)
);

OAI31xp33_ASAP7_75t_L g7973 ( 
.A1(n_7631),
.A2(n_7410),
.A3(n_7049),
.B(n_7040),
.Y(n_7973)
);

OAI211xp5_ASAP7_75t_SL g7974 ( 
.A1(n_7715),
.A2(n_7384),
.B(n_7385),
.C(n_7377),
.Y(n_7974)
);

INVx2_ASAP7_75t_L g7975 ( 
.A(n_7578),
.Y(n_7975)
);

OA211x2_ASAP7_75t_L g7976 ( 
.A1(n_7721),
.A2(n_6597),
.B(n_6535),
.C(n_6237),
.Y(n_7976)
);

NAND3xp33_ASAP7_75t_L g7977 ( 
.A(n_7531),
.B(n_7393),
.C(n_7389),
.Y(n_7977)
);

INVx1_ASAP7_75t_SL g7978 ( 
.A(n_7566),
.Y(n_7978)
);

NAND2x1_ASAP7_75t_L g7979 ( 
.A(n_7682),
.B(n_7306),
.Y(n_7979)
);

INVx2_ASAP7_75t_L g7980 ( 
.A(n_7563),
.Y(n_7980)
);

NOR2xp33_ASAP7_75t_L g7981 ( 
.A(n_7462),
.B(n_7343),
.Y(n_7981)
);

NAND2xp5_ASAP7_75t_L g7982 ( 
.A(n_7736),
.B(n_7412),
.Y(n_7982)
);

NAND3xp33_ASAP7_75t_L g7983 ( 
.A(n_7539),
.B(n_7401),
.C(n_7396),
.Y(n_7983)
);

AND2x2_ASAP7_75t_L g7984 ( 
.A(n_7767),
.B(n_7388),
.Y(n_7984)
);

NAND3xp33_ASAP7_75t_L g7985 ( 
.A(n_7539),
.B(n_7411),
.C(n_7409),
.Y(n_7985)
);

AND2x2_ASAP7_75t_L g7986 ( 
.A(n_7566),
.B(n_7254),
.Y(n_7986)
);

AOI22xp33_ASAP7_75t_L g7987 ( 
.A1(n_7628),
.A2(n_7634),
.B1(n_7640),
.B2(n_7633),
.Y(n_7987)
);

NOR3xp33_ASAP7_75t_L g7988 ( 
.A(n_7591),
.B(n_7293),
.C(n_7292),
.Y(n_7988)
);

NOR2xp33_ASAP7_75t_L g7989 ( 
.A(n_7462),
.B(n_7306),
.Y(n_7989)
);

OR2x2_ASAP7_75t_L g7990 ( 
.A(n_7517),
.B(n_7314),
.Y(n_7990)
);

NOR2xp33_ASAP7_75t_L g7991 ( 
.A(n_7462),
.B(n_7312),
.Y(n_7991)
);

AOI22xp33_ASAP7_75t_L g7992 ( 
.A1(n_7642),
.A2(n_7418),
.B1(n_7419),
.B2(n_7415),
.Y(n_7992)
);

AND2x4_ASAP7_75t_L g7993 ( 
.A(n_7777),
.B(n_7256),
.Y(n_7993)
);

NOR3xp33_ASAP7_75t_L g7994 ( 
.A(n_7591),
.B(n_7305),
.C(n_7302),
.Y(n_7994)
);

NAND3xp33_ASAP7_75t_L g7995 ( 
.A(n_7689),
.B(n_7669),
.C(n_7663),
.Y(n_7995)
);

NAND3xp33_ASAP7_75t_L g7996 ( 
.A(n_7689),
.B(n_7481),
.C(n_7563),
.Y(n_7996)
);

AND2x2_ASAP7_75t_L g7997 ( 
.A(n_7735),
.B(n_7254),
.Y(n_7997)
);

INVx2_ASAP7_75t_L g7998 ( 
.A(n_7563),
.Y(n_7998)
);

NAND2xp5_ASAP7_75t_L g7999 ( 
.A(n_7684),
.B(n_7348),
.Y(n_7999)
);

BUFx2_ASAP7_75t_L g8000 ( 
.A(n_7469),
.Y(n_8000)
);

AOI22xp33_ASAP7_75t_L g8001 ( 
.A1(n_7646),
.A2(n_7650),
.B1(n_7653),
.B2(n_7648),
.Y(n_8001)
);

AND2x2_ASAP7_75t_L g8002 ( 
.A(n_7737),
.B(n_7312),
.Y(n_8002)
);

AND2x2_ASAP7_75t_L g8003 ( 
.A(n_7488),
.B(n_6150),
.Y(n_8003)
);

NAND3xp33_ASAP7_75t_L g8004 ( 
.A(n_7605),
.B(n_7305),
.C(n_7302),
.Y(n_8004)
);

INVx1_ASAP7_75t_L g8005 ( 
.A(n_7554),
.Y(n_8005)
);

AND2x2_ASAP7_75t_L g8006 ( 
.A(n_7574),
.B(n_6180),
.Y(n_8006)
);

NAND3xp33_ASAP7_75t_L g8007 ( 
.A(n_7607),
.B(n_7616),
.C(n_7609),
.Y(n_8007)
);

OR2x2_ASAP7_75t_L g8008 ( 
.A(n_7530),
.B(n_7001),
.Y(n_8008)
);

NAND3xp33_ASAP7_75t_L g8009 ( 
.A(n_7617),
.B(n_7310),
.C(n_7308),
.Y(n_8009)
);

NOR2xp33_ASAP7_75t_L g8010 ( 
.A(n_7487),
.B(n_4774),
.Y(n_8010)
);

OR2x2_ASAP7_75t_L g8011 ( 
.A(n_7657),
.B(n_7002),
.Y(n_8011)
);

AOI22xp5_ASAP7_75t_L g8012 ( 
.A1(n_7672),
.A2(n_7419),
.B1(n_7423),
.B2(n_7418),
.Y(n_8012)
);

INVx2_ASAP7_75t_SL g8013 ( 
.A(n_7534),
.Y(n_8013)
);

INVx1_ASAP7_75t_L g8014 ( 
.A(n_7568),
.Y(n_8014)
);

NOR3xp33_ASAP7_75t_L g8015 ( 
.A(n_7659),
.B(n_7310),
.C(n_7308),
.Y(n_8015)
);

NOR2xp33_ASAP7_75t_L g8016 ( 
.A(n_7487),
.B(n_4874),
.Y(n_8016)
);

AOI221xp5_ASAP7_75t_L g8017 ( 
.A1(n_7794),
.A2(n_7444),
.B1(n_7428),
.B2(n_7423),
.C(n_7445),
.Y(n_8017)
);

AND2x2_ASAP7_75t_L g8018 ( 
.A(n_7820),
.B(n_6180),
.Y(n_8018)
);

AOI22xp33_ASAP7_75t_L g8019 ( 
.A1(n_7673),
.A2(n_7753),
.B1(n_7757),
.B2(n_7752),
.Y(n_8019)
);

NAND3xp33_ASAP7_75t_L g8020 ( 
.A(n_7476),
.B(n_7444),
.C(n_7428),
.Y(n_8020)
);

AO21x2_ASAP7_75t_L g8021 ( 
.A1(n_7453),
.A2(n_7445),
.B(n_7337),
.Y(n_8021)
);

NAND2xp5_ASAP7_75t_L g8022 ( 
.A(n_7477),
.B(n_6267),
.Y(n_8022)
);

OR2x2_ASAP7_75t_L g8023 ( 
.A(n_7725),
.B(n_7571),
.Y(n_8023)
);

NOR2xp33_ASAP7_75t_L g8024 ( 
.A(n_7487),
.B(n_4887),
.Y(n_8024)
);

NAND2xp5_ASAP7_75t_L g8025 ( 
.A(n_7564),
.B(n_6271),
.Y(n_8025)
);

NOR3xp33_ASAP7_75t_L g8026 ( 
.A(n_7659),
.B(n_7346),
.C(n_7344),
.Y(n_8026)
);

AND2x2_ASAP7_75t_L g8027 ( 
.A(n_7629),
.B(n_6187),
.Y(n_8027)
);

AND2x2_ASAP7_75t_L g8028 ( 
.A(n_7629),
.B(n_7792),
.Y(n_8028)
);

AOI22xp33_ASAP7_75t_SL g8029 ( 
.A1(n_7561),
.A2(n_6928),
.B1(n_7007),
.B2(n_7322),
.Y(n_8029)
);

AND2x2_ASAP7_75t_L g8030 ( 
.A(n_7792),
.B(n_7680),
.Y(n_8030)
);

NAND4xp25_ASAP7_75t_L g8031 ( 
.A(n_7511),
.B(n_6371),
.C(n_6407),
.D(n_6368),
.Y(n_8031)
);

AND2x2_ASAP7_75t_L g8032 ( 
.A(n_7701),
.B(n_6187),
.Y(n_8032)
);

HB1xp67_ASAP7_75t_L g8033 ( 
.A(n_7807),
.Y(n_8033)
);

INVx1_ASAP7_75t_L g8034 ( 
.A(n_7568),
.Y(n_8034)
);

NAND2xp5_ASAP7_75t_L g8035 ( 
.A(n_7720),
.B(n_7534),
.Y(n_8035)
);

OR2x2_ASAP7_75t_L g8036 ( 
.A(n_7678),
.B(n_6276),
.Y(n_8036)
);

NOR3xp33_ASAP7_75t_L g8037 ( 
.A(n_7706),
.B(n_7337),
.C(n_7322),
.Y(n_8037)
);

NAND4xp75_ASAP7_75t_L g8038 ( 
.A(n_7712),
.B(n_7060),
.C(n_7062),
.D(n_7059),
.Y(n_8038)
);

AO21x2_ASAP7_75t_L g8039 ( 
.A1(n_7453),
.A2(n_7344),
.B(n_7342),
.Y(n_8039)
);

NAND4xp75_ASAP7_75t_L g8040 ( 
.A(n_7770),
.B(n_7065),
.C(n_7066),
.D(n_7063),
.Y(n_8040)
);

NOR3xp33_ASAP7_75t_L g8041 ( 
.A(n_7706),
.B(n_7346),
.C(n_7342),
.Y(n_8041)
);

OAI211xp5_ASAP7_75t_L g8042 ( 
.A1(n_7722),
.A2(n_6440),
.B(n_6476),
.C(n_6407),
.Y(n_8042)
);

BUFx2_ASAP7_75t_L g8043 ( 
.A(n_7469),
.Y(n_8043)
);

INVx1_ASAP7_75t_L g8044 ( 
.A(n_7495),
.Y(n_8044)
);

AND2x2_ASAP7_75t_L g8045 ( 
.A(n_7805),
.B(n_6440),
.Y(n_8045)
);

NAND2xp5_ASAP7_75t_L g8046 ( 
.A(n_7501),
.B(n_6273),
.Y(n_8046)
);

AND2x2_ASAP7_75t_L g8047 ( 
.A(n_7807),
.B(n_6440),
.Y(n_8047)
);

AND2x4_ASAP7_75t_L g8048 ( 
.A(n_7454),
.B(n_6476),
.Y(n_8048)
);

HB1xp67_ASAP7_75t_L g8049 ( 
.A(n_7613),
.Y(n_8049)
);

AND2x2_ASAP7_75t_L g8050 ( 
.A(n_7532),
.B(n_6476),
.Y(n_8050)
);

AOI221xp5_ASAP7_75t_L g8051 ( 
.A1(n_7747),
.A2(n_7350),
.B1(n_7066),
.B2(n_7068),
.C(n_7065),
.Y(n_8051)
);

OR2x2_ASAP7_75t_L g8052 ( 
.A(n_7704),
.B(n_6279),
.Y(n_8052)
);

NOR3xp33_ASAP7_75t_L g8053 ( 
.A(n_7738),
.B(n_7350),
.C(n_7068),
.Y(n_8053)
);

AOI21x1_ASAP7_75t_L g8054 ( 
.A1(n_7455),
.A2(n_7070),
.B(n_7063),
.Y(n_8054)
);

OR2x2_ASAP7_75t_L g8055 ( 
.A(n_7758),
.B(n_6295),
.Y(n_8055)
);

NAND2xp33_ASAP7_75t_SL g8056 ( 
.A(n_7759),
.B(n_4917),
.Y(n_8056)
);

NOR2x1_ASAP7_75t_L g8057 ( 
.A(n_7592),
.B(n_7119),
.Y(n_8057)
);

NAND3xp33_ASAP7_75t_L g8058 ( 
.A(n_7619),
.B(n_7071),
.C(n_7070),
.Y(n_8058)
);

AND2x2_ASAP7_75t_L g8059 ( 
.A(n_7559),
.B(n_7460),
.Y(n_8059)
);

NAND2xp5_ASAP7_75t_L g8060 ( 
.A(n_7513),
.B(n_6274),
.Y(n_8060)
);

AOI21x1_ASAP7_75t_L g8061 ( 
.A1(n_7455),
.A2(n_7101),
.B(n_7071),
.Y(n_8061)
);

AND2x2_ASAP7_75t_L g8062 ( 
.A(n_7622),
.B(n_6516),
.Y(n_8062)
);

AOI22xp33_ASAP7_75t_L g8063 ( 
.A1(n_7752),
.A2(n_7101),
.B1(n_7119),
.B2(n_7108),
.Y(n_8063)
);

OR2x2_ASAP7_75t_L g8064 ( 
.A(n_7811),
.B(n_6323),
.Y(n_8064)
);

NAND2xp5_ASAP7_75t_L g8065 ( 
.A(n_7516),
.B(n_6285),
.Y(n_8065)
);

NAND2xp5_ASAP7_75t_L g8066 ( 
.A(n_7525),
.B(n_6288),
.Y(n_8066)
);

INVx2_ASAP7_75t_L g8067 ( 
.A(n_7738),
.Y(n_8067)
);

INVx1_ASAP7_75t_L g8068 ( 
.A(n_7498),
.Y(n_8068)
);

AND2x4_ASAP7_75t_L g8069 ( 
.A(n_7454),
.B(n_6516),
.Y(n_8069)
);

NOR3xp33_ASAP7_75t_L g8070 ( 
.A(n_7769),
.B(n_7126),
.C(n_7108),
.Y(n_8070)
);

NOR2xp33_ASAP7_75t_L g8071 ( 
.A(n_7452),
.B(n_6516),
.Y(n_8071)
);

NAND3xp33_ASAP7_75t_SL g8072 ( 
.A(n_7763),
.B(n_7128),
.C(n_7126),
.Y(n_8072)
);

AOI221xp5_ASAP7_75t_L g8073 ( 
.A1(n_7776),
.A2(n_7135),
.B1(n_7138),
.B2(n_7129),
.C(n_7128),
.Y(n_8073)
);

NAND2xp5_ASAP7_75t_SL g8074 ( 
.A(n_7497),
.B(n_6535),
.Y(n_8074)
);

AND2x2_ASAP7_75t_L g8075 ( 
.A(n_7624),
.B(n_6543),
.Y(n_8075)
);

NOR2x1_ASAP7_75t_L g8076 ( 
.A(n_7597),
.B(n_7129),
.Y(n_8076)
);

OAI211xp5_ASAP7_75t_L g8077 ( 
.A1(n_7529),
.A2(n_6543),
.B(n_5084),
.C(n_5136),
.Y(n_8077)
);

AOI22xp33_ASAP7_75t_L g8078 ( 
.A1(n_7753),
.A2(n_7135),
.B1(n_7139),
.B2(n_7138),
.Y(n_8078)
);

HB1xp67_ASAP7_75t_L g8079 ( 
.A(n_7625),
.Y(n_8079)
);

AND2x2_ASAP7_75t_L g8080 ( 
.A(n_7627),
.B(n_6543),
.Y(n_8080)
);

INVxp67_ASAP7_75t_SL g8081 ( 
.A(n_7791),
.Y(n_8081)
);

AO21x2_ASAP7_75t_L g8082 ( 
.A1(n_7641),
.A2(n_7140),
.B(n_7139),
.Y(n_8082)
);

AND2x2_ASAP7_75t_L g8083 ( 
.A(n_7636),
.B(n_5716),
.Y(n_8083)
);

NAND4xp75_ASAP7_75t_L g8084 ( 
.A(n_7783),
.B(n_7142),
.C(n_7140),
.D(n_6621),
.Y(n_8084)
);

NOR3xp33_ASAP7_75t_L g8085 ( 
.A(n_7472),
.B(n_7142),
.C(n_6623),
.Y(n_8085)
);

OR2x2_ASAP7_75t_L g8086 ( 
.A(n_7745),
.B(n_6334),
.Y(n_8086)
);

AND2x2_ASAP7_75t_L g8087 ( 
.A(n_7647),
.B(n_5718),
.Y(n_8087)
);

AOI22xp33_ASAP7_75t_L g8088 ( 
.A1(n_7757),
.A2(n_7184),
.B1(n_6420),
.B2(n_6928),
.Y(n_8088)
);

INVx1_ASAP7_75t_L g8089 ( 
.A(n_7503),
.Y(n_8089)
);

AND2x2_ASAP7_75t_L g8090 ( 
.A(n_7661),
.B(n_5718),
.Y(n_8090)
);

OAI211xp5_ASAP7_75t_SL g8091 ( 
.A1(n_7727),
.A2(n_5767),
.B(n_5789),
.C(n_5724),
.Y(n_8091)
);

AND2x2_ASAP7_75t_L g8092 ( 
.A(n_7670),
.B(n_5724),
.Y(n_8092)
);

NAND2xp5_ASAP7_75t_L g8093 ( 
.A(n_7527),
.B(n_6297),
.Y(n_8093)
);

AND2x2_ASAP7_75t_L g8094 ( 
.A(n_7671),
.B(n_5724),
.Y(n_8094)
);

AND2x2_ASAP7_75t_L g8095 ( 
.A(n_7683),
.B(n_5767),
.Y(n_8095)
);

AND2x4_ASAP7_75t_L g8096 ( 
.A(n_7496),
.B(n_6393),
.Y(n_8096)
);

AO21x2_ASAP7_75t_L g8097 ( 
.A1(n_7621),
.A2(n_7184),
.B(n_6629),
.Y(n_8097)
);

INVx1_ASAP7_75t_SL g8098 ( 
.A(n_7596),
.Y(n_8098)
);

OR2x2_ASAP7_75t_L g8099 ( 
.A(n_7786),
.B(n_6361),
.Y(n_8099)
);

AOI22xp33_ASAP7_75t_L g8100 ( 
.A1(n_7761),
.A2(n_6420),
.B1(n_6928),
.B2(n_6629),
.Y(n_8100)
);

NAND2xp5_ASAP7_75t_L g8101 ( 
.A(n_7551),
.B(n_7569),
.Y(n_8101)
);

NOR3xp33_ASAP7_75t_L g8102 ( 
.A(n_7482),
.B(n_6632),
.C(n_6617),
.Y(n_8102)
);

NOR2xp33_ASAP7_75t_L g8103 ( 
.A(n_7502),
.B(n_6393),
.Y(n_8103)
);

NAND2xp5_ASAP7_75t_L g8104 ( 
.A(n_7594),
.B(n_6544),
.Y(n_8104)
);

NAND3xp33_ASAP7_75t_L g8105 ( 
.A(n_7598),
.B(n_6663),
.C(n_6643),
.Y(n_8105)
);

NAND3xp33_ASAP7_75t_L g8106 ( 
.A(n_7601),
.B(n_6663),
.C(n_6643),
.Y(n_8106)
);

INVx1_ASAP7_75t_L g8107 ( 
.A(n_7504),
.Y(n_8107)
);

OR2x2_ASAP7_75t_L g8108 ( 
.A(n_7544),
.B(n_6401),
.Y(n_8108)
);

NAND2xp5_ASAP7_75t_L g8109 ( 
.A(n_7732),
.B(n_6548),
.Y(n_8109)
);

AND2x2_ASAP7_75t_L g8110 ( 
.A(n_7694),
.B(n_5767),
.Y(n_8110)
);

OR2x2_ASAP7_75t_L g8111 ( 
.A(n_7556),
.B(n_6298),
.Y(n_8111)
);

AND2x2_ASAP7_75t_L g8112 ( 
.A(n_7496),
.B(n_5789),
.Y(n_8112)
);

AOI221xp5_ASAP7_75t_L g8113 ( 
.A1(n_7788),
.A2(n_6649),
.B1(n_6632),
.B2(n_6449),
.C(n_6489),
.Y(n_8113)
);

AND2x2_ASAP7_75t_L g8114 ( 
.A(n_7819),
.B(n_5789),
.Y(n_8114)
);

NAND2xp5_ASAP7_75t_L g8115 ( 
.A(n_7821),
.B(n_7596),
.Y(n_8115)
);

NOR2x1_ASAP7_75t_R g8116 ( 
.A(n_7658),
.B(n_6535),
.Y(n_8116)
);

AND2x2_ASAP7_75t_L g8117 ( 
.A(n_7548),
.B(n_5791),
.Y(n_8117)
);

OR2x2_ASAP7_75t_L g8118 ( 
.A(n_7557),
.B(n_6301),
.Y(n_8118)
);

OR2x2_ASAP7_75t_L g8119 ( 
.A(n_7760),
.B(n_6333),
.Y(n_8119)
);

OR2x2_ASAP7_75t_L g8120 ( 
.A(n_7782),
.B(n_6339),
.Y(n_8120)
);

AOI22xp33_ASAP7_75t_L g8121 ( 
.A1(n_7761),
.A2(n_7771),
.B1(n_7768),
.B2(n_7685),
.Y(n_8121)
);

INVx1_ASAP7_75t_L g8122 ( 
.A(n_7512),
.Y(n_8122)
);

HB1xp67_ASAP7_75t_L g8123 ( 
.A(n_7773),
.Y(n_8123)
);

INVx2_ASAP7_75t_L g8124 ( 
.A(n_7484),
.Y(n_8124)
);

AOI22xp5_ASAP7_75t_L g8125 ( 
.A1(n_7561),
.A2(n_6649),
.B1(n_5252),
.B2(n_5070),
.Y(n_8125)
);

NAND2xp5_ASAP7_75t_L g8126 ( 
.A(n_7790),
.B(n_6533),
.Y(n_8126)
);

AND2x2_ASAP7_75t_L g8127 ( 
.A(n_7677),
.B(n_5791),
.Y(n_8127)
);

AO21x2_ASAP7_75t_L g8128 ( 
.A1(n_7494),
.A2(n_6185),
.B(n_6184),
.Y(n_8128)
);

BUFx2_ASAP7_75t_L g8129 ( 
.A(n_7469),
.Y(n_8129)
);

NAND4xp75_ASAP7_75t_L g8130 ( 
.A(n_7784),
.B(n_6536),
.C(n_6211),
.D(n_6395),
.Y(n_8130)
);

OR2x2_ASAP7_75t_L g8131 ( 
.A(n_7711),
.B(n_6341),
.Y(n_8131)
);

OR2x2_ASAP7_75t_SL g8132 ( 
.A(n_7798),
.B(n_5964),
.Y(n_8132)
);

AND2x2_ASAP7_75t_L g8133 ( 
.A(n_7728),
.B(n_5791),
.Y(n_8133)
);

OAI22xp5_ASAP7_75t_L g8134 ( 
.A1(n_7810),
.A2(n_6408),
.B1(n_6518),
.B2(n_5810),
.Y(n_8134)
);

NAND3xp33_ASAP7_75t_L g8135 ( 
.A(n_7806),
.B(n_6110),
.C(n_6106),
.Y(n_8135)
);

INVx2_ASAP7_75t_L g8136 ( 
.A(n_7573),
.Y(n_8136)
);

BUFx3_ASAP7_75t_L g8137 ( 
.A(n_7497),
.Y(n_8137)
);

AOI22xp33_ASAP7_75t_L g8138 ( 
.A1(n_7768),
.A2(n_6420),
.B1(n_6185),
.B2(n_6186),
.Y(n_8138)
);

OR2x2_ASAP7_75t_L g8139 ( 
.A(n_7541),
.B(n_6352),
.Y(n_8139)
);

NAND4xp75_ASAP7_75t_L g8140 ( 
.A(n_7789),
.B(n_6536),
.C(n_6211),
.D(n_6395),
.Y(n_8140)
);

XOR2x2_ASAP7_75t_L g8141 ( 
.A(n_7741),
.B(n_5347),
.Y(n_8141)
);

AND2x2_ASAP7_75t_L g8142 ( 
.A(n_7645),
.B(n_5808),
.Y(n_8142)
);

NOR3xp33_ASAP7_75t_L g8143 ( 
.A(n_7708),
.B(n_6110),
.C(n_6106),
.Y(n_8143)
);

INVx2_ASAP7_75t_SL g8144 ( 
.A(n_7810),
.Y(n_8144)
);

INVx4_ASAP7_75t_L g8145 ( 
.A(n_7658),
.Y(n_8145)
);

NAND3xp33_ASAP7_75t_L g8146 ( 
.A(n_7515),
.B(n_6102),
.C(n_6195),
.Y(n_8146)
);

AND2x2_ASAP7_75t_L g8147 ( 
.A(n_7847),
.B(n_7849),
.Y(n_8147)
);

AND2x2_ASAP7_75t_L g8148 ( 
.A(n_7921),
.B(n_7802),
.Y(n_8148)
);

INVx2_ASAP7_75t_L g8149 ( 
.A(n_8082),
.Y(n_8149)
);

AND2x2_ASAP7_75t_L g8150 ( 
.A(n_7924),
.B(n_7655),
.Y(n_8150)
);

INVx2_ASAP7_75t_L g8151 ( 
.A(n_8082),
.Y(n_8151)
);

AO21x2_ASAP7_75t_L g8152 ( 
.A1(n_7892),
.A2(n_7577),
.B(n_7518),
.Y(n_8152)
);

INVx2_ASAP7_75t_L g8153 ( 
.A(n_7993),
.Y(n_8153)
);

INVx2_ASAP7_75t_L g8154 ( 
.A(n_7993),
.Y(n_8154)
);

INVx1_ASAP7_75t_SL g8155 ( 
.A(n_7823),
.Y(n_8155)
);

OAI22xp5_ASAP7_75t_SL g8156 ( 
.A1(n_7833),
.A2(n_7662),
.B1(n_7690),
.B2(n_7560),
.Y(n_8156)
);

INVx3_ASAP7_75t_L g8157 ( 
.A(n_7859),
.Y(n_8157)
);

AOI21xp33_ASAP7_75t_SL g8158 ( 
.A1(n_7892),
.A2(n_7538),
.B(n_7536),
.Y(n_8158)
);

INVx2_ASAP7_75t_L g8159 ( 
.A(n_7858),
.Y(n_8159)
);

INVx1_ASAP7_75t_L g8160 ( 
.A(n_7841),
.Y(n_8160)
);

NAND2xp5_ASAP7_75t_SL g8161 ( 
.A(n_7859),
.B(n_6535),
.Y(n_8161)
);

OAI31xp33_ASAP7_75t_L g8162 ( 
.A1(n_7973),
.A2(n_7804),
.A3(n_7716),
.B(n_7681),
.Y(n_8162)
);

BUFx3_ASAP7_75t_L g8163 ( 
.A(n_7916),
.Y(n_8163)
);

INVx1_ASAP7_75t_SL g8164 ( 
.A(n_8059),
.Y(n_8164)
);

NAND2xp5_ASAP7_75t_L g8165 ( 
.A(n_8081),
.B(n_7817),
.Y(n_8165)
);

AND2x2_ASAP7_75t_L g8166 ( 
.A(n_7879),
.B(n_7603),
.Y(n_8166)
);

AND2x2_ASAP7_75t_L g8167 ( 
.A(n_7889),
.B(n_7611),
.Y(n_8167)
);

BUFx2_ASAP7_75t_L g8168 ( 
.A(n_7926),
.Y(n_8168)
);

OR2x6_ASAP7_75t_L g8169 ( 
.A(n_7964),
.B(n_7709),
.Y(n_8169)
);

INVx1_ASAP7_75t_L g8170 ( 
.A(n_7841),
.Y(n_8170)
);

INVx1_ASAP7_75t_L g8171 ( 
.A(n_7880),
.Y(n_8171)
);

OAI31xp33_ASAP7_75t_L g8172 ( 
.A1(n_7895),
.A2(n_7695),
.A3(n_7696),
.B(n_7676),
.Y(n_8172)
);

INVx1_ASAP7_75t_L g8173 ( 
.A(n_7880),
.Y(n_8173)
);

INVx1_ASAP7_75t_L g8174 ( 
.A(n_8021),
.Y(n_8174)
);

AND2x4_ASAP7_75t_L g8175 ( 
.A(n_7986),
.B(n_7658),
.Y(n_8175)
);

INVx2_ASAP7_75t_L g8176 ( 
.A(n_7826),
.Y(n_8176)
);

OA21x2_ASAP7_75t_L g8177 ( 
.A1(n_7828),
.A2(n_7793),
.B(n_7702),
.Y(n_8177)
);

OR2x2_ASAP7_75t_L g8178 ( 
.A(n_7870),
.B(n_8023),
.Y(n_8178)
);

OAI31xp33_ASAP7_75t_L g8179 ( 
.A1(n_7871),
.A2(n_7700),
.A3(n_7699),
.B(n_7771),
.Y(n_8179)
);

INVxp67_ASAP7_75t_L g8180 ( 
.A(n_8033),
.Y(n_8180)
);

AND2x2_ASAP7_75t_L g8181 ( 
.A(n_7869),
.B(n_7514),
.Y(n_8181)
);

NAND2xp5_ASAP7_75t_L g8182 ( 
.A(n_7934),
.B(n_7579),
.Y(n_8182)
);

AND2x2_ASAP7_75t_L g8183 ( 
.A(n_7886),
.B(n_7514),
.Y(n_8183)
);

NAND2xp5_ASAP7_75t_L g8184 ( 
.A(n_7967),
.B(n_7580),
.Y(n_8184)
);

HB1xp67_ASAP7_75t_L g8185 ( 
.A(n_8021),
.Y(n_8185)
);

BUFx2_ASAP7_75t_L g8186 ( 
.A(n_7929),
.Y(n_8186)
);

BUFx2_ASAP7_75t_L g8187 ( 
.A(n_7856),
.Y(n_8187)
);

INVx1_ASAP7_75t_L g8188 ( 
.A(n_8039),
.Y(n_8188)
);

INVx1_ASAP7_75t_L g8189 ( 
.A(n_8039),
.Y(n_8189)
);

NAND2xp5_ASAP7_75t_L g8190 ( 
.A(n_7978),
.B(n_7587),
.Y(n_8190)
);

INVxp67_ASAP7_75t_L g8191 ( 
.A(n_8016),
.Y(n_8191)
);

AND2x2_ASAP7_75t_L g8192 ( 
.A(n_7959),
.B(n_7610),
.Y(n_8192)
);

AND2x4_ASAP7_75t_L g8193 ( 
.A(n_8028),
.B(n_7597),
.Y(n_8193)
);

AND2x4_ASAP7_75t_SL g8194 ( 
.A(n_7839),
.B(n_7652),
.Y(n_8194)
);

OAI22xp33_ASAP7_75t_L g8195 ( 
.A1(n_7900),
.A2(n_7643),
.B1(n_6408),
.B2(n_7698),
.Y(n_8195)
);

OR2x2_ASAP7_75t_L g8196 ( 
.A(n_7912),
.B(n_7724),
.Y(n_8196)
);

INVx2_ASAP7_75t_L g8197 ( 
.A(n_7915),
.Y(n_8197)
);

AND2x2_ASAP7_75t_L g8198 ( 
.A(n_7935),
.B(n_7588),
.Y(n_8198)
);

INVx2_ASAP7_75t_L g8199 ( 
.A(n_8030),
.Y(n_8199)
);

AND2x2_ASAP7_75t_L g8200 ( 
.A(n_7927),
.B(n_7652),
.Y(n_8200)
);

OR2x2_ASAP7_75t_L g8201 ( 
.A(n_7899),
.B(n_7746),
.Y(n_8201)
);

INVx1_ASAP7_75t_L g8202 ( 
.A(n_8097),
.Y(n_8202)
);

INVx1_ASAP7_75t_L g8203 ( 
.A(n_8097),
.Y(n_8203)
);

AND2x4_ASAP7_75t_L g8204 ( 
.A(n_7918),
.B(n_7567),
.Y(n_8204)
);

AND2x2_ASAP7_75t_L g8205 ( 
.A(n_7894),
.B(n_7457),
.Y(n_8205)
);

OAI221xp5_ASAP7_75t_L g8206 ( 
.A1(n_7863),
.A2(n_7643),
.B1(n_7586),
.B2(n_7565),
.C(n_7674),
.Y(n_8206)
);

INVx1_ASAP7_75t_L g8207 ( 
.A(n_8054),
.Y(n_8207)
);

INVx1_ASAP7_75t_L g8208 ( 
.A(n_8061),
.Y(n_8208)
);

OR2x2_ASAP7_75t_L g8209 ( 
.A(n_7990),
.B(n_7703),
.Y(n_8209)
);

INVx2_ASAP7_75t_L g8210 ( 
.A(n_7855),
.Y(n_8210)
);

INVxp67_ASAP7_75t_L g8211 ( 
.A(n_8024),
.Y(n_8211)
);

INVx1_ASAP7_75t_L g8212 ( 
.A(n_8123),
.Y(n_8212)
);

NAND2xp5_ASAP7_75t_L g8213 ( 
.A(n_7968),
.B(n_7714),
.Y(n_8213)
);

NAND3xp33_ASAP7_75t_SL g8214 ( 
.A(n_7863),
.B(n_7719),
.C(n_7714),
.Y(n_8214)
);

INVxp67_ASAP7_75t_L g8215 ( 
.A(n_7836),
.Y(n_8215)
);

NAND2xp5_ASAP7_75t_L g8216 ( 
.A(n_7971),
.B(n_7719),
.Y(n_8216)
);

OAI211xp5_ASAP7_75t_L g8217 ( 
.A1(n_7833),
.A2(n_7593),
.B(n_7774),
.C(n_7772),
.Y(n_8217)
);

INVx1_ASAP7_75t_L g8218 ( 
.A(n_8049),
.Y(n_8218)
);

HB1xp67_ASAP7_75t_L g8219 ( 
.A(n_8013),
.Y(n_8219)
);

AND2x2_ASAP7_75t_L g8220 ( 
.A(n_7997),
.B(n_7589),
.Y(n_8220)
);

AND2x2_ASAP7_75t_L g8221 ( 
.A(n_7944),
.B(n_7742),
.Y(n_8221)
);

AOI33xp33_ASAP7_75t_L g8222 ( 
.A1(n_7911),
.A2(n_7795),
.A3(n_7774),
.B1(n_7799),
.B2(n_7778),
.B3(n_7772),
.Y(n_8222)
);

INVx2_ASAP7_75t_L g8223 ( 
.A(n_7946),
.Y(n_8223)
);

NAND2xp5_ASAP7_75t_SL g8224 ( 
.A(n_7942),
.B(n_6535),
.Y(n_8224)
);

NAND2xp5_ASAP7_75t_L g8225 ( 
.A(n_8098),
.B(n_7744),
.Y(n_8225)
);

AND2x2_ASAP7_75t_L g8226 ( 
.A(n_7896),
.B(n_7742),
.Y(n_8226)
);

INVx1_ASAP7_75t_SL g8227 ( 
.A(n_7979),
.Y(n_8227)
);

AND2x2_ASAP7_75t_L g8228 ( 
.A(n_7887),
.B(n_7743),
.Y(n_8228)
);

INVx1_ASAP7_75t_L g8229 ( 
.A(n_8079),
.Y(n_8229)
);

AND2x2_ASAP7_75t_L g8230 ( 
.A(n_7888),
.B(n_7743),
.Y(n_8230)
);

INVx2_ASAP7_75t_L g8231 ( 
.A(n_8137),
.Y(n_8231)
);

AOI211xp5_ASAP7_75t_L g8232 ( 
.A1(n_7834),
.A2(n_7860),
.B(n_7865),
.C(n_7866),
.Y(n_8232)
);

INVx4_ASAP7_75t_L g8233 ( 
.A(n_8145),
.Y(n_8233)
);

NAND3xp33_ASAP7_75t_L g8234 ( 
.A(n_7837),
.B(n_7795),
.C(n_7778),
.Y(n_8234)
);

AND2x2_ASAP7_75t_L g8235 ( 
.A(n_8002),
.B(n_7984),
.Y(n_8235)
);

INVxp67_ASAP7_75t_SL g8236 ( 
.A(n_7867),
.Y(n_8236)
);

INVx2_ASAP7_75t_L g8237 ( 
.A(n_7938),
.Y(n_8237)
);

INVx1_ASAP7_75t_L g8238 ( 
.A(n_7822),
.Y(n_8238)
);

INVx1_ASAP7_75t_SL g8239 ( 
.A(n_8056),
.Y(n_8239)
);

BUFx2_ASAP7_75t_L g8240 ( 
.A(n_7940),
.Y(n_8240)
);

AND2x2_ASAP7_75t_L g8241 ( 
.A(n_8003),
.B(n_7744),
.Y(n_8241)
);

AND2x2_ASAP7_75t_L g8242 ( 
.A(n_8027),
.B(n_7749),
.Y(n_8242)
);

NAND2xp5_ASAP7_75t_L g8243 ( 
.A(n_8050),
.B(n_7751),
.Y(n_8243)
);

NAND2xp5_ASAP7_75t_L g8244 ( 
.A(n_7825),
.B(n_7751),
.Y(n_8244)
);

NAND2xp5_ASAP7_75t_L g8245 ( 
.A(n_7846),
.B(n_7749),
.Y(n_8245)
);

HB1xp67_ASAP7_75t_L g8246 ( 
.A(n_8057),
.Y(n_8246)
);

INVx1_ASAP7_75t_L g8247 ( 
.A(n_7843),
.Y(n_8247)
);

INVx1_ASAP7_75t_SL g8248 ( 
.A(n_7897),
.Y(n_8248)
);

INVx1_ASAP7_75t_L g8249 ( 
.A(n_7932),
.Y(n_8249)
);

INVx1_ASAP7_75t_L g8250 ( 
.A(n_7930),
.Y(n_8250)
);

AND2x2_ASAP7_75t_L g8251 ( 
.A(n_8032),
.B(n_7750),
.Y(n_8251)
);

NAND3xp33_ASAP7_75t_L g8252 ( 
.A(n_7911),
.B(n_7801),
.C(n_7799),
.Y(n_8252)
);

NAND5xp2_ASAP7_75t_L g8253 ( 
.A(n_7844),
.B(n_7750),
.C(n_7801),
.D(n_7818),
.E(n_7808),
.Y(n_8253)
);

NAND2xp5_ASAP7_75t_L g8254 ( 
.A(n_7848),
.B(n_7818),
.Y(n_8254)
);

OAI221xp5_ASAP7_75t_L g8255 ( 
.A1(n_8029),
.A2(n_7586),
.B1(n_7565),
.B2(n_7674),
.C(n_6408),
.Y(n_8255)
);

INVx2_ASAP7_75t_L g8256 ( 
.A(n_7914),
.Y(n_8256)
);

INVx1_ASAP7_75t_L g8257 ( 
.A(n_7913),
.Y(n_8257)
);

INVx1_ASAP7_75t_L g8258 ( 
.A(n_7913),
.Y(n_8258)
);

INVx3_ASAP7_75t_L g8259 ( 
.A(n_8048),
.Y(n_8259)
);

AND2x4_ASAP7_75t_L g8260 ( 
.A(n_8067),
.B(n_7623),
.Y(n_8260)
);

OAI33xp33_ASAP7_75t_L g8261 ( 
.A1(n_7827),
.A2(n_7974),
.A3(n_7854),
.B1(n_8007),
.B2(n_7851),
.B3(n_7909),
.Y(n_8261)
);

INVx4_ASAP7_75t_SL g8262 ( 
.A(n_8000),
.Y(n_8262)
);

AOI211xp5_ASAP7_75t_L g8263 ( 
.A1(n_7830),
.A2(n_7651),
.B(n_5975),
.C(n_6121),
.Y(n_8263)
);

INVx2_ASAP7_75t_L g8264 ( 
.A(n_8043),
.Y(n_8264)
);

HB1xp67_ASAP7_75t_L g8265 ( 
.A(n_7857),
.Y(n_8265)
);

NOR3xp33_ASAP7_75t_L g8266 ( 
.A(n_7995),
.B(n_7687),
.C(n_7656),
.Y(n_8266)
);

BUFx2_ASAP7_75t_L g8267 ( 
.A(n_8048),
.Y(n_8267)
);

AND2x2_ASAP7_75t_L g8268 ( 
.A(n_8006),
.B(n_5810),
.Y(n_8268)
);

OAI321xp33_ASAP7_75t_L g8269 ( 
.A1(n_7900),
.A2(n_6189),
.A3(n_6186),
.B1(n_6184),
.B2(n_6246),
.C(n_6224),
.Y(n_8269)
);

NAND2xp5_ASAP7_75t_L g8270 ( 
.A(n_7850),
.B(n_7688),
.Y(n_8270)
);

INVx1_ASAP7_75t_L g8271 ( 
.A(n_7882),
.Y(n_8271)
);

OR2x2_ASAP7_75t_L g8272 ( 
.A(n_7947),
.B(n_6552),
.Y(n_8272)
);

AND2x2_ASAP7_75t_L g8273 ( 
.A(n_8136),
.B(n_8018),
.Y(n_8273)
);

INVx2_ASAP7_75t_L g8274 ( 
.A(n_8129),
.Y(n_8274)
);

NAND4xp25_ASAP7_75t_SL g8275 ( 
.A(n_7906),
.B(n_6113),
.C(n_6128),
.D(n_6121),
.Y(n_8275)
);

INVx2_ASAP7_75t_L g8276 ( 
.A(n_8047),
.Y(n_8276)
);

AOI22xp33_ASAP7_75t_L g8277 ( 
.A1(n_7852),
.A2(n_7739),
.B1(n_7785),
.B2(n_7754),
.Y(n_8277)
);

AND2x2_ASAP7_75t_L g8278 ( 
.A(n_8117),
.B(n_5810),
.Y(n_8278)
);

OAI221xp5_ASAP7_75t_L g8279 ( 
.A1(n_8113),
.A2(n_7739),
.B1(n_7785),
.B2(n_7754),
.C(n_7765),
.Y(n_8279)
);

AOI221xp5_ASAP7_75t_L g8280 ( 
.A1(n_8004),
.A2(n_6189),
.B1(n_6432),
.B2(n_6446),
.C(n_6449),
.Y(n_8280)
);

INVx2_ASAP7_75t_L g8281 ( 
.A(n_8069),
.Y(n_8281)
);

NAND2x1_ASAP7_75t_SL g8282 ( 
.A(n_8069),
.B(n_5808),
.Y(n_8282)
);

AND2x4_ASAP7_75t_L g8283 ( 
.A(n_7907),
.B(n_5808),
.Y(n_8283)
);

INVx1_ASAP7_75t_SL g8284 ( 
.A(n_7922),
.Y(n_8284)
);

NAND2xp5_ASAP7_75t_L g8285 ( 
.A(n_7904),
.B(n_6314),
.Y(n_8285)
);

OR2x2_ASAP7_75t_L g8286 ( 
.A(n_7931),
.B(n_6526),
.Y(n_8286)
);

AND2x2_ASAP7_75t_L g8287 ( 
.A(n_7989),
.B(n_5913),
.Y(n_8287)
);

AND2x2_ASAP7_75t_L g8288 ( 
.A(n_7991),
.B(n_5913),
.Y(n_8288)
);

INVx3_ASAP7_75t_L g8289 ( 
.A(n_8096),
.Y(n_8289)
);

OAI31xp33_ASAP7_75t_L g8290 ( 
.A1(n_8146),
.A2(n_6198),
.A3(n_6207),
.B(n_6194),
.Y(n_8290)
);

NAND2xp5_ASAP7_75t_L g8291 ( 
.A(n_7919),
.B(n_6322),
.Y(n_8291)
);

AOI21xp33_ASAP7_75t_L g8292 ( 
.A1(n_8124),
.A2(n_7765),
.B(n_7797),
.Y(n_8292)
);

INVx2_ASAP7_75t_L g8293 ( 
.A(n_7878),
.Y(n_8293)
);

INVx5_ASAP7_75t_L g8294 ( 
.A(n_8145),
.Y(n_8294)
);

OAI33xp33_ASAP7_75t_L g8295 ( 
.A1(n_8007),
.A2(n_6357),
.A3(n_6344),
.B1(n_6377),
.B2(n_6353),
.B3(n_6326),
.Y(n_8295)
);

AND2x2_ASAP7_75t_L g8296 ( 
.A(n_8045),
.B(n_5913),
.Y(n_8296)
);

AOI22xp33_ASAP7_75t_L g8297 ( 
.A1(n_7908),
.A2(n_7797),
.B1(n_6375),
.B2(n_6370),
.Y(n_8297)
);

BUFx3_ASAP7_75t_L g8298 ( 
.A(n_8035),
.Y(n_8298)
);

INVx1_ASAP7_75t_L g8299 ( 
.A(n_8011),
.Y(n_8299)
);

INVx1_ASAP7_75t_L g8300 ( 
.A(n_7873),
.Y(n_8300)
);

OAI21x1_ASAP7_75t_L g8301 ( 
.A1(n_7960),
.A2(n_6409),
.B(n_6406),
.Y(n_8301)
);

AND2x2_ASAP7_75t_L g8302 ( 
.A(n_7831),
.B(n_8010),
.Y(n_8302)
);

INVx1_ASAP7_75t_L g8303 ( 
.A(n_7864),
.Y(n_8303)
);

INVx1_ASAP7_75t_L g8304 ( 
.A(n_7872),
.Y(n_8304)
);

INVx2_ASAP7_75t_L g8305 ( 
.A(n_8084),
.Y(n_8305)
);

AND2x2_ASAP7_75t_L g8306 ( 
.A(n_7941),
.B(n_5818),
.Y(n_8306)
);

INVx2_ASAP7_75t_L g8307 ( 
.A(n_7853),
.Y(n_8307)
);

INVx1_ASAP7_75t_L g8308 ( 
.A(n_7933),
.Y(n_8308)
);

AND2x2_ASAP7_75t_L g8309 ( 
.A(n_7963),
.B(n_5818),
.Y(n_8309)
);

AND2x2_ASAP7_75t_L g8310 ( 
.A(n_7981),
.B(n_7936),
.Y(n_8310)
);

AND2x2_ASAP7_75t_L g8311 ( 
.A(n_8133),
.B(n_8062),
.Y(n_8311)
);

INVxp67_ASAP7_75t_L g8312 ( 
.A(n_7838),
.Y(n_8312)
);

OAI21xp5_ASAP7_75t_L g8313 ( 
.A1(n_7845),
.A2(n_6128),
.B(n_6113),
.Y(n_8313)
);

INVx3_ASAP7_75t_L g8314 ( 
.A(n_8096),
.Y(n_8314)
);

INVx2_ASAP7_75t_L g8315 ( 
.A(n_7874),
.Y(n_8315)
);

OAI221xp5_ASAP7_75t_L g8316 ( 
.A1(n_8121),
.A2(n_8019),
.B1(n_8001),
.B2(n_7987),
.C(n_8088),
.Y(n_8316)
);

INVx1_ASAP7_75t_L g8317 ( 
.A(n_7937),
.Y(n_8317)
);

INVx5_ASAP7_75t_L g8318 ( 
.A(n_7890),
.Y(n_8318)
);

NAND2xp5_ASAP7_75t_SL g8319 ( 
.A(n_7842),
.B(n_6535),
.Y(n_8319)
);

INVx2_ASAP7_75t_L g8320 ( 
.A(n_7948),
.Y(n_8320)
);

AND2x2_ASAP7_75t_L g8321 ( 
.A(n_8075),
.B(n_8080),
.Y(n_8321)
);

OA211x2_ASAP7_75t_L g8322 ( 
.A1(n_7928),
.A2(n_6535),
.B(n_5151),
.C(n_4550),
.Y(n_8322)
);

OAI21xp5_ASAP7_75t_L g8323 ( 
.A1(n_7961),
.A2(n_6134),
.B(n_6131),
.Y(n_8323)
);

OAI22xp5_ASAP7_75t_L g8324 ( 
.A1(n_7862),
.A2(n_6518),
.B1(n_6246),
.B2(n_6282),
.Y(n_8324)
);

AND2x4_ASAP7_75t_L g8325 ( 
.A(n_7996),
.B(n_5818),
.Y(n_8325)
);

INVx1_ASAP7_75t_L g8326 ( 
.A(n_8004),
.Y(n_8326)
);

AND2x2_ASAP7_75t_L g8327 ( 
.A(n_7832),
.B(n_5971),
.Y(n_8327)
);

INVx1_ASAP7_75t_L g8328 ( 
.A(n_8009),
.Y(n_8328)
);

OAI211xp5_ASAP7_75t_L g8329 ( 
.A1(n_7905),
.A2(n_5084),
.B(n_5136),
.C(n_5126),
.Y(n_8329)
);

INVx2_ASAP7_75t_SL g8330 ( 
.A(n_8112),
.Y(n_8330)
);

INVx1_ASAP7_75t_L g8331 ( 
.A(n_8009),
.Y(n_8331)
);

INVx1_ASAP7_75t_L g8332 ( 
.A(n_8058),
.Y(n_8332)
);

OR2x2_ASAP7_75t_L g8333 ( 
.A(n_7999),
.B(n_6534),
.Y(n_8333)
);

AND2x4_ASAP7_75t_L g8334 ( 
.A(n_7824),
.B(n_5824),
.Y(n_8334)
);

AOI221xp5_ASAP7_75t_L g8335 ( 
.A1(n_8072),
.A2(n_6446),
.B1(n_6432),
.B2(n_6465),
.C(n_6449),
.Y(n_8335)
);

AND2x2_ASAP7_75t_L g8336 ( 
.A(n_8114),
.B(n_5824),
.Y(n_8336)
);

BUFx3_ASAP7_75t_L g8337 ( 
.A(n_7861),
.Y(n_8337)
);

NAND2xp5_ASAP7_75t_L g8338 ( 
.A(n_7835),
.B(n_6410),
.Y(n_8338)
);

INVx1_ASAP7_75t_L g8339 ( 
.A(n_8105),
.Y(n_8339)
);

AND2x4_ASAP7_75t_SL g8340 ( 
.A(n_7840),
.B(n_5975),
.Y(n_8340)
);

OAI31xp33_ASAP7_75t_L g8341 ( 
.A1(n_8146),
.A2(n_6207),
.A3(n_6215),
.B(n_6198),
.Y(n_8341)
);

AOI33xp33_ASAP7_75t_L g8342 ( 
.A1(n_8144),
.A2(n_6141),
.A3(n_6131),
.B1(n_6143),
.B2(n_6139),
.B3(n_6134),
.Y(n_8342)
);

HB1xp67_ASAP7_75t_L g8343 ( 
.A(n_8038),
.Y(n_8343)
);

INVx1_ASAP7_75t_L g8344 ( 
.A(n_8105),
.Y(n_8344)
);

NAND2xp5_ASAP7_75t_L g8345 ( 
.A(n_7962),
.B(n_6411),
.Y(n_8345)
);

OAI221xp5_ASAP7_75t_L g8346 ( 
.A1(n_7875),
.A2(n_6246),
.B1(n_6300),
.B2(n_6282),
.C(n_6224),
.Y(n_8346)
);

INVx1_ASAP7_75t_L g8347 ( 
.A(n_8106),
.Y(n_8347)
);

INVx1_ASAP7_75t_L g8348 ( 
.A(n_8106),
.Y(n_8348)
);

INVx2_ASAP7_75t_L g8349 ( 
.A(n_7975),
.Y(n_8349)
);

INVx1_ASAP7_75t_L g8350 ( 
.A(n_7920),
.Y(n_8350)
);

AND2x2_ASAP7_75t_L g8351 ( 
.A(n_8083),
.B(n_5824),
.Y(n_8351)
);

OAI221xp5_ASAP7_75t_SL g8352 ( 
.A1(n_8108),
.A2(n_6518),
.B1(n_6300),
.B2(n_6246),
.C(n_6282),
.Y(n_8352)
);

AND2x2_ASAP7_75t_L g8353 ( 
.A(n_8087),
.B(n_5921),
.Y(n_8353)
);

INVx3_ASAP7_75t_L g8354 ( 
.A(n_7980),
.Y(n_8354)
);

HB1xp67_ASAP7_75t_L g8355 ( 
.A(n_8115),
.Y(n_8355)
);

INVx1_ASAP7_75t_L g8356 ( 
.A(n_7920),
.Y(n_8356)
);

INVx4_ASAP7_75t_L g8357 ( 
.A(n_7998),
.Y(n_8357)
);

NOR2xp33_ASAP7_75t_L g8358 ( 
.A(n_7868),
.B(n_5964),
.Y(n_8358)
);

OR2x2_ASAP7_75t_L g8359 ( 
.A(n_7982),
.B(n_8008),
.Y(n_8359)
);

INVx1_ASAP7_75t_L g8360 ( 
.A(n_7925),
.Y(n_8360)
);

NOR3xp33_ASAP7_75t_L g8361 ( 
.A(n_7891),
.B(n_6141),
.C(n_6139),
.Y(n_8361)
);

AND2x2_ASAP7_75t_L g8362 ( 
.A(n_8090),
.B(n_5921),
.Y(n_8362)
);

OAI22xp5_ASAP7_75t_L g8363 ( 
.A1(n_7883),
.A2(n_6518),
.B1(n_6282),
.B2(n_6300),
.Y(n_8363)
);

INVx1_ASAP7_75t_L g8364 ( 
.A(n_7925),
.Y(n_8364)
);

INVx1_ASAP7_75t_L g8365 ( 
.A(n_7966),
.Y(n_8365)
);

INVx1_ASAP7_75t_L g8366 ( 
.A(n_7966),
.Y(n_8366)
);

INVx1_ASAP7_75t_L g8367 ( 
.A(n_7969),
.Y(n_8367)
);

NOR3xp33_ASAP7_75t_SL g8368 ( 
.A(n_7977),
.B(n_4820),
.C(n_5332),
.Y(n_8368)
);

INVx2_ASAP7_75t_L g8369 ( 
.A(n_8132),
.Y(n_8369)
);

BUFx2_ASAP7_75t_L g8370 ( 
.A(n_8092),
.Y(n_8370)
);

OAI221xp5_ASAP7_75t_L g8371 ( 
.A1(n_8070),
.A2(n_6355),
.B1(n_6359),
.B2(n_6300),
.C(n_6224),
.Y(n_8371)
);

INVx1_ASAP7_75t_L g8372 ( 
.A(n_8036),
.Y(n_8372)
);

BUFx6f_ASAP7_75t_L g8373 ( 
.A(n_8101),
.Y(n_8373)
);

OR2x2_ASAP7_75t_L g8374 ( 
.A(n_7901),
.B(n_6537),
.Y(n_8374)
);

HB1xp67_ASAP7_75t_L g8375 ( 
.A(n_8076),
.Y(n_8375)
);

OAI221xp5_ASAP7_75t_SL g8376 ( 
.A1(n_8119),
.A2(n_6355),
.B1(n_6359),
.B2(n_6224),
.C(n_6477),
.Y(n_8376)
);

NAND2xp5_ASAP7_75t_L g8377 ( 
.A(n_7957),
.B(n_6463),
.Y(n_8377)
);

NOR3xp33_ASAP7_75t_SL g8378 ( 
.A(n_7898),
.B(n_4820),
.C(n_5332),
.Y(n_8378)
);

NAND2xp5_ASAP7_75t_L g8379 ( 
.A(n_7877),
.B(n_6471),
.Y(n_8379)
);

INVx2_ASAP7_75t_L g8380 ( 
.A(n_8052),
.Y(n_8380)
);

AO21x2_ASAP7_75t_L g8381 ( 
.A1(n_7945),
.A2(n_6383),
.B(n_6378),
.Y(n_8381)
);

OAI21xp5_ASAP7_75t_L g8382 ( 
.A1(n_7885),
.A2(n_6144),
.B(n_6143),
.Y(n_8382)
);

AOI22xp5_ASAP7_75t_L g8383 ( 
.A1(n_8130),
.A2(n_6359),
.B1(n_6355),
.B2(n_6215),
.Y(n_8383)
);

INVx1_ASAP7_75t_L g8384 ( 
.A(n_8055),
.Y(n_8384)
);

AND2x2_ASAP7_75t_L g8385 ( 
.A(n_8094),
.B(n_5921),
.Y(n_8385)
);

AND2x2_ASAP7_75t_L g8386 ( 
.A(n_8095),
.B(n_5971),
.Y(n_8386)
);

INVx2_ASAP7_75t_L g8387 ( 
.A(n_8064),
.Y(n_8387)
);

INVx5_ASAP7_75t_L g8388 ( 
.A(n_8141),
.Y(n_8388)
);

INVx2_ASAP7_75t_L g8389 ( 
.A(n_8086),
.Y(n_8389)
);

INVx1_ASAP7_75t_SL g8390 ( 
.A(n_8110),
.Y(n_8390)
);

NOR3xp33_ASAP7_75t_L g8391 ( 
.A(n_8020),
.B(n_6145),
.C(n_6144),
.Y(n_8391)
);

NAND2x1p5_ASAP7_75t_L g8392 ( 
.A(n_8074),
.B(n_5975),
.Y(n_8392)
);

NAND2xp5_ASAP7_75t_L g8393 ( 
.A(n_8085),
.B(n_6472),
.Y(n_8393)
);

OAI31xp33_ASAP7_75t_L g8394 ( 
.A1(n_8100),
.A2(n_6223),
.A3(n_6225),
.B(n_6220),
.Y(n_8394)
);

AND2x2_ASAP7_75t_L g8395 ( 
.A(n_8142),
.B(n_5971),
.Y(n_8395)
);

OAI221xp5_ASAP7_75t_L g8396 ( 
.A1(n_7970),
.A2(n_6359),
.B1(n_6355),
.B2(n_6477),
.C(n_6329),
.Y(n_8396)
);

AND2x2_ASAP7_75t_L g8397 ( 
.A(n_8127),
.B(n_5991),
.Y(n_8397)
);

NOR2xp33_ASAP7_75t_L g8398 ( 
.A(n_8031),
.B(n_5964),
.Y(n_8398)
);

NAND2xp5_ASAP7_75t_L g8399 ( 
.A(n_8102),
.B(n_6482),
.Y(n_8399)
);

HB1xp67_ASAP7_75t_L g8400 ( 
.A(n_7829),
.Y(n_8400)
);

OR2x2_ASAP7_75t_L g8401 ( 
.A(n_8109),
.B(n_6521),
.Y(n_8401)
);

INVxp67_ASAP7_75t_SL g8402 ( 
.A(n_8116),
.Y(n_8402)
);

OAI31xp33_ASAP7_75t_L g8403 ( 
.A1(n_7903),
.A2(n_8015),
.A3(n_8037),
.B(n_8026),
.Y(n_8403)
);

OR2x2_ASAP7_75t_L g8404 ( 
.A(n_8111),
.B(n_6539),
.Y(n_8404)
);

AND2x2_ASAP7_75t_L g8405 ( 
.A(n_8103),
.B(n_5991),
.Y(n_8405)
);

NAND2xp5_ASAP7_75t_SL g8406 ( 
.A(n_8134),
.B(n_5975),
.Y(n_8406)
);

AND2x4_ASAP7_75t_L g8407 ( 
.A(n_7902),
.B(n_5991),
.Y(n_8407)
);

OR2x2_ASAP7_75t_L g8408 ( 
.A(n_8118),
.B(n_6547),
.Y(n_8408)
);

OAI33xp33_ASAP7_75t_L g8409 ( 
.A1(n_7969),
.A2(n_7985),
.A3(n_7983),
.B1(n_7923),
.B2(n_7951),
.B3(n_8044),
.Y(n_8409)
);

INVx1_ASAP7_75t_SL g8410 ( 
.A(n_8040),
.Y(n_8410)
);

AOI221xp5_ASAP7_75t_L g8411 ( 
.A1(n_7972),
.A2(n_6446),
.B1(n_6432),
.B2(n_6489),
.C(n_6465),
.Y(n_8411)
);

OR2x2_ASAP7_75t_L g8412 ( 
.A(n_8099),
.B(n_6483),
.Y(n_8412)
);

AND2x4_ASAP7_75t_SL g8413 ( 
.A(n_8071),
.B(n_8068),
.Y(n_8413)
);

HB1xp67_ASAP7_75t_L g8414 ( 
.A(n_7876),
.Y(n_8414)
);

INVx3_ASAP7_75t_L g8415 ( 
.A(n_8140),
.Y(n_8415)
);

AND2x2_ASAP7_75t_L g8416 ( 
.A(n_8089),
.B(n_5679),
.Y(n_8416)
);

INVx1_ASAP7_75t_L g8417 ( 
.A(n_7983),
.Y(n_8417)
);

AND2x2_ASAP7_75t_L g8418 ( 
.A(n_8107),
.B(n_5679),
.Y(n_8418)
);

INVxp67_ASAP7_75t_L g8419 ( 
.A(n_8116),
.Y(n_8419)
);

HB1xp67_ASAP7_75t_L g8420 ( 
.A(n_7881),
.Y(n_8420)
);

INVx2_ASAP7_75t_L g8421 ( 
.A(n_8131),
.Y(n_8421)
);

INVx1_ASAP7_75t_L g8422 ( 
.A(n_7910),
.Y(n_8422)
);

INVx1_ASAP7_75t_L g8423 ( 
.A(n_7949),
.Y(n_8423)
);

OR2x2_ASAP7_75t_L g8424 ( 
.A(n_8139),
.B(n_6488),
.Y(n_8424)
);

HB1xp67_ASAP7_75t_L g8425 ( 
.A(n_7952),
.Y(n_8425)
);

AND2x2_ASAP7_75t_L g8426 ( 
.A(n_8122),
.B(n_5683),
.Y(n_8426)
);

AND2x2_ASAP7_75t_L g8427 ( 
.A(n_7953),
.B(n_5683),
.Y(n_8427)
);

INVx2_ASAP7_75t_L g8428 ( 
.A(n_8128),
.Y(n_8428)
);

AND2x2_ASAP7_75t_L g8429 ( 
.A(n_7955),
.B(n_7965),
.Y(n_8429)
);

INVx1_ASAP7_75t_L g8430 ( 
.A(n_8005),
.Y(n_8430)
);

NAND2xp5_ASAP7_75t_L g8431 ( 
.A(n_7950),
.B(n_6494),
.Y(n_8431)
);

HB1xp67_ASAP7_75t_L g8432 ( 
.A(n_8014),
.Y(n_8432)
);

AND2x2_ASAP7_75t_L g8433 ( 
.A(n_8034),
.B(n_5689),
.Y(n_8433)
);

AND2x2_ASAP7_75t_SL g8434 ( 
.A(n_8041),
.B(n_5975),
.Y(n_8434)
);

AND2x2_ASAP7_75t_L g8435 ( 
.A(n_8143),
.B(n_5689),
.Y(n_8435)
);

AOI221xp5_ASAP7_75t_L g8436 ( 
.A1(n_7988),
.A2(n_6489),
.B1(n_6465),
.B2(n_6375),
.C(n_6514),
.Y(n_8436)
);

NAND2xp5_ASAP7_75t_L g8437 ( 
.A(n_7994),
.B(n_6497),
.Y(n_8437)
);

INVx1_ASAP7_75t_L g8438 ( 
.A(n_7985),
.Y(n_8438)
);

NAND2x1p5_ASAP7_75t_L g8439 ( 
.A(n_8022),
.B(n_5081),
.Y(n_8439)
);

INVx4_ASAP7_75t_L g8440 ( 
.A(n_8120),
.Y(n_8440)
);

OR2x2_ASAP7_75t_L g8441 ( 
.A(n_7893),
.B(n_8025),
.Y(n_8441)
);

AOI21xp5_ASAP7_75t_L g8442 ( 
.A1(n_7939),
.A2(n_6505),
.B(n_6499),
.Y(n_8442)
);

INVx2_ASAP7_75t_L g8443 ( 
.A(n_8128),
.Y(n_8443)
);

NOR2xp67_ASAP7_75t_L g8444 ( 
.A(n_8042),
.B(n_5126),
.Y(n_8444)
);

NOR2xp67_ASAP7_75t_L g8445 ( 
.A(n_7958),
.B(n_5126),
.Y(n_8445)
);

AND2x2_ASAP7_75t_L g8446 ( 
.A(n_8126),
.B(n_5715),
.Y(n_8446)
);

INVx1_ASAP7_75t_L g8447 ( 
.A(n_8185),
.Y(n_8447)
);

INVx1_ASAP7_75t_L g8448 ( 
.A(n_8160),
.Y(n_8448)
);

AND2x2_ASAP7_75t_L g8449 ( 
.A(n_8235),
.B(n_8046),
.Y(n_8449)
);

AND2x2_ASAP7_75t_L g8450 ( 
.A(n_8187),
.B(n_8060),
.Y(n_8450)
);

INVx1_ASAP7_75t_L g8451 ( 
.A(n_8160),
.Y(n_8451)
);

INVxp67_ASAP7_75t_L g8452 ( 
.A(n_8186),
.Y(n_8452)
);

INVx1_ASAP7_75t_L g8453 ( 
.A(n_8202),
.Y(n_8453)
);

INVx2_ASAP7_75t_L g8454 ( 
.A(n_8163),
.Y(n_8454)
);

INVx1_ASAP7_75t_L g8455 ( 
.A(n_8202),
.Y(n_8455)
);

NOR2xp33_ASAP7_75t_L g8456 ( 
.A(n_8373),
.B(n_8091),
.Y(n_8456)
);

INVx1_ASAP7_75t_L g8457 ( 
.A(n_8203),
.Y(n_8457)
);

NAND2xp5_ASAP7_75t_L g8458 ( 
.A(n_8164),
.B(n_8053),
.Y(n_8458)
);

NAND2xp5_ASAP7_75t_L g8459 ( 
.A(n_8226),
.B(n_7884),
.Y(n_8459)
);

AND2x2_ASAP7_75t_SL g8460 ( 
.A(n_8178),
.B(n_8065),
.Y(n_8460)
);

OA21x2_ASAP7_75t_L g8461 ( 
.A1(n_8174),
.A2(n_7917),
.B(n_8017),
.Y(n_8461)
);

NAND2x1_ASAP7_75t_L g8462 ( 
.A(n_8157),
.B(n_8135),
.Y(n_8462)
);

INVx2_ASAP7_75t_L g8463 ( 
.A(n_8157),
.Y(n_8463)
);

INVx1_ASAP7_75t_L g8464 ( 
.A(n_8188),
.Y(n_8464)
);

AND2x2_ASAP7_75t_L g8465 ( 
.A(n_8147),
.B(n_8198),
.Y(n_8465)
);

OR2x2_ASAP7_75t_L g8466 ( 
.A(n_8155),
.B(n_7954),
.Y(n_8466)
);

NAND2xp5_ASAP7_75t_L g8467 ( 
.A(n_8373),
.B(n_8066),
.Y(n_8467)
);

INVx1_ASAP7_75t_L g8468 ( 
.A(n_8189),
.Y(n_8468)
);

AND2x2_ASAP7_75t_L g8469 ( 
.A(n_8167),
.B(n_8093),
.Y(n_8469)
);

HB1xp67_ASAP7_75t_L g8470 ( 
.A(n_8152),
.Y(n_8470)
);

OR2x2_ASAP7_75t_L g8471 ( 
.A(n_8196),
.B(n_8104),
.Y(n_8471)
);

INVx1_ASAP7_75t_L g8472 ( 
.A(n_8170),
.Y(n_8472)
);

NAND2xp5_ASAP7_75t_L g8473 ( 
.A(n_8373),
.B(n_8073),
.Y(n_8473)
);

AND2x2_ASAP7_75t_L g8474 ( 
.A(n_8183),
.B(n_8077),
.Y(n_8474)
);

AOI22xp5_ASAP7_75t_L g8475 ( 
.A1(n_8415),
.A2(n_7976),
.B1(n_8051),
.B2(n_8012),
.Y(n_8475)
);

INVx1_ASAP7_75t_L g8476 ( 
.A(n_8171),
.Y(n_8476)
);

OR2x6_ASAP7_75t_L g8477 ( 
.A(n_8169),
.B(n_6477),
.Y(n_8477)
);

INVx1_ASAP7_75t_L g8478 ( 
.A(n_8173),
.Y(n_8478)
);

OAI32xp33_ASAP7_75t_L g8479 ( 
.A1(n_8326),
.A2(n_7992),
.A3(n_7956),
.B1(n_7976),
.B2(n_8063),
.Y(n_8479)
);

INVx1_ASAP7_75t_L g8480 ( 
.A(n_8219),
.Y(n_8480)
);

INVx1_ASAP7_75t_L g8481 ( 
.A(n_8228),
.Y(n_8481)
);

NAND2xp5_ASAP7_75t_L g8482 ( 
.A(n_8248),
.B(n_8012),
.Y(n_8482)
);

AND2x2_ASAP7_75t_L g8483 ( 
.A(n_8166),
.B(n_5715),
.Y(n_8483)
);

AND2x2_ASAP7_75t_L g8484 ( 
.A(n_8221),
.B(n_5726),
.Y(n_8484)
);

AND2x2_ASAP7_75t_SL g8485 ( 
.A(n_8168),
.B(n_7943),
.Y(n_8485)
);

INVx1_ASAP7_75t_L g8486 ( 
.A(n_8230),
.Y(n_8486)
);

INVx3_ASAP7_75t_L g8487 ( 
.A(n_8204),
.Y(n_8487)
);

NOR2x1_ASAP7_75t_L g8488 ( 
.A(n_8350),
.B(n_5081),
.Y(n_8488)
);

AND2x2_ASAP7_75t_L g8489 ( 
.A(n_8159),
.B(n_5726),
.Y(n_8489)
);

INVx1_ASAP7_75t_L g8490 ( 
.A(n_8241),
.Y(n_8490)
);

HB1xp67_ASAP7_75t_L g8491 ( 
.A(n_8262),
.Y(n_8491)
);

INVx1_ASAP7_75t_L g8492 ( 
.A(n_8251),
.Y(n_8492)
);

NAND2xp5_ASAP7_75t_L g8493 ( 
.A(n_8370),
.B(n_8078),
.Y(n_8493)
);

AND2x2_ASAP7_75t_L g8494 ( 
.A(n_8169),
.B(n_5745),
.Y(n_8494)
);

NAND2xp5_ASAP7_75t_L g8495 ( 
.A(n_8242),
.B(n_8138),
.Y(n_8495)
);

OR2x2_ASAP7_75t_L g8496 ( 
.A(n_8284),
.B(n_6500),
.Y(n_8496)
);

INVx1_ASAP7_75t_L g8497 ( 
.A(n_8355),
.Y(n_8497)
);

NOR2xp33_ASAP7_75t_L g8498 ( 
.A(n_8289),
.B(n_5964),
.Y(n_8498)
);

OR2x2_ASAP7_75t_L g8499 ( 
.A(n_8244),
.B(n_6510),
.Y(n_8499)
);

INVx1_ASAP7_75t_L g8500 ( 
.A(n_8203),
.Y(n_8500)
);

OR2x2_ASAP7_75t_L g8501 ( 
.A(n_8326),
.B(n_6512),
.Y(n_8501)
);

INVxp67_ASAP7_75t_L g8502 ( 
.A(n_8240),
.Y(n_8502)
);

NAND2xp5_ASAP7_75t_L g8503 ( 
.A(n_8210),
.B(n_6513),
.Y(n_8503)
);

INVx1_ASAP7_75t_L g8504 ( 
.A(n_8149),
.Y(n_8504)
);

HB1xp67_ASAP7_75t_L g8505 ( 
.A(n_8262),
.Y(n_8505)
);

INVx1_ASAP7_75t_L g8506 ( 
.A(n_8151),
.Y(n_8506)
);

AND2x2_ASAP7_75t_L g8507 ( 
.A(n_8197),
.B(n_8199),
.Y(n_8507)
);

INVx2_ASAP7_75t_L g8508 ( 
.A(n_8282),
.Y(n_8508)
);

INVx3_ASAP7_75t_L g8509 ( 
.A(n_8204),
.Y(n_8509)
);

INVxp67_ASAP7_75t_SL g8510 ( 
.A(n_8328),
.Y(n_8510)
);

INVx1_ASAP7_75t_L g8511 ( 
.A(n_8265),
.Y(n_8511)
);

INVx1_ASAP7_75t_L g8512 ( 
.A(n_8328),
.Y(n_8512)
);

NOR2x1_ASAP7_75t_L g8513 ( 
.A(n_8350),
.B(n_5081),
.Y(n_8513)
);

INVx1_ASAP7_75t_L g8514 ( 
.A(n_8331),
.Y(n_8514)
);

AND2x2_ASAP7_75t_L g8515 ( 
.A(n_8176),
.B(n_5745),
.Y(n_8515)
);

CKINVDCx5p33_ASAP7_75t_R g8516 ( 
.A(n_8194),
.Y(n_8516)
);

INVx1_ASAP7_75t_SL g8517 ( 
.A(n_8227),
.Y(n_8517)
);

HB1xp67_ASAP7_75t_L g8518 ( 
.A(n_8331),
.Y(n_8518)
);

OR2x2_ASAP7_75t_L g8519 ( 
.A(n_8213),
.B(n_8216),
.Y(n_8519)
);

INVx1_ASAP7_75t_L g8520 ( 
.A(n_8359),
.Y(n_8520)
);

INVx1_ASAP7_75t_L g8521 ( 
.A(n_8184),
.Y(n_8521)
);

INVx2_ASAP7_75t_L g8522 ( 
.A(n_8259),
.Y(n_8522)
);

INVx2_ASAP7_75t_SL g8523 ( 
.A(n_8318),
.Y(n_8523)
);

AND2x2_ASAP7_75t_L g8524 ( 
.A(n_8321),
.B(n_5847),
.Y(n_8524)
);

AND2x2_ASAP7_75t_L g8525 ( 
.A(n_8337),
.B(n_5847),
.Y(n_8525)
);

NAND2xp5_ASAP7_75t_L g8526 ( 
.A(n_8390),
.B(n_6515),
.Y(n_8526)
);

INVx1_ASAP7_75t_L g8527 ( 
.A(n_8428),
.Y(n_8527)
);

OAI21xp33_ASAP7_75t_L g8528 ( 
.A1(n_8253),
.A2(n_5122),
.B(n_5120),
.Y(n_8528)
);

INVx1_ASAP7_75t_L g8529 ( 
.A(n_8212),
.Y(n_8529)
);

NOR2xp33_ASAP7_75t_L g8530 ( 
.A(n_8289),
.B(n_6145),
.Y(n_8530)
);

AND2x4_ASAP7_75t_L g8531 ( 
.A(n_8153),
.B(n_6149),
.Y(n_8531)
);

AND2x2_ASAP7_75t_L g8532 ( 
.A(n_8192),
.B(n_8310),
.Y(n_8532)
);

INVx2_ASAP7_75t_L g8533 ( 
.A(n_8259),
.Y(n_8533)
);

INVx2_ASAP7_75t_L g8534 ( 
.A(n_8267),
.Y(n_8534)
);

AND2x2_ASAP7_75t_L g8535 ( 
.A(n_8205),
.B(n_5853),
.Y(n_8535)
);

NAND2x1p5_ASAP7_75t_L g8536 ( 
.A(n_8314),
.B(n_5120),
.Y(n_8536)
);

INVx1_ASAP7_75t_L g8537 ( 
.A(n_8190),
.Y(n_8537)
);

INVx1_ASAP7_75t_L g8538 ( 
.A(n_8182),
.Y(n_8538)
);

INVx2_ASAP7_75t_L g8539 ( 
.A(n_8314),
.Y(n_8539)
);

INVx1_ASAP7_75t_L g8540 ( 
.A(n_8225),
.Y(n_8540)
);

OR2x2_ASAP7_75t_L g8541 ( 
.A(n_8209),
.B(n_6517),
.Y(n_8541)
);

INVx1_ASAP7_75t_L g8542 ( 
.A(n_8400),
.Y(n_8542)
);

NAND2xp5_ASAP7_75t_L g8543 ( 
.A(n_8223),
.B(n_6149),
.Y(n_8543)
);

INVx2_ASAP7_75t_L g8544 ( 
.A(n_8260),
.Y(n_8544)
);

INVx1_ASAP7_75t_SL g8545 ( 
.A(n_8220),
.Y(n_8545)
);

NAND2xp5_ASAP7_75t_L g8546 ( 
.A(n_8298),
.B(n_6163),
.Y(n_8546)
);

NAND2xp5_ASAP7_75t_L g8547 ( 
.A(n_8308),
.B(n_6163),
.Y(n_8547)
);

INVxp67_ASAP7_75t_L g8548 ( 
.A(n_8246),
.Y(n_8548)
);

INVx1_ASAP7_75t_L g8549 ( 
.A(n_8414),
.Y(n_8549)
);

OR2x2_ASAP7_75t_L g8550 ( 
.A(n_8214),
.B(n_6174),
.Y(n_8550)
);

INVx2_ASAP7_75t_L g8551 ( 
.A(n_8260),
.Y(n_8551)
);

INVx2_ASAP7_75t_SL g8552 ( 
.A(n_8318),
.Y(n_8552)
);

INVxp67_ASAP7_75t_L g8553 ( 
.A(n_8148),
.Y(n_8553)
);

INVx1_ASAP7_75t_L g8554 ( 
.A(n_8443),
.Y(n_8554)
);

OR2x2_ASAP7_75t_L g8555 ( 
.A(n_8218),
.B(n_6174),
.Y(n_8555)
);

OR2x6_ASAP7_75t_L g8556 ( 
.A(n_8231),
.B(n_6477),
.Y(n_8556)
);

OR2x6_ASAP7_75t_L g8557 ( 
.A(n_8315),
.B(n_5629),
.Y(n_8557)
);

OR2x2_ASAP7_75t_L g8558 ( 
.A(n_8229),
.B(n_6171),
.Y(n_8558)
);

INVx2_ASAP7_75t_SL g8559 ( 
.A(n_8318),
.Y(n_8559)
);

OAI21xp33_ASAP7_75t_L g8560 ( 
.A1(n_8368),
.A2(n_5122),
.B(n_5120),
.Y(n_8560)
);

INVx1_ASAP7_75t_L g8561 ( 
.A(n_8420),
.Y(n_8561)
);

OR2x2_ASAP7_75t_L g8562 ( 
.A(n_8356),
.B(n_6171),
.Y(n_8562)
);

INVx1_ASAP7_75t_L g8563 ( 
.A(n_8425),
.Y(n_8563)
);

NAND2xp5_ASAP7_75t_L g8564 ( 
.A(n_8354),
.B(n_6172),
.Y(n_8564)
);

OAI21xp5_ASAP7_75t_L g8565 ( 
.A1(n_8356),
.A2(n_8125),
.B(n_6173),
.Y(n_8565)
);

NAND2xp5_ASAP7_75t_L g8566 ( 
.A(n_8354),
.B(n_6172),
.Y(n_8566)
);

INVx1_ASAP7_75t_L g8567 ( 
.A(n_8432),
.Y(n_8567)
);

OR2x2_ASAP7_75t_L g8568 ( 
.A(n_8360),
.B(n_6173),
.Y(n_8568)
);

INVx1_ASAP7_75t_L g8569 ( 
.A(n_8360),
.Y(n_8569)
);

NAND2xp5_ASAP7_75t_L g8570 ( 
.A(n_8421),
.B(n_5575),
.Y(n_8570)
);

INVx1_ASAP7_75t_L g8571 ( 
.A(n_8364),
.Y(n_8571)
);

AND2x2_ASAP7_75t_L g8572 ( 
.A(n_8154),
.B(n_5853),
.Y(n_8572)
);

AND2x2_ASAP7_75t_L g8573 ( 
.A(n_8200),
.B(n_5917),
.Y(n_8573)
);

INVx1_ASAP7_75t_L g8574 ( 
.A(n_8364),
.Y(n_8574)
);

OR2x2_ASAP7_75t_L g8575 ( 
.A(n_8365),
.B(n_5576),
.Y(n_8575)
);

NOR3xp33_ASAP7_75t_L g8576 ( 
.A(n_8365),
.B(n_8125),
.C(n_6278),
.Y(n_8576)
);

INVx1_ASAP7_75t_L g8577 ( 
.A(n_8366),
.Y(n_8577)
);

INVx1_ASAP7_75t_L g8578 ( 
.A(n_8366),
.Y(n_8578)
);

NAND2xp5_ASAP7_75t_L g8579 ( 
.A(n_8299),
.B(n_5576),
.Y(n_8579)
);

NAND2xp5_ASAP7_75t_L g8580 ( 
.A(n_8380),
.B(n_5577),
.Y(n_8580)
);

INVx2_ASAP7_75t_L g8581 ( 
.A(n_8175),
.Y(n_8581)
);

INVx2_ASAP7_75t_SL g8582 ( 
.A(n_8181),
.Y(n_8582)
);

INVx1_ASAP7_75t_L g8583 ( 
.A(n_8367),
.Y(n_8583)
);

INVx1_ASAP7_75t_SL g8584 ( 
.A(n_8302),
.Y(n_8584)
);

AND2x2_ASAP7_75t_L g8585 ( 
.A(n_8311),
.B(n_5857),
.Y(n_8585)
);

INVx1_ASAP7_75t_L g8586 ( 
.A(n_8367),
.Y(n_8586)
);

OR2x2_ASAP7_75t_L g8587 ( 
.A(n_8417),
.B(n_5577),
.Y(n_8587)
);

INVx1_ASAP7_75t_SL g8588 ( 
.A(n_8175),
.Y(n_8588)
);

BUFx3_ASAP7_75t_L g8589 ( 
.A(n_8193),
.Y(n_8589)
);

NOR2xp33_ASAP7_75t_L g8590 ( 
.A(n_8409),
.B(n_8357),
.Y(n_8590)
);

INVx2_ASAP7_75t_L g8591 ( 
.A(n_8294),
.Y(n_8591)
);

INVx1_ASAP7_75t_L g8592 ( 
.A(n_8417),
.Y(n_8592)
);

OR2x2_ASAP7_75t_L g8593 ( 
.A(n_8438),
.B(n_5580),
.Y(n_8593)
);

INVx1_ASAP7_75t_L g8594 ( 
.A(n_8438),
.Y(n_8594)
);

AND2x2_ASAP7_75t_L g8595 ( 
.A(n_8334),
.B(n_5857),
.Y(n_8595)
);

INVxp67_ASAP7_75t_L g8596 ( 
.A(n_8343),
.Y(n_8596)
);

INVx1_ASAP7_75t_L g8597 ( 
.A(n_8339),
.Y(n_8597)
);

INVx2_ASAP7_75t_L g8598 ( 
.A(n_8294),
.Y(n_8598)
);

NOR2xp33_ASAP7_75t_L g8599 ( 
.A(n_8357),
.B(n_5122),
.Y(n_8599)
);

NAND2xp5_ASAP7_75t_SL g8600 ( 
.A(n_8232),
.B(n_5134),
.Y(n_8600)
);

AND2x2_ASAP7_75t_L g8601 ( 
.A(n_8334),
.B(n_5865),
.Y(n_8601)
);

NAND2xp5_ASAP7_75t_L g8602 ( 
.A(n_8372),
.B(n_5580),
.Y(n_8602)
);

INVx1_ASAP7_75t_L g8603 ( 
.A(n_8339),
.Y(n_8603)
);

AOI21xp5_ASAP7_75t_L g8604 ( 
.A1(n_8162),
.A2(n_8347),
.B(n_8344),
.Y(n_8604)
);

NAND2xp5_ASAP7_75t_SL g8605 ( 
.A(n_8388),
.B(n_5134),
.Y(n_8605)
);

INVx1_ASAP7_75t_L g8606 ( 
.A(n_8344),
.Y(n_8606)
);

INVxp33_ASAP7_75t_L g8607 ( 
.A(n_8237),
.Y(n_8607)
);

INVx1_ASAP7_75t_L g8608 ( 
.A(n_8347),
.Y(n_8608)
);

INVx1_ASAP7_75t_L g8609 ( 
.A(n_8348),
.Y(n_8609)
);

OR2x2_ASAP7_75t_L g8610 ( 
.A(n_8243),
.B(n_5581),
.Y(n_8610)
);

INVx1_ASAP7_75t_L g8611 ( 
.A(n_8348),
.Y(n_8611)
);

INVx2_ASAP7_75t_L g8612 ( 
.A(n_8294),
.Y(n_8612)
);

AND2x2_ASAP7_75t_L g8613 ( 
.A(n_8150),
.B(n_5865),
.Y(n_8613)
);

INVx1_ASAP7_75t_L g8614 ( 
.A(n_8165),
.Y(n_8614)
);

AND2x2_ASAP7_75t_L g8615 ( 
.A(n_8193),
.B(n_5917),
.Y(n_8615)
);

NOR2x1p5_ASAP7_75t_SL g8616 ( 
.A(n_8207),
.B(n_6220),
.Y(n_8616)
);

AND2x2_ASAP7_75t_L g8617 ( 
.A(n_8273),
.B(n_5932),
.Y(n_8617)
);

OR2x2_ASAP7_75t_L g8618 ( 
.A(n_8201),
.B(n_5581),
.Y(n_8618)
);

OR2x2_ASAP7_75t_L g8619 ( 
.A(n_8332),
.B(n_5585),
.Y(n_8619)
);

INVx1_ASAP7_75t_L g8620 ( 
.A(n_8429),
.Y(n_8620)
);

NAND2xp5_ASAP7_75t_L g8621 ( 
.A(n_8387),
.B(n_5585),
.Y(n_8621)
);

INVx2_ASAP7_75t_L g8622 ( 
.A(n_8439),
.Y(n_8622)
);

AND2x2_ASAP7_75t_L g8623 ( 
.A(n_8306),
.B(n_5932),
.Y(n_8623)
);

OR2x2_ASAP7_75t_L g8624 ( 
.A(n_8332),
.B(n_5590),
.Y(n_8624)
);

AND2x4_ASAP7_75t_L g8625 ( 
.A(n_8281),
.B(n_5134),
.Y(n_8625)
);

OR2x2_ASAP7_75t_L g8626 ( 
.A(n_8389),
.B(n_5590),
.Y(n_8626)
);

AND2x2_ASAP7_75t_L g8627 ( 
.A(n_8309),
.B(n_5955),
.Y(n_8627)
);

NAND2xp5_ASAP7_75t_L g8628 ( 
.A(n_8158),
.B(n_5595),
.Y(n_8628)
);

AND2x2_ASAP7_75t_L g8629 ( 
.A(n_8287),
.B(n_5955),
.Y(n_8629)
);

INVx2_ASAP7_75t_L g8630 ( 
.A(n_8233),
.Y(n_8630)
);

O2A1O1Ixp33_ASAP7_75t_L g8631 ( 
.A1(n_8206),
.A2(n_6223),
.B(n_6231),
.C(n_6225),
.Y(n_8631)
);

OR2x2_ASAP7_75t_L g8632 ( 
.A(n_8441),
.B(n_5595),
.Y(n_8632)
);

INVx1_ASAP7_75t_L g8633 ( 
.A(n_8286),
.Y(n_8633)
);

HB1xp67_ASAP7_75t_L g8634 ( 
.A(n_8177),
.Y(n_8634)
);

BUFx2_ASAP7_75t_L g8635 ( 
.A(n_8215),
.Y(n_8635)
);

INVx1_ASAP7_75t_L g8636 ( 
.A(n_8180),
.Y(n_8636)
);

INVx1_ASAP7_75t_L g8637 ( 
.A(n_8207),
.Y(n_8637)
);

NAND2xp33_ASAP7_75t_L g8638 ( 
.A(n_8239),
.B(n_4928),
.Y(n_8638)
);

AND2x4_ASAP7_75t_L g8639 ( 
.A(n_8330),
.B(n_5164),
.Y(n_8639)
);

OR2x2_ASAP7_75t_L g8640 ( 
.A(n_8384),
.B(n_5597),
.Y(n_8640)
);

INVx2_ASAP7_75t_L g8641 ( 
.A(n_8233),
.Y(n_8641)
);

INVx1_ASAP7_75t_L g8642 ( 
.A(n_8208),
.Y(n_8642)
);

INVx1_ASAP7_75t_L g8643 ( 
.A(n_8208),
.Y(n_8643)
);

INVx2_ASAP7_75t_SL g8644 ( 
.A(n_8413),
.Y(n_8644)
);

NAND2xp5_ASAP7_75t_L g8645 ( 
.A(n_8427),
.B(n_5597),
.Y(n_8645)
);

INVx1_ASAP7_75t_L g8646 ( 
.A(n_8272),
.Y(n_8646)
);

INVx2_ASAP7_75t_L g8647 ( 
.A(n_8407),
.Y(n_8647)
);

AND2x2_ASAP7_75t_L g8648 ( 
.A(n_8288),
.B(n_5973),
.Y(n_8648)
);

INVx2_ASAP7_75t_L g8649 ( 
.A(n_8407),
.Y(n_8649)
);

AND2x2_ASAP7_75t_L g8650 ( 
.A(n_8433),
.B(n_5973),
.Y(n_8650)
);

INVx1_ASAP7_75t_L g8651 ( 
.A(n_8222),
.Y(n_8651)
);

OR2x2_ASAP7_75t_L g8652 ( 
.A(n_8247),
.B(n_5598),
.Y(n_8652)
);

NAND4xp75_ASAP7_75t_L g8653 ( 
.A(n_8322),
.B(n_6211),
.C(n_6536),
.D(n_6245),
.Y(n_8653)
);

NAND2xp5_ASAP7_75t_L g8654 ( 
.A(n_8403),
.B(n_5598),
.Y(n_8654)
);

INVx2_ASAP7_75t_L g8655 ( 
.A(n_8283),
.Y(n_8655)
);

INVx1_ASAP7_75t_L g8656 ( 
.A(n_8401),
.Y(n_8656)
);

AND2x2_ASAP7_75t_L g8657 ( 
.A(n_8416),
.B(n_5980),
.Y(n_8657)
);

INVxp67_ASAP7_75t_SL g8658 ( 
.A(n_8177),
.Y(n_8658)
);

INVx1_ASAP7_75t_L g8659 ( 
.A(n_8245),
.Y(n_8659)
);

INVx1_ASAP7_75t_L g8660 ( 
.A(n_8254),
.Y(n_8660)
);

NAND2xp5_ASAP7_75t_L g8661 ( 
.A(n_8317),
.B(n_8418),
.Y(n_8661)
);

INVx2_ASAP7_75t_SL g8662 ( 
.A(n_8283),
.Y(n_8662)
);

INVx2_ASAP7_75t_L g8663 ( 
.A(n_8268),
.Y(n_8663)
);

HB1xp67_ASAP7_75t_L g8664 ( 
.A(n_8375),
.Y(n_8664)
);

OAI222xp33_ASAP7_75t_L g8665 ( 
.A1(n_8410),
.A2(n_5242),
.B1(n_5629),
.B2(n_6238),
.C1(n_6234),
.C2(n_6231),
.Y(n_8665)
);

INVx2_ASAP7_75t_L g8666 ( 
.A(n_8381),
.Y(n_8666)
);

AND2x2_ASAP7_75t_L g8667 ( 
.A(n_8426),
.B(n_5980),
.Y(n_8667)
);

INVx3_ASAP7_75t_L g8668 ( 
.A(n_8325),
.Y(n_8668)
);

INVx1_ASAP7_75t_L g8669 ( 
.A(n_8424),
.Y(n_8669)
);

INVxp67_ASAP7_75t_L g8670 ( 
.A(n_8236),
.Y(n_8670)
);

AND2x2_ASAP7_75t_L g8671 ( 
.A(n_8327),
.B(n_6000),
.Y(n_8671)
);

AND2x2_ASAP7_75t_L g8672 ( 
.A(n_8388),
.B(n_6000),
.Y(n_8672)
);

OR2x2_ASAP7_75t_L g8673 ( 
.A(n_8271),
.B(n_5599),
.Y(n_8673)
);

INVx2_ASAP7_75t_L g8674 ( 
.A(n_8296),
.Y(n_8674)
);

AND2x2_ASAP7_75t_L g8675 ( 
.A(n_8388),
.B(n_5747),
.Y(n_8675)
);

INVx1_ASAP7_75t_L g8676 ( 
.A(n_8404),
.Y(n_8676)
);

AND2x2_ASAP7_75t_L g8677 ( 
.A(n_8446),
.B(n_8276),
.Y(n_8677)
);

INVx1_ASAP7_75t_L g8678 ( 
.A(n_8408),
.Y(n_8678)
);

NAND2xp5_ASAP7_75t_L g8679 ( 
.A(n_8256),
.B(n_5599),
.Y(n_8679)
);

AND2x2_ASAP7_75t_L g8680 ( 
.A(n_8405),
.B(n_5747),
.Y(n_8680)
);

NAND2x1p5_ASAP7_75t_L g8681 ( 
.A(n_8238),
.B(n_5164),
.Y(n_8681)
);

NAND2xp5_ASAP7_75t_L g8682 ( 
.A(n_8264),
.B(n_5605),
.Y(n_8682)
);

NAND2xp5_ASAP7_75t_L g8683 ( 
.A(n_8274),
.B(n_5605),
.Y(n_8683)
);

AND2x4_ASAP7_75t_L g8684 ( 
.A(n_8320),
.B(n_5164),
.Y(n_8684)
);

INVx2_ASAP7_75t_L g8685 ( 
.A(n_8434),
.Y(n_8685)
);

INVx2_ASAP7_75t_L g8686 ( 
.A(n_8301),
.Y(n_8686)
);

OAI211xp5_ASAP7_75t_SL g8687 ( 
.A1(n_8415),
.A2(n_5214),
.B(n_5300),
.C(n_5159),
.Y(n_8687)
);

AND2x4_ASAP7_75t_L g8688 ( 
.A(n_8349),
.B(n_8369),
.Y(n_8688)
);

OR2x6_ASAP7_75t_L g8689 ( 
.A(n_8191),
.B(n_5203),
.Y(n_8689)
);

INVx1_ASAP7_75t_L g8690 ( 
.A(n_8270),
.Y(n_8690)
);

NAND2xp5_ASAP7_75t_L g8691 ( 
.A(n_8300),
.B(n_5606),
.Y(n_8691)
);

AO22x1_ASAP7_75t_L g8692 ( 
.A1(n_8266),
.A2(n_5203),
.B1(n_5256),
.B2(n_5217),
.Y(n_8692)
);

OR2x2_ASAP7_75t_L g8693 ( 
.A(n_8303),
.B(n_5606),
.Y(n_8693)
);

INVx1_ASAP7_75t_L g8694 ( 
.A(n_8234),
.Y(n_8694)
);

OR2x2_ASAP7_75t_L g8695 ( 
.A(n_8304),
.B(n_5611),
.Y(n_8695)
);

INVx2_ASAP7_75t_L g8696 ( 
.A(n_8336),
.Y(n_8696)
);

OAI21xp5_ASAP7_75t_L g8697 ( 
.A1(n_8252),
.A2(n_6383),
.B(n_6378),
.Y(n_8697)
);

A2O1A1Ixp33_ASAP7_75t_L g8698 ( 
.A1(n_8255),
.A2(n_6492),
.B(n_6507),
.C(n_6484),
.Y(n_8698)
);

O2A1O1Ixp33_ASAP7_75t_L g8699 ( 
.A1(n_8261),
.A2(n_6234),
.B(n_6243),
.C(n_6238),
.Y(n_8699)
);

INVx1_ASAP7_75t_L g8700 ( 
.A(n_8257),
.Y(n_8700)
);

AND2x2_ASAP7_75t_L g8701 ( 
.A(n_8293),
.B(n_5785),
.Y(n_8701)
);

INVxp67_ASAP7_75t_L g8702 ( 
.A(n_8358),
.Y(n_8702)
);

AND2x2_ASAP7_75t_L g8703 ( 
.A(n_8532),
.B(n_8465),
.Y(n_8703)
);

INVx1_ASAP7_75t_L g8704 ( 
.A(n_8470),
.Y(n_8704)
);

INVx1_ASAP7_75t_L g8705 ( 
.A(n_8634),
.Y(n_8705)
);

INVx2_ASAP7_75t_L g8706 ( 
.A(n_8487),
.Y(n_8706)
);

OR2x2_ASAP7_75t_L g8707 ( 
.A(n_8584),
.B(n_8249),
.Y(n_8707)
);

NAND2xp5_ASAP7_75t_L g8708 ( 
.A(n_8460),
.B(n_8305),
.Y(n_8708)
);

INVx2_ASAP7_75t_L g8709 ( 
.A(n_8487),
.Y(n_8709)
);

INVx2_ASAP7_75t_SL g8710 ( 
.A(n_8589),
.Y(n_8710)
);

INVx1_ASAP7_75t_L g8711 ( 
.A(n_8658),
.Y(n_8711)
);

OAI21xp5_ASAP7_75t_L g8712 ( 
.A1(n_8604),
.A2(n_8217),
.B(n_8316),
.Y(n_8712)
);

INVx1_ASAP7_75t_SL g8713 ( 
.A(n_8635),
.Y(n_8713)
);

INVxp67_ASAP7_75t_L g8714 ( 
.A(n_8491),
.Y(n_8714)
);

AND2x2_ASAP7_75t_L g8715 ( 
.A(n_8672),
.B(n_8340),
.Y(n_8715)
);

INVx1_ASAP7_75t_L g8716 ( 
.A(n_8482),
.Y(n_8716)
);

NAND2xp5_ASAP7_75t_L g8717 ( 
.A(n_8469),
.B(n_8250),
.Y(n_8717)
);

NOR2xp33_ASAP7_75t_SL g8718 ( 
.A(n_8516),
.B(n_8440),
.Y(n_8718)
);

NAND3xp33_ASAP7_75t_L g8719 ( 
.A(n_8518),
.B(n_8172),
.C(n_8179),
.Y(n_8719)
);

AOI322xp5_ASAP7_75t_L g8720 ( 
.A1(n_8510),
.A2(n_8258),
.A3(n_8277),
.B1(n_8297),
.B2(n_8292),
.C1(n_8307),
.C2(n_8335),
.Y(n_8720)
);

INVx1_ASAP7_75t_L g8721 ( 
.A(n_8616),
.Y(n_8721)
);

INVx1_ASAP7_75t_L g8722 ( 
.A(n_8463),
.Y(n_8722)
);

INVx1_ASAP7_75t_L g8723 ( 
.A(n_8539),
.Y(n_8723)
);

INVx1_ASAP7_75t_L g8724 ( 
.A(n_8450),
.Y(n_8724)
);

NAND2xp5_ASAP7_75t_L g8725 ( 
.A(n_8449),
.B(n_8312),
.Y(n_8725)
);

INVx1_ASAP7_75t_L g8726 ( 
.A(n_8507),
.Y(n_8726)
);

INVx1_ASAP7_75t_L g8727 ( 
.A(n_8466),
.Y(n_8727)
);

AOI22xp5_ASAP7_75t_L g8728 ( 
.A1(n_8461),
.A2(n_8596),
.B1(n_8666),
.B2(n_8279),
.Y(n_8728)
);

OR2x2_ASAP7_75t_L g8729 ( 
.A(n_8517),
.B(n_8440),
.Y(n_8729)
);

AND2x2_ASAP7_75t_L g8730 ( 
.A(n_8675),
.B(n_8395),
.Y(n_8730)
);

INVx1_ASAP7_75t_L g8731 ( 
.A(n_8534),
.Y(n_8731)
);

INVx2_ASAP7_75t_L g8732 ( 
.A(n_8509),
.Y(n_8732)
);

INVx1_ASAP7_75t_L g8733 ( 
.A(n_8544),
.Y(n_8733)
);

AND2x2_ASAP7_75t_L g8734 ( 
.A(n_8525),
.B(n_8351),
.Y(n_8734)
);

NAND2xp5_ASAP7_75t_L g8735 ( 
.A(n_8505),
.B(n_8342),
.Y(n_8735)
);

NOR2xp33_ASAP7_75t_L g8736 ( 
.A(n_8553),
.B(n_8352),
.Y(n_8736)
);

INVx1_ASAP7_75t_L g8737 ( 
.A(n_8551),
.Y(n_8737)
);

AOI32xp33_ASAP7_75t_L g8738 ( 
.A1(n_8694),
.A2(n_8377),
.A3(n_8431),
.B1(n_8430),
.B2(n_8423),
.Y(n_8738)
);

INVx1_ASAP7_75t_L g8739 ( 
.A(n_8664),
.Y(n_8739)
);

INVx1_ASAP7_75t_L g8740 ( 
.A(n_8471),
.Y(n_8740)
);

INVx1_ASAP7_75t_L g8741 ( 
.A(n_8509),
.Y(n_8741)
);

NOR3xp33_ASAP7_75t_L g8742 ( 
.A(n_8473),
.B(n_8694),
.C(n_8590),
.Y(n_8742)
);

AOI222xp33_ASAP7_75t_L g8743 ( 
.A1(n_8700),
.A2(n_8156),
.B1(n_8436),
.B2(n_8280),
.C1(n_8411),
.C2(n_8269),
.Y(n_8743)
);

AND2x4_ASAP7_75t_L g8744 ( 
.A(n_8582),
.B(n_8211),
.Y(n_8744)
);

OAI21xp5_ASAP7_75t_L g8745 ( 
.A1(n_8485),
.A2(n_8323),
.B(n_8378),
.Y(n_8745)
);

AND2x2_ASAP7_75t_L g8746 ( 
.A(n_8545),
.B(n_8353),
.Y(n_8746)
);

AOI221xp5_ASAP7_75t_L g8747 ( 
.A1(n_8631),
.A2(n_8479),
.B1(n_8606),
.B2(n_8603),
.C(n_8597),
.Y(n_8747)
);

INVx1_ASAP7_75t_L g8748 ( 
.A(n_8522),
.Y(n_8748)
);

INVx1_ASAP7_75t_L g8749 ( 
.A(n_8533),
.Y(n_8749)
);

AO22x1_ASAP7_75t_L g8750 ( 
.A1(n_8569),
.A2(n_8402),
.B1(n_8422),
.B2(n_8325),
.Y(n_8750)
);

NAND2xp5_ASAP7_75t_L g8751 ( 
.A(n_8523),
.B(n_8442),
.Y(n_8751)
);

INVx1_ASAP7_75t_L g8752 ( 
.A(n_8481),
.Y(n_8752)
);

NAND2xp5_ASAP7_75t_L g8753 ( 
.A(n_8552),
.B(n_8412),
.Y(n_8753)
);

HB1xp67_ASAP7_75t_L g8754 ( 
.A(n_8559),
.Y(n_8754)
);

OAI32xp33_ASAP7_75t_L g8755 ( 
.A1(n_8651),
.A2(n_8577),
.A3(n_8578),
.B1(n_8574),
.B2(n_8571),
.Y(n_8755)
);

OAI32xp33_ASAP7_75t_L g8756 ( 
.A1(n_8583),
.A2(n_8437),
.A3(n_8393),
.B1(n_8399),
.B2(n_8391),
.Y(n_8756)
);

INVx1_ASAP7_75t_L g8757 ( 
.A(n_8486),
.Y(n_8757)
);

INVx1_ASAP7_75t_L g8758 ( 
.A(n_8458),
.Y(n_8758)
);

NAND2xp5_ASAP7_75t_L g8759 ( 
.A(n_8490),
.B(n_8445),
.Y(n_8759)
);

INVx1_ASAP7_75t_L g8760 ( 
.A(n_8492),
.Y(n_8760)
);

AOI21xp5_ASAP7_75t_SL g8761 ( 
.A1(n_8467),
.A2(n_8419),
.B(n_8224),
.Y(n_8761)
);

NAND2xp5_ASAP7_75t_L g8762 ( 
.A(n_8688),
.B(n_8374),
.Y(n_8762)
);

INVx1_ASAP7_75t_L g8763 ( 
.A(n_8519),
.Y(n_8763)
);

NAND3xp33_ASAP7_75t_L g8764 ( 
.A(n_8461),
.B(n_8263),
.C(n_8290),
.Y(n_8764)
);

NAND2xp5_ASAP7_75t_L g8765 ( 
.A(n_8688),
.B(n_8285),
.Y(n_8765)
);

INVx1_ASAP7_75t_L g8766 ( 
.A(n_8520),
.Y(n_8766)
);

NAND2xp5_ASAP7_75t_L g8767 ( 
.A(n_8588),
.B(n_8291),
.Y(n_8767)
);

INVx1_ASAP7_75t_L g8768 ( 
.A(n_8493),
.Y(n_8768)
);

INVx1_ASAP7_75t_L g8769 ( 
.A(n_8452),
.Y(n_8769)
);

NOR2x1_ASAP7_75t_L g8770 ( 
.A(n_8608),
.B(n_8275),
.Y(n_8770)
);

NAND2xp5_ASAP7_75t_L g8771 ( 
.A(n_8677),
.B(n_8345),
.Y(n_8771)
);

HB1xp67_ASAP7_75t_L g8772 ( 
.A(n_8462),
.Y(n_8772)
);

INVx3_ASAP7_75t_SL g8773 ( 
.A(n_8644),
.Y(n_8773)
);

AND2x2_ASAP7_75t_L g8774 ( 
.A(n_8483),
.B(n_8362),
.Y(n_8774)
);

XOR2x2_ASAP7_75t_L g8775 ( 
.A(n_8459),
.B(n_8376),
.Y(n_8775)
);

INVx1_ASAP7_75t_L g8776 ( 
.A(n_8454),
.Y(n_8776)
);

INVx1_ASAP7_75t_L g8777 ( 
.A(n_8480),
.Y(n_8777)
);

INVx1_ASAP7_75t_L g8778 ( 
.A(n_8620),
.Y(n_8778)
);

AOI222xp33_ASAP7_75t_L g8779 ( 
.A1(n_8700),
.A2(n_8295),
.B1(n_8313),
.B2(n_8382),
.C1(n_8379),
.C2(n_8195),
.Y(n_8779)
);

NAND2xp67_ASAP7_75t_L g8780 ( 
.A(n_8647),
.B(n_8338),
.Y(n_8780)
);

NAND4xp25_ASAP7_75t_L g8781 ( 
.A(n_8456),
.B(n_8398),
.C(n_8444),
.D(n_8329),
.Y(n_8781)
);

OAI22xp5_ASAP7_75t_L g8782 ( 
.A1(n_8475),
.A2(n_8435),
.B1(n_8406),
.B2(n_8333),
.Y(n_8782)
);

AND2x2_ASAP7_75t_L g8783 ( 
.A(n_8494),
.B(n_8385),
.Y(n_8783)
);

INVxp67_ASAP7_75t_L g8784 ( 
.A(n_8599),
.Y(n_8784)
);

INVx2_ASAP7_75t_L g8785 ( 
.A(n_8536),
.Y(n_8785)
);

NOR2x1_ASAP7_75t_L g8786 ( 
.A(n_8609),
.B(n_8161),
.Y(n_8786)
);

INVx2_ASAP7_75t_L g8787 ( 
.A(n_8477),
.Y(n_8787)
);

NAND2xp5_ASAP7_75t_L g8788 ( 
.A(n_8524),
.B(n_8361),
.Y(n_8788)
);

AOI22xp5_ASAP7_75t_L g8789 ( 
.A1(n_8576),
.A2(n_8383),
.B1(n_8363),
.B2(n_8324),
.Y(n_8789)
);

NOR3xp33_ASAP7_75t_L g8790 ( 
.A(n_8479),
.B(n_8670),
.C(n_8537),
.Y(n_8790)
);

HB1xp67_ASAP7_75t_L g8791 ( 
.A(n_8488),
.Y(n_8791)
);

NAND2xp5_ASAP7_75t_SL g8792 ( 
.A(n_8508),
.B(n_8341),
.Y(n_8792)
);

OR2x2_ASAP7_75t_L g8793 ( 
.A(n_8497),
.B(n_8386),
.Y(n_8793)
);

INVx2_ASAP7_75t_L g8794 ( 
.A(n_8477),
.Y(n_8794)
);

O2A1O1Ixp33_ASAP7_75t_L g8795 ( 
.A1(n_8611),
.A2(n_8319),
.B(n_8394),
.C(n_8346),
.Y(n_8795)
);

NAND2xp5_ASAP7_75t_L g8796 ( 
.A(n_8617),
.B(n_8278),
.Y(n_8796)
);

INVx1_ASAP7_75t_L g8797 ( 
.A(n_8661),
.Y(n_8797)
);

OAI21xp33_ASAP7_75t_SL g8798 ( 
.A1(n_8512),
.A2(n_8397),
.B(n_6469),
.Y(n_8798)
);

NAND2xp5_ASAP7_75t_L g8799 ( 
.A(n_8585),
.B(n_8392),
.Y(n_8799)
);

NOR2xp33_ASAP7_75t_L g8800 ( 
.A(n_8528),
.B(n_8371),
.Y(n_8800)
);

AND2x2_ASAP7_75t_L g8801 ( 
.A(n_8484),
.B(n_5785),
.Y(n_8801)
);

NAND2xp5_ASAP7_75t_L g8802 ( 
.A(n_8656),
.B(n_8396),
.Y(n_8802)
);

AOI22xp5_ASAP7_75t_L g8803 ( 
.A1(n_8607),
.A2(n_6243),
.B1(n_6253),
.B2(n_6250),
.Y(n_8803)
);

AOI22xp33_ASAP7_75t_L g8804 ( 
.A1(n_8514),
.A2(n_6375),
.B1(n_6370),
.B2(n_6358),
.Y(n_8804)
);

INVx1_ASAP7_75t_L g8805 ( 
.A(n_8541),
.Y(n_8805)
);

INVx1_ASAP7_75t_L g8806 ( 
.A(n_8511),
.Y(n_8806)
);

NAND2xp5_ASAP7_75t_L g8807 ( 
.A(n_8668),
.B(n_5611),
.Y(n_8807)
);

INVx1_ASAP7_75t_L g8808 ( 
.A(n_8562),
.Y(n_8808)
);

INVx1_ASAP7_75t_SL g8809 ( 
.A(n_8684),
.Y(n_8809)
);

INVx1_ASAP7_75t_L g8810 ( 
.A(n_8568),
.Y(n_8810)
);

HB1xp67_ASAP7_75t_L g8811 ( 
.A(n_8513),
.Y(n_8811)
);

CKINVDCx20_ASAP7_75t_R g8812 ( 
.A(n_8495),
.Y(n_8812)
);

INVx1_ASAP7_75t_L g8813 ( 
.A(n_8618),
.Y(n_8813)
);

INVx2_ASAP7_75t_SL g8814 ( 
.A(n_8684),
.Y(n_8814)
);

INVx1_ASAP7_75t_L g8815 ( 
.A(n_8633),
.Y(n_8815)
);

INVx1_ASAP7_75t_L g8816 ( 
.A(n_8646),
.Y(n_8816)
);

OAI22xp5_ASAP7_75t_L g8817 ( 
.A1(n_8586),
.A2(n_5203),
.B1(n_5256),
.B2(n_5217),
.Y(n_8817)
);

INVx1_ASAP7_75t_L g8818 ( 
.A(n_8496),
.Y(n_8818)
);

AND2x2_ASAP7_75t_L g8819 ( 
.A(n_8573),
.B(n_8615),
.Y(n_8819)
);

OA222x2_ASAP7_75t_L g8820 ( 
.A1(n_8592),
.A2(n_8594),
.B1(n_8550),
.B2(n_8628),
.C1(n_8502),
.C2(n_8548),
.Y(n_8820)
);

OAI22xp33_ASAP7_75t_L g8821 ( 
.A1(n_8697),
.A2(n_6253),
.B1(n_6268),
.B2(n_6250),
.Y(n_8821)
);

AND2x4_ASAP7_75t_L g8822 ( 
.A(n_8581),
.B(n_5217),
.Y(n_8822)
);

OR2x2_ASAP7_75t_L g8823 ( 
.A(n_8546),
.B(n_5246),
.Y(n_8823)
);

OAI21xp33_ASAP7_75t_L g8824 ( 
.A1(n_8560),
.A2(n_8498),
.B(n_8474),
.Y(n_8824)
);

NAND2x1p5_ASAP7_75t_L g8825 ( 
.A(n_8605),
.B(n_5256),
.Y(n_8825)
);

INVx2_ASAP7_75t_SL g8826 ( 
.A(n_8625),
.Y(n_8826)
);

OAI32xp33_ASAP7_75t_L g8827 ( 
.A1(n_8542),
.A2(n_5753),
.A3(n_5836),
.B1(n_5588),
.B2(n_5136),
.Y(n_8827)
);

OAI21xp5_ASAP7_75t_L g8828 ( 
.A1(n_8600),
.A2(n_6469),
.B(n_6439),
.Y(n_8828)
);

NAND2x1p5_ASAP7_75t_L g8829 ( 
.A(n_8636),
.B(n_4836),
.Y(n_8829)
);

INVx1_ASAP7_75t_L g8830 ( 
.A(n_8549),
.Y(n_8830)
);

NAND2xp5_ASAP7_75t_L g8831 ( 
.A(n_8668),
.B(n_5612),
.Y(n_8831)
);

INVx2_ASAP7_75t_L g8832 ( 
.A(n_8535),
.Y(n_8832)
);

AOI21xp33_ASAP7_75t_L g8833 ( 
.A1(n_8699),
.A2(n_6270),
.B(n_6268),
.Y(n_8833)
);

AOI22xp5_ASAP7_75t_L g8834 ( 
.A1(n_8637),
.A2(n_8642),
.B1(n_8643),
.B2(n_8690),
.Y(n_8834)
);

INVx2_ASAP7_75t_L g8835 ( 
.A(n_8657),
.Y(n_8835)
);

INVx1_ASAP7_75t_L g8836 ( 
.A(n_8561),
.Y(n_8836)
);

AND2x2_ASAP7_75t_L g8837 ( 
.A(n_8572),
.B(n_5803),
.Y(n_8837)
);

OAI221xp5_ASAP7_75t_L g8838 ( 
.A1(n_8565),
.A2(n_8698),
.B1(n_8447),
.B2(n_8686),
.C(n_8685),
.Y(n_8838)
);

INVx1_ASAP7_75t_L g8839 ( 
.A(n_8563),
.Y(n_8839)
);

AND2x2_ASAP7_75t_L g8840 ( 
.A(n_8515),
.B(n_5803),
.Y(n_8840)
);

INVxp67_ASAP7_75t_L g8841 ( 
.A(n_8530),
.Y(n_8841)
);

INVx2_ASAP7_75t_L g8842 ( 
.A(n_8667),
.Y(n_8842)
);

BUFx2_ASAP7_75t_L g8843 ( 
.A(n_8689),
.Y(n_8843)
);

INVx1_ASAP7_75t_L g8844 ( 
.A(n_8567),
.Y(n_8844)
);

NAND3xp33_ASAP7_75t_L g8845 ( 
.A(n_8649),
.B(n_8540),
.C(n_8638),
.Y(n_8845)
);

OR2x2_ASAP7_75t_L g8846 ( 
.A(n_8669),
.B(n_5358),
.Y(n_8846)
);

NAND2xp5_ASAP7_75t_L g8847 ( 
.A(n_8531),
.B(n_5612),
.Y(n_8847)
);

INVx1_ASAP7_75t_L g8848 ( 
.A(n_8676),
.Y(n_8848)
);

HB1xp67_ASAP7_75t_L g8849 ( 
.A(n_8689),
.Y(n_8849)
);

INVx1_ASAP7_75t_L g8850 ( 
.A(n_8678),
.Y(n_8850)
);

INVx3_ASAP7_75t_L g8851 ( 
.A(n_8625),
.Y(n_8851)
);

A2O1A1Ixp33_ASAP7_75t_L g8852 ( 
.A1(n_8504),
.A2(n_8506),
.B(n_8451),
.C(n_8448),
.Y(n_8852)
);

INVx1_ASAP7_75t_L g8853 ( 
.A(n_8499),
.Y(n_8853)
);

NOR4xp25_ASAP7_75t_SL g8854 ( 
.A(n_8659),
.B(n_5246),
.C(n_5358),
.D(n_5127),
.Y(n_8854)
);

OAI21xp33_ASAP7_75t_L g8855 ( 
.A1(n_8701),
.A2(n_6439),
.B(n_4846),
.Y(n_8855)
);

INVx1_ASAP7_75t_SL g8856 ( 
.A(n_8639),
.Y(n_8856)
);

NOR3xp33_ASAP7_75t_L g8857 ( 
.A(n_8692),
.B(n_6278),
.C(n_6270),
.Y(n_8857)
);

AND2x2_ASAP7_75t_L g8858 ( 
.A(n_8613),
.B(n_8489),
.Y(n_8858)
);

HB1xp67_ASAP7_75t_L g8859 ( 
.A(n_8639),
.Y(n_8859)
);

INVxp67_ASAP7_75t_L g8860 ( 
.A(n_8674),
.Y(n_8860)
);

AND2x2_ASAP7_75t_L g8861 ( 
.A(n_8663),
.B(n_5813),
.Y(n_8861)
);

INVx1_ASAP7_75t_L g8862 ( 
.A(n_8564),
.Y(n_8862)
);

NOR2xp67_ASAP7_75t_SL g8863 ( 
.A(n_8529),
.B(n_5106),
.Y(n_8863)
);

OAI22xp33_ASAP7_75t_L g8864 ( 
.A1(n_8501),
.A2(n_6280),
.B1(n_6286),
.B2(n_6284),
.Y(n_8864)
);

OR2x2_ASAP7_75t_L g8865 ( 
.A(n_8521),
.B(n_5127),
.Y(n_8865)
);

INVx1_ASAP7_75t_L g8866 ( 
.A(n_8566),
.Y(n_8866)
);

NAND2xp33_ASAP7_75t_SL g8867 ( 
.A(n_8662),
.B(n_5813),
.Y(n_8867)
);

INVx2_ASAP7_75t_L g8868 ( 
.A(n_8650),
.Y(n_8868)
);

OR2x2_ASAP7_75t_L g8869 ( 
.A(n_8538),
.B(n_5613),
.Y(n_8869)
);

NAND2xp5_ASAP7_75t_L g8870 ( 
.A(n_8531),
.B(n_5613),
.Y(n_8870)
);

AOI21xp33_ASAP7_75t_L g8871 ( 
.A1(n_8575),
.A2(n_6284),
.B(n_6280),
.Y(n_8871)
);

INVx1_ASAP7_75t_L g8872 ( 
.A(n_8632),
.Y(n_8872)
);

OAI22xp5_ASAP7_75t_L g8873 ( 
.A1(n_8622),
.A2(n_5615),
.B1(n_5630),
.B2(n_5623),
.Y(n_8873)
);

OAI21xp33_ASAP7_75t_L g8874 ( 
.A1(n_8671),
.A2(n_4846),
.B(n_4826),
.Y(n_8874)
);

INVx1_ASAP7_75t_L g8875 ( 
.A(n_8660),
.Y(n_8875)
);

NAND2x1_ASAP7_75t_L g8876 ( 
.A(n_8655),
.B(n_8696),
.Y(n_8876)
);

NAND2xp5_ASAP7_75t_SL g8877 ( 
.A(n_8630),
.B(n_5838),
.Y(n_8877)
);

NOR2xp33_ASAP7_75t_L g8878 ( 
.A(n_8681),
.B(n_3886),
.Y(n_8878)
);

AND2x4_ASAP7_75t_L g8879 ( 
.A(n_8641),
.B(n_4826),
.Y(n_8879)
);

INVx1_ASAP7_75t_L g8880 ( 
.A(n_8610),
.Y(n_8880)
);

AOI32xp33_ASAP7_75t_L g8881 ( 
.A1(n_8614),
.A2(n_5192),
.A3(n_6292),
.B1(n_6289),
.B2(n_6286),
.Y(n_8881)
);

AND2x2_ASAP7_75t_L g8882 ( 
.A(n_8595),
.B(n_4922),
.Y(n_8882)
);

INVx1_ASAP7_75t_SL g8883 ( 
.A(n_8555),
.Y(n_8883)
);

AOI22xp5_ASAP7_75t_L g8884 ( 
.A1(n_8527),
.A2(n_6289),
.B1(n_6303),
.B2(n_6292),
.Y(n_8884)
);

INVx1_ASAP7_75t_L g8885 ( 
.A(n_8558),
.Y(n_8885)
);

NOR3xp33_ASAP7_75t_L g8886 ( 
.A(n_8692),
.B(n_6308),
.C(n_6303),
.Y(n_8886)
);

AND2x2_ASAP7_75t_L g8887 ( 
.A(n_8601),
.B(n_4922),
.Y(n_8887)
);

NAND4xp75_ASAP7_75t_SL g8888 ( 
.A(n_8680),
.B(n_6195),
.C(n_4736),
.D(n_4689),
.Y(n_8888)
);

NAND2xp5_ASAP7_75t_SL g8889 ( 
.A(n_8591),
.B(n_5838),
.Y(n_8889)
);

NAND2xp5_ASAP7_75t_L g8890 ( 
.A(n_8598),
.B(n_5615),
.Y(n_8890)
);

NOR2x1_ASAP7_75t_L g8891 ( 
.A(n_8448),
.B(n_5139),
.Y(n_8891)
);

INVx1_ASAP7_75t_L g8892 ( 
.A(n_8626),
.Y(n_8892)
);

AND2x2_ASAP7_75t_L g8893 ( 
.A(n_8623),
.B(n_5133),
.Y(n_8893)
);

INVx1_ASAP7_75t_L g8894 ( 
.A(n_8587),
.Y(n_8894)
);

AND2x2_ASAP7_75t_L g8895 ( 
.A(n_8627),
.B(n_5133),
.Y(n_8895)
);

INVx1_ASAP7_75t_L g8896 ( 
.A(n_8593),
.Y(n_8896)
);

INVx2_ASAP7_75t_L g8897 ( 
.A(n_8557),
.Y(n_8897)
);

NAND3xp33_ASAP7_75t_SL g8898 ( 
.A(n_8702),
.B(n_5272),
.C(n_5588),
.Y(n_8898)
);

INVx2_ASAP7_75t_L g8899 ( 
.A(n_8557),
.Y(n_8899)
);

AND2x2_ASAP7_75t_L g8900 ( 
.A(n_8629),
.B(n_5143),
.Y(n_8900)
);

AOI32xp33_ASAP7_75t_L g8901 ( 
.A1(n_8654),
.A2(n_6312),
.A3(n_6329),
.B1(n_6315),
.B2(n_6308),
.Y(n_8901)
);

NOR2xp67_ASAP7_75t_L g8902 ( 
.A(n_8612),
.B(n_4836),
.Y(n_8902)
);

NAND2xp5_ASAP7_75t_L g8903 ( 
.A(n_8526),
.B(n_8645),
.Y(n_8903)
);

NOR2x1_ASAP7_75t_L g8904 ( 
.A(n_8451),
.B(n_5139),
.Y(n_8904)
);

INVx3_ASAP7_75t_L g8905 ( 
.A(n_8640),
.Y(n_8905)
);

AOI21xp5_ASAP7_75t_L g8906 ( 
.A1(n_8547),
.A2(n_6195),
.B(n_6102),
.Y(n_8906)
);

INVx1_ASAP7_75t_L g8907 ( 
.A(n_8652),
.Y(n_8907)
);

INVx2_ASAP7_75t_L g8908 ( 
.A(n_8648),
.Y(n_8908)
);

INVx1_ASAP7_75t_L g8909 ( 
.A(n_8619),
.Y(n_8909)
);

INVx2_ASAP7_75t_L g8910 ( 
.A(n_8556),
.Y(n_8910)
);

INVx2_ASAP7_75t_L g8911 ( 
.A(n_8556),
.Y(n_8911)
);

INVx1_ASAP7_75t_L g8912 ( 
.A(n_8624),
.Y(n_8912)
);

INVx1_ASAP7_75t_L g8913 ( 
.A(n_8543),
.Y(n_8913)
);

AOI22xp5_ASAP7_75t_L g8914 ( 
.A1(n_8527),
.A2(n_6312),
.B1(n_6350),
.B2(n_6315),
.Y(n_8914)
);

OAI22xp33_ASAP7_75t_L g8915 ( 
.A1(n_8453),
.A2(n_6350),
.B1(n_6362),
.B2(n_6360),
.Y(n_8915)
);

NAND2xp5_ASAP7_75t_L g8916 ( 
.A(n_8570),
.B(n_5623),
.Y(n_8916)
);

NAND4xp25_ASAP7_75t_L g8917 ( 
.A(n_8503),
.B(n_4836),
.C(n_4889),
.D(n_4849),
.Y(n_8917)
);

INVx2_ASAP7_75t_L g8918 ( 
.A(n_8653),
.Y(n_8918)
);

O2A1O1Ixp33_ASAP7_75t_L g8919 ( 
.A1(n_8500),
.A2(n_6102),
.B(n_6362),
.C(n_6360),
.Y(n_8919)
);

INVx1_ASAP7_75t_L g8920 ( 
.A(n_8693),
.Y(n_8920)
);

OAI32xp33_ASAP7_75t_L g8921 ( 
.A1(n_8580),
.A2(n_5836),
.A3(n_5753),
.B1(n_5588),
.B2(n_5351),
.Y(n_8921)
);

AOI211xp5_ASAP7_75t_L g8922 ( 
.A1(n_8687),
.A2(n_4920),
.B(n_5176),
.C(n_4913),
.Y(n_8922)
);

INVxp67_ASAP7_75t_L g8923 ( 
.A(n_8673),
.Y(n_8923)
);

NAND3xp33_ASAP7_75t_L g8924 ( 
.A(n_8554),
.B(n_6384),
.C(n_6374),
.Y(n_8924)
);

OAI22xp33_ASAP7_75t_L g8925 ( 
.A1(n_8453),
.A2(n_8457),
.B1(n_8455),
.B2(n_8554),
.Y(n_8925)
);

OAI221xp5_ASAP7_75t_L g8926 ( 
.A1(n_8455),
.A2(n_6520),
.B1(n_6522),
.B2(n_6514),
.C(n_6507),
.Y(n_8926)
);

HB1xp67_ASAP7_75t_L g8927 ( 
.A(n_8695),
.Y(n_8927)
);

OAI221xp5_ASAP7_75t_SL g8928 ( 
.A1(n_8679),
.A2(n_5272),
.B1(n_5104),
.B2(n_5250),
.C(n_6399),
.Y(n_8928)
);

INVx1_ASAP7_75t_L g8929 ( 
.A(n_8621),
.Y(n_8929)
);

AND2x2_ASAP7_75t_L g8930 ( 
.A(n_8682),
.B(n_5143),
.Y(n_8930)
);

INVx1_ASAP7_75t_L g8931 ( 
.A(n_8683),
.Y(n_8931)
);

AND2x2_ASAP7_75t_L g8932 ( 
.A(n_8579),
.B(n_8602),
.Y(n_8932)
);

OAI21xp33_ASAP7_75t_L g8933 ( 
.A1(n_8691),
.A2(n_5855),
.B(n_5838),
.Y(n_8933)
);

INVx1_ASAP7_75t_L g8934 ( 
.A(n_8464),
.Y(n_8934)
);

OAI32xp33_ASAP7_75t_L g8935 ( 
.A1(n_8457),
.A2(n_5836),
.A3(n_5753),
.B1(n_5351),
.B2(n_5300),
.Y(n_8935)
);

INVx1_ASAP7_75t_L g8936 ( 
.A(n_8468),
.Y(n_8936)
);

AOI221xp5_ASAP7_75t_L g8937 ( 
.A1(n_8472),
.A2(n_6370),
.B1(n_6384),
.B2(n_6385),
.C(n_6374),
.Y(n_8937)
);

CKINVDCx5p33_ASAP7_75t_R g8938 ( 
.A(n_8773),
.Y(n_8938)
);

INVx1_ASAP7_75t_L g8939 ( 
.A(n_8703),
.Y(n_8939)
);

AND2x4_ASAP7_75t_L g8940 ( 
.A(n_8744),
.B(n_8476),
.Y(n_8940)
);

NAND2x1_ASAP7_75t_L g8941 ( 
.A(n_8744),
.B(n_8478),
.Y(n_8941)
);

INVxp67_ASAP7_75t_SL g8942 ( 
.A(n_8772),
.Y(n_8942)
);

NAND2xp5_ASAP7_75t_L g8943 ( 
.A(n_8713),
.B(n_6385),
.Y(n_8943)
);

AOI22xp33_ASAP7_75t_L g8944 ( 
.A1(n_8918),
.A2(n_8728),
.B1(n_8711),
.B2(n_8764),
.Y(n_8944)
);

INVx1_ASAP7_75t_L g8945 ( 
.A(n_8859),
.Y(n_8945)
);

AND2x2_ASAP7_75t_L g8946 ( 
.A(n_8858),
.B(n_5168),
.Y(n_8946)
);

OR2x2_ASAP7_75t_L g8947 ( 
.A(n_8762),
.B(n_5630),
.Y(n_8947)
);

NAND2xp5_ASAP7_75t_L g8948 ( 
.A(n_8851),
.B(n_6388),
.Y(n_8948)
);

NAND3xp33_ASAP7_75t_L g8949 ( 
.A(n_8712),
.B(n_8665),
.C(n_6389),
.Y(n_8949)
);

AOI221xp5_ASAP7_75t_L g8950 ( 
.A1(n_8747),
.A2(n_6389),
.B1(n_6396),
.B2(n_6391),
.C(n_6388),
.Y(n_8950)
);

NAND2xp5_ASAP7_75t_L g8951 ( 
.A(n_8851),
.B(n_6391),
.Y(n_8951)
);

AND2x2_ASAP7_75t_L g8952 ( 
.A(n_8730),
.B(n_5168),
.Y(n_8952)
);

INVxp33_ASAP7_75t_L g8953 ( 
.A(n_8718),
.Y(n_8953)
);

OR2x2_ASAP7_75t_L g8954 ( 
.A(n_8729),
.B(n_5635),
.Y(n_8954)
);

OR2x2_ASAP7_75t_L g8955 ( 
.A(n_8876),
.B(n_5635),
.Y(n_8955)
);

OR2x2_ASAP7_75t_L g8956 ( 
.A(n_8765),
.B(n_5640),
.Y(n_8956)
);

INVx1_ASAP7_75t_L g8957 ( 
.A(n_8707),
.Y(n_8957)
);

AND2x2_ASAP7_75t_L g8958 ( 
.A(n_8746),
.B(n_5838),
.Y(n_8958)
);

INVx2_ASAP7_75t_L g8959 ( 
.A(n_8812),
.Y(n_8959)
);

AOI21xp5_ASAP7_75t_L g8960 ( 
.A1(n_8745),
.A2(n_6399),
.B(n_6396),
.Y(n_8960)
);

INVx1_ASAP7_75t_L g8961 ( 
.A(n_8780),
.Y(n_8961)
);

INVx1_ASAP7_75t_L g8962 ( 
.A(n_8754),
.Y(n_8962)
);

INVx1_ASAP7_75t_L g8963 ( 
.A(n_8706),
.Y(n_8963)
);

AND2x2_ASAP7_75t_L g8964 ( 
.A(n_8820),
.B(n_5855),
.Y(n_8964)
);

INVx3_ASAP7_75t_L g8965 ( 
.A(n_8822),
.Y(n_8965)
);

INVx1_ASAP7_75t_L g8966 ( 
.A(n_8709),
.Y(n_8966)
);

INVx1_ASAP7_75t_SL g8967 ( 
.A(n_8809),
.Y(n_8967)
);

INVx1_ASAP7_75t_L g8968 ( 
.A(n_8732),
.Y(n_8968)
);

NAND2xp5_ASAP7_75t_L g8969 ( 
.A(n_8710),
.B(n_8763),
.Y(n_8969)
);

OR2x2_ASAP7_75t_L g8970 ( 
.A(n_8883),
.B(n_5640),
.Y(n_8970)
);

INVx1_ASAP7_75t_SL g8971 ( 
.A(n_8856),
.Y(n_8971)
);

AND2x2_ASAP7_75t_L g8972 ( 
.A(n_8774),
.B(n_8819),
.Y(n_8972)
);

INVx1_ASAP7_75t_L g8973 ( 
.A(n_8721),
.Y(n_8973)
);

NOR2xp33_ASAP7_75t_L g8974 ( 
.A(n_8826),
.B(n_6416),
.Y(n_8974)
);

OR2x2_ASAP7_75t_L g8975 ( 
.A(n_8726),
.B(n_5641),
.Y(n_8975)
);

INVx1_ASAP7_75t_L g8976 ( 
.A(n_8725),
.Y(n_8976)
);

OR2x2_ASAP7_75t_L g8977 ( 
.A(n_8771),
.B(n_5641),
.Y(n_8977)
);

CKINVDCx16_ASAP7_75t_R g8978 ( 
.A(n_8727),
.Y(n_8978)
);

AOI22xp5_ASAP7_75t_L g8979 ( 
.A1(n_8742),
.A2(n_6417),
.B1(n_6423),
.B2(n_6416),
.Y(n_8979)
);

INVx2_ASAP7_75t_L g8980 ( 
.A(n_8905),
.Y(n_8980)
);

INVx1_ASAP7_75t_L g8981 ( 
.A(n_8927),
.Y(n_8981)
);

INVx2_ASAP7_75t_SL g8982 ( 
.A(n_8734),
.Y(n_8982)
);

AND2x2_ASAP7_75t_L g8983 ( 
.A(n_8783),
.B(n_5855),
.Y(n_8983)
);

AND2x2_ASAP7_75t_L g8984 ( 
.A(n_8861),
.B(n_5855),
.Y(n_8984)
);

OR2x2_ASAP7_75t_L g8985 ( 
.A(n_8767),
.B(n_5642),
.Y(n_8985)
);

INVx1_ASAP7_75t_L g8986 ( 
.A(n_8717),
.Y(n_8986)
);

AND2x2_ASAP7_75t_L g8987 ( 
.A(n_8715),
.B(n_5895),
.Y(n_8987)
);

INVx1_ASAP7_75t_L g8988 ( 
.A(n_8716),
.Y(n_8988)
);

AND2x2_ASAP7_75t_L g8989 ( 
.A(n_8837),
.B(n_5895),
.Y(n_8989)
);

AND2x2_ASAP7_75t_L g8990 ( 
.A(n_8840),
.B(n_5895),
.Y(n_8990)
);

NAND2xp5_ASAP7_75t_L g8991 ( 
.A(n_8740),
.B(n_6417),
.Y(n_8991)
);

INVx2_ASAP7_75t_L g8992 ( 
.A(n_8905),
.Y(n_8992)
);

INVx2_ASAP7_75t_SL g8993 ( 
.A(n_8822),
.Y(n_8993)
);

AOI22xp5_ASAP7_75t_L g8994 ( 
.A1(n_8708),
.A2(n_6433),
.B1(n_6435),
.B2(n_6423),
.Y(n_8994)
);

NAND2xp5_ASAP7_75t_L g8995 ( 
.A(n_8814),
.B(n_6433),
.Y(n_8995)
);

INVx2_ASAP7_75t_L g8996 ( 
.A(n_8825),
.Y(n_8996)
);

AND2x2_ASAP7_75t_L g8997 ( 
.A(n_8832),
.B(n_5895),
.Y(n_8997)
);

NAND2xp5_ASAP7_75t_L g8998 ( 
.A(n_8724),
.B(n_6435),
.Y(n_8998)
);

INVxp67_ASAP7_75t_L g8999 ( 
.A(n_8791),
.Y(n_8999)
);

OR2x2_ASAP7_75t_L g9000 ( 
.A(n_8793),
.B(n_5642),
.Y(n_9000)
);

AND2x2_ASAP7_75t_L g9001 ( 
.A(n_8860),
.B(n_5912),
.Y(n_9001)
);

AND2x2_ASAP7_75t_L g9002 ( 
.A(n_8835),
.B(n_5912),
.Y(n_9002)
);

INVx1_ASAP7_75t_SL g9003 ( 
.A(n_8843),
.Y(n_9003)
);

INVx1_ASAP7_75t_SL g9004 ( 
.A(n_8796),
.Y(n_9004)
);

OR2x2_ASAP7_75t_L g9005 ( 
.A(n_8741),
.B(n_5646),
.Y(n_9005)
);

NOR2xp33_ASAP7_75t_L g9006 ( 
.A(n_8714),
.B(n_6436),
.Y(n_9006)
);

INVx1_ASAP7_75t_SL g9007 ( 
.A(n_8753),
.Y(n_9007)
);

INVx1_ASAP7_75t_L g9008 ( 
.A(n_8705),
.Y(n_9008)
);

CKINVDCx16_ASAP7_75t_R g9009 ( 
.A(n_8768),
.Y(n_9009)
);

OR2x2_ASAP7_75t_L g9010 ( 
.A(n_8842),
.B(n_5646),
.Y(n_9010)
);

AND2x2_ASAP7_75t_L g9011 ( 
.A(n_8868),
.B(n_8908),
.Y(n_9011)
);

INVx1_ASAP7_75t_L g9012 ( 
.A(n_8808),
.Y(n_9012)
);

AND2x2_ASAP7_75t_L g9013 ( 
.A(n_8731),
.B(n_5912),
.Y(n_9013)
);

INVx1_ASAP7_75t_L g9014 ( 
.A(n_8810),
.Y(n_9014)
);

INVxp67_ASAP7_75t_SL g9015 ( 
.A(n_8770),
.Y(n_9015)
);

INVx2_ASAP7_75t_L g9016 ( 
.A(n_8801),
.Y(n_9016)
);

AND2x2_ASAP7_75t_L g9017 ( 
.A(n_8776),
.B(n_5912),
.Y(n_9017)
);

INVx1_ASAP7_75t_L g9018 ( 
.A(n_8733),
.Y(n_9018)
);

NAND2xp5_ASAP7_75t_L g9019 ( 
.A(n_8750),
.B(n_6436),
.Y(n_9019)
);

AND2x2_ASAP7_75t_L g9020 ( 
.A(n_8930),
.B(n_8882),
.Y(n_9020)
);

NOR2xp33_ASAP7_75t_L g9021 ( 
.A(n_8811),
.B(n_6458),
.Y(n_9021)
);

AND2x4_ASAP7_75t_L g9022 ( 
.A(n_8722),
.B(n_6458),
.Y(n_9022)
);

AND2x2_ASAP7_75t_L g9023 ( 
.A(n_8887),
.B(n_4928),
.Y(n_9023)
);

NAND2xp5_ASAP7_75t_L g9024 ( 
.A(n_8909),
.B(n_6468),
.Y(n_9024)
);

HB1xp67_ASAP7_75t_L g9025 ( 
.A(n_8770),
.Y(n_9025)
);

OAI21xp33_ASAP7_75t_L g9026 ( 
.A1(n_8736),
.A2(n_5300),
.B(n_5214),
.Y(n_9026)
);

AND2x2_ASAP7_75t_L g9027 ( 
.A(n_8723),
.B(n_5022),
.Y(n_9027)
);

AND2x4_ASAP7_75t_L g9028 ( 
.A(n_8748),
.B(n_6468),
.Y(n_9028)
);

INVx1_ASAP7_75t_L g9029 ( 
.A(n_8737),
.Y(n_9029)
);

INVx1_ASAP7_75t_SL g9030 ( 
.A(n_8865),
.Y(n_9030)
);

NAND4xp75_ASAP7_75t_L g9031 ( 
.A(n_8786),
.B(n_6395),
.C(n_6460),
.D(n_6245),
.Y(n_9031)
);

AND2x2_ASAP7_75t_L g9032 ( 
.A(n_8749),
.B(n_5022),
.Y(n_9032)
);

BUFx3_ASAP7_75t_L g9033 ( 
.A(n_8766),
.Y(n_9033)
);

INVx2_ASAP7_75t_SL g9034 ( 
.A(n_8846),
.Y(n_9034)
);

NAND2xp5_ASAP7_75t_L g9035 ( 
.A(n_8912),
.B(n_6470),
.Y(n_9035)
);

INVx1_ASAP7_75t_SL g9036 ( 
.A(n_8932),
.Y(n_9036)
);

AND2x2_ASAP7_75t_L g9037 ( 
.A(n_8797),
.B(n_8829),
.Y(n_9037)
);

NOR2x1_ASAP7_75t_L g9038 ( 
.A(n_8719),
.B(n_5157),
.Y(n_9038)
);

AND2x2_ASAP7_75t_L g9039 ( 
.A(n_8790),
.B(n_8893),
.Y(n_9039)
);

HB1xp67_ASAP7_75t_L g9040 ( 
.A(n_8891),
.Y(n_9040)
);

BUFx3_ASAP7_75t_L g9041 ( 
.A(n_8815),
.Y(n_9041)
);

INVx1_ASAP7_75t_SL g9042 ( 
.A(n_8849),
.Y(n_9042)
);

INVx1_ASAP7_75t_L g9043 ( 
.A(n_8885),
.Y(n_9043)
);

INVx1_ASAP7_75t_SL g9044 ( 
.A(n_8788),
.Y(n_9044)
);

OAI22xp5_ASAP7_75t_L g9045 ( 
.A1(n_8845),
.A2(n_6484),
.B1(n_6492),
.B2(n_6470),
.Y(n_9045)
);

AND2x2_ASAP7_75t_L g9046 ( 
.A(n_8895),
.B(n_5109),
.Y(n_9046)
);

INVx1_ASAP7_75t_L g9047 ( 
.A(n_8739),
.Y(n_9047)
);

NAND2xp5_ASAP7_75t_SL g9048 ( 
.A(n_8779),
.B(n_6522),
.Y(n_9048)
);

AND2x2_ASAP7_75t_L g9049 ( 
.A(n_8900),
.B(n_5109),
.Y(n_9049)
);

INVx4_ASAP7_75t_L g9050 ( 
.A(n_8769),
.Y(n_9050)
);

INVx1_ASAP7_75t_SL g9051 ( 
.A(n_8775),
.Y(n_9051)
);

INVx3_ASAP7_75t_L g9052 ( 
.A(n_8879),
.Y(n_9052)
);

INVx1_ASAP7_75t_L g9053 ( 
.A(n_8704),
.Y(n_9053)
);

OR2x2_ASAP7_75t_L g9054 ( 
.A(n_8805),
.B(n_5647),
.Y(n_9054)
);

INVx1_ASAP7_75t_L g9055 ( 
.A(n_8894),
.Y(n_9055)
);

NOR2xp33_ASAP7_75t_L g9056 ( 
.A(n_8841),
.B(n_6520),
.Y(n_9056)
);

OR2x2_ASAP7_75t_L g9057 ( 
.A(n_8818),
.B(n_5647),
.Y(n_9057)
);

AOI22x1_ASAP7_75t_L g9058 ( 
.A1(n_8816),
.A2(n_5157),
.B1(n_5313),
.B2(n_5274),
.Y(n_9058)
);

CKINVDCx20_ASAP7_75t_L g9059 ( 
.A(n_8761),
.Y(n_9059)
);

INVx1_ASAP7_75t_L g9060 ( 
.A(n_8896),
.Y(n_9060)
);

INVx2_ASAP7_75t_L g9061 ( 
.A(n_8853),
.Y(n_9061)
);

INVx1_ASAP7_75t_L g9062 ( 
.A(n_8903),
.Y(n_9062)
);

AND2x2_ASAP7_75t_L g9063 ( 
.A(n_8878),
.B(n_5198),
.Y(n_9063)
);

INVx2_ASAP7_75t_L g9064 ( 
.A(n_8892),
.Y(n_9064)
);

INVx2_ASAP7_75t_L g9065 ( 
.A(n_8872),
.Y(n_9065)
);

NAND2xp5_ASAP7_75t_L g9066 ( 
.A(n_8907),
.B(n_6523),
.Y(n_9066)
);

OR2x2_ASAP7_75t_L g9067 ( 
.A(n_8848),
.B(n_5654),
.Y(n_9067)
);

INVx2_ASAP7_75t_SL g9068 ( 
.A(n_8879),
.Y(n_9068)
);

INVx2_ASAP7_75t_L g9069 ( 
.A(n_8920),
.Y(n_9069)
);

NOR2xp33_ASAP7_75t_L g9070 ( 
.A(n_8923),
.B(n_6523),
.Y(n_9070)
);

INVx1_ASAP7_75t_L g9071 ( 
.A(n_8813),
.Y(n_9071)
);

AND2x2_ASAP7_75t_L g9072 ( 
.A(n_8785),
.B(n_8850),
.Y(n_9072)
);

NAND3xp33_ASAP7_75t_L g9073 ( 
.A(n_8720),
.B(n_6540),
.C(n_6524),
.Y(n_9073)
);

OR2x2_ASAP7_75t_L g9074 ( 
.A(n_8751),
.B(n_8735),
.Y(n_9074)
);

NOR2x1p5_ASAP7_75t_L g9075 ( 
.A(n_8799),
.B(n_4810),
.Y(n_9075)
);

AND2x2_ASAP7_75t_L g9076 ( 
.A(n_8778),
.B(n_5198),
.Y(n_9076)
);

INVx1_ASAP7_75t_SL g9077 ( 
.A(n_8867),
.Y(n_9077)
);

AOI222xp33_ASAP7_75t_L g9078 ( 
.A1(n_8798),
.A2(n_6551),
.B1(n_6540),
.B2(n_6541),
.C1(n_6524),
.C2(n_5462),
.Y(n_9078)
);

INVx1_ASAP7_75t_L g9079 ( 
.A(n_8925),
.Y(n_9079)
);

INVx2_ASAP7_75t_L g9080 ( 
.A(n_8880),
.Y(n_9080)
);

AND2x2_ASAP7_75t_L g9081 ( 
.A(n_8752),
.B(n_5199),
.Y(n_9081)
);

AO22x1_ASAP7_75t_L g9082 ( 
.A1(n_8891),
.A2(n_4836),
.B1(n_4889),
.B2(n_4849),
.Y(n_9082)
);

NOR2x1_ASAP7_75t_L g9083 ( 
.A(n_8786),
.B(n_4849),
.Y(n_9083)
);

OAI22xp5_ASAP7_75t_L g9084 ( 
.A1(n_8757),
.A2(n_6551),
.B1(n_6541),
.B2(n_5657),
.Y(n_9084)
);

INVx1_ASAP7_75t_L g9085 ( 
.A(n_8852),
.Y(n_9085)
);

INVx1_ASAP7_75t_L g9086 ( 
.A(n_8847),
.Y(n_9086)
);

HB1xp67_ASAP7_75t_L g9087 ( 
.A(n_8904),
.Y(n_9087)
);

AND2x2_ASAP7_75t_L g9088 ( 
.A(n_8760),
.B(n_5199),
.Y(n_9088)
);

INVx1_ASAP7_75t_L g9089 ( 
.A(n_8870),
.Y(n_9089)
);

OR2x2_ASAP7_75t_L g9090 ( 
.A(n_8777),
.B(n_5654),
.Y(n_9090)
);

AND2x2_ASAP7_75t_L g9091 ( 
.A(n_8902),
.B(n_8806),
.Y(n_9091)
);

INVx1_ASAP7_75t_L g9092 ( 
.A(n_8869),
.Y(n_9092)
);

NAND2xp5_ASAP7_75t_L g9093 ( 
.A(n_8913),
.B(n_5657),
.Y(n_9093)
);

INVxp67_ASAP7_75t_L g9094 ( 
.A(n_8863),
.Y(n_9094)
);

AND2x2_ASAP7_75t_L g9095 ( 
.A(n_8784),
.B(n_5273),
.Y(n_9095)
);

NOR2x1_ASAP7_75t_L g9096 ( 
.A(n_8830),
.B(n_4849),
.Y(n_9096)
);

OR2x2_ASAP7_75t_L g9097 ( 
.A(n_8823),
.B(n_5658),
.Y(n_9097)
);

NOR2x1_ASAP7_75t_L g9098 ( 
.A(n_8836),
.B(n_4889),
.Y(n_9098)
);

INVx2_ASAP7_75t_L g9099 ( 
.A(n_8758),
.Y(n_9099)
);

INVx1_ASAP7_75t_L g9100 ( 
.A(n_8875),
.Y(n_9100)
);

AOI22xp33_ASAP7_75t_L g9101 ( 
.A1(n_8743),
.A2(n_6382),
.B1(n_6418),
.B2(n_6245),
.Y(n_9101)
);

INVx1_ASAP7_75t_SL g9102 ( 
.A(n_8792),
.Y(n_9102)
);

NAND3xp33_ASAP7_75t_L g9103 ( 
.A(n_8738),
.B(n_4898),
.C(n_4893),
.Y(n_9103)
);

AND2x2_ASAP7_75t_L g9104 ( 
.A(n_8854),
.B(n_5273),
.Y(n_9104)
);

AOI22xp5_ASAP7_75t_L g9105 ( 
.A1(n_8800),
.A2(n_5624),
.B1(n_5625),
.B2(n_5622),
.Y(n_9105)
);

INVx1_ASAP7_75t_L g9106 ( 
.A(n_8807),
.Y(n_9106)
);

NAND3xp33_ASAP7_75t_SL g9107 ( 
.A(n_8738),
.B(n_5312),
.C(n_4918),
.Y(n_9107)
);

INVx1_ASAP7_75t_SL g9108 ( 
.A(n_8759),
.Y(n_9108)
);

INVx1_ASAP7_75t_SL g9109 ( 
.A(n_8802),
.Y(n_9109)
);

INVx1_ASAP7_75t_L g9110 ( 
.A(n_8831),
.Y(n_9110)
);

AND2x2_ASAP7_75t_L g9111 ( 
.A(n_8839),
.B(n_5364),
.Y(n_9111)
);

INVx1_ASAP7_75t_L g9112 ( 
.A(n_8931),
.Y(n_9112)
);

AND2x2_ASAP7_75t_L g9113 ( 
.A(n_8844),
.B(n_5364),
.Y(n_9113)
);

INVxp67_ASAP7_75t_L g9114 ( 
.A(n_8838),
.Y(n_9114)
);

AND2x2_ASAP7_75t_L g9115 ( 
.A(n_8877),
.B(n_4889),
.Y(n_9115)
);

AND2x2_ASAP7_75t_L g9116 ( 
.A(n_8929),
.B(n_4942),
.Y(n_9116)
);

NAND2xp5_ASAP7_75t_L g9117 ( 
.A(n_8901),
.B(n_5658),
.Y(n_9117)
);

OR2x2_ASAP7_75t_L g9118 ( 
.A(n_8862),
.B(n_5659),
.Y(n_9118)
);

NAND2x1_ASAP7_75t_L g9119 ( 
.A(n_8866),
.B(n_8934),
.Y(n_9119)
);

INVx1_ASAP7_75t_L g9120 ( 
.A(n_8834),
.Y(n_9120)
);

BUFx6f_ASAP7_75t_L g9121 ( 
.A(n_8936),
.Y(n_9121)
);

INVx1_ASAP7_75t_L g9122 ( 
.A(n_8916),
.Y(n_9122)
);

INVx2_ASAP7_75t_L g9123 ( 
.A(n_8889),
.Y(n_9123)
);

AND2x4_ASAP7_75t_L g9124 ( 
.A(n_8787),
.B(n_4810),
.Y(n_9124)
);

INVx1_ASAP7_75t_L g9125 ( 
.A(n_8890),
.Y(n_9125)
);

HB1xp67_ASAP7_75t_L g9126 ( 
.A(n_8817),
.Y(n_9126)
);

CKINVDCx16_ASAP7_75t_R g9127 ( 
.A(n_8782),
.Y(n_9127)
);

INVx1_ASAP7_75t_L g9128 ( 
.A(n_8755),
.Y(n_9128)
);

AOI22xp33_ASAP7_75t_L g9129 ( 
.A1(n_8906),
.A2(n_6382),
.B1(n_6418),
.B2(n_6460),
.Y(n_9129)
);

AND2x4_ASAP7_75t_L g9130 ( 
.A(n_8959),
.B(n_8794),
.Y(n_9130)
);

INVx2_ASAP7_75t_L g9131 ( 
.A(n_8972),
.Y(n_9131)
);

AND2x2_ASAP7_75t_L g9132 ( 
.A(n_8939),
.B(n_8964),
.Y(n_9132)
);

INVxp67_ASAP7_75t_L g9133 ( 
.A(n_9025),
.Y(n_9133)
);

INVx1_ASAP7_75t_L g9134 ( 
.A(n_8939),
.Y(n_9134)
);

OAI211xp5_ASAP7_75t_L g9135 ( 
.A1(n_9015),
.A2(n_8824),
.B(n_8756),
.C(n_8781),
.Y(n_9135)
);

NAND4xp75_ASAP7_75t_L g9136 ( 
.A(n_9039),
.B(n_8789),
.C(n_8911),
.D(n_8910),
.Y(n_9136)
);

OAI211xp5_ASAP7_75t_L g9137 ( 
.A1(n_8944),
.A2(n_8795),
.B(n_8917),
.C(n_8874),
.Y(n_9137)
);

INVxp67_ASAP7_75t_SL g9138 ( 
.A(n_8942),
.Y(n_9138)
);

NOR2xp33_ASAP7_75t_SL g9139 ( 
.A(n_8938),
.B(n_8897),
.Y(n_9139)
);

NAND3x1_ASAP7_75t_L g9140 ( 
.A(n_9052),
.B(n_8828),
.C(n_8937),
.Y(n_9140)
);

INVx2_ASAP7_75t_L g9141 ( 
.A(n_9059),
.Y(n_9141)
);

NAND2xp5_ASAP7_75t_SL g9142 ( 
.A(n_9127),
.B(n_8901),
.Y(n_9142)
);

INVxp67_ASAP7_75t_SL g9143 ( 
.A(n_9052),
.Y(n_9143)
);

AOI21xp33_ASAP7_75t_L g9144 ( 
.A1(n_9051),
.A2(n_8899),
.B(n_8919),
.Y(n_9144)
);

INVx1_ASAP7_75t_SL g9145 ( 
.A(n_9102),
.Y(n_9145)
);

OAI21xp33_ASAP7_75t_SL g9146 ( 
.A1(n_9128),
.A2(n_8888),
.B(n_8881),
.Y(n_9146)
);

AND2x2_ASAP7_75t_L g9147 ( 
.A(n_8978),
.B(n_8933),
.Y(n_9147)
);

INVx1_ASAP7_75t_L g9148 ( 
.A(n_8941),
.Y(n_9148)
);

A2O1A1Ixp33_ASAP7_75t_L g9149 ( 
.A1(n_9085),
.A2(n_8833),
.B(n_8881),
.C(n_8804),
.Y(n_9149)
);

NAND2xp5_ASAP7_75t_L g9150 ( 
.A(n_9009),
.B(n_9036),
.Y(n_9150)
);

OAI221xp5_ASAP7_75t_SL g9151 ( 
.A1(n_9101),
.A2(n_8821),
.B1(n_8855),
.B2(n_8803),
.C(n_8857),
.Y(n_9151)
);

INVxp67_ASAP7_75t_L g9152 ( 
.A(n_8982),
.Y(n_9152)
);

NAND2xp5_ASAP7_75t_SL g9153 ( 
.A(n_9121),
.B(n_8915),
.Y(n_9153)
);

OAI21xp33_ASAP7_75t_L g9154 ( 
.A1(n_8953),
.A2(n_8898),
.B(n_8928),
.Y(n_9154)
);

INVx2_ASAP7_75t_L g9155 ( 
.A(n_9121),
.Y(n_9155)
);

INVx1_ASAP7_75t_L g9156 ( 
.A(n_9011),
.Y(n_9156)
);

AOI21xp33_ASAP7_75t_R g9157 ( 
.A1(n_8962),
.A2(n_8873),
.B(n_8827),
.Y(n_9157)
);

NAND3xp33_ASAP7_75t_L g9158 ( 
.A(n_9085),
.B(n_8924),
.C(n_8886),
.Y(n_9158)
);

NAND2x1_ASAP7_75t_L g9159 ( 
.A(n_9083),
.B(n_8884),
.Y(n_9159)
);

INVx2_ASAP7_75t_L g9160 ( 
.A(n_9121),
.Y(n_9160)
);

AND2x2_ASAP7_75t_L g9161 ( 
.A(n_8958),
.B(n_8922),
.Y(n_9161)
);

INVx1_ASAP7_75t_L g9162 ( 
.A(n_8965),
.Y(n_9162)
);

NAND2xp33_ASAP7_75t_SL g9163 ( 
.A(n_9119),
.B(n_4942),
.Y(n_9163)
);

NAND2xp5_ASAP7_75t_L g9164 ( 
.A(n_8965),
.B(n_8864),
.Y(n_9164)
);

INVx1_ASAP7_75t_L g9165 ( 
.A(n_9079),
.Y(n_9165)
);

INVx1_ASAP7_75t_L g9166 ( 
.A(n_9079),
.Y(n_9166)
);

AOI22xp5_ASAP7_75t_L g9167 ( 
.A1(n_9048),
.A2(n_8914),
.B1(n_8871),
.B2(n_8926),
.Y(n_9167)
);

INVx1_ASAP7_75t_L g9168 ( 
.A(n_8940),
.Y(n_9168)
);

INVx1_ASAP7_75t_L g9169 ( 
.A(n_8940),
.Y(n_9169)
);

INVx1_ASAP7_75t_L g9170 ( 
.A(n_8957),
.Y(n_9170)
);

INVx1_ASAP7_75t_L g9171 ( 
.A(n_8945),
.Y(n_9171)
);

INVx1_ASAP7_75t_L g9172 ( 
.A(n_8980),
.Y(n_9172)
);

INVx1_ASAP7_75t_L g9173 ( 
.A(n_8992),
.Y(n_9173)
);

AOI21xp33_ASAP7_75t_L g9174 ( 
.A1(n_9114),
.A2(n_8921),
.B(n_8935),
.Y(n_9174)
);

INVx1_ASAP7_75t_L g9175 ( 
.A(n_8969),
.Y(n_9175)
);

INVx1_ASAP7_75t_L g9176 ( 
.A(n_8955),
.Y(n_9176)
);

A2O1A1Ixp33_ASAP7_75t_L g9177 ( 
.A1(n_9021),
.A2(n_5624),
.B(n_5625),
.C(n_5622),
.Y(n_9177)
);

INVx1_ASAP7_75t_L g9178 ( 
.A(n_9033),
.Y(n_9178)
);

AND2x2_ASAP7_75t_L g9179 ( 
.A(n_8983),
.B(n_8967),
.Y(n_9179)
);

O2A1O1Ixp5_ASAP7_75t_L g9180 ( 
.A1(n_9128),
.A2(n_5300),
.B(n_5351),
.C(n_5214),
.Y(n_9180)
);

INVx2_ASAP7_75t_L g9181 ( 
.A(n_8946),
.Y(n_9181)
);

OAI32xp33_ASAP7_75t_L g9182 ( 
.A1(n_9003),
.A2(n_5351),
.A3(n_5319),
.B1(n_4285),
.B2(n_4338),
.Y(n_9182)
);

INVxp67_ASAP7_75t_SL g9183 ( 
.A(n_9087),
.Y(n_9183)
);

INVx2_ASAP7_75t_L g9184 ( 
.A(n_9041),
.Y(n_9184)
);

AND2x2_ASAP7_75t_L g9185 ( 
.A(n_8971),
.B(n_4942),
.Y(n_9185)
);

AOI22xp5_ASAP7_75t_L g9186 ( 
.A1(n_9042),
.A2(n_5632),
.B1(n_5648),
.B2(n_5631),
.Y(n_9186)
);

OAI21xp5_ASAP7_75t_SL g9187 ( 
.A1(n_9007),
.A2(n_5673),
.B(n_5669),
.Y(n_9187)
);

NAND2xp5_ASAP7_75t_L g9188 ( 
.A(n_9004),
.B(n_5631),
.Y(n_9188)
);

A2O1A1Ixp33_ASAP7_75t_L g9189 ( 
.A1(n_9074),
.A2(n_5648),
.B(n_5652),
.C(n_5632),
.Y(n_9189)
);

NAND2xp5_ASAP7_75t_L g9190 ( 
.A(n_8993),
.B(n_9068),
.Y(n_9190)
);

OA21x2_ASAP7_75t_L g9191 ( 
.A1(n_9120),
.A2(n_5823),
.B(n_5786),
.Y(n_9191)
);

AOI22xp5_ASAP7_75t_L g9192 ( 
.A1(n_9044),
.A2(n_5656),
.B1(n_5666),
.B2(n_5652),
.Y(n_9192)
);

OR2x2_ASAP7_75t_L g9193 ( 
.A(n_9016),
.B(n_5659),
.Y(n_9193)
);

INVx2_ASAP7_75t_L g9194 ( 
.A(n_8952),
.Y(n_9194)
);

HB1xp67_ASAP7_75t_L g9195 ( 
.A(n_9040),
.Y(n_9195)
);

AND2x2_ASAP7_75t_L g9196 ( 
.A(n_9013),
.B(n_4942),
.Y(n_9196)
);

INVx1_ASAP7_75t_L g9197 ( 
.A(n_9019),
.Y(n_9197)
);

INVx1_ASAP7_75t_L g9198 ( 
.A(n_8981),
.Y(n_9198)
);

OAI22xp5_ASAP7_75t_L g9199 ( 
.A1(n_8963),
.A2(n_3955),
.B1(n_5676),
.B2(n_5663),
.Y(n_9199)
);

INVx2_ASAP7_75t_SL g9200 ( 
.A(n_9017),
.Y(n_9200)
);

INVx1_ASAP7_75t_L g9201 ( 
.A(n_8966),
.Y(n_9201)
);

INVx1_ASAP7_75t_L g9202 ( 
.A(n_8968),
.Y(n_9202)
);

INVx1_ASAP7_75t_L g9203 ( 
.A(n_9018),
.Y(n_9203)
);

INVx2_ASAP7_75t_L g9204 ( 
.A(n_9020),
.Y(n_9204)
);

NAND2xp5_ASAP7_75t_L g9205 ( 
.A(n_8986),
.B(n_5656),
.Y(n_9205)
);

OAI22xp33_ASAP7_75t_L g9206 ( 
.A1(n_8943),
.A2(n_5668),
.B1(n_5681),
.B2(n_5666),
.Y(n_9206)
);

AOI321xp33_ASAP7_75t_L g9207 ( 
.A1(n_9038),
.A2(n_4896),
.A3(n_4856),
.B1(n_4892),
.B2(n_5341),
.C(n_4729),
.Y(n_9207)
);

NAND3xp33_ASAP7_75t_SL g9208 ( 
.A(n_9109),
.B(n_5681),
.C(n_5668),
.Y(n_9208)
);

OR2x2_ASAP7_75t_L g9209 ( 
.A(n_9030),
.B(n_5663),
.Y(n_9209)
);

INVx2_ASAP7_75t_L g9210 ( 
.A(n_9099),
.Y(n_9210)
);

AND2x2_ASAP7_75t_L g9211 ( 
.A(n_8984),
.B(n_4948),
.Y(n_9211)
);

INVx1_ASAP7_75t_L g9212 ( 
.A(n_9029),
.Y(n_9212)
);

AOI22xp5_ASAP7_75t_L g9213 ( 
.A1(n_8973),
.A2(n_5691),
.B1(n_5703),
.B2(n_5685),
.Y(n_9213)
);

OR2x2_ASAP7_75t_L g9214 ( 
.A(n_9050),
.B(n_5667),
.Y(n_9214)
);

INVx1_ASAP7_75t_L g9215 ( 
.A(n_8948),
.Y(n_9215)
);

NAND2xp5_ASAP7_75t_L g9216 ( 
.A(n_9050),
.B(n_5685),
.Y(n_9216)
);

AOI22xp5_ASAP7_75t_L g9217 ( 
.A1(n_9108),
.A2(n_5703),
.B1(n_5704),
.B2(n_5691),
.Y(n_9217)
);

INVx1_ASAP7_75t_L g9218 ( 
.A(n_8951),
.Y(n_9218)
);

AOI322xp5_ASAP7_75t_L g9219 ( 
.A1(n_9008),
.A2(n_5704),
.A3(n_5475),
.B1(n_5478),
.B2(n_5462),
.C1(n_5483),
.C2(n_5482),
.Y(n_9219)
);

NAND2xp5_ASAP7_75t_L g9220 ( 
.A(n_8976),
.B(n_5667),
.Y(n_9220)
);

NAND2xp33_ASAP7_75t_SL g9221 ( 
.A(n_9034),
.B(n_4948),
.Y(n_9221)
);

INVx1_ASAP7_75t_L g9222 ( 
.A(n_9072),
.Y(n_9222)
);

OAI22xp5_ASAP7_75t_L g9223 ( 
.A1(n_9061),
.A2(n_3955),
.B1(n_5723),
.B2(n_5693),
.Y(n_9223)
);

INVx1_ASAP7_75t_SL g9224 ( 
.A(n_9077),
.Y(n_9224)
);

OAI21xp33_ASAP7_75t_L g9225 ( 
.A1(n_9123),
.A2(n_4313),
.B(n_4285),
.Y(n_9225)
);

INVxp67_ASAP7_75t_L g9226 ( 
.A(n_9126),
.Y(n_9226)
);

NOR2xp33_ASAP7_75t_L g9227 ( 
.A(n_8999),
.B(n_5458),
.Y(n_9227)
);

AND2x2_ASAP7_75t_L g9228 ( 
.A(n_9001),
.B(n_4948),
.Y(n_9228)
);

INVxp67_ASAP7_75t_SL g9229 ( 
.A(n_9065),
.Y(n_9229)
);

INVx1_ASAP7_75t_L g9230 ( 
.A(n_8988),
.Y(n_9230)
);

INVx1_ASAP7_75t_L g9231 ( 
.A(n_9080),
.Y(n_9231)
);

OAI22xp5_ASAP7_75t_L g9232 ( 
.A1(n_9069),
.A2(n_5731),
.B1(n_5756),
.B2(n_5697),
.Y(n_9232)
);

AOI22xp5_ASAP7_75t_L g9233 ( 
.A1(n_9064),
.A2(n_5463),
.B1(n_5475),
.B2(n_5458),
.Y(n_9233)
);

HB1xp67_ASAP7_75t_L g9234 ( 
.A(n_9096),
.Y(n_9234)
);

INVx2_ASAP7_75t_L g9235 ( 
.A(n_8989),
.Y(n_9235)
);

INVx1_ASAP7_75t_L g9236 ( 
.A(n_9022),
.Y(n_9236)
);

AND2x2_ASAP7_75t_L g9237 ( 
.A(n_8997),
.B(n_4948),
.Y(n_9237)
);

A2O1A1Ixp33_ASAP7_75t_SL g9238 ( 
.A1(n_9008),
.A2(n_5676),
.B(n_5680),
.C(n_5675),
.Y(n_9238)
);

NOR2xp67_ASAP7_75t_L g9239 ( 
.A(n_9012),
.B(n_4988),
.Y(n_9239)
);

NAND3xp33_ASAP7_75t_L g9240 ( 
.A(n_8961),
.B(n_6493),
.C(n_6460),
.Y(n_9240)
);

NAND2xp5_ASAP7_75t_L g9241 ( 
.A(n_9022),
.B(n_5675),
.Y(n_9241)
);

OAI222xp33_ASAP7_75t_L g9242 ( 
.A1(n_8994),
.A2(n_4914),
.B1(n_4924),
.B2(n_4957),
.C1(n_4925),
.C2(n_4898),
.Y(n_9242)
);

AOI211xp5_ASAP7_75t_L g9243 ( 
.A1(n_9006),
.A2(n_9053),
.B(n_9091),
.C(n_9047),
.Y(n_9243)
);

NAND2xp5_ASAP7_75t_L g9244 ( 
.A(n_9028),
.B(n_5680),
.Y(n_9244)
);

AOI32xp33_ASAP7_75t_L g9245 ( 
.A1(n_9043),
.A2(n_5823),
.A3(n_5786),
.B1(n_5764),
.B2(n_5776),
.Y(n_9245)
);

INVx1_ASAP7_75t_L g9246 ( 
.A(n_9028),
.Y(n_9246)
);

OAI21xp5_ASAP7_75t_L g9247 ( 
.A1(n_9098),
.A2(n_6493),
.B(n_5554),
.Y(n_9247)
);

INVx1_ASAP7_75t_SL g9248 ( 
.A(n_9037),
.Y(n_9248)
);

NOR2xp33_ASAP7_75t_L g9249 ( 
.A(n_9092),
.B(n_5463),
.Y(n_9249)
);

AND2x2_ASAP7_75t_L g9250 ( 
.A(n_9002),
.B(n_4988),
.Y(n_9250)
);

INVx1_ASAP7_75t_L g9251 ( 
.A(n_9062),
.Y(n_9251)
);

NAND2xp5_ASAP7_75t_L g9252 ( 
.A(n_9104),
.B(n_5688),
.Y(n_9252)
);

INVx1_ASAP7_75t_L g9253 ( 
.A(n_8949),
.Y(n_9253)
);

INVxp67_ASAP7_75t_L g9254 ( 
.A(n_8974),
.Y(n_9254)
);

OR2x2_ASAP7_75t_L g9255 ( 
.A(n_9014),
.B(n_5688),
.Y(n_9255)
);

AOI222xp33_ASAP7_75t_L g9256 ( 
.A1(n_9073),
.A2(n_5482),
.B1(n_5478),
.B2(n_5490),
.C1(n_5486),
.C2(n_5483),
.Y(n_9256)
);

INVx1_ASAP7_75t_L g9257 ( 
.A(n_9000),
.Y(n_9257)
);

NAND2xp5_ASAP7_75t_SL g9258 ( 
.A(n_8996),
.B(n_5486),
.Y(n_9258)
);

AND2x2_ASAP7_75t_L g9259 ( 
.A(n_8987),
.B(n_4988),
.Y(n_9259)
);

INVx1_ASAP7_75t_L g9260 ( 
.A(n_8995),
.Y(n_9260)
);

OAI22xp33_ASAP7_75t_L g9261 ( 
.A1(n_8991),
.A2(n_5490),
.B1(n_5520),
.B2(n_5499),
.Y(n_9261)
);

AND2x2_ASAP7_75t_L g9262 ( 
.A(n_8990),
.B(n_4988),
.Y(n_9262)
);

INVx1_ASAP7_75t_L g9263 ( 
.A(n_9071),
.Y(n_9263)
);

INVx2_ASAP7_75t_L g9264 ( 
.A(n_9031),
.Y(n_9264)
);

AOI221xp5_ASAP7_75t_L g9265 ( 
.A1(n_9129),
.A2(n_6382),
.B1(n_6418),
.B2(n_5524),
.C(n_5538),
.Y(n_9265)
);

AOI21xp33_ASAP7_75t_L g9266 ( 
.A1(n_9056),
.A2(n_6493),
.B(n_6506),
.Y(n_9266)
);

INVx1_ASAP7_75t_SL g9267 ( 
.A(n_9124),
.Y(n_9267)
);

OAI21xp5_ASAP7_75t_SL g9268 ( 
.A1(n_9094),
.A2(n_5673),
.B(n_5669),
.Y(n_9268)
);

AOI21xp33_ASAP7_75t_L g9269 ( 
.A1(n_9070),
.A2(n_8998),
.B(n_9100),
.Y(n_9269)
);

NAND2xp5_ASAP7_75t_L g9270 ( 
.A(n_9116),
.B(n_5693),
.Y(n_9270)
);

INVx2_ASAP7_75t_L g9271 ( 
.A(n_9058),
.Y(n_9271)
);

NOR3xp33_ASAP7_75t_L g9272 ( 
.A(n_9055),
.B(n_5520),
.C(n_5499),
.Y(n_9272)
);

NOR2xp33_ASAP7_75t_L g9273 ( 
.A(n_9060),
.B(n_5524),
.Y(n_9273)
);

OAI21xp5_ASAP7_75t_L g9274 ( 
.A1(n_8960),
.A2(n_5541),
.B(n_5538),
.Y(n_9274)
);

INVx1_ASAP7_75t_L g9275 ( 
.A(n_8977),
.Y(n_9275)
);

AOI22xp5_ASAP7_75t_L g9276 ( 
.A1(n_9078),
.A2(n_5541),
.B1(n_5554),
.B2(n_6506),
.Y(n_9276)
);

OAI22xp5_ASAP7_75t_L g9277 ( 
.A1(n_9112),
.A2(n_5748),
.B1(n_5765),
.B2(n_5723),
.Y(n_9277)
);

AND2x2_ASAP7_75t_L g9278 ( 
.A(n_9115),
.B(n_4994),
.Y(n_9278)
);

OAI321xp33_ASAP7_75t_L g9279 ( 
.A1(n_9026),
.A2(n_9107),
.A3(n_9066),
.B1(n_9035),
.B2(n_9024),
.C(n_8979),
.Y(n_9279)
);

OAI222xp33_ASAP7_75t_L g9280 ( 
.A1(n_9045),
.A2(n_4957),
.B1(n_4924),
.B2(n_4962),
.C1(n_4925),
.C2(n_4914),
.Y(n_9280)
);

NAND2xp5_ASAP7_75t_L g9281 ( 
.A(n_9027),
.B(n_9032),
.Y(n_9281)
);

INVx1_ASAP7_75t_L g9282 ( 
.A(n_8985),
.Y(n_9282)
);

AOI22x1_ASAP7_75t_L g9283 ( 
.A1(n_9075),
.A2(n_5274),
.B1(n_5313),
.B2(n_5697),
.Y(n_9283)
);

AOI221xp5_ASAP7_75t_L g9284 ( 
.A1(n_9125),
.A2(n_6555),
.B1(n_6542),
.B2(n_6506),
.C(n_4925),
.Y(n_9284)
);

OAI21xp33_ASAP7_75t_SL g9285 ( 
.A1(n_9076),
.A2(n_5764),
.B(n_5784),
.Y(n_9285)
);

NAND2xp5_ASAP7_75t_L g9286 ( 
.A(n_9122),
.B(n_5698),
.Y(n_9286)
);

NAND2xp5_ASAP7_75t_SL g9287 ( 
.A(n_9124),
.B(n_5669),
.Y(n_9287)
);

AOI221x1_ASAP7_75t_L g9288 ( 
.A1(n_9106),
.A2(n_5972),
.B1(n_5701),
.B2(n_5702),
.C(n_5700),
.Y(n_9288)
);

NAND2xp5_ASAP7_75t_L g9289 ( 
.A(n_9081),
.B(n_5698),
.Y(n_9289)
);

AND2x2_ASAP7_75t_L g9290 ( 
.A(n_9095),
.B(n_4994),
.Y(n_9290)
);

INVx1_ASAP7_75t_L g9291 ( 
.A(n_8970),
.Y(n_9291)
);

INVx2_ASAP7_75t_L g9292 ( 
.A(n_9058),
.Y(n_9292)
);

NOR2x1_ASAP7_75t_L g9293 ( 
.A(n_9110),
.B(n_5422),
.Y(n_9293)
);

OAI22xp5_ASAP7_75t_L g9294 ( 
.A1(n_9010),
.A2(n_5759),
.B1(n_5774),
.B2(n_5736),
.Y(n_9294)
);

INVx1_ASAP7_75t_L g9295 ( 
.A(n_9088),
.Y(n_9295)
);

AOI22xp5_ASAP7_75t_L g9296 ( 
.A1(n_9086),
.A2(n_6555),
.B1(n_6542),
.B2(n_5626),
.Y(n_9296)
);

O2A1O1Ixp33_ASAP7_75t_L g9297 ( 
.A1(n_9089),
.A2(n_5798),
.B(n_5999),
.C(n_5834),
.Y(n_9297)
);

INVx1_ASAP7_75t_L g9298 ( 
.A(n_9111),
.Y(n_9298)
);

NAND2xp5_ASAP7_75t_SL g9299 ( 
.A(n_9113),
.B(n_5669),
.Y(n_9299)
);

OAI22xp5_ASAP7_75t_L g9300 ( 
.A1(n_8947),
.A2(n_5737),
.B1(n_5760),
.B2(n_5700),
.Y(n_9300)
);

OAI22xp5_ASAP7_75t_L g9301 ( 
.A1(n_9057),
.A2(n_5738),
.B1(n_5761),
.B2(n_5701),
.Y(n_9301)
);

O2A1O1Ixp33_ASAP7_75t_L g9302 ( 
.A1(n_9117),
.A2(n_5798),
.B(n_5999),
.C(n_5834),
.Y(n_9302)
);

AND2x2_ASAP7_75t_L g9303 ( 
.A(n_9023),
.B(n_4994),
.Y(n_9303)
);

NAND2x1p5_ASAP7_75t_L g9304 ( 
.A(n_8954),
.B(n_8956),
.Y(n_9304)
);

AOI222xp33_ASAP7_75t_L g9305 ( 
.A1(n_8950),
.A2(n_5781),
.B1(n_5778),
.B2(n_5796),
.C1(n_5795),
.C2(n_5794),
.Y(n_9305)
);

OAI22xp5_ASAP7_75t_L g9306 ( 
.A1(n_9054),
.A2(n_5707),
.B1(n_5768),
.B2(n_5748),
.Y(n_9306)
);

OR2x2_ASAP7_75t_L g9307 ( 
.A(n_8975),
.B(n_5702),
.Y(n_9307)
);

OAI21xp33_ASAP7_75t_L g9308 ( 
.A1(n_9063),
.A2(n_4338),
.B(n_4313),
.Y(n_9308)
);

NAND2x1_ASAP7_75t_L g9309 ( 
.A(n_9067),
.B(n_5180),
.Y(n_9309)
);

OAI22xp5_ASAP7_75t_L g9310 ( 
.A1(n_9090),
.A2(n_5759),
.B1(n_5774),
.B2(n_5732),
.Y(n_9310)
);

NAND2xp5_ASAP7_75t_L g9311 ( 
.A(n_9145),
.B(n_9046),
.Y(n_9311)
);

NAND2xp5_ASAP7_75t_L g9312 ( 
.A(n_9132),
.B(n_9143),
.Y(n_9312)
);

AOI21xp5_ASAP7_75t_L g9313 ( 
.A1(n_9150),
.A2(n_9093),
.B(n_9005),
.Y(n_9313)
);

AND2x2_ASAP7_75t_L g9314 ( 
.A(n_9131),
.B(n_9049),
.Y(n_9314)
);

NOR3xp33_ASAP7_75t_SL g9315 ( 
.A(n_9135),
.B(n_9084),
.C(n_9103),
.Y(n_9315)
);

NAND3xp33_ASAP7_75t_L g9316 ( 
.A(n_9226),
.B(n_9118),
.C(n_9097),
.Y(n_9316)
);

INVx1_ASAP7_75t_L g9317 ( 
.A(n_9138),
.Y(n_9317)
);

INVx2_ASAP7_75t_SL g9318 ( 
.A(n_9179),
.Y(n_9318)
);

OAI22xp5_ASAP7_75t_L g9319 ( 
.A1(n_9229),
.A2(n_9105),
.B1(n_9082),
.B2(n_5728),
.Y(n_9319)
);

INVx1_ASAP7_75t_L g9320 ( 
.A(n_9195),
.Y(n_9320)
);

NOR3xp33_ASAP7_75t_L g9321 ( 
.A(n_9144),
.B(n_4918),
.C(n_5249),
.Y(n_9321)
);

INVx2_ASAP7_75t_SL g9322 ( 
.A(n_9204),
.Y(n_9322)
);

NAND3xp33_ASAP7_75t_L g9323 ( 
.A(n_9243),
.B(n_4924),
.C(n_4914),
.Y(n_9323)
);

INVx1_ASAP7_75t_L g9324 ( 
.A(n_9183),
.Y(n_9324)
);

AOI22xp5_ASAP7_75t_L g9325 ( 
.A1(n_9264),
.A2(n_6555),
.B1(n_6542),
.B2(n_5626),
.Y(n_9325)
);

AOI21xp33_ASAP7_75t_SL g9326 ( 
.A1(n_9142),
.A2(n_4736),
.B(n_4689),
.Y(n_9326)
);

INVx1_ASAP7_75t_SL g9327 ( 
.A(n_9248),
.Y(n_9327)
);

NAND2xp5_ASAP7_75t_L g9328 ( 
.A(n_9168),
.B(n_9169),
.Y(n_9328)
);

NOR3xp33_ASAP7_75t_SL g9329 ( 
.A(n_9153),
.B(n_4920),
.C(n_4913),
.Y(n_9329)
);

INVx1_ASAP7_75t_L g9330 ( 
.A(n_9156),
.Y(n_9330)
);

NOR2xp33_ASAP7_75t_L g9331 ( 
.A(n_9267),
.B(n_5534),
.Y(n_9331)
);

OAI22xp33_ASAP7_75t_SL g9332 ( 
.A1(n_9159),
.A2(n_5781),
.B1(n_5794),
.B2(n_5778),
.Y(n_9332)
);

O2A1O1Ixp33_ASAP7_75t_L g9333 ( 
.A1(n_9149),
.A2(n_5798),
.B(n_5534),
.C(n_5626),
.Y(n_9333)
);

AOI21xp5_ASAP7_75t_L g9334 ( 
.A1(n_9163),
.A2(n_9190),
.B(n_9133),
.Y(n_9334)
);

HB1xp67_ASAP7_75t_L g9335 ( 
.A(n_9239),
.Y(n_9335)
);

INVx1_ASAP7_75t_L g9336 ( 
.A(n_9222),
.Y(n_9336)
);

OAI21xp5_ASAP7_75t_SL g9337 ( 
.A1(n_9224),
.A2(n_5673),
.B(n_5674),
.Y(n_9337)
);

INVxp67_ASAP7_75t_SL g9338 ( 
.A(n_9304),
.Y(n_9338)
);

AOI22xp33_ASAP7_75t_L g9339 ( 
.A1(n_9197),
.A2(n_5626),
.B1(n_5534),
.B2(n_4962),
.Y(n_9339)
);

AND2x2_ASAP7_75t_L g9340 ( 
.A(n_9185),
.B(n_4879),
.Y(n_9340)
);

OAI211xp5_ASAP7_75t_SL g9341 ( 
.A1(n_9146),
.A2(n_5707),
.B(n_5731),
.C(n_5728),
.Y(n_9341)
);

OAI22xp33_ASAP7_75t_SL g9342 ( 
.A1(n_9253),
.A2(n_5796),
.B1(n_5805),
.B2(n_5795),
.Y(n_9342)
);

INVx1_ASAP7_75t_L g9343 ( 
.A(n_9165),
.Y(n_9343)
);

AOI22xp5_ASAP7_75t_L g9344 ( 
.A1(n_9140),
.A2(n_5534),
.B1(n_5999),
.B2(n_5834),
.Y(n_9344)
);

AND2x2_ASAP7_75t_L g9345 ( 
.A(n_9200),
.B(n_4879),
.Y(n_9345)
);

OAI322xp33_ASAP7_75t_L g9346 ( 
.A1(n_9139),
.A2(n_4974),
.A3(n_4957),
.B1(n_4978),
.B2(n_4982),
.C1(n_4971),
.C2(n_4962),
.Y(n_9346)
);

OR2x2_ASAP7_75t_L g9347 ( 
.A(n_9148),
.B(n_5732),
.Y(n_9347)
);

NAND2xp5_ASAP7_75t_L g9348 ( 
.A(n_9130),
.B(n_5736),
.Y(n_9348)
);

INVx1_ASAP7_75t_L g9349 ( 
.A(n_9166),
.Y(n_9349)
);

INVx1_ASAP7_75t_L g9350 ( 
.A(n_9134),
.Y(n_9350)
);

NAND2xp5_ASAP7_75t_SL g9351 ( 
.A(n_9130),
.B(n_9155),
.Y(n_9351)
);

OR2x2_ASAP7_75t_L g9352 ( 
.A(n_9160),
.B(n_5737),
.Y(n_9352)
);

NAND2xp5_ASAP7_75t_L g9353 ( 
.A(n_9239),
.B(n_5738),
.Y(n_9353)
);

AOI322xp5_ASAP7_75t_L g9354 ( 
.A1(n_9154),
.A2(n_4971),
.A3(n_4974),
.B1(n_4983),
.B2(n_4982),
.C1(n_4978),
.C2(n_5805),
.Y(n_9354)
);

INVx1_ASAP7_75t_L g9355 ( 
.A(n_9162),
.Y(n_9355)
);

NAND2xp5_ASAP7_75t_L g9356 ( 
.A(n_9152),
.B(n_5746),
.Y(n_9356)
);

AOI21xp5_ASAP7_75t_L g9357 ( 
.A1(n_9281),
.A2(n_5752),
.B(n_5746),
.Y(n_9357)
);

INVx1_ASAP7_75t_L g9358 ( 
.A(n_9231),
.Y(n_9358)
);

OAI22xp5_ASAP7_75t_L g9359 ( 
.A1(n_9172),
.A2(n_5756),
.B1(n_5757),
.B2(n_5752),
.Y(n_9359)
);

OR2x2_ASAP7_75t_L g9360 ( 
.A(n_9210),
.B(n_5757),
.Y(n_9360)
);

NOR2xp33_ASAP7_75t_L g9361 ( 
.A(n_9236),
.B(n_4971),
.Y(n_9361)
);

INVx1_ASAP7_75t_L g9362 ( 
.A(n_9164),
.Y(n_9362)
);

OAI22xp5_ASAP7_75t_L g9363 ( 
.A1(n_9173),
.A2(n_5761),
.B1(n_5765),
.B2(n_5760),
.Y(n_9363)
);

AND2x2_ASAP7_75t_L g9364 ( 
.A(n_9235),
.B(n_4879),
.Y(n_9364)
);

INVx2_ASAP7_75t_L g9365 ( 
.A(n_9136),
.Y(n_9365)
);

AOI21xp5_ASAP7_75t_L g9366 ( 
.A1(n_9216),
.A2(n_5769),
.B(n_5768),
.Y(n_9366)
);

INVx1_ASAP7_75t_L g9367 ( 
.A(n_9184),
.Y(n_9367)
);

INVx1_ASAP7_75t_L g9368 ( 
.A(n_9170),
.Y(n_9368)
);

OAI21xp5_ASAP7_75t_SL g9369 ( 
.A1(n_9137),
.A2(n_5673),
.B(n_5674),
.Y(n_9369)
);

AND2x4_ASAP7_75t_L g9370 ( 
.A(n_9181),
.B(n_4810),
.Y(n_9370)
);

INVx1_ASAP7_75t_L g9371 ( 
.A(n_9246),
.Y(n_9371)
);

AOI221xp5_ASAP7_75t_L g9372 ( 
.A1(n_9269),
.A2(n_4978),
.B1(n_4983),
.B2(n_4982),
.C(n_4974),
.Y(n_9372)
);

INVx2_ASAP7_75t_L g9373 ( 
.A(n_9259),
.Y(n_9373)
);

INVx1_ASAP7_75t_L g9374 ( 
.A(n_9178),
.Y(n_9374)
);

NAND2xp5_ASAP7_75t_L g9375 ( 
.A(n_9175),
.B(n_9275),
.Y(n_9375)
);

NOR2x1_ASAP7_75t_L g9376 ( 
.A(n_9201),
.B(n_5422),
.Y(n_9376)
);

INVx1_ASAP7_75t_L g9377 ( 
.A(n_9202),
.Y(n_9377)
);

INVxp67_ASAP7_75t_L g9378 ( 
.A(n_9234),
.Y(n_9378)
);

OAI21xp5_ASAP7_75t_L g9379 ( 
.A1(n_9158),
.A2(n_5798),
.B(n_5834),
.Y(n_9379)
);

AOI322xp5_ASAP7_75t_L g9380 ( 
.A1(n_9167),
.A2(n_4983),
.A3(n_5830),
.B1(n_5819),
.B2(n_5837),
.C1(n_5822),
.C2(n_5821),
.Y(n_9380)
);

INVx1_ASAP7_75t_L g9381 ( 
.A(n_9194),
.Y(n_9381)
);

OAI21xp33_ASAP7_75t_L g9382 ( 
.A1(n_9225),
.A2(n_5770),
.B(n_5769),
.Y(n_9382)
);

OAI31xp33_ASAP7_75t_L g9383 ( 
.A1(n_9151),
.A2(n_5821),
.A3(n_5822),
.B(n_5819),
.Y(n_9383)
);

INVx1_ASAP7_75t_L g9384 ( 
.A(n_9188),
.Y(n_9384)
);

AOI32xp33_ASAP7_75t_L g9385 ( 
.A1(n_9147),
.A2(n_5784),
.A3(n_4831),
.B1(n_5674),
.B2(n_4822),
.Y(n_9385)
);

NOR2x1_ASAP7_75t_L g9386 ( 
.A(n_9141),
.B(n_4882),
.Y(n_9386)
);

AOI21xp33_ASAP7_75t_L g9387 ( 
.A1(n_9254),
.A2(n_9227),
.B(n_9291),
.Y(n_9387)
);

AND2x2_ASAP7_75t_L g9388 ( 
.A(n_9303),
.B(n_4879),
.Y(n_9388)
);

AOI221x1_ASAP7_75t_L g9389 ( 
.A1(n_9171),
.A2(n_5968),
.B1(n_5969),
.B2(n_5965),
.C(n_5962),
.Y(n_9389)
);

OAI22xp5_ASAP7_75t_L g9390 ( 
.A1(n_9198),
.A2(n_5773),
.B1(n_5777),
.B2(n_5770),
.Y(n_9390)
);

AND2x2_ASAP7_75t_L g9391 ( 
.A(n_9196),
.B(n_4906),
.Y(n_9391)
);

INVx1_ASAP7_75t_L g9392 ( 
.A(n_9176),
.Y(n_9392)
);

INVx1_ASAP7_75t_L g9393 ( 
.A(n_9263),
.Y(n_9393)
);

INVx2_ASAP7_75t_L g9394 ( 
.A(n_9237),
.Y(n_9394)
);

NAND2xp33_ASAP7_75t_SL g9395 ( 
.A(n_9271),
.B(n_5773),
.Y(n_9395)
);

OAI21xp5_ASAP7_75t_SL g9396 ( 
.A1(n_9174),
.A2(n_5674),
.B(n_5020),
.Y(n_9396)
);

OAI22xp5_ASAP7_75t_L g9397 ( 
.A1(n_9251),
.A2(n_5788),
.B1(n_5800),
.B2(n_5777),
.Y(n_9397)
);

NAND2xp5_ASAP7_75t_L g9398 ( 
.A(n_9282),
.B(n_5788),
.Y(n_9398)
);

NAND2xp5_ASAP7_75t_L g9399 ( 
.A(n_9257),
.B(n_5800),
.Y(n_9399)
);

OAI32xp33_ASAP7_75t_L g9400 ( 
.A1(n_9203),
.A2(n_5825),
.A3(n_5826),
.B1(n_5815),
.B2(n_5807),
.Y(n_9400)
);

OA21x2_ASAP7_75t_L g9401 ( 
.A1(n_9292),
.A2(n_5815),
.B(n_5807),
.Y(n_9401)
);

OAI21xp33_ASAP7_75t_L g9402 ( 
.A1(n_9187),
.A2(n_5826),
.B(n_5825),
.Y(n_9402)
);

INVx1_ASAP7_75t_L g9403 ( 
.A(n_9214),
.Y(n_9403)
);

AND2x2_ASAP7_75t_L g9404 ( 
.A(n_9290),
.B(n_9250),
.Y(n_9404)
);

NOR2xp33_ASAP7_75t_L g9405 ( 
.A(n_9279),
.B(n_5827),
.Y(n_9405)
);

OR2x2_ASAP7_75t_L g9406 ( 
.A(n_9209),
.B(n_5827),
.Y(n_9406)
);

AOI21xp5_ASAP7_75t_L g9407 ( 
.A1(n_9221),
.A2(n_5833),
.B(n_5828),
.Y(n_9407)
);

INVx1_ASAP7_75t_L g9408 ( 
.A(n_9212),
.Y(n_9408)
);

INVx1_ASAP7_75t_L g9409 ( 
.A(n_9307),
.Y(n_9409)
);

INVx1_ASAP7_75t_L g9410 ( 
.A(n_9230),
.Y(n_9410)
);

AOI222xp33_ASAP7_75t_L g9411 ( 
.A1(n_9208),
.A2(n_9240),
.B1(n_9265),
.B2(n_9285),
.C1(n_9293),
.C2(n_9284),
.Y(n_9411)
);

OAI22x1_ASAP7_75t_L g9412 ( 
.A1(n_9283),
.A2(n_6009),
.B1(n_6010),
.B2(n_6008),
.Y(n_9412)
);

NOR2xp33_ASAP7_75t_L g9413 ( 
.A(n_9287),
.B(n_9295),
.Y(n_9413)
);

OAI21xp5_ASAP7_75t_SL g9414 ( 
.A1(n_9161),
.A2(n_5020),
.B(n_5312),
.Y(n_9414)
);

AOI22xp33_ASAP7_75t_L g9415 ( 
.A1(n_9260),
.A2(n_5999),
.B1(n_5252),
.B2(n_5070),
.Y(n_9415)
);

AND2x2_ASAP7_75t_L g9416 ( 
.A(n_9262),
.B(n_9211),
.Y(n_9416)
);

NAND2xp5_ASAP7_75t_L g9417 ( 
.A(n_9298),
.B(n_5828),
.Y(n_9417)
);

INVx1_ASAP7_75t_L g9418 ( 
.A(n_9252),
.Y(n_9418)
);

AOI221xp5_ASAP7_75t_L g9419 ( 
.A1(n_9157),
.A2(n_5860),
.B1(n_5863),
.B2(n_5837),
.C(n_5830),
.Y(n_9419)
);

INVx1_ASAP7_75t_L g9420 ( 
.A(n_9193),
.Y(n_9420)
);

OAI32xp33_ASAP7_75t_L g9421 ( 
.A1(n_9205),
.A2(n_5843),
.A3(n_5844),
.B1(n_5835),
.B2(n_5833),
.Y(n_9421)
);

NOR2x1_ASAP7_75t_L g9422 ( 
.A(n_9215),
.B(n_4882),
.Y(n_9422)
);

O2A1O1Ixp33_ASAP7_75t_L g9423 ( 
.A1(n_9218),
.A2(n_4689),
.B(n_5863),
.C(n_5860),
.Y(n_9423)
);

INVx1_ASAP7_75t_SL g9424 ( 
.A(n_9220),
.Y(n_9424)
);

INVx1_ASAP7_75t_L g9425 ( 
.A(n_9255),
.Y(n_9425)
);

INVx2_ASAP7_75t_L g9426 ( 
.A(n_9309),
.Y(n_9426)
);

INVx2_ASAP7_75t_L g9427 ( 
.A(n_9228),
.Y(n_9427)
);

AOI221xp5_ASAP7_75t_L g9428 ( 
.A1(n_9157),
.A2(n_5889),
.B1(n_5890),
.B2(n_5883),
.C(n_5874),
.Y(n_9428)
);

AOI21xp5_ASAP7_75t_L g9429 ( 
.A1(n_9286),
.A2(n_5843),
.B(n_5835),
.Y(n_9429)
);

INVx1_ASAP7_75t_L g9430 ( 
.A(n_9241),
.Y(n_9430)
);

OAI321xp33_ASAP7_75t_L g9431 ( 
.A1(n_9258),
.A2(n_5311),
.A3(n_4809),
.B1(n_5059),
.B2(n_4808),
.C(n_4726),
.Y(n_9431)
);

NAND2xp5_ASAP7_75t_L g9432 ( 
.A(n_9273),
.B(n_5844),
.Y(n_9432)
);

INVxp67_ASAP7_75t_SL g9433 ( 
.A(n_9249),
.Y(n_9433)
);

AOI221xp5_ASAP7_75t_L g9434 ( 
.A1(n_9266),
.A2(n_5889),
.B1(n_5890),
.B2(n_5883),
.C(n_5874),
.Y(n_9434)
);

AOI21xp5_ASAP7_75t_L g9435 ( 
.A1(n_9299),
.A2(n_5846),
.B(n_5845),
.Y(n_9435)
);

INVx1_ASAP7_75t_L g9436 ( 
.A(n_9244),
.Y(n_9436)
);

INVx1_ASAP7_75t_L g9437 ( 
.A(n_9289),
.Y(n_9437)
);

OAI211xp5_ASAP7_75t_L g9438 ( 
.A1(n_9268),
.A2(n_9293),
.B(n_9308),
.C(n_9182),
.Y(n_9438)
);

AOI221x1_ASAP7_75t_L g9439 ( 
.A1(n_9272),
.A2(n_5962),
.B1(n_5965),
.B2(n_5961),
.C(n_5959),
.Y(n_9439)
);

NOR2xp33_ASAP7_75t_L g9440 ( 
.A(n_9270),
.B(n_5845),
.Y(n_9440)
);

AND2x2_ASAP7_75t_L g9441 ( 
.A(n_9278),
.B(n_4906),
.Y(n_9441)
);

OAI32xp33_ASAP7_75t_L g9442 ( 
.A1(n_9285),
.A2(n_5852),
.A3(n_5854),
.B1(n_5851),
.B2(n_5846),
.Y(n_9442)
);

INVx2_ASAP7_75t_L g9443 ( 
.A(n_9191),
.Y(n_9443)
);

O2A1O1Ixp33_ASAP7_75t_L g9444 ( 
.A1(n_9238),
.A2(n_5896),
.B(n_5901),
.C(n_5900),
.Y(n_9444)
);

INVx1_ASAP7_75t_L g9445 ( 
.A(n_9288),
.Y(n_9445)
);

AOI32xp33_ASAP7_75t_L g9446 ( 
.A1(n_9199),
.A2(n_4831),
.A3(n_4822),
.B1(n_5969),
.B2(n_5968),
.Y(n_9446)
);

A2O1A1Ixp33_ASAP7_75t_L g9447 ( 
.A1(n_9180),
.A2(n_5902),
.B(n_5900),
.C(n_5901),
.Y(n_9447)
);

OAI22xp33_ASAP7_75t_L g9448 ( 
.A1(n_9186),
.A2(n_5896),
.B1(n_5906),
.B2(n_5902),
.Y(n_9448)
);

INVx2_ASAP7_75t_SL g9449 ( 
.A(n_9223),
.Y(n_9449)
);

INVx1_ASAP7_75t_L g9450 ( 
.A(n_9232),
.Y(n_9450)
);

AO21x1_ASAP7_75t_L g9451 ( 
.A1(n_9277),
.A2(n_5852),
.B(n_5851),
.Y(n_9451)
);

AOI32xp33_ASAP7_75t_L g9452 ( 
.A1(n_9294),
.A2(n_5954),
.A3(n_5957),
.B1(n_5953),
.B2(n_5950),
.Y(n_9452)
);

OAI221xp5_ASAP7_75t_L g9453 ( 
.A1(n_9245),
.A2(n_5422),
.B1(n_5574),
.B2(n_5449),
.C(n_4885),
.Y(n_9453)
);

INVx1_ASAP7_75t_L g9454 ( 
.A(n_9276),
.Y(n_9454)
);

AOI221xp5_ASAP7_75t_L g9455 ( 
.A1(n_9247),
.A2(n_5910),
.B1(n_5911),
.B2(n_5908),
.C(n_5906),
.Y(n_9455)
);

OAI221xp5_ASAP7_75t_SL g9456 ( 
.A1(n_9296),
.A2(n_5275),
.B1(n_5304),
.B2(n_5291),
.C(n_5287),
.Y(n_9456)
);

INVx1_ASAP7_75t_L g9457 ( 
.A(n_9191),
.Y(n_9457)
);

NAND2xp5_ASAP7_75t_L g9458 ( 
.A(n_9217),
.B(n_5854),
.Y(n_9458)
);

INVx1_ASAP7_75t_L g9459 ( 
.A(n_9192),
.Y(n_9459)
);

INVx1_ASAP7_75t_L g9460 ( 
.A(n_9338),
.Y(n_9460)
);

NAND2xp5_ASAP7_75t_L g9461 ( 
.A(n_9318),
.B(n_9327),
.Y(n_9461)
);

NAND2xp5_ASAP7_75t_L g9462 ( 
.A(n_9365),
.B(n_9233),
.Y(n_9462)
);

NAND2xp5_ASAP7_75t_L g9463 ( 
.A(n_9322),
.B(n_9189),
.Y(n_9463)
);

INVx2_ASAP7_75t_L g9464 ( 
.A(n_9312),
.Y(n_9464)
);

HB1xp67_ASAP7_75t_L g9465 ( 
.A(n_9351),
.Y(n_9465)
);

NAND2xp33_ASAP7_75t_L g9466 ( 
.A(n_9324),
.B(n_9300),
.Y(n_9466)
);

NAND2xp5_ASAP7_75t_L g9467 ( 
.A(n_9314),
.B(n_9274),
.Y(n_9467)
);

INVxp67_ASAP7_75t_L g9468 ( 
.A(n_9311),
.Y(n_9468)
);

NAND2xp5_ASAP7_75t_L g9469 ( 
.A(n_9424),
.B(n_9219),
.Y(n_9469)
);

AND2x4_ASAP7_75t_L g9470 ( 
.A(n_9381),
.B(n_9213),
.Y(n_9470)
);

AND2x2_ASAP7_75t_L g9471 ( 
.A(n_9329),
.B(n_9301),
.Y(n_9471)
);

AND2x2_ASAP7_75t_L g9472 ( 
.A(n_9404),
.B(n_9306),
.Y(n_9472)
);

NAND2xp5_ASAP7_75t_L g9473 ( 
.A(n_9433),
.B(n_9206),
.Y(n_9473)
);

INVx1_ASAP7_75t_L g9474 ( 
.A(n_9335),
.Y(n_9474)
);

NAND2x1_ASAP7_75t_L g9475 ( 
.A(n_9370),
.B(n_9320),
.Y(n_9475)
);

INVx2_ASAP7_75t_L g9476 ( 
.A(n_9401),
.Y(n_9476)
);

NAND2xp5_ASAP7_75t_L g9477 ( 
.A(n_9362),
.B(n_9261),
.Y(n_9477)
);

OAI31xp33_ASAP7_75t_SL g9478 ( 
.A1(n_9438),
.A2(n_9310),
.A3(n_9302),
.B(n_9297),
.Y(n_9478)
);

INVx1_ASAP7_75t_L g9479 ( 
.A(n_9328),
.Y(n_9479)
);

INVx1_ASAP7_75t_L g9480 ( 
.A(n_9457),
.Y(n_9480)
);

AND2x2_ASAP7_75t_L g9481 ( 
.A(n_9370),
.B(n_9177),
.Y(n_9481)
);

NAND2xp5_ASAP7_75t_L g9482 ( 
.A(n_9343),
.B(n_9256),
.Y(n_9482)
);

AND2x2_ASAP7_75t_L g9483 ( 
.A(n_9367),
.B(n_9305),
.Y(n_9483)
);

AND2x2_ASAP7_75t_L g9484 ( 
.A(n_9386),
.B(n_4906),
.Y(n_9484)
);

INVx1_ASAP7_75t_L g9485 ( 
.A(n_9443),
.Y(n_9485)
);

NOR2xp33_ASAP7_75t_L g9486 ( 
.A(n_9317),
.B(n_9280),
.Y(n_9486)
);

AND2x2_ASAP7_75t_L g9487 ( 
.A(n_9416),
.B(n_4906),
.Y(n_9487)
);

AND2x2_ASAP7_75t_L g9488 ( 
.A(n_9330),
.B(n_9336),
.Y(n_9488)
);

OR2x2_ASAP7_75t_L g9489 ( 
.A(n_9349),
.B(n_5856),
.Y(n_9489)
);

INVx2_ASAP7_75t_L g9490 ( 
.A(n_9401),
.Y(n_9490)
);

NAND2xp5_ASAP7_75t_L g9491 ( 
.A(n_9425),
.B(n_9420),
.Y(n_9491)
);

AOI22xp5_ASAP7_75t_L g9492 ( 
.A1(n_9331),
.A2(n_9207),
.B1(n_5910),
.B2(n_5911),
.Y(n_9492)
);

NOR3xp33_ASAP7_75t_L g9493 ( 
.A(n_9378),
.B(n_9242),
.C(n_4975),
.Y(n_9493)
);

INVx1_ASAP7_75t_L g9494 ( 
.A(n_9445),
.Y(n_9494)
);

OAI22xp5_ASAP7_75t_L g9495 ( 
.A1(n_9316),
.A2(n_5864),
.B1(n_5866),
.B2(n_5856),
.Y(n_9495)
);

OAI22xp5_ASAP7_75t_L g9496 ( 
.A1(n_9368),
.A2(n_5866),
.B1(n_5870),
.B2(n_5864),
.Y(n_9496)
);

OAI22xp5_ASAP7_75t_L g9497 ( 
.A1(n_9355),
.A2(n_5871),
.B1(n_5872),
.B2(n_5870),
.Y(n_9497)
);

AND2x2_ASAP7_75t_L g9498 ( 
.A(n_9364),
.B(n_4934),
.Y(n_9498)
);

INVx1_ASAP7_75t_L g9499 ( 
.A(n_9375),
.Y(n_9499)
);

AND2x2_ASAP7_75t_L g9500 ( 
.A(n_9345),
.B(n_9358),
.Y(n_9500)
);

INVx1_ASAP7_75t_L g9501 ( 
.A(n_9348),
.Y(n_9501)
);

AND2x2_ASAP7_75t_SL g9502 ( 
.A(n_9413),
.B(n_4885),
.Y(n_9502)
);

AND2x4_ASAP7_75t_L g9503 ( 
.A(n_9422),
.B(n_4882),
.Y(n_9503)
);

AND2x2_ASAP7_75t_L g9504 ( 
.A(n_9394),
.B(n_4934),
.Y(n_9504)
);

NOR2x1_ASAP7_75t_R g9505 ( 
.A(n_9377),
.B(n_5342),
.Y(n_9505)
);

INVx1_ASAP7_75t_L g9506 ( 
.A(n_9350),
.Y(n_9506)
);

NOR2xp33_ASAP7_75t_L g9507 ( 
.A(n_9396),
.B(n_5908),
.Y(n_9507)
);

CKINVDCx20_ASAP7_75t_R g9508 ( 
.A(n_9315),
.Y(n_9508)
);

INVx2_ASAP7_75t_L g9509 ( 
.A(n_9360),
.Y(n_9509)
);

NAND2xp5_ASAP7_75t_L g9510 ( 
.A(n_9313),
.B(n_5871),
.Y(n_9510)
);

INVx2_ASAP7_75t_L g9511 ( 
.A(n_9406),
.Y(n_9511)
);

NOR2x1_ASAP7_75t_L g9512 ( 
.A(n_9392),
.B(n_4894),
.Y(n_9512)
);

INVx1_ASAP7_75t_L g9513 ( 
.A(n_9371),
.Y(n_9513)
);

INVx1_ASAP7_75t_SL g9514 ( 
.A(n_9393),
.Y(n_9514)
);

NAND2xp5_ASAP7_75t_L g9515 ( 
.A(n_9409),
.B(n_5872),
.Y(n_9515)
);

NAND2xp5_ASAP7_75t_L g9516 ( 
.A(n_9403),
.B(n_5873),
.Y(n_9516)
);

INVx1_ASAP7_75t_L g9517 ( 
.A(n_9408),
.Y(n_9517)
);

AOI22xp33_ASAP7_75t_L g9518 ( 
.A1(n_9384),
.A2(n_5924),
.B1(n_5928),
.B2(n_5918),
.Y(n_9518)
);

OR2x2_ASAP7_75t_L g9519 ( 
.A(n_9410),
.B(n_5873),
.Y(n_9519)
);

NOR2xp33_ASAP7_75t_L g9520 ( 
.A(n_9341),
.B(n_5918),
.Y(n_9520)
);

AOI22xp33_ASAP7_75t_L g9521 ( 
.A1(n_9454),
.A2(n_5928),
.B1(n_5929),
.B2(n_5924),
.Y(n_9521)
);

NAND2xp5_ASAP7_75t_L g9522 ( 
.A(n_9426),
.B(n_5875),
.Y(n_9522)
);

OAI222xp33_ASAP7_75t_L g9523 ( 
.A1(n_9334),
.A2(n_5312),
.B1(n_5885),
.B2(n_5886),
.C1(n_5876),
.C2(n_5875),
.Y(n_9523)
);

NAND2x1_ASAP7_75t_L g9524 ( 
.A(n_9374),
.B(n_5180),
.Y(n_9524)
);

NAND2xp5_ASAP7_75t_L g9525 ( 
.A(n_9437),
.B(n_5876),
.Y(n_9525)
);

NAND2xp5_ASAP7_75t_L g9526 ( 
.A(n_9427),
.B(n_5885),
.Y(n_9526)
);

INVxp67_ASAP7_75t_SL g9527 ( 
.A(n_9373),
.Y(n_9527)
);

NAND2xp5_ASAP7_75t_L g9528 ( 
.A(n_9337),
.B(n_5886),
.Y(n_9528)
);

NAND2xp5_ASAP7_75t_L g9529 ( 
.A(n_9440),
.B(n_5887),
.Y(n_9529)
);

AND2x2_ASAP7_75t_L g9530 ( 
.A(n_9441),
.B(n_4934),
.Y(n_9530)
);

INVx1_ASAP7_75t_L g9531 ( 
.A(n_9376),
.Y(n_9531)
);

INVx2_ASAP7_75t_L g9532 ( 
.A(n_9352),
.Y(n_9532)
);

INVx1_ASAP7_75t_L g9533 ( 
.A(n_9376),
.Y(n_9533)
);

NOR2xp33_ASAP7_75t_SL g9534 ( 
.A(n_9387),
.B(n_4894),
.Y(n_9534)
);

AND2x4_ASAP7_75t_L g9535 ( 
.A(n_9430),
.B(n_4894),
.Y(n_9535)
);

NAND2xp5_ASAP7_75t_L g9536 ( 
.A(n_9369),
.B(n_5887),
.Y(n_9536)
);

NAND2xp5_ASAP7_75t_L g9537 ( 
.A(n_9418),
.B(n_5888),
.Y(n_9537)
);

INVx2_ASAP7_75t_SL g9538 ( 
.A(n_9347),
.Y(n_9538)
);

INVx1_ASAP7_75t_L g9539 ( 
.A(n_9353),
.Y(n_9539)
);

INVx1_ASAP7_75t_L g9540 ( 
.A(n_9432),
.Y(n_9540)
);

INVx2_ASAP7_75t_L g9541 ( 
.A(n_9388),
.Y(n_9541)
);

INVx1_ASAP7_75t_L g9542 ( 
.A(n_9398),
.Y(n_9542)
);

AND2x2_ASAP7_75t_L g9543 ( 
.A(n_9340),
.B(n_4934),
.Y(n_9543)
);

INVx1_ASAP7_75t_SL g9544 ( 
.A(n_9395),
.Y(n_9544)
);

OAI221xp5_ASAP7_75t_L g9545 ( 
.A1(n_9405),
.A2(n_5422),
.B1(n_5574),
.B2(n_5449),
.C(n_4885),
.Y(n_9545)
);

OAI221xp5_ASAP7_75t_L g9546 ( 
.A1(n_9383),
.A2(n_5449),
.B1(n_5574),
.B2(n_4885),
.C(n_4740),
.Y(n_9546)
);

INVx1_ASAP7_75t_SL g9547 ( 
.A(n_9356),
.Y(n_9547)
);

INVx1_ASAP7_75t_L g9548 ( 
.A(n_9399),
.Y(n_9548)
);

INVx1_ASAP7_75t_L g9549 ( 
.A(n_9417),
.Y(n_9549)
);

AND2x2_ASAP7_75t_L g9550 ( 
.A(n_9391),
.B(n_4996),
.Y(n_9550)
);

INVx1_ASAP7_75t_L g9551 ( 
.A(n_9319),
.Y(n_9551)
);

INVx1_ASAP7_75t_L g9552 ( 
.A(n_9459),
.Y(n_9552)
);

AND2x2_ASAP7_75t_L g9553 ( 
.A(n_9449),
.B(n_4996),
.Y(n_9553)
);

INVx1_ASAP7_75t_L g9554 ( 
.A(n_9436),
.Y(n_9554)
);

INVx1_ASAP7_75t_L g9555 ( 
.A(n_9450),
.Y(n_9555)
);

NOR2xp33_ASAP7_75t_L g9556 ( 
.A(n_9332),
.B(n_5929),
.Y(n_9556)
);

INVx1_ASAP7_75t_SL g9557 ( 
.A(n_9412),
.Y(n_9557)
);

NAND2xp5_ASAP7_75t_L g9558 ( 
.A(n_9357),
.B(n_5888),
.Y(n_9558)
);

AND2x4_ASAP7_75t_L g9559 ( 
.A(n_9389),
.B(n_4931),
.Y(n_9559)
);

NAND2xp5_ASAP7_75t_L g9560 ( 
.A(n_9435),
.B(n_5892),
.Y(n_9560)
);

NOR2xp33_ASAP7_75t_L g9561 ( 
.A(n_9361),
.B(n_5937),
.Y(n_9561)
);

INVx1_ASAP7_75t_L g9562 ( 
.A(n_9458),
.Y(n_9562)
);

NAND2xp5_ASAP7_75t_L g9563 ( 
.A(n_9429),
.B(n_5892),
.Y(n_9563)
);

HB1xp67_ASAP7_75t_L g9564 ( 
.A(n_9411),
.Y(n_9564)
);

INVx1_ASAP7_75t_L g9565 ( 
.A(n_9451),
.Y(n_9565)
);

NAND2xp5_ASAP7_75t_L g9566 ( 
.A(n_9321),
.B(n_5893),
.Y(n_9566)
);

NOR2xp33_ASAP7_75t_L g9567 ( 
.A(n_9442),
.B(n_5937),
.Y(n_9567)
);

NAND2xp5_ASAP7_75t_L g9568 ( 
.A(n_9402),
.B(n_9439),
.Y(n_9568)
);

OAI22xp5_ASAP7_75t_L g9569 ( 
.A1(n_9456),
.A2(n_5894),
.B1(n_5907),
.B2(n_5893),
.Y(n_9569)
);

INVx2_ASAP7_75t_L g9570 ( 
.A(n_9344),
.Y(n_9570)
);

NAND2xp5_ASAP7_75t_L g9571 ( 
.A(n_9366),
.B(n_5894),
.Y(n_9571)
);

NAND2xp5_ASAP7_75t_L g9572 ( 
.A(n_9452),
.B(n_5899),
.Y(n_9572)
);

AND2x2_ASAP7_75t_L g9573 ( 
.A(n_9414),
.B(n_4996),
.Y(n_9573)
);

INVx1_ASAP7_75t_L g9574 ( 
.A(n_9333),
.Y(n_9574)
);

NAND2xp5_ASAP7_75t_L g9575 ( 
.A(n_9385),
.B(n_5899),
.Y(n_9575)
);

INVx1_ASAP7_75t_L g9576 ( 
.A(n_9342),
.Y(n_9576)
);

INVx1_ASAP7_75t_L g9577 ( 
.A(n_9400),
.Y(n_9577)
);

NAND2xp5_ASAP7_75t_L g9578 ( 
.A(n_9407),
.B(n_5907),
.Y(n_9578)
);

OR2x2_ASAP7_75t_L g9579 ( 
.A(n_9323),
.B(n_5914),
.Y(n_9579)
);

AND2x2_ASAP7_75t_L g9580 ( 
.A(n_9382),
.B(n_4996),
.Y(n_9580)
);

OAI221xp5_ASAP7_75t_L g9581 ( 
.A1(n_9325),
.A2(n_5574),
.B1(n_5449),
.B2(n_4740),
.C(n_4807),
.Y(n_9581)
);

NOR4xp25_ASAP7_75t_L g9582 ( 
.A(n_9485),
.B(n_9431),
.C(n_9379),
.D(n_9423),
.Y(n_9582)
);

OAI21xp33_ASAP7_75t_SL g9583 ( 
.A1(n_9461),
.A2(n_9446),
.B(n_9363),
.Y(n_9583)
);

INVx1_ASAP7_75t_L g9584 ( 
.A(n_9465),
.Y(n_9584)
);

NAND5xp2_ASAP7_75t_L g9585 ( 
.A(n_9534),
.B(n_9380),
.C(n_9428),
.D(n_9419),
.E(n_9339),
.Y(n_9585)
);

AOI222xp33_ASAP7_75t_L g9586 ( 
.A1(n_9564),
.A2(n_9448),
.B1(n_9434),
.B2(n_9415),
.C1(n_9421),
.C2(n_9455),
.Y(n_9586)
);

NOR3xp33_ASAP7_75t_L g9587 ( 
.A(n_9475),
.B(n_9326),
.C(n_9359),
.Y(n_9587)
);

NOR3x1_ASAP7_75t_L g9588 ( 
.A(n_9527),
.B(n_9397),
.C(n_9390),
.Y(n_9588)
);

NOR3xp33_ASAP7_75t_L g9589 ( 
.A(n_9468),
.B(n_9474),
.C(n_9479),
.Y(n_9589)
);

INVx1_ASAP7_75t_L g9590 ( 
.A(n_9488),
.Y(n_9590)
);

AND2x2_ASAP7_75t_L g9591 ( 
.A(n_9464),
.B(n_9444),
.Y(n_9591)
);

INVx2_ASAP7_75t_L g9592 ( 
.A(n_9559),
.Y(n_9592)
);

AOI22xp5_ASAP7_75t_L g9593 ( 
.A1(n_9508),
.A2(n_9453),
.B1(n_9372),
.B2(n_9447),
.Y(n_9593)
);

INVx1_ASAP7_75t_L g9594 ( 
.A(n_9460),
.Y(n_9594)
);

OAI21xp5_ASAP7_75t_SL g9595 ( 
.A1(n_9514),
.A2(n_9354),
.B(n_9346),
.Y(n_9595)
);

AOI21xp5_ASAP7_75t_L g9596 ( 
.A1(n_9466),
.A2(n_5953),
.B(n_5930),
.Y(n_9596)
);

NAND2xp5_ASAP7_75t_SL g9597 ( 
.A(n_9470),
.B(n_5986),
.Y(n_9597)
);

NAND2xp5_ASAP7_75t_SL g9598 ( 
.A(n_9470),
.B(n_5987),
.Y(n_9598)
);

INVx2_ASAP7_75t_L g9599 ( 
.A(n_9559),
.Y(n_9599)
);

INVx1_ASAP7_75t_L g9600 ( 
.A(n_9476),
.Y(n_9600)
);

INVx1_ASAP7_75t_L g9601 ( 
.A(n_9490),
.Y(n_9601)
);

INVx2_ASAP7_75t_L g9602 ( 
.A(n_9472),
.Y(n_9602)
);

NAND3xp33_ASAP7_75t_L g9603 ( 
.A(n_9494),
.B(n_9576),
.C(n_9480),
.Y(n_9603)
);

AOI21xp5_ASAP7_75t_L g9604 ( 
.A1(n_9568),
.A2(n_5954),
.B(n_5930),
.Y(n_9604)
);

NAND2x1_ASAP7_75t_L g9605 ( 
.A(n_9503),
.B(n_5180),
.Y(n_9605)
);

NOR3x1_ASAP7_75t_L g9606 ( 
.A(n_9538),
.B(n_5915),
.C(n_5914),
.Y(n_9606)
);

NOR2xp33_ASAP7_75t_L g9607 ( 
.A(n_9544),
.B(n_5946),
.Y(n_9607)
);

NAND2xp5_ASAP7_75t_L g9608 ( 
.A(n_9512),
.B(n_5946),
.Y(n_9608)
);

NOR3xp33_ASAP7_75t_L g9609 ( 
.A(n_9491),
.B(n_9513),
.C(n_9499),
.Y(n_9609)
);

NAND2xp5_ASAP7_75t_SL g9610 ( 
.A(n_9503),
.B(n_5948),
.Y(n_9610)
);

INVx1_ASAP7_75t_L g9611 ( 
.A(n_9512),
.Y(n_9611)
);

NOR3x1_ASAP7_75t_L g9612 ( 
.A(n_9467),
.B(n_5916),
.C(n_5915),
.Y(n_9612)
);

AND2x2_ASAP7_75t_L g9613 ( 
.A(n_9487),
.B(n_5191),
.Y(n_9613)
);

INVx1_ASAP7_75t_L g9614 ( 
.A(n_9531),
.Y(n_9614)
);

INVx1_ASAP7_75t_L g9615 ( 
.A(n_9533),
.Y(n_9615)
);

NOR2xp33_ASAP7_75t_L g9616 ( 
.A(n_9557),
.B(n_5949),
.Y(n_9616)
);

NAND4xp25_ASAP7_75t_L g9617 ( 
.A(n_9462),
.B(n_4972),
.C(n_4931),
.D(n_5116),
.Y(n_9617)
);

NAND4xp25_ASAP7_75t_L g9618 ( 
.A(n_9555),
.B(n_4972),
.C(n_4931),
.D(n_5335),
.Y(n_9618)
);

NAND2xp5_ASAP7_75t_L g9619 ( 
.A(n_9547),
.B(n_5949),
.Y(n_9619)
);

INVx1_ASAP7_75t_L g9620 ( 
.A(n_9552),
.Y(n_9620)
);

OA22x2_ASAP7_75t_L g9621 ( 
.A1(n_9524),
.A2(n_5925),
.B1(n_5926),
.B2(n_5916),
.Y(n_9621)
);

A2O1A1Ixp33_ASAP7_75t_SL g9622 ( 
.A1(n_9517),
.A2(n_9506),
.B(n_9554),
.C(n_9532),
.Y(n_9622)
);

AOI221xp5_ASAP7_75t_SL g9623 ( 
.A1(n_9565),
.A2(n_5935),
.B1(n_5942),
.B2(n_5926),
.C(n_5925),
.Y(n_9623)
);

NOR2xp33_ASAP7_75t_L g9624 ( 
.A(n_9509),
.B(n_5951),
.Y(n_9624)
);

INVx1_ASAP7_75t_SL g9625 ( 
.A(n_9500),
.Y(n_9625)
);

NAND4xp25_ASAP7_75t_L g9626 ( 
.A(n_9469),
.B(n_4972),
.C(n_5335),
.D(n_5088),
.Y(n_9626)
);

OAI21xp33_ASAP7_75t_SL g9627 ( 
.A1(n_9484),
.A2(n_5942),
.B(n_5935),
.Y(n_9627)
);

INVx1_ASAP7_75t_L g9628 ( 
.A(n_9463),
.Y(n_9628)
);

INVx1_ASAP7_75t_L g9629 ( 
.A(n_9471),
.Y(n_9629)
);

AND2x2_ASAP7_75t_L g9630 ( 
.A(n_9553),
.B(n_5191),
.Y(n_9630)
);

NOR2xp33_ASAP7_75t_SL g9631 ( 
.A(n_9541),
.B(n_5274),
.Y(n_9631)
);

NOR2xp33_ASAP7_75t_L g9632 ( 
.A(n_9511),
.B(n_5951),
.Y(n_9632)
);

NAND2xp5_ASAP7_75t_L g9633 ( 
.A(n_9481),
.B(n_5956),
.Y(n_9633)
);

NAND2x1_ASAP7_75t_L g9634 ( 
.A(n_9535),
.B(n_5180),
.Y(n_9634)
);

NAND4xp25_ASAP7_75t_L g9635 ( 
.A(n_9477),
.B(n_5078),
.C(n_5213),
.D(n_4975),
.Y(n_9635)
);

AOI22x1_ASAP7_75t_L g9636 ( 
.A1(n_9577),
.A2(n_5313),
.B1(n_5950),
.B2(n_5948),
.Y(n_9636)
);

NOR3x1_ASAP7_75t_L g9637 ( 
.A(n_9482),
.B(n_5959),
.C(n_5957),
.Y(n_9637)
);

NAND2xp5_ASAP7_75t_L g9638 ( 
.A(n_9483),
.B(n_5956),
.Y(n_9638)
);

NAND4xp25_ASAP7_75t_L g9639 ( 
.A(n_9486),
.B(n_4663),
.C(n_5329),
.D(n_5317),
.Y(n_9639)
);

OAI21xp5_ASAP7_75t_SL g9640 ( 
.A1(n_9478),
.A2(n_5307),
.B(n_5237),
.Y(n_9640)
);

NOR2x1_ASAP7_75t_L g9641 ( 
.A(n_9551),
.B(n_5961),
.Y(n_9641)
);

AOI21xp5_ASAP7_75t_L g9642 ( 
.A1(n_9510),
.A2(n_5972),
.B(n_5970),
.Y(n_9642)
);

NAND2xp5_ASAP7_75t_SL g9643 ( 
.A(n_9535),
.B(n_5987),
.Y(n_9643)
);

NOR4xp25_ASAP7_75t_L g9644 ( 
.A(n_9473),
.B(n_5970),
.C(n_6008),
.D(n_5979),
.Y(n_9644)
);

AOI221xp5_ASAP7_75t_L g9645 ( 
.A1(n_9574),
.A2(n_5966),
.B1(n_4788),
.B2(n_4702),
.C(n_4703),
.Y(n_9645)
);

INVx1_ASAP7_75t_L g9646 ( 
.A(n_9519),
.Y(n_9646)
);

OAI321xp33_ASAP7_75t_L g9647 ( 
.A1(n_9570),
.A2(n_4726),
.A3(n_4744),
.B1(n_4711),
.B2(n_5966),
.C(n_4771),
.Y(n_9647)
);

AND2x2_ASAP7_75t_L g9648 ( 
.A(n_9504),
.B(n_5244),
.Y(n_9648)
);

OAI21xp5_ASAP7_75t_L g9649 ( 
.A1(n_9562),
.A2(n_5056),
.B(n_4740),
.Y(n_9649)
);

AOI21xp5_ASAP7_75t_L g9650 ( 
.A1(n_9542),
.A2(n_4740),
.B(n_4907),
.Y(n_9650)
);

OAI21xp33_ASAP7_75t_L g9651 ( 
.A1(n_9548),
.A2(n_5220),
.B(n_5219),
.Y(n_9651)
);

AO21x1_ASAP7_75t_L g9652 ( 
.A1(n_9549),
.A2(n_5357),
.B(n_5355),
.Y(n_9652)
);

AOI22xp5_ASAP7_75t_L g9653 ( 
.A1(n_9539),
.A2(n_4780),
.B1(n_4833),
.B2(n_4807),
.Y(n_9653)
);

NAND3xp33_ASAP7_75t_SL g9654 ( 
.A(n_9501),
.B(n_4726),
.C(n_4711),
.Y(n_9654)
);

NAND4xp25_ASAP7_75t_L g9655 ( 
.A(n_9493),
.B(n_4663),
.C(n_4939),
.D(n_5119),
.Y(n_9655)
);

NAND2xp5_ASAP7_75t_L g9656 ( 
.A(n_9492),
.B(n_4993),
.Y(n_9656)
);

INVxp67_ASAP7_75t_L g9657 ( 
.A(n_9540),
.Y(n_9657)
);

AOI221xp5_ASAP7_75t_L g9658 ( 
.A1(n_9567),
.A2(n_4702),
.B1(n_4703),
.B2(n_5019),
.C(n_4993),
.Y(n_9658)
);

AOI21xp33_ASAP7_75t_SL g9659 ( 
.A1(n_9489),
.A2(n_5347),
.B(n_4744),
.Y(n_9659)
);

INVx1_ASAP7_75t_L g9660 ( 
.A(n_9558),
.Y(n_9660)
);

INVx1_ASAP7_75t_L g9661 ( 
.A(n_9563),
.Y(n_9661)
);

NAND2xp5_ASAP7_75t_L g9662 ( 
.A(n_9520),
.B(n_4993),
.Y(n_9662)
);

NOR3xp33_ASAP7_75t_L g9663 ( 
.A(n_9505),
.B(n_9526),
.C(n_9516),
.Y(n_9663)
);

NAND3xp33_ASAP7_75t_L g9664 ( 
.A(n_9507),
.B(n_4703),
.C(n_4702),
.Y(n_9664)
);

AOI211xp5_ASAP7_75t_L g9665 ( 
.A1(n_9505),
.A2(n_5347),
.B(n_5047),
.C(n_4860),
.Y(n_9665)
);

NAND2xp5_ASAP7_75t_L g9666 ( 
.A(n_9556),
.B(n_4993),
.Y(n_9666)
);

OA22x2_ASAP7_75t_L g9667 ( 
.A1(n_9536),
.A2(n_9575),
.B1(n_9528),
.B2(n_9522),
.Y(n_9667)
);

NAND4xp25_ASAP7_75t_L g9668 ( 
.A(n_9525),
.B(n_5187),
.C(n_5058),
.D(n_4834),
.Y(n_9668)
);

AOI22xp5_ASAP7_75t_SL g9669 ( 
.A1(n_9515),
.A2(n_5263),
.B1(n_4180),
.B2(n_4225),
.Y(n_9669)
);

NOR2xp33_ASAP7_75t_L g9670 ( 
.A(n_9537),
.B(n_3842),
.Y(n_9670)
);

NAND2xp5_ASAP7_75t_L g9671 ( 
.A(n_9529),
.B(n_9560),
.Y(n_9671)
);

NOR3xp33_ASAP7_75t_L g9672 ( 
.A(n_9569),
.B(n_4393),
.C(n_4619),
.Y(n_9672)
);

NAND3xp33_ASAP7_75t_L g9673 ( 
.A(n_9561),
.B(n_5182),
.C(n_5171),
.Y(n_9673)
);

NAND3xp33_ASAP7_75t_L g9674 ( 
.A(n_9566),
.B(n_5182),
.C(n_5171),
.Y(n_9674)
);

NAND2xp5_ASAP7_75t_L g9675 ( 
.A(n_9571),
.B(n_5019),
.Y(n_9675)
);

AOI21xp5_ASAP7_75t_SL g9676 ( 
.A1(n_9578),
.A2(n_4442),
.B(n_5244),
.Y(n_9676)
);

NAND4xp75_ASAP7_75t_L g9677 ( 
.A(n_9573),
.B(n_4904),
.C(n_4427),
.D(n_4461),
.Y(n_9677)
);

NAND4xp25_ASAP7_75t_L g9678 ( 
.A(n_9572),
.B(n_4751),
.C(n_5210),
.D(n_5202),
.Y(n_9678)
);

NOR2x1_ASAP7_75t_L g9679 ( 
.A(n_9579),
.B(n_5263),
.Y(n_9679)
);

NAND4xp25_ASAP7_75t_L g9680 ( 
.A(n_9580),
.B(n_5338),
.C(n_4963),
.D(n_4940),
.Y(n_9680)
);

NAND2xp5_ASAP7_75t_L g9681 ( 
.A(n_9495),
.B(n_5019),
.Y(n_9681)
);

AOI21xp5_ASAP7_75t_L g9682 ( 
.A1(n_9523),
.A2(n_4907),
.B(n_5220),
.Y(n_9682)
);

INVx1_ASAP7_75t_L g9683 ( 
.A(n_9496),
.Y(n_9683)
);

AND2x2_ASAP7_75t_L g9684 ( 
.A(n_9498),
.B(n_5283),
.Y(n_9684)
);

AOI211xp5_ASAP7_75t_L g9685 ( 
.A1(n_9581),
.A2(n_4860),
.B(n_4868),
.C(n_4859),
.Y(n_9685)
);

AOI211xp5_ASAP7_75t_L g9686 ( 
.A1(n_9545),
.A2(n_4860),
.B(n_4868),
.C(n_4859),
.Y(n_9686)
);

NAND2xp5_ASAP7_75t_L g9687 ( 
.A(n_9502),
.B(n_5019),
.Y(n_9687)
);

NAND2xp5_ASAP7_75t_L g9688 ( 
.A(n_9543),
.B(n_5070),
.Y(n_9688)
);

BUFx2_ASAP7_75t_L g9689 ( 
.A(n_9550),
.Y(n_9689)
);

AOI221xp5_ASAP7_75t_L g9690 ( 
.A1(n_9546),
.A2(n_3891),
.B1(n_3874),
.B2(n_5226),
.C(n_5222),
.Y(n_9690)
);

INVx1_ASAP7_75t_L g9691 ( 
.A(n_9497),
.Y(n_9691)
);

NAND5xp2_ASAP7_75t_L g9692 ( 
.A(n_9530),
.B(n_4711),
.C(n_4744),
.D(n_5208),
.E(n_4181),
.Y(n_9692)
);

AND2x2_ASAP7_75t_L g9693 ( 
.A(n_9584),
.B(n_9521),
.Y(n_9693)
);

NAND2xp5_ASAP7_75t_SL g9694 ( 
.A(n_9602),
.B(n_9518),
.Y(n_9694)
);

INVx1_ASAP7_75t_L g9695 ( 
.A(n_9592),
.Y(n_9695)
);

AND2x2_ASAP7_75t_L g9696 ( 
.A(n_9625),
.B(n_5283),
.Y(n_9696)
);

NAND2xp5_ASAP7_75t_L g9697 ( 
.A(n_9599),
.B(n_9590),
.Y(n_9697)
);

OR2x2_ASAP7_75t_L g9698 ( 
.A(n_9582),
.B(n_4501),
.Y(n_9698)
);

AOI221xp5_ASAP7_75t_L g9699 ( 
.A1(n_9603),
.A2(n_3891),
.B1(n_3874),
.B2(n_5343),
.C(n_5337),
.Y(n_9699)
);

INVx1_ASAP7_75t_L g9700 ( 
.A(n_9620),
.Y(n_9700)
);

AND2x2_ASAP7_75t_L g9701 ( 
.A(n_9609),
.B(n_5293),
.Y(n_9701)
);

INVx1_ASAP7_75t_L g9702 ( 
.A(n_9591),
.Y(n_9702)
);

INVx1_ASAP7_75t_L g9703 ( 
.A(n_9689),
.Y(n_9703)
);

NAND2xp5_ASAP7_75t_L g9704 ( 
.A(n_9629),
.B(n_5252),
.Y(n_9704)
);

OAI321xp33_ASAP7_75t_L g9705 ( 
.A1(n_9593),
.A2(n_4839),
.A3(n_4976),
.B1(n_4181),
.B2(n_4168),
.C(n_5237),
.Y(n_9705)
);

NOR3xp33_ASAP7_75t_L g9706 ( 
.A(n_9589),
.B(n_9594),
.C(n_9614),
.Y(n_9706)
);

NOR2xp33_ASAP7_75t_L g9707 ( 
.A(n_9595),
.B(n_4780),
.Y(n_9707)
);

HB1xp67_ASAP7_75t_L g9708 ( 
.A(n_9600),
.Y(n_9708)
);

NAND4xp25_ASAP7_75t_L g9709 ( 
.A(n_9622),
.B(n_4813),
.C(n_5015),
.D(n_4815),
.Y(n_9709)
);

AOI211xp5_ASAP7_75t_L g9710 ( 
.A1(n_9601),
.A2(n_4860),
.B(n_4868),
.C(n_4859),
.Y(n_9710)
);

AOI211xp5_ASAP7_75t_L g9711 ( 
.A1(n_9587),
.A2(n_4860),
.B(n_4868),
.C(n_4859),
.Y(n_9711)
);

NAND2xp5_ASAP7_75t_SL g9712 ( 
.A(n_9583),
.B(n_4868),
.Y(n_9712)
);

NOR3xp33_ASAP7_75t_L g9713 ( 
.A(n_9615),
.B(n_9657),
.C(n_9628),
.Y(n_9713)
);

NOR3xp33_ASAP7_75t_L g9714 ( 
.A(n_9611),
.B(n_4112),
.C(n_4086),
.Y(n_9714)
);

INVx1_ASAP7_75t_L g9715 ( 
.A(n_9608),
.Y(n_9715)
);

INVx1_ASAP7_75t_L g9716 ( 
.A(n_9652),
.Y(n_9716)
);

NAND2xp5_ASAP7_75t_L g9717 ( 
.A(n_9646),
.B(n_5314),
.Y(n_9717)
);

AOI21xp5_ASAP7_75t_L g9718 ( 
.A1(n_9671),
.A2(n_4180),
.B(n_4907),
.Y(n_9718)
);

NOR3xp33_ASAP7_75t_L g9719 ( 
.A(n_9663),
.B(n_4125),
.C(n_5013),
.Y(n_9719)
);

INVx1_ASAP7_75t_SL g9720 ( 
.A(n_9660),
.Y(n_9720)
);

O2A1O1Ixp33_ASAP7_75t_L g9721 ( 
.A1(n_9661),
.A2(n_4530),
.B(n_4168),
.C(n_5237),
.Y(n_9721)
);

CKINVDCx20_ASAP7_75t_R g9722 ( 
.A(n_9683),
.Y(n_9722)
);

INVx1_ASAP7_75t_L g9723 ( 
.A(n_9597),
.Y(n_9723)
);

NAND3xp33_ASAP7_75t_L g9724 ( 
.A(n_9691),
.B(n_5182),
.C(n_5171),
.Y(n_9724)
);

NOR2x1_ASAP7_75t_L g9725 ( 
.A(n_9641),
.B(n_9585),
.Y(n_9725)
);

NAND2xp5_ASAP7_75t_SL g9726 ( 
.A(n_9631),
.B(n_5037),
.Y(n_9726)
);

OR2x2_ASAP7_75t_L g9727 ( 
.A(n_9626),
.B(n_4501),
.Y(n_9727)
);

NAND5xp2_ASAP7_75t_L g9728 ( 
.A(n_9586),
.B(n_5208),
.C(n_5307),
.D(n_4847),
.E(n_4855),
.Y(n_9728)
);

AND2x2_ASAP7_75t_L g9729 ( 
.A(n_9630),
.B(n_5293),
.Y(n_9729)
);

O2A1O1Ixp5_ASAP7_75t_L g9730 ( 
.A1(n_9598),
.A2(n_5226),
.B(n_5227),
.C(n_5222),
.Y(n_9730)
);

NOR2xp33_ASAP7_75t_L g9731 ( 
.A(n_9638),
.B(n_4780),
.Y(n_9731)
);

NOR2xp33_ASAP7_75t_L g9732 ( 
.A(n_9633),
.B(n_4780),
.Y(n_9732)
);

OAI21xp5_ASAP7_75t_L g9733 ( 
.A1(n_9616),
.A2(n_4198),
.B(n_4508),
.Y(n_9733)
);

XOR2xp5_ASAP7_75t_L g9734 ( 
.A(n_9667),
.B(n_4741),
.Y(n_9734)
);

INVx1_ASAP7_75t_L g9735 ( 
.A(n_9588),
.Y(n_9735)
);

NOR2xp33_ASAP7_75t_L g9736 ( 
.A(n_9619),
.B(n_4780),
.Y(n_9736)
);

NOR2xp33_ASAP7_75t_L g9737 ( 
.A(n_9607),
.B(n_4807),
.Y(n_9737)
);

AOI332xp33_ASAP7_75t_L g9738 ( 
.A1(n_9636),
.A2(n_5236),
.A3(n_5230),
.B1(n_5264),
.B2(n_5253),
.B3(n_5270),
.C1(n_5234),
.C2(n_5227),
.Y(n_9738)
);

INVx1_ASAP7_75t_L g9739 ( 
.A(n_9612),
.Y(n_9739)
);

NAND3xp33_ASAP7_75t_L g9740 ( 
.A(n_9624),
.B(n_5188),
.C(n_5184),
.Y(n_9740)
);

INVx1_ASAP7_75t_L g9741 ( 
.A(n_9637),
.Y(n_9741)
);

OR2x2_ASAP7_75t_L g9742 ( 
.A(n_9639),
.B(n_4508),
.Y(n_9742)
);

OAI21xp5_ASAP7_75t_L g9743 ( 
.A1(n_9604),
.A2(n_4198),
.B(n_4515),
.Y(n_9743)
);

INVx1_ASAP7_75t_L g9744 ( 
.A(n_9632),
.Y(n_9744)
);

NOR3xp33_ASAP7_75t_L g9745 ( 
.A(n_9605),
.B(n_5013),
.C(n_4427),
.Y(n_9745)
);

INVx1_ASAP7_75t_L g9746 ( 
.A(n_9606),
.Y(n_9746)
);

AOI211xp5_ASAP7_75t_L g9747 ( 
.A1(n_9640),
.A2(n_4859),
.B(n_4868),
.C(n_4860),
.Y(n_9747)
);

AND2x2_ASAP7_75t_L g9748 ( 
.A(n_9648),
.B(n_5297),
.Y(n_9748)
);

INVx1_ASAP7_75t_L g9749 ( 
.A(n_9610),
.Y(n_9749)
);

INVx1_ASAP7_75t_L g9750 ( 
.A(n_9621),
.Y(n_9750)
);

NAND2xp5_ASAP7_75t_SL g9751 ( 
.A(n_9679),
.B(n_5251),
.Y(n_9751)
);

INVx1_ASAP7_75t_L g9752 ( 
.A(n_9643),
.Y(n_9752)
);

NOR3xp33_ASAP7_75t_L g9753 ( 
.A(n_9670),
.B(n_5013),
.C(n_4590),
.Y(n_9753)
);

NAND4xp25_ASAP7_75t_L g9754 ( 
.A(n_9665),
.B(n_4757),
.C(n_4461),
.D(n_4446),
.Y(n_9754)
);

NAND2xp5_ASAP7_75t_L g9755 ( 
.A(n_9644),
.B(n_5209),
.Y(n_9755)
);

NOR2xp33_ASAP7_75t_L g9756 ( 
.A(n_9627),
.B(n_4807),
.Y(n_9756)
);

OAI22xp5_ASAP7_75t_L g9757 ( 
.A1(n_9653),
.A2(n_4807),
.B1(n_4953),
.B2(n_4833),
.Y(n_9757)
);

NAND2xp5_ASAP7_75t_L g9758 ( 
.A(n_9623),
.B(n_5216),
.Y(n_9758)
);

NOR3xp33_ASAP7_75t_L g9759 ( 
.A(n_9656),
.B(n_4589),
.C(n_4515),
.Y(n_9759)
);

AND2x2_ASAP7_75t_L g9760 ( 
.A(n_9613),
.B(n_5297),
.Y(n_9760)
);

NAND3xp33_ASAP7_75t_L g9761 ( 
.A(n_9686),
.B(n_5188),
.C(n_5184),
.Y(n_9761)
);

NOR3xp33_ASAP7_75t_L g9762 ( 
.A(n_9634),
.B(n_4762),
.C(n_4749),
.Y(n_9762)
);

NOR2xp33_ASAP7_75t_L g9763 ( 
.A(n_9675),
.B(n_4833),
.Y(n_9763)
);

NOR3xp33_ASAP7_75t_L g9764 ( 
.A(n_9666),
.B(n_4762),
.C(n_4749),
.Y(n_9764)
);

NOR4xp25_ASAP7_75t_SL g9765 ( 
.A(n_9651),
.B(n_4256),
.C(n_4336),
.D(n_4186),
.Y(n_9765)
);

AND2x2_ASAP7_75t_L g9766 ( 
.A(n_9684),
.B(n_5303),
.Y(n_9766)
);

NAND3xp33_ASAP7_75t_SL g9767 ( 
.A(n_9685),
.B(n_4756),
.C(n_4742),
.Y(n_9767)
);

AOI22xp5_ASAP7_75t_L g9768 ( 
.A1(n_9688),
.A2(n_4953),
.B1(n_4833),
.B2(n_5342),
.Y(n_9768)
);

NAND2xp5_ASAP7_75t_L g9769 ( 
.A(n_9642),
.B(n_5207),
.Y(n_9769)
);

NAND2xp5_ASAP7_75t_L g9770 ( 
.A(n_9596),
.B(n_5207),
.Y(n_9770)
);

O2A1O1Ixp33_ASAP7_75t_L g9771 ( 
.A1(n_9681),
.A2(n_5307),
.B(n_4334),
.C(n_4225),
.Y(n_9771)
);

NOR2xp33_ASAP7_75t_L g9772 ( 
.A(n_9662),
.B(n_4833),
.Y(n_9772)
);

NAND2xp5_ASAP7_75t_L g9773 ( 
.A(n_9651),
.B(n_5209),
.Y(n_9773)
);

NAND2xp5_ASAP7_75t_SL g9774 ( 
.A(n_9658),
.B(n_4859),
.Y(n_9774)
);

NOR2xp33_ASAP7_75t_L g9775 ( 
.A(n_9664),
.B(n_4953),
.Y(n_9775)
);

NOR4xp25_ASAP7_75t_L g9776 ( 
.A(n_9687),
.B(n_5367),
.C(n_5365),
.D(n_5234),
.Y(n_9776)
);

NAND3xp33_ASAP7_75t_SL g9777 ( 
.A(n_9672),
.B(n_4819),
.C(n_5208),
.Y(n_9777)
);

AND2x2_ASAP7_75t_L g9778 ( 
.A(n_9676),
.B(n_5303),
.Y(n_9778)
);

OAI21xp5_ASAP7_75t_L g9779 ( 
.A1(n_9650),
.A2(n_4198),
.B(n_4187),
.Y(n_9779)
);

AND2x2_ASAP7_75t_L g9780 ( 
.A(n_9682),
.B(n_5316),
.Y(n_9780)
);

OAI221xp5_ASAP7_75t_SL g9781 ( 
.A1(n_9690),
.A2(n_9618),
.B1(n_9617),
.B2(n_9645),
.C(n_9635),
.Y(n_9781)
);

NAND3xp33_ASAP7_75t_L g9782 ( 
.A(n_9674),
.B(n_5188),
.C(n_5184),
.Y(n_9782)
);

OR2x2_ASAP7_75t_L g9783 ( 
.A(n_9655),
.B(n_4634),
.Y(n_9783)
);

AND2x2_ASAP7_75t_L g9784 ( 
.A(n_9659),
.B(n_5316),
.Y(n_9784)
);

NAND2xp5_ASAP7_75t_L g9785 ( 
.A(n_9649),
.B(n_5259),
.Y(n_9785)
);

NAND4xp75_ASAP7_75t_L g9786 ( 
.A(n_9677),
.B(n_9654),
.C(n_9647),
.D(n_9678),
.Y(n_9786)
);

NAND3xp33_ASAP7_75t_L g9787 ( 
.A(n_9673),
.B(n_5209),
.C(n_5207),
.Y(n_9787)
);

NOR2xp33_ASAP7_75t_L g9788 ( 
.A(n_9668),
.B(n_4953),
.Y(n_9788)
);

AOI22xp5_ASAP7_75t_L g9789 ( 
.A1(n_9680),
.A2(n_4953),
.B1(n_5342),
.B2(n_4198),
.Y(n_9789)
);

OR2x2_ASAP7_75t_L g9790 ( 
.A(n_9692),
.B(n_9669),
.Y(n_9790)
);

INVx1_ASAP7_75t_SL g9791 ( 
.A(n_9669),
.Y(n_9791)
);

NAND3xp33_ASAP7_75t_L g9792 ( 
.A(n_9584),
.B(n_5218),
.C(n_5216),
.Y(n_9792)
);

INVx1_ASAP7_75t_L g9793 ( 
.A(n_9584),
.Y(n_9793)
);

NAND3xp33_ASAP7_75t_L g9794 ( 
.A(n_9584),
.B(n_5218),
.C(n_5216),
.Y(n_9794)
);

NAND5xp2_ASAP7_75t_L g9795 ( 
.A(n_9584),
.B(n_4854),
.C(n_4855),
.D(n_4847),
.E(n_4827),
.Y(n_9795)
);

AOI221xp5_ASAP7_75t_L g9796 ( 
.A1(n_9582),
.A2(n_3891),
.B1(n_3874),
.B2(n_5357),
.C(n_5355),
.Y(n_9796)
);

INVx2_ASAP7_75t_L g9797 ( 
.A(n_9602),
.Y(n_9797)
);

NAND2xp33_ASAP7_75t_SL g9798 ( 
.A(n_9584),
.B(n_4869),
.Y(n_9798)
);

INVx1_ASAP7_75t_L g9799 ( 
.A(n_9584),
.Y(n_9799)
);

INVx1_ASAP7_75t_L g9800 ( 
.A(n_9584),
.Y(n_9800)
);

OAI21xp33_ASAP7_75t_L g9801 ( 
.A1(n_9584),
.A2(n_3755),
.B(n_3754),
.Y(n_9801)
);

NAND2xp5_ASAP7_75t_L g9802 ( 
.A(n_9592),
.B(n_5232),
.Y(n_9802)
);

AOI211xp5_ASAP7_75t_L g9803 ( 
.A1(n_9625),
.A2(n_4961),
.B(n_5037),
.C(n_4869),
.Y(n_9803)
);

OR2x2_ASAP7_75t_L g9804 ( 
.A(n_9698),
.B(n_4634),
.Y(n_9804)
);

AOI21xp5_ASAP7_75t_L g9805 ( 
.A1(n_9708),
.A2(n_4198),
.B(n_4907),
.Y(n_9805)
);

OAI22xp5_ASAP7_75t_L g9806 ( 
.A1(n_9703),
.A2(n_5289),
.B1(n_5180),
.B2(n_4961),
.Y(n_9806)
);

XNOR2x1_ASAP7_75t_L g9807 ( 
.A(n_9725),
.B(n_9797),
.Y(n_9807)
);

XOR2xp5_ASAP7_75t_L g9808 ( 
.A(n_9722),
.B(n_4817),
.Y(n_9808)
);

INVx1_ASAP7_75t_SL g9809 ( 
.A(n_9697),
.Y(n_9809)
);

INVx1_ASAP7_75t_L g9810 ( 
.A(n_9695),
.Y(n_9810)
);

XNOR2xp5_ASAP7_75t_L g9811 ( 
.A(n_9734),
.B(n_4827),
.Y(n_9811)
);

AND2x2_ASAP7_75t_L g9812 ( 
.A(n_9701),
.B(n_5073),
.Y(n_9812)
);

AOI22xp5_ASAP7_75t_L g9813 ( 
.A1(n_9700),
.A2(n_5289),
.B1(n_4187),
.B2(n_4961),
.Y(n_9813)
);

NOR2xp33_ASAP7_75t_L g9814 ( 
.A(n_9702),
.B(n_3690),
.Y(n_9814)
);

INVx1_ASAP7_75t_L g9815 ( 
.A(n_9793),
.Y(n_9815)
);

NAND2x1p5_ASAP7_75t_L g9816 ( 
.A(n_9799),
.B(n_3635),
.Y(n_9816)
);

XNOR2x1_ASAP7_75t_L g9817 ( 
.A(n_9735),
.B(n_4827),
.Y(n_9817)
);

OAI22xp5_ASAP7_75t_L g9818 ( 
.A1(n_9800),
.A2(n_5289),
.B1(n_4961),
.B2(n_5037),
.Y(n_9818)
);

AOI31xp33_ASAP7_75t_L g9819 ( 
.A1(n_9720),
.A2(n_4503),
.A3(n_4442),
.B(n_4606),
.Y(n_9819)
);

XOR2x2_ASAP7_75t_L g9820 ( 
.A(n_9706),
.B(n_4847),
.Y(n_9820)
);

NOR3xp33_ASAP7_75t_L g9821 ( 
.A(n_9713),
.B(n_4021),
.C(n_4017),
.Y(n_9821)
);

INVx1_ASAP7_75t_L g9822 ( 
.A(n_9696),
.Y(n_9822)
);

OAI211xp5_ASAP7_75t_L g9823 ( 
.A1(n_9712),
.A2(n_9741),
.B(n_9746),
.C(n_9739),
.Y(n_9823)
);

AOI22xp5_ASAP7_75t_L g9824 ( 
.A1(n_9707),
.A2(n_5289),
.B1(n_4187),
.B2(n_4961),
.Y(n_9824)
);

INVx1_ASAP7_75t_SL g9825 ( 
.A(n_9693),
.Y(n_9825)
);

AND2x2_ASAP7_75t_L g9826 ( 
.A(n_9778),
.B(n_9748),
.Y(n_9826)
);

INVx1_ASAP7_75t_L g9827 ( 
.A(n_9694),
.Y(n_9827)
);

O2A1O1Ixp33_ASAP7_75t_L g9828 ( 
.A1(n_9716),
.A2(n_4334),
.B(n_4976),
.C(n_4839),
.Y(n_9828)
);

NAND2xp5_ASAP7_75t_SL g9829 ( 
.A(n_9723),
.B(n_4869),
.Y(n_9829)
);

INVx1_ASAP7_75t_L g9830 ( 
.A(n_9790),
.Y(n_9830)
);

CKINVDCx5p33_ASAP7_75t_R g9831 ( 
.A(n_9744),
.Y(n_9831)
);

AOI22xp5_ASAP7_75t_L g9832 ( 
.A1(n_9791),
.A2(n_5289),
.B1(n_4187),
.B2(n_4961),
.Y(n_9832)
);

OR2x2_ASAP7_75t_L g9833 ( 
.A(n_9709),
.B(n_4242),
.Y(n_9833)
);

XOR2xp5_ASAP7_75t_L g9834 ( 
.A(n_9786),
.B(n_4797),
.Y(n_9834)
);

INVx1_ASAP7_75t_L g9835 ( 
.A(n_9715),
.Y(n_9835)
);

AOI322xp5_ASAP7_75t_L g9836 ( 
.A1(n_9788),
.A2(n_4470),
.A3(n_4346),
.B1(n_5361),
.B2(n_5346),
.C1(n_5232),
.C2(n_5218),
.Y(n_9836)
);

INVxp67_ASAP7_75t_SL g9837 ( 
.A(n_9752),
.Y(n_9837)
);

AOI222xp33_ASAP7_75t_L g9838 ( 
.A1(n_9798),
.A2(n_5261),
.B1(n_5223),
.B2(n_5262),
.C1(n_5259),
.C2(n_5232),
.Y(n_9838)
);

AOI21xp5_ASAP7_75t_L g9839 ( 
.A1(n_9750),
.A2(n_4907),
.B(n_4187),
.Y(n_9839)
);

AOI22xp33_ASAP7_75t_SL g9840 ( 
.A1(n_9772),
.A2(n_5286),
.B1(n_4838),
.B2(n_5090),
.Y(n_9840)
);

INVx1_ASAP7_75t_L g9841 ( 
.A(n_9755),
.Y(n_9841)
);

INVxp67_ASAP7_75t_SL g9842 ( 
.A(n_9749),
.Y(n_9842)
);

AND2x2_ASAP7_75t_L g9843 ( 
.A(n_9729),
.B(n_4457),
.Y(n_9843)
);

INVxp67_ASAP7_75t_L g9844 ( 
.A(n_9704),
.Y(n_9844)
);

OAI21xp5_ASAP7_75t_SL g9845 ( 
.A1(n_9763),
.A2(n_4446),
.B(n_4503),
.Y(n_9845)
);

INVx1_ASAP7_75t_L g9846 ( 
.A(n_9802),
.Y(n_9846)
);

NAND2xp5_ASAP7_75t_L g9847 ( 
.A(n_9756),
.B(n_4191),
.Y(n_9847)
);

AOI21xp5_ASAP7_75t_L g9848 ( 
.A1(n_9751),
.A2(n_4301),
.B(n_4269),
.Y(n_9848)
);

NAND4xp25_ASAP7_75t_L g9849 ( 
.A(n_9728),
.B(n_5345),
.C(n_5039),
.D(n_5035),
.Y(n_9849)
);

BUFx3_ASAP7_75t_L g9850 ( 
.A(n_9731),
.Y(n_9850)
);

INVx2_ASAP7_75t_SL g9851 ( 
.A(n_9726),
.Y(n_9851)
);

NAND3xp33_ASAP7_75t_L g9852 ( 
.A(n_9711),
.B(n_5259),
.C(n_5223),
.Y(n_9852)
);

INVx1_ASAP7_75t_L g9853 ( 
.A(n_9727),
.Y(n_9853)
);

NOR2x1_ASAP7_75t_L g9854 ( 
.A(n_9737),
.B(n_4976),
.Y(n_9854)
);

NOR2xp33_ASAP7_75t_L g9855 ( 
.A(n_9781),
.B(n_9732),
.Y(n_9855)
);

AND2x2_ASAP7_75t_L g9856 ( 
.A(n_9760),
.B(n_4457),
.Y(n_9856)
);

AOI21xp5_ASAP7_75t_L g9857 ( 
.A1(n_9774),
.A2(n_4301),
.B(n_4269),
.Y(n_9857)
);

AND2x2_ASAP7_75t_L g9858 ( 
.A(n_9766),
.B(n_4463),
.Y(n_9858)
);

NAND2xp5_ASAP7_75t_L g9859 ( 
.A(n_9736),
.B(n_4191),
.Y(n_9859)
);

NAND2xp5_ASAP7_75t_L g9860 ( 
.A(n_9775),
.B(n_4191),
.Y(n_9860)
);

INVx1_ASAP7_75t_L g9861 ( 
.A(n_9758),
.Y(n_9861)
);

CKINVDCx20_ASAP7_75t_R g9862 ( 
.A(n_9783),
.Y(n_9862)
);

NAND2xp5_ASAP7_75t_SL g9863 ( 
.A(n_9796),
.B(n_4869),
.Y(n_9863)
);

HB1xp67_ASAP7_75t_L g9864 ( 
.A(n_9717),
.Y(n_9864)
);

INVx1_ASAP7_75t_L g9865 ( 
.A(n_9742),
.Y(n_9865)
);

NAND2xp5_ASAP7_75t_L g9866 ( 
.A(n_9747),
.B(n_4191),
.Y(n_9866)
);

INVx1_ASAP7_75t_L g9867 ( 
.A(n_9769),
.Y(n_9867)
);

INVx2_ASAP7_75t_L g9868 ( 
.A(n_9780),
.Y(n_9868)
);

INVx1_ASAP7_75t_L g9869 ( 
.A(n_9770),
.Y(n_9869)
);

INVx1_ASAP7_75t_L g9870 ( 
.A(n_9784),
.Y(n_9870)
);

XOR2x2_ASAP7_75t_L g9871 ( 
.A(n_9777),
.B(n_4854),
.Y(n_9871)
);

AOI221x1_ASAP7_75t_L g9872 ( 
.A1(n_9801),
.A2(n_5253),
.B1(n_5264),
.B2(n_5236),
.C(n_5230),
.Y(n_9872)
);

AOI31xp33_ASAP7_75t_L g9873 ( 
.A1(n_9710),
.A2(n_4503),
.A3(n_4639),
.B(n_4606),
.Y(n_9873)
);

INVx2_ASAP7_75t_SL g9874 ( 
.A(n_9792),
.Y(n_9874)
);

INVx1_ASAP7_75t_L g9875 ( 
.A(n_9714),
.Y(n_9875)
);

INVx1_ASAP7_75t_L g9876 ( 
.A(n_9773),
.Y(n_9876)
);

INVx1_ASAP7_75t_L g9877 ( 
.A(n_9730),
.Y(n_9877)
);

NAND2xp5_ASAP7_75t_L g9878 ( 
.A(n_9776),
.B(n_4191),
.Y(n_9878)
);

INVx1_ASAP7_75t_SL g9879 ( 
.A(n_9785),
.Y(n_9879)
);

AOI22xp33_ASAP7_75t_SL g9880 ( 
.A1(n_9794),
.A2(n_5286),
.B1(n_4838),
.B2(n_5090),
.Y(n_9880)
);

OR2x2_ASAP7_75t_L g9881 ( 
.A(n_9767),
.B(n_4242),
.Y(n_9881)
);

NAND2xp5_ASAP7_75t_L g9882 ( 
.A(n_9759),
.B(n_4191),
.Y(n_9882)
);

NAND4xp75_ASAP7_75t_L g9883 ( 
.A(n_9699),
.B(n_4904),
.C(n_4389),
.D(n_5112),
.Y(n_9883)
);

OAI21xp5_ASAP7_75t_L g9884 ( 
.A1(n_9718),
.A2(n_5064),
.B(n_5030),
.Y(n_9884)
);

AOI22xp5_ASAP7_75t_L g9885 ( 
.A1(n_9764),
.A2(n_4205),
.B1(n_5204),
.B2(n_5089),
.Y(n_9885)
);

NOR4xp25_ASAP7_75t_L g9886 ( 
.A(n_9809),
.B(n_9771),
.C(n_9724),
.D(n_9733),
.Y(n_9886)
);

NOR2x1_ASAP7_75t_L g9887 ( 
.A(n_9807),
.B(n_9754),
.Y(n_9887)
);

AOI22xp5_ASAP7_75t_L g9888 ( 
.A1(n_9830),
.A2(n_9789),
.B1(n_9768),
.B2(n_9745),
.Y(n_9888)
);

AOI22xp5_ASAP7_75t_L g9889 ( 
.A1(n_9825),
.A2(n_9719),
.B1(n_9710),
.B2(n_9753),
.Y(n_9889)
);

OAI22xp5_ASAP7_75t_L g9890 ( 
.A1(n_9837),
.A2(n_9842),
.B1(n_9851),
.B2(n_9822),
.Y(n_9890)
);

INVx1_ASAP7_75t_L g9891 ( 
.A(n_9827),
.Y(n_9891)
);

NOR2x1p5_ASAP7_75t_L g9892 ( 
.A(n_9815),
.B(n_9765),
.Y(n_9892)
);

AOI22xp5_ASAP7_75t_L g9893 ( 
.A1(n_9870),
.A2(n_9862),
.B1(n_9826),
.B2(n_9823),
.Y(n_9893)
);

INVx1_ASAP7_75t_L g9894 ( 
.A(n_9810),
.Y(n_9894)
);

NOR2x1_ASAP7_75t_L g9895 ( 
.A(n_9850),
.B(n_9757),
.Y(n_9895)
);

OAI22xp33_ASAP7_75t_L g9896 ( 
.A1(n_9877),
.A2(n_9743),
.B1(n_9761),
.B2(n_9740),
.Y(n_9896)
);

INVx1_ASAP7_75t_L g9897 ( 
.A(n_9808),
.Y(n_9897)
);

NOR4xp25_ASAP7_75t_L g9898 ( 
.A(n_9835),
.B(n_9705),
.C(n_9782),
.D(n_9787),
.Y(n_9898)
);

OAI22xp33_ASAP7_75t_L g9899 ( 
.A1(n_9868),
.A2(n_9779),
.B1(n_9803),
.B2(n_9738),
.Y(n_9899)
);

OAI22xp5_ASAP7_75t_SL g9900 ( 
.A1(n_9855),
.A2(n_9803),
.B1(n_9721),
.B2(n_9795),
.Y(n_9900)
);

OA22x2_ASAP7_75t_L g9901 ( 
.A1(n_9834),
.A2(n_9762),
.B1(n_5277),
.B2(n_5278),
.Y(n_9901)
);

AOI22xp5_ASAP7_75t_L g9902 ( 
.A1(n_9831),
.A2(n_4869),
.B1(n_5071),
.B2(n_5037),
.Y(n_9902)
);

INVxp67_ASAP7_75t_SL g9903 ( 
.A(n_9864),
.Y(n_9903)
);

NOR4xp25_ASAP7_75t_L g9904 ( 
.A(n_9841),
.B(n_5277),
.C(n_5278),
.D(n_5270),
.Y(n_9904)
);

INVx1_ASAP7_75t_L g9905 ( 
.A(n_9804),
.Y(n_9905)
);

INVx2_ASAP7_75t_L g9906 ( 
.A(n_9816),
.Y(n_9906)
);

AOI22xp33_ASAP7_75t_SL g9907 ( 
.A1(n_9874),
.A2(n_9861),
.B1(n_9865),
.B2(n_9879),
.Y(n_9907)
);

AOI22xp5_ASAP7_75t_L g9908 ( 
.A1(n_9853),
.A2(n_4869),
.B1(n_5071),
.B2(n_5037),
.Y(n_9908)
);

INVx1_ASAP7_75t_L g9909 ( 
.A(n_9820),
.Y(n_9909)
);

BUFx2_ASAP7_75t_L g9910 ( 
.A(n_9817),
.Y(n_9910)
);

AOI22xp5_ASAP7_75t_L g9911 ( 
.A1(n_9875),
.A2(n_5037),
.B1(n_5085),
.B2(n_5071),
.Y(n_9911)
);

AOI22xp5_ASAP7_75t_L g9912 ( 
.A1(n_9811),
.A2(n_9876),
.B1(n_9844),
.B2(n_9814),
.Y(n_9912)
);

NAND2xp5_ASAP7_75t_L g9913 ( 
.A(n_9867),
.B(n_5223),
.Y(n_9913)
);

AOI22xp5_ASAP7_75t_L g9914 ( 
.A1(n_9869),
.A2(n_5071),
.B1(n_5089),
.B2(n_5085),
.Y(n_9914)
);

NOR4xp25_ASAP7_75t_L g9915 ( 
.A(n_9846),
.B(n_5282),
.C(n_5284),
.D(n_5281),
.Y(n_9915)
);

INVx1_ASAP7_75t_L g9916 ( 
.A(n_9829),
.Y(n_9916)
);

INVx1_ASAP7_75t_L g9917 ( 
.A(n_9833),
.Y(n_9917)
);

AOI22xp33_ASAP7_75t_SL g9918 ( 
.A1(n_9812),
.A2(n_4838),
.B1(n_5286),
.B2(n_5090),
.Y(n_9918)
);

INVx1_ASAP7_75t_L g9919 ( 
.A(n_9881),
.Y(n_9919)
);

O2A1O1Ixp33_ASAP7_75t_L g9920 ( 
.A1(n_9821),
.A2(n_9863),
.B(n_9847),
.C(n_9878),
.Y(n_9920)
);

A2O1A1Ixp33_ASAP7_75t_SL g9921 ( 
.A1(n_9857),
.A2(n_5282),
.B(n_5284),
.C(n_5281),
.Y(n_9921)
);

INVx1_ASAP7_75t_L g9922 ( 
.A(n_9871),
.Y(n_9922)
);

INVx1_ASAP7_75t_L g9923 ( 
.A(n_9859),
.Y(n_9923)
);

INVx1_ASAP7_75t_L g9924 ( 
.A(n_9860),
.Y(n_9924)
);

AOI22xp5_ASAP7_75t_L g9925 ( 
.A1(n_9866),
.A2(n_5071),
.B1(n_5089),
.B2(n_5085),
.Y(n_9925)
);

INVx1_ASAP7_75t_L g9926 ( 
.A(n_9843),
.Y(n_9926)
);

OA22x2_ASAP7_75t_L g9927 ( 
.A1(n_9806),
.A2(n_5298),
.B1(n_5305),
.B2(n_5296),
.Y(n_9927)
);

AOI22xp5_ASAP7_75t_L g9928 ( 
.A1(n_9839),
.A2(n_5071),
.B1(n_5089),
.B2(n_5085),
.Y(n_9928)
);

NOR2x1_ASAP7_75t_L g9929 ( 
.A(n_9854),
.B(n_4976),
.Y(n_9929)
);

INVx1_ASAP7_75t_L g9930 ( 
.A(n_9856),
.Y(n_9930)
);

AOI22xp5_ASAP7_75t_L g9931 ( 
.A1(n_9818),
.A2(n_5085),
.B1(n_5113),
.B2(n_5089),
.Y(n_9931)
);

INVx1_ASAP7_75t_L g9932 ( 
.A(n_9858),
.Y(n_9932)
);

NOR2xp33_ASAP7_75t_L g9933 ( 
.A(n_9882),
.B(n_3690),
.Y(n_9933)
);

NAND2xp5_ASAP7_75t_L g9934 ( 
.A(n_9885),
.B(n_5261),
.Y(n_9934)
);

INVx2_ASAP7_75t_L g9935 ( 
.A(n_9854),
.Y(n_9935)
);

INVx1_ASAP7_75t_L g9936 ( 
.A(n_9872),
.Y(n_9936)
);

NAND2xp5_ASAP7_75t_L g9937 ( 
.A(n_9885),
.B(n_5261),
.Y(n_9937)
);

INVx1_ASAP7_75t_L g9938 ( 
.A(n_9848),
.Y(n_9938)
);

NAND2xp5_ASAP7_75t_L g9939 ( 
.A(n_9832),
.B(n_5262),
.Y(n_9939)
);

AOI22xp5_ASAP7_75t_L g9940 ( 
.A1(n_9883),
.A2(n_5085),
.B1(n_5113),
.B2(n_5089),
.Y(n_9940)
);

INVx1_ASAP7_75t_L g9941 ( 
.A(n_9852),
.Y(n_9941)
);

NOR2xp33_ASAP7_75t_L g9942 ( 
.A(n_9845),
.B(n_3690),
.Y(n_9942)
);

NOR2x1_ASAP7_75t_L g9943 ( 
.A(n_9828),
.B(n_3636),
.Y(n_9943)
);

OAI22xp5_ASAP7_75t_L g9944 ( 
.A1(n_9824),
.A2(n_5204),
.B1(n_5221),
.B2(n_5113),
.Y(n_9944)
);

AOI22xp5_ASAP7_75t_L g9945 ( 
.A1(n_9880),
.A2(n_5204),
.B1(n_5221),
.B2(n_5113),
.Y(n_9945)
);

NOR2x1_ASAP7_75t_L g9946 ( 
.A(n_9819),
.B(n_3642),
.Y(n_9946)
);

INVx1_ASAP7_75t_L g9947 ( 
.A(n_9805),
.Y(n_9947)
);

AOI22xp5_ASAP7_75t_L g9948 ( 
.A1(n_9884),
.A2(n_4205),
.B1(n_5204),
.B2(n_5113),
.Y(n_9948)
);

AOI22xp5_ASAP7_75t_L g9949 ( 
.A1(n_9840),
.A2(n_5113),
.B1(n_5221),
.B2(n_5204),
.Y(n_9949)
);

NOR2x1_ASAP7_75t_L g9950 ( 
.A(n_9849),
.B(n_3676),
.Y(n_9950)
);

INVx2_ASAP7_75t_L g9951 ( 
.A(n_9813),
.Y(n_9951)
);

NOR4xp25_ASAP7_75t_L g9952 ( 
.A(n_9873),
.B(n_5298),
.C(n_5305),
.D(n_5296),
.Y(n_9952)
);

NAND2xp5_ASAP7_75t_L g9953 ( 
.A(n_9836),
.B(n_5262),
.Y(n_9953)
);

INVx1_ASAP7_75t_L g9954 ( 
.A(n_9838),
.Y(n_9954)
);

INVx1_ASAP7_75t_L g9955 ( 
.A(n_9903),
.Y(n_9955)
);

INVx1_ASAP7_75t_L g9956 ( 
.A(n_9891),
.Y(n_9956)
);

NAND2xp5_ASAP7_75t_L g9957 ( 
.A(n_9893),
.B(n_4271),
.Y(n_9957)
);

NOR2x1_ASAP7_75t_L g9958 ( 
.A(n_9890),
.B(n_4623),
.Y(n_9958)
);

NOR2x1p5_ASAP7_75t_L g9959 ( 
.A(n_9894),
.B(n_3644),
.Y(n_9959)
);

NOR2x1_ASAP7_75t_L g9960 ( 
.A(n_9892),
.B(n_4623),
.Y(n_9960)
);

NAND2xp5_ASAP7_75t_L g9961 ( 
.A(n_9935),
.B(n_4271),
.Y(n_9961)
);

NAND2xp5_ASAP7_75t_SL g9962 ( 
.A(n_9907),
.B(n_5055),
.Y(n_9962)
);

A2O1A1Ixp33_ASAP7_75t_L g9963 ( 
.A1(n_9920),
.A2(n_5320),
.B(n_5326),
.C(n_5318),
.Y(n_9963)
);

NOR3xp33_ASAP7_75t_L g9964 ( 
.A(n_9897),
.B(n_3698),
.C(n_3676),
.Y(n_9964)
);

INVxp33_ASAP7_75t_L g9965 ( 
.A(n_9887),
.Y(n_9965)
);

OAI22xp33_ASAP7_75t_L g9966 ( 
.A1(n_9888),
.A2(n_5221),
.B1(n_5225),
.B2(n_5204),
.Y(n_9966)
);

AOI311xp33_ASAP7_75t_L g9967 ( 
.A1(n_9900),
.A2(n_9922),
.A3(n_9909),
.B(n_9899),
.C(n_9916),
.Y(n_9967)
);

AOI222xp33_ASAP7_75t_L g9968 ( 
.A1(n_9919),
.A2(n_5320),
.B1(n_5326),
.B2(n_5334),
.C1(n_5327),
.C2(n_5318),
.Y(n_9968)
);

INVx2_ASAP7_75t_L g9969 ( 
.A(n_9905),
.Y(n_9969)
);

AND2x4_ASAP7_75t_L g9970 ( 
.A(n_9895),
.B(n_5221),
.Y(n_9970)
);

OR2x2_ASAP7_75t_L g9971 ( 
.A(n_9917),
.B(n_4271),
.Y(n_9971)
);

INVx1_ASAP7_75t_L g9972 ( 
.A(n_9936),
.Y(n_9972)
);

INVx1_ASAP7_75t_SL g9973 ( 
.A(n_9926),
.Y(n_9973)
);

NAND4xp75_ASAP7_75t_L g9974 ( 
.A(n_9912),
.B(n_4904),
.C(n_4320),
.D(n_5112),
.Y(n_9974)
);

AND2x2_ASAP7_75t_L g9975 ( 
.A(n_9929),
.B(n_4463),
.Y(n_9975)
);

INVx2_ASAP7_75t_L g9976 ( 
.A(n_9906),
.Y(n_9976)
);

INVx1_ASAP7_75t_L g9977 ( 
.A(n_9930),
.Y(n_9977)
);

NAND2xp5_ASAP7_75t_L g9978 ( 
.A(n_9910),
.B(n_4271),
.Y(n_9978)
);

INVx1_ASAP7_75t_L g9979 ( 
.A(n_9932),
.Y(n_9979)
);

NAND2x1p5_ASAP7_75t_L g9980 ( 
.A(n_9924),
.B(n_3676),
.Y(n_9980)
);

INVxp67_ASAP7_75t_L g9981 ( 
.A(n_9954),
.Y(n_9981)
);

INVx2_ASAP7_75t_L g9982 ( 
.A(n_9901),
.Y(n_9982)
);

NAND2xp33_ASAP7_75t_L g9983 ( 
.A(n_9951),
.B(n_5221),
.Y(n_9983)
);

AND2x2_ASAP7_75t_L g9984 ( 
.A(n_9950),
.B(n_4781),
.Y(n_9984)
);

NOR3xp33_ASAP7_75t_L g9985 ( 
.A(n_9923),
.B(n_3698),
.C(n_3676),
.Y(n_9985)
);

INVx1_ASAP7_75t_SL g9986 ( 
.A(n_9941),
.Y(n_9986)
);

OAI21xp5_ASAP7_75t_L g9987 ( 
.A1(n_9898),
.A2(n_5064),
.B(n_5030),
.Y(n_9987)
);

NAND2xp5_ASAP7_75t_L g9988 ( 
.A(n_9886),
.B(n_4271),
.Y(n_9988)
);

BUFx4f_ASAP7_75t_SL g9989 ( 
.A(n_9947),
.Y(n_9989)
);

OAI21xp33_ASAP7_75t_L g9990 ( 
.A1(n_9889),
.A2(n_5251),
.B(n_5225),
.Y(n_9990)
);

NAND3xp33_ASAP7_75t_L g9991 ( 
.A(n_9938),
.B(n_5090),
.C(n_5055),
.Y(n_9991)
);

NAND2xp5_ASAP7_75t_L g9992 ( 
.A(n_9896),
.B(n_4271),
.Y(n_9992)
);

AND2x2_ASAP7_75t_L g9993 ( 
.A(n_9946),
.B(n_4781),
.Y(n_9993)
);

INVx3_ASAP7_75t_SL g9994 ( 
.A(n_9927),
.Y(n_9994)
);

AOI21xp5_ASAP7_75t_L g9995 ( 
.A1(n_9921),
.A2(n_4301),
.B(n_4269),
.Y(n_9995)
);

INVx1_ASAP7_75t_L g9996 ( 
.A(n_9913),
.Y(n_9996)
);

AND2x2_ASAP7_75t_L g9997 ( 
.A(n_9943),
.B(n_4781),
.Y(n_9997)
);

NAND2xp5_ASAP7_75t_L g9998 ( 
.A(n_9933),
.B(n_5694),
.Y(n_9998)
);

INVxp67_ASAP7_75t_L g9999 ( 
.A(n_9953),
.Y(n_9999)
);

NAND2xp33_ASAP7_75t_L g10000 ( 
.A(n_9902),
.B(n_9908),
.Y(n_10000)
);

NAND3x1_ASAP7_75t_SL g10001 ( 
.A(n_9952),
.B(n_3690),
.C(n_4965),
.Y(n_10001)
);

AND2x4_ASAP7_75t_L g10002 ( 
.A(n_9942),
.B(n_9914),
.Y(n_10002)
);

AOI22xp5_ASAP7_75t_L g10003 ( 
.A1(n_9939),
.A2(n_5225),
.B1(n_5251),
.B2(n_4205),
.Y(n_10003)
);

INVx1_ASAP7_75t_L g10004 ( 
.A(n_9934),
.Y(n_10004)
);

NOR2xp33_ASAP7_75t_L g10005 ( 
.A(n_9937),
.B(n_5225),
.Y(n_10005)
);

OAI21xp33_ASAP7_75t_L g10006 ( 
.A1(n_9911),
.A2(n_9925),
.B(n_9918),
.Y(n_10006)
);

NOR2x1_ASAP7_75t_L g10007 ( 
.A(n_9944),
.B(n_4623),
.Y(n_10007)
);

XNOR2x1_ASAP7_75t_L g10008 ( 
.A(n_9928),
.B(n_4854),
.Y(n_10008)
);

NAND2xp33_ASAP7_75t_SL g10009 ( 
.A(n_9904),
.B(n_5225),
.Y(n_10009)
);

NAND2xp5_ASAP7_75t_L g10010 ( 
.A(n_9915),
.B(n_5694),
.Y(n_10010)
);

AOI22x1_ASAP7_75t_L g10011 ( 
.A1(n_9955),
.A2(n_9940),
.B1(n_9949),
.B2(n_9945),
.Y(n_10011)
);

NOR2x1_ASAP7_75t_L g10012 ( 
.A(n_9956),
.B(n_9948),
.Y(n_10012)
);

NOR3xp33_ASAP7_75t_SL g10013 ( 
.A(n_9972),
.B(n_9948),
.C(n_9931),
.Y(n_10013)
);

AND2x4_ASAP7_75t_L g10014 ( 
.A(n_9970),
.B(n_5225),
.Y(n_10014)
);

XNOR2xp5_ASAP7_75t_L g10015 ( 
.A(n_9965),
.B(n_9973),
.Y(n_10015)
);

INVx1_ASAP7_75t_L g10016 ( 
.A(n_9970),
.Y(n_10016)
);

INVx1_ASAP7_75t_SL g10017 ( 
.A(n_9986),
.Y(n_10017)
);

AND2x4_ASAP7_75t_L g10018 ( 
.A(n_9975),
.B(n_5251),
.Y(n_10018)
);

INVx1_ASAP7_75t_L g10019 ( 
.A(n_9969),
.Y(n_10019)
);

AND4x1_ASAP7_75t_L g10020 ( 
.A(n_9967),
.B(n_4616),
.C(n_4489),
.D(n_4526),
.Y(n_10020)
);

INVx1_ASAP7_75t_L g10021 ( 
.A(n_9976),
.Y(n_10021)
);

NOR2xp33_ASAP7_75t_L g10022 ( 
.A(n_9981),
.B(n_9989),
.Y(n_10022)
);

NAND4xp25_ASAP7_75t_L g10023 ( 
.A(n_9977),
.B(n_4655),
.C(n_4666),
.D(n_3698),
.Y(n_10023)
);

NAND3xp33_ASAP7_75t_SL g10024 ( 
.A(n_9979),
.B(n_4862),
.C(n_4855),
.Y(n_10024)
);

NOR3xp33_ASAP7_75t_SL g10025 ( 
.A(n_9996),
.B(n_4616),
.C(n_4489),
.Y(n_10025)
);

NOR3xp33_ASAP7_75t_L g10026 ( 
.A(n_9999),
.B(n_3698),
.C(n_4017),
.Y(n_10026)
);

INVx1_ASAP7_75t_L g10027 ( 
.A(n_9960),
.Y(n_10027)
);

AND2x4_ASAP7_75t_L g10028 ( 
.A(n_9959),
.B(n_5251),
.Y(n_10028)
);

INVx1_ASAP7_75t_L g10029 ( 
.A(n_9988),
.Y(n_10029)
);

NAND4xp25_ASAP7_75t_L g10030 ( 
.A(n_9962),
.B(n_3755),
.C(n_3756),
.D(n_3754),
.Y(n_10030)
);

NOR2x1_ASAP7_75t_L g10031 ( 
.A(n_9982),
.B(n_4623),
.Y(n_10031)
);

OR2x2_ASAP7_75t_L g10032 ( 
.A(n_9980),
.B(n_5694),
.Y(n_10032)
);

NAND3xp33_ASAP7_75t_L g10033 ( 
.A(n_10004),
.B(n_9983),
.C(n_10000),
.Y(n_10033)
);

NOR2x1_ASAP7_75t_L g10034 ( 
.A(n_10002),
.B(n_5308),
.Y(n_10034)
);

NOR2x1p5_ASAP7_75t_L g10035 ( 
.A(n_9957),
.B(n_3644),
.Y(n_10035)
);

AOI211xp5_ASAP7_75t_SL g10036 ( 
.A1(n_10006),
.A2(n_4071),
.B(n_4090),
.C(n_4331),
.Y(n_10036)
);

NAND2xp5_ASAP7_75t_L g10037 ( 
.A(n_10005),
.B(n_5694),
.Y(n_10037)
);

NOR4xp25_ASAP7_75t_L g10038 ( 
.A(n_9978),
.B(n_5309),
.C(n_5306),
.D(n_5327),
.Y(n_10038)
);

NOR4xp25_ASAP7_75t_L g10039 ( 
.A(n_9992),
.B(n_5309),
.C(n_5306),
.D(n_5334),
.Y(n_10039)
);

NAND3xp33_ASAP7_75t_L g10040 ( 
.A(n_10002),
.B(n_5090),
.C(n_5055),
.Y(n_10040)
);

NAND3xp33_ASAP7_75t_SL g10041 ( 
.A(n_9961),
.B(n_4926),
.C(n_4862),
.Y(n_10041)
);

AOI22xp5_ASAP7_75t_L g10042 ( 
.A1(n_9984),
.A2(n_5251),
.B1(n_4965),
.B2(n_4269),
.Y(n_10042)
);

INVx1_ASAP7_75t_L g10043 ( 
.A(n_9958),
.Y(n_10043)
);

NOR3xp33_ASAP7_75t_L g10044 ( 
.A(n_10001),
.B(n_4021),
.C(n_4017),
.Y(n_10044)
);

NOR3xp33_ASAP7_75t_L g10045 ( 
.A(n_9993),
.B(n_4021),
.C(n_4017),
.Y(n_10045)
);

NAND4xp25_ASAP7_75t_L g10046 ( 
.A(n_9990),
.B(n_3755),
.C(n_3756),
.D(n_3754),
.Y(n_10046)
);

NOR2x1_ASAP7_75t_L g10047 ( 
.A(n_9997),
.B(n_5308),
.Y(n_10047)
);

AND2x4_ASAP7_75t_L g10048 ( 
.A(n_9964),
.B(n_3756),
.Y(n_10048)
);

OAI211xp5_ASAP7_75t_L g10049 ( 
.A1(n_10009),
.A2(n_3800),
.B(n_3889),
.C(n_4256),
.Y(n_10049)
);

NAND2xp5_ASAP7_75t_L g10050 ( 
.A(n_9994),
.B(n_5694),
.Y(n_10050)
);

AOI221xp5_ASAP7_75t_L g10051 ( 
.A1(n_9966),
.A2(n_10010),
.B1(n_9998),
.B2(n_9987),
.C(n_9991),
.Y(n_10051)
);

NOR2xp67_ASAP7_75t_L g10052 ( 
.A(n_9971),
.B(n_5055),
.Y(n_10052)
);

NOR3xp33_ASAP7_75t_L g10053 ( 
.A(n_10007),
.B(n_4038),
.C(n_4021),
.Y(n_10053)
);

NOR2xp33_ASAP7_75t_L g10054 ( 
.A(n_10008),
.B(n_9963),
.Y(n_10054)
);

NOR2xp33_ASAP7_75t_L g10055 ( 
.A(n_10003),
.B(n_4965),
.Y(n_10055)
);

NOR3xp33_ASAP7_75t_L g10056 ( 
.A(n_9985),
.B(n_4038),
.C(n_3719),
.Y(n_10056)
);

OAI211xp5_ASAP7_75t_L g10057 ( 
.A1(n_9995),
.A2(n_3800),
.B(n_4368),
.C(n_4336),
.Y(n_10057)
);

NOR2xp67_ASAP7_75t_L g10058 ( 
.A(n_9968),
.B(n_5090),
.Y(n_10058)
);

BUFx3_ASAP7_75t_L g10059 ( 
.A(n_9974),
.Y(n_10059)
);

NAND5xp2_ASAP7_75t_L g10060 ( 
.A(n_10022),
.B(n_5040),
.C(n_5046),
.D(n_4926),
.E(n_4862),
.Y(n_10060)
);

NOR3xp33_ASAP7_75t_SL g10061 ( 
.A(n_10015),
.B(n_4526),
.C(n_5336),
.Y(n_10061)
);

NAND4xp75_ASAP7_75t_L g10062 ( 
.A(n_10012),
.B(n_4320),
.C(n_4904),
.D(n_5112),
.Y(n_10062)
);

AND3x2_ASAP7_75t_L g10063 ( 
.A(n_10021),
.B(n_4394),
.C(n_4368),
.Y(n_10063)
);

BUFx6f_ASAP7_75t_L g10064 ( 
.A(n_10019),
.Y(n_10064)
);

NAND3x1_ASAP7_75t_L g10065 ( 
.A(n_10016),
.B(n_5337),
.C(n_5336),
.Y(n_10065)
);

AND2x2_ASAP7_75t_SL g10066 ( 
.A(n_10029),
.B(n_4320),
.Y(n_10066)
);

INVx1_ASAP7_75t_L g10067 ( 
.A(n_10017),
.Y(n_10067)
);

AO22x1_ASAP7_75t_L g10068 ( 
.A1(n_10027),
.A2(n_3793),
.B1(n_5344),
.B2(n_5343),
.Y(n_10068)
);

NAND2x1p5_ASAP7_75t_L g10069 ( 
.A(n_10043),
.B(n_3789),
.Y(n_10069)
);

INVxp33_ASAP7_75t_SL g10070 ( 
.A(n_10033),
.Y(n_10070)
);

NAND2xp5_ASAP7_75t_L g10071 ( 
.A(n_10014),
.B(n_5280),
.Y(n_10071)
);

AOI21xp33_ASAP7_75t_L g10072 ( 
.A1(n_10011),
.A2(n_5290),
.B(n_5280),
.Y(n_10072)
);

NOR2xp33_ASAP7_75t_L g10073 ( 
.A(n_10050),
.B(n_4965),
.Y(n_10073)
);

AND2x2_ASAP7_75t_L g10074 ( 
.A(n_10047),
.B(n_5224),
.Y(n_10074)
);

OAI322xp33_ASAP7_75t_L g10075 ( 
.A1(n_10054),
.A2(n_5365),
.A3(n_5367),
.B1(n_5344),
.B2(n_4537),
.C1(n_4487),
.C2(n_4559),
.Y(n_10075)
);

NAND4xp75_ASAP7_75t_L g10076 ( 
.A(n_10013),
.B(n_4320),
.C(n_5112),
.D(n_4254),
.Y(n_10076)
);

AND2x2_ASAP7_75t_L g10077 ( 
.A(n_10034),
.B(n_5224),
.Y(n_10077)
);

AND3x4_ASAP7_75t_L g10078 ( 
.A(n_10020),
.B(n_10059),
.C(n_10028),
.Y(n_10078)
);

INVx1_ASAP7_75t_L g10079 ( 
.A(n_10035),
.Y(n_10079)
);

OAI21xp5_ASAP7_75t_SL g10080 ( 
.A1(n_10051),
.A2(n_4926),
.B(n_5040),
.Y(n_10080)
);

XNOR2x1_ASAP7_75t_SL g10081 ( 
.A(n_10039),
.B(n_4606),
.Y(n_10081)
);

NOR2xp33_ASAP7_75t_L g10082 ( 
.A(n_10018),
.B(n_10052),
.Y(n_10082)
);

OAI221xp5_ASAP7_75t_L g10083 ( 
.A1(n_10044),
.A2(n_4394),
.B1(n_3757),
.B2(n_3793),
.C(n_4458),
.Y(n_10083)
);

NAND2xp5_ASAP7_75t_L g10084 ( 
.A(n_10037),
.B(n_5290),
.Y(n_10084)
);

INVx1_ASAP7_75t_L g10085 ( 
.A(n_10032),
.Y(n_10085)
);

INVxp67_ASAP7_75t_L g10086 ( 
.A(n_10055),
.Y(n_10086)
);

INVxp67_ASAP7_75t_L g10087 ( 
.A(n_10031),
.Y(n_10087)
);

NAND4xp25_ASAP7_75t_L g10088 ( 
.A(n_10045),
.B(n_3757),
.C(n_4495),
.D(n_4038),
.Y(n_10088)
);

INVx2_ASAP7_75t_L g10089 ( 
.A(n_10048),
.Y(n_10089)
);

HB1xp67_ASAP7_75t_L g10090 ( 
.A(n_10058),
.Y(n_10090)
);

NAND2xp33_ASAP7_75t_SL g10091 ( 
.A(n_10048),
.B(n_3793),
.Y(n_10091)
);

INVxp67_ASAP7_75t_SL g10092 ( 
.A(n_10053),
.Y(n_10092)
);

AND2x2_ASAP7_75t_L g10093 ( 
.A(n_10026),
.B(n_5224),
.Y(n_10093)
);

NAND2x1p5_ASAP7_75t_L g10094 ( 
.A(n_10042),
.B(n_4038),
.Y(n_10094)
);

NOR2x1_ASAP7_75t_L g10095 ( 
.A(n_10057),
.B(n_5308),
.Y(n_10095)
);

AND2x4_ASAP7_75t_L g10096 ( 
.A(n_10067),
.B(n_10056),
.Y(n_10096)
);

OR2x2_ASAP7_75t_L g10097 ( 
.A(n_10064),
.B(n_10038),
.Y(n_10097)
);

INVxp67_ASAP7_75t_L g10098 ( 
.A(n_10064),
.Y(n_10098)
);

OR2x2_ASAP7_75t_L g10099 ( 
.A(n_10064),
.B(n_10041),
.Y(n_10099)
);

OR4x2_ASAP7_75t_L g10100 ( 
.A(n_10070),
.B(n_10024),
.C(n_10049),
.D(n_10036),
.Y(n_10100)
);

NOR2x1_ASAP7_75t_L g10101 ( 
.A(n_10078),
.B(n_10040),
.Y(n_10101)
);

NOR2xp33_ASAP7_75t_L g10102 ( 
.A(n_10090),
.B(n_10085),
.Y(n_10102)
);

NAND2xp5_ASAP7_75t_L g10103 ( 
.A(n_10082),
.B(n_10030),
.Y(n_10103)
);

BUFx2_ASAP7_75t_L g10104 ( 
.A(n_10087),
.Y(n_10104)
);

INVx1_ASAP7_75t_L g10105 ( 
.A(n_10069),
.Y(n_10105)
);

OR2x6_ASAP7_75t_L g10106 ( 
.A(n_10089),
.B(n_10046),
.Y(n_10106)
);

NOR2xp33_ASAP7_75t_L g10107 ( 
.A(n_10079),
.B(n_10023),
.Y(n_10107)
);

INVx2_ASAP7_75t_L g10108 ( 
.A(n_10074),
.Y(n_10108)
);

NAND3x1_ASAP7_75t_SL g10109 ( 
.A(n_10095),
.B(n_10025),
.C(n_3644),
.Y(n_10109)
);

INVx2_ASAP7_75t_L g10110 ( 
.A(n_10077),
.Y(n_10110)
);

HB1xp67_ASAP7_75t_L g10111 ( 
.A(n_10092),
.Y(n_10111)
);

INVx1_ASAP7_75t_L g10112 ( 
.A(n_10073),
.Y(n_10112)
);

AO22x1_ASAP7_75t_L g10113 ( 
.A1(n_10086),
.A2(n_3757),
.B1(n_3696),
.B2(n_4107),
.Y(n_10113)
);

BUFx3_ASAP7_75t_L g10114 ( 
.A(n_10094),
.Y(n_10114)
);

INVxp33_ASAP7_75t_L g10115 ( 
.A(n_10081),
.Y(n_10115)
);

NOR3xp33_ASAP7_75t_L g10116 ( 
.A(n_10091),
.B(n_10084),
.C(n_10093),
.Y(n_10116)
);

INVx1_ASAP7_75t_L g10117 ( 
.A(n_10071),
.Y(n_10117)
);

INVx4_ASAP7_75t_L g10118 ( 
.A(n_10063),
.Y(n_10118)
);

INVx1_ASAP7_75t_L g10119 ( 
.A(n_10061),
.Y(n_10119)
);

INVx1_ASAP7_75t_L g10120 ( 
.A(n_10066),
.Y(n_10120)
);

AND3x4_ASAP7_75t_L g10121 ( 
.A(n_10072),
.B(n_4422),
.C(n_4178),
.Y(n_10121)
);

NOR2xp33_ASAP7_75t_L g10122 ( 
.A(n_10080),
.B(n_5224),
.Y(n_10122)
);

NOR2x1_ASAP7_75t_L g10123 ( 
.A(n_10088),
.B(n_4320),
.Y(n_10123)
);

INVx1_ASAP7_75t_L g10124 ( 
.A(n_10111),
.Y(n_10124)
);

INVx2_ASAP7_75t_L g10125 ( 
.A(n_10104),
.Y(n_10125)
);

AOI22xp5_ASAP7_75t_L g10126 ( 
.A1(n_10098),
.A2(n_10065),
.B1(n_10083),
.B2(n_10076),
.Y(n_10126)
);

INVx1_ASAP7_75t_L g10127 ( 
.A(n_10102),
.Y(n_10127)
);

AND2x4_ASAP7_75t_SL g10128 ( 
.A(n_10108),
.B(n_10068),
.Y(n_10128)
);

INVx2_ASAP7_75t_L g10129 ( 
.A(n_10097),
.Y(n_10129)
);

CKINVDCx20_ASAP7_75t_R g10130 ( 
.A(n_10110),
.Y(n_10130)
);

INVx1_ASAP7_75t_L g10131 ( 
.A(n_10118),
.Y(n_10131)
);

INVx1_ASAP7_75t_L g10132 ( 
.A(n_10099),
.Y(n_10132)
);

NAND2xp5_ASAP7_75t_L g10133 ( 
.A(n_10120),
.B(n_10062),
.Y(n_10133)
);

OAI22xp5_ASAP7_75t_L g10134 ( 
.A1(n_10115),
.A2(n_10075),
.B1(n_10060),
.B2(n_4473),
.Y(n_10134)
);

INVx1_ASAP7_75t_L g10135 ( 
.A(n_10105),
.Y(n_10135)
);

NAND2xp5_ASAP7_75t_L g10136 ( 
.A(n_10119),
.B(n_4838),
.Y(n_10136)
);

HB1xp67_ASAP7_75t_L g10137 ( 
.A(n_10101),
.Y(n_10137)
);

CKINVDCx20_ASAP7_75t_R g10138 ( 
.A(n_10103),
.Y(n_10138)
);

AOI222xp33_ASAP7_75t_L g10139 ( 
.A1(n_10114),
.A2(n_5228),
.B1(n_4552),
.B2(n_5290),
.C1(n_5299),
.C2(n_5280),
.Y(n_10139)
);

CKINVDCx20_ASAP7_75t_R g10140 ( 
.A(n_10106),
.Y(n_10140)
);

NAND2xp5_ASAP7_75t_L g10141 ( 
.A(n_10117),
.B(n_4838),
.Y(n_10141)
);

NAND2xp5_ASAP7_75t_L g10142 ( 
.A(n_10116),
.B(n_4838),
.Y(n_10142)
);

HB1xp67_ASAP7_75t_L g10143 ( 
.A(n_10106),
.Y(n_10143)
);

OAI21xp5_ASAP7_75t_L g10144 ( 
.A1(n_10107),
.A2(n_4762),
.B(n_4749),
.Y(n_10144)
);

NAND2xp5_ASAP7_75t_L g10145 ( 
.A(n_10112),
.B(n_4838),
.Y(n_10145)
);

OAI22xp5_ASAP7_75t_L g10146 ( 
.A1(n_10096),
.A2(n_4473),
.B1(n_4543),
.B2(n_4402),
.Y(n_10146)
);

AOI211x1_ASAP7_75t_L g10147 ( 
.A1(n_10109),
.A2(n_4652),
.B(n_4653),
.C(n_4651),
.Y(n_10147)
);

AND3x1_ASAP7_75t_L g10148 ( 
.A(n_10122),
.B(n_5314),
.C(n_5299),
.Y(n_10148)
);

INVx2_ASAP7_75t_L g10149 ( 
.A(n_10125),
.Y(n_10149)
);

INVx1_ASAP7_75t_SL g10150 ( 
.A(n_10137),
.Y(n_10150)
);

INVx2_ASAP7_75t_L g10151 ( 
.A(n_10124),
.Y(n_10151)
);

AND2x2_ASAP7_75t_L g10152 ( 
.A(n_10143),
.B(n_10123),
.Y(n_10152)
);

INVx2_ASAP7_75t_L g10153 ( 
.A(n_10140),
.Y(n_10153)
);

INVx2_ASAP7_75t_SL g10154 ( 
.A(n_10127),
.Y(n_10154)
);

INVx1_ASAP7_75t_L g10155 ( 
.A(n_10130),
.Y(n_10155)
);

XOR2xp5_ASAP7_75t_L g10156 ( 
.A(n_10138),
.B(n_10100),
.Y(n_10156)
);

OAI22xp5_ASAP7_75t_SL g10157 ( 
.A1(n_10131),
.A2(n_10121),
.B1(n_10113),
.B2(n_5040),
.Y(n_10157)
);

INVxp67_ASAP7_75t_L g10158 ( 
.A(n_10132),
.Y(n_10158)
);

INVx2_ASAP7_75t_SL g10159 ( 
.A(n_10135),
.Y(n_10159)
);

AOI22xp5_ASAP7_75t_L g10160 ( 
.A1(n_10129),
.A2(n_3759),
.B1(n_3763),
.B2(n_3760),
.Y(n_10160)
);

AOI22xp5_ASAP7_75t_L g10161 ( 
.A1(n_10134),
.A2(n_3759),
.B1(n_3763),
.B2(n_3760),
.Y(n_10161)
);

INVx1_ASAP7_75t_L g10162 ( 
.A(n_10128),
.Y(n_10162)
);

AOI22x1_ASAP7_75t_L g10163 ( 
.A1(n_10133),
.A2(n_3760),
.B1(n_3763),
.B2(n_3759),
.Y(n_10163)
);

INVx1_ASAP7_75t_L g10164 ( 
.A(n_10126),
.Y(n_10164)
);

INVx1_ASAP7_75t_L g10165 ( 
.A(n_10142),
.Y(n_10165)
);

NAND2xp5_ASAP7_75t_SL g10166 ( 
.A(n_10145),
.B(n_5228),
.Y(n_10166)
);

INVx1_ASAP7_75t_L g10167 ( 
.A(n_10141),
.Y(n_10167)
);

INVx1_ASAP7_75t_L g10168 ( 
.A(n_10136),
.Y(n_10168)
);

INVx1_ASAP7_75t_L g10169 ( 
.A(n_10148),
.Y(n_10169)
);

INVx2_ASAP7_75t_SL g10170 ( 
.A(n_10146),
.Y(n_10170)
);

INVx1_ASAP7_75t_L g10171 ( 
.A(n_10147),
.Y(n_10171)
);

OR2x2_ASAP7_75t_L g10172 ( 
.A(n_10150),
.B(n_10144),
.Y(n_10172)
);

OAI21x1_ASAP7_75t_SL g10173 ( 
.A1(n_10156),
.A2(n_10139),
.B(n_4604),
.Y(n_10173)
);

CKINVDCx20_ASAP7_75t_R g10174 ( 
.A(n_10153),
.Y(n_10174)
);

AOI22xp33_ASAP7_75t_L g10175 ( 
.A1(n_10159),
.A2(n_5286),
.B1(n_4838),
.B2(n_3891),
.Y(n_10175)
);

NAND2xp5_ASAP7_75t_L g10176 ( 
.A(n_10158),
.B(n_4838),
.Y(n_10176)
);

AOI22xp33_ASAP7_75t_L g10177 ( 
.A1(n_10149),
.A2(n_5286),
.B1(n_4838),
.B2(n_3891),
.Y(n_10177)
);

HB1xp67_ASAP7_75t_L g10178 ( 
.A(n_10155),
.Y(n_10178)
);

NOR3xp33_ASAP7_75t_L g10179 ( 
.A(n_10151),
.B(n_3719),
.C(n_3709),
.Y(n_10179)
);

NAND2xp5_ASAP7_75t_L g10180 ( 
.A(n_10154),
.B(n_5286),
.Y(n_10180)
);

HB1xp67_ASAP7_75t_L g10181 ( 
.A(n_10152),
.Y(n_10181)
);

AOI22xp33_ASAP7_75t_L g10182 ( 
.A1(n_10162),
.A2(n_5286),
.B1(n_3891),
.B2(n_3874),
.Y(n_10182)
);

AOI22xp5_ASAP7_75t_L g10183 ( 
.A1(n_10164),
.A2(n_3784),
.B1(n_3812),
.B2(n_3810),
.Y(n_10183)
);

OAI22xp33_ASAP7_75t_L g10184 ( 
.A1(n_10171),
.A2(n_3786),
.B1(n_3810),
.B2(n_3784),
.Y(n_10184)
);

AND2x4_ASAP7_75t_L g10185 ( 
.A(n_10169),
.B(n_5308),
.Y(n_10185)
);

INVx1_ASAP7_75t_L g10186 ( 
.A(n_10168),
.Y(n_10186)
);

INVx1_ASAP7_75t_L g10187 ( 
.A(n_10178),
.Y(n_10187)
);

INVx1_ASAP7_75t_L g10188 ( 
.A(n_10174),
.Y(n_10188)
);

OR2x2_ASAP7_75t_L g10189 ( 
.A(n_10181),
.B(n_10167),
.Y(n_10189)
);

INVx3_ASAP7_75t_L g10190 ( 
.A(n_10186),
.Y(n_10190)
);

INVx1_ASAP7_75t_L g10191 ( 
.A(n_10172),
.Y(n_10191)
);

INVx1_ASAP7_75t_L g10192 ( 
.A(n_10180),
.Y(n_10192)
);

HB1xp67_ASAP7_75t_L g10193 ( 
.A(n_10176),
.Y(n_10193)
);

INVx1_ASAP7_75t_L g10194 ( 
.A(n_10173),
.Y(n_10194)
);

INVx1_ASAP7_75t_L g10195 ( 
.A(n_10183),
.Y(n_10195)
);

INVx1_ASAP7_75t_L g10196 ( 
.A(n_10184),
.Y(n_10196)
);

INVx1_ASAP7_75t_L g10197 ( 
.A(n_10179),
.Y(n_10197)
);

INVx1_ASAP7_75t_L g10198 ( 
.A(n_10182),
.Y(n_10198)
);

INVx1_ASAP7_75t_L g10199 ( 
.A(n_10187),
.Y(n_10199)
);

AOI21xp5_ASAP7_75t_L g10200 ( 
.A1(n_10188),
.A2(n_10165),
.B(n_10170),
.Y(n_10200)
);

INVx2_ASAP7_75t_L g10201 ( 
.A(n_10189),
.Y(n_10201)
);

OAI21xp33_ASAP7_75t_L g10202 ( 
.A1(n_10191),
.A2(n_10160),
.B(n_10166),
.Y(n_10202)
);

OAI21xp5_ASAP7_75t_L g10203 ( 
.A1(n_10190),
.A2(n_10161),
.B(n_10163),
.Y(n_10203)
);

NAND2xp5_ASAP7_75t_SL g10204 ( 
.A(n_10194),
.B(n_10157),
.Y(n_10204)
);

INVx1_ASAP7_75t_L g10205 ( 
.A(n_10201),
.Y(n_10205)
);

OAI22x1_ASAP7_75t_L g10206 ( 
.A1(n_10199),
.A2(n_10196),
.B1(n_10192),
.B2(n_10193),
.Y(n_10206)
);

OA21x2_ASAP7_75t_L g10207 ( 
.A1(n_10200),
.A2(n_10204),
.B(n_10202),
.Y(n_10207)
);

NAND3xp33_ASAP7_75t_L g10208 ( 
.A(n_10203),
.B(n_10195),
.C(n_10198),
.Y(n_10208)
);

INVx1_ASAP7_75t_L g10209 ( 
.A(n_10205),
.Y(n_10209)
);

OAI21xp5_ASAP7_75t_L g10210 ( 
.A1(n_10208),
.A2(n_10197),
.B(n_10175),
.Y(n_10210)
);

OAI22xp5_ASAP7_75t_SL g10211 ( 
.A1(n_10209),
.A2(n_10207),
.B1(n_10206),
.B2(n_10177),
.Y(n_10211)
);

AOI22xp33_ASAP7_75t_SL g10212 ( 
.A1(n_10211),
.A2(n_10210),
.B1(n_10185),
.B2(n_3784),
.Y(n_10212)
);

AO21x2_ASAP7_75t_L g10213 ( 
.A1(n_10212),
.A2(n_10185),
.B(n_4604),
.Y(n_10213)
);

INVx1_ASAP7_75t_L g10214 ( 
.A(n_10213),
.Y(n_10214)
);

OAI221xp5_ASAP7_75t_R g10215 ( 
.A1(n_10214),
.A2(n_4502),
.B1(n_3952),
.B2(n_3916),
.C(n_5228),
.Y(n_10215)
);

AOI21xp5_ASAP7_75t_L g10216 ( 
.A1(n_10215),
.A2(n_4051),
.B(n_4592),
.Y(n_10216)
);

AOI211xp5_ASAP7_75t_L g10217 ( 
.A1(n_10216),
.A2(n_4111),
.B(n_4107),
.C(n_3844),
.Y(n_10217)
);


endmodule