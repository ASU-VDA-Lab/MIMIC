module fake_ariane_545_n_1864 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1864);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1864;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx2_ASAP7_75t_L g188 ( 
.A(n_29),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_128),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_132),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_176),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_104),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_158),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_89),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_99),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_40),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_64),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_36),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_168),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_75),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_11),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_50),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_138),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_111),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_80),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_2),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_3),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_129),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_103),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_160),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_77),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_4),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_43),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_134),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_177),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_60),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_48),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_180),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_30),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_39),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_137),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_48),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_24),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_47),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_156),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_0),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_30),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_49),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_167),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_65),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_155),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_87),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_0),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_165),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_10),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_92),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_88),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_171),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_23),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_10),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_101),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_17),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_82),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_127),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_100),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_27),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_93),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_121),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_115),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_31),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_110),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_108),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_68),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_72),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_3),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_94),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_122),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_105),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_36),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_120),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_13),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_12),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_26),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_56),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_29),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_107),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_1),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_98),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_146),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_182),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_140),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_84),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_73),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_76),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_56),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_169),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_43),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_37),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_28),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_159),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_179),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_7),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_97),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_183),
.Y(n_285)
);

CKINVDCx6p67_ASAP7_75t_R g286 ( 
.A(n_150),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_50),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_45),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_145),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_112),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_14),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_144),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_62),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_42),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_9),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_147),
.Y(n_296)
);

BUFx5_ASAP7_75t_L g297 ( 
.A(n_67),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_109),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_106),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_172),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_86),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_61),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_123),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_17),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g305 ( 
.A(n_96),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_20),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_118),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_139),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_131),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_157),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_178),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_46),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_59),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_58),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_31),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_38),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_25),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_27),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_164),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_63),
.Y(n_320)
);

BUFx5_ASAP7_75t_L g321 ( 
.A(n_148),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_59),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_46),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_22),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_143),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_53),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_154),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_11),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_78),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_14),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_130),
.Y(n_331)
);

BUFx10_ASAP7_75t_L g332 ( 
.A(n_37),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_44),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_7),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_85),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_173),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_166),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_24),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_35),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_52),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_32),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_162),
.Y(n_342)
);

BUFx10_ASAP7_75t_L g343 ( 
.A(n_170),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_133),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_61),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_60),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_114),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_22),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_5),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_83),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_5),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_12),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_151),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_66),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_136),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_58),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_42),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_81),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_18),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_54),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_153),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_135),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_181),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_23),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_113),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_53),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_71),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_21),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_15),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_119),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_49),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_184),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_116),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_90),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_16),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_161),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_34),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_234),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_234),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_234),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_234),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_247),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_247),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_288),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_283),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_262),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_194),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_247),
.Y(n_388)
);

INVxp33_ASAP7_75t_L g389 ( 
.A(n_198),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_247),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_263),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_262),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_286),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_368),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_368),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_333),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_211),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_206),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_286),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_368),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_368),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_211),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_203),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_215),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_188),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_333),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_202),
.Y(n_407)
);

INVxp33_ASAP7_75t_L g408 ( 
.A(n_201),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_188),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_215),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_217),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_291),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_218),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_237),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_291),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_323),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_323),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_263),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_364),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_224),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_364),
.Y(n_421)
);

INVxp33_ASAP7_75t_L g422 ( 
.A(n_220),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_225),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_248),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_248),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_362),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_228),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_362),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_269),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_221),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_223),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_227),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_240),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_229),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_241),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_206),
.Y(n_436)
);

CKINVDCx14_ASAP7_75t_R g437 ( 
.A(n_191),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_264),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_265),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_250),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_236),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_250),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_268),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_276),
.Y(n_444)
);

BUFx6f_ASAP7_75t_SL g445 ( 
.A(n_269),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_237),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_279),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_271),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_263),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_251),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_256),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_280),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_294),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_260),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_204),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_243),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_314),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_316),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_207),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_317),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_322),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_328),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_338),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_208),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_339),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_340),
.Y(n_466)
);

INVxp33_ASAP7_75t_SL g467 ( 
.A(n_208),
.Y(n_467)
);

INVxp33_ASAP7_75t_SL g468 ( 
.A(n_213),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_231),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_341),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_356),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_360),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_232),
.Y(n_473)
);

INVx6_ASAP7_75t_L g474 ( 
.A(n_387),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_424),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_429),
.B(n_226),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_437),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_440),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_393),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_395),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_430),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_429),
.B(n_235),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_440),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_429),
.B(n_396),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_424),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_406),
.B(n_242),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_399),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_389),
.B(n_332),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_425),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_425),
.Y(n_490)
);

OA21x2_ASAP7_75t_L g491 ( 
.A1(n_426),
.A2(n_254),
.B(n_252),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_440),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_426),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_440),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_440),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_432),
.B(n_444),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_387),
.B(n_226),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_397),
.A2(n_243),
.B1(n_315),
.B2(n_290),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_398),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_442),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_407),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_384),
.Y(n_502)
);

NAND2xp33_ASAP7_75t_L g503 ( 
.A(n_411),
.B(n_377),
.Y(n_503)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_413),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_402),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_430),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_455),
.B(n_253),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_442),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_442),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_431),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_455),
.B(n_459),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_420),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_408),
.B(n_422),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_428),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_431),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_433),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_423),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_404),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_385),
.B(n_212),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_442),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_442),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_428),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_459),
.B(n_253),
.Y(n_523)
);

CKINVDCx8_ASAP7_75t_R g524 ( 
.A(n_391),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_473),
.B(n_212),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_395),
.Y(n_526)
);

NAND3xp33_ASAP7_75t_L g527 ( 
.A(n_386),
.B(n_214),
.C(n_213),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_400),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_400),
.Y(n_529)
);

CKINVDCx8_ASAP7_75t_R g530 ( 
.A(n_418),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_392),
.B(n_332),
.Y(n_531)
);

AOI22x1_ASAP7_75t_SL g532 ( 
.A1(n_410),
.A2(n_315),
.B1(n_214),
.B2(n_366),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_467),
.B(n_212),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_401),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_473),
.B(n_255),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_401),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_433),
.B(n_332),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_403),
.B(n_258),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_378),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_378),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_403),
.B(n_274),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_469),
.B(n_259),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_379),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_469),
.B(n_435),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_468),
.B(n_259),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_379),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_380),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_472),
.B(n_259),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_427),
.B(n_269),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_380),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_381),
.Y(n_551)
);

OR2x6_ASAP7_75t_L g552 ( 
.A(n_449),
.B(n_271),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_381),
.Y(n_553)
);

NAND2xp33_ASAP7_75t_L g554 ( 
.A(n_501),
.B(n_512),
.Y(n_554)
);

BUFx10_ASAP7_75t_L g555 ( 
.A(n_533),
.Y(n_555)
);

INVx11_ASAP7_75t_L g556 ( 
.A(n_524),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_545),
.B(n_434),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_484),
.B(n_445),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_476),
.B(n_441),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_539),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_547),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_537),
.A2(n_445),
.B1(n_464),
.B2(n_436),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_499),
.A2(n_369),
.B1(n_366),
.B2(n_266),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_537),
.A2(n_273),
.B1(n_298),
.B2(n_290),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_547),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_474),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_539),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_513),
.A2(n_445),
.B1(n_273),
.B2(n_303),
.Y(n_568)
);

BUFx10_ASAP7_75t_L g569 ( 
.A(n_501),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_547),
.Y(n_570)
);

NAND2xp33_ASAP7_75t_L g571 ( 
.A(n_512),
.B(n_450),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_513),
.B(n_435),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_474),
.Y(n_573)
);

CKINVDCx6p67_ASAP7_75t_R g574 ( 
.A(n_504),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_540),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_517),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_476),
.B(n_451),
.Y(n_577)
);

AND2x6_ASAP7_75t_L g578 ( 
.A(n_525),
.B(n_488),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_519),
.B(n_454),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_526),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_543),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_543),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_550),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_476),
.B(n_382),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_496),
.B(n_438),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_540),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_550),
.Y(n_587)
);

AO21x2_ASAP7_75t_L g588 ( 
.A1(n_482),
.A2(n_285),
.B(n_277),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_517),
.B(n_205),
.Y(n_589)
);

INVxp67_ASAP7_75t_L g590 ( 
.A(n_488),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_511),
.B(n_438),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_526),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_526),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_526),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_526),
.Y(n_595)
);

OR2x6_ASAP7_75t_L g596 ( 
.A(n_552),
.B(n_439),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_553),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_546),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_511),
.B(n_382),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_511),
.B(n_383),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_546),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_553),
.Y(n_602)
);

NAND2xp33_ASAP7_75t_L g603 ( 
.A(n_477),
.B(n_205),
.Y(n_603)
);

BUFx10_ASAP7_75t_L g604 ( 
.A(n_477),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_544),
.B(n_439),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_534),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_474),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_497),
.B(n_383),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_544),
.B(n_443),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_544),
.A2(n_325),
.B1(n_298),
.B2(n_303),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_551),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_504),
.B(n_210),
.Y(n_612)
);

INVxp33_ASAP7_75t_SL g613 ( 
.A(n_479),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_548),
.B(n_443),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_481),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_497),
.A2(n_308),
.B1(n_325),
.B2(n_331),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_531),
.B(n_479),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_531),
.B(n_210),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_475),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_497),
.B(n_507),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_487),
.B(n_507),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_548),
.B(n_447),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_551),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_507),
.B(n_388),
.Y(n_624)
);

OAI22xp33_ASAP7_75t_L g625 ( 
.A1(n_552),
.A2(n_527),
.B1(n_196),
.B2(n_487),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_551),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_551),
.Y(n_627)
);

INVx1_ASAP7_75t_SL g628 ( 
.A(n_502),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_525),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_523),
.B(n_388),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_551),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_525),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_523),
.B(n_390),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_483),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_483),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_478),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_523),
.Y(n_637)
);

NAND3xp33_ASAP7_75t_L g638 ( 
.A(n_491),
.B(n_219),
.C(n_289),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_494),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_494),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_495),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_495),
.Y(n_642)
);

INVx1_ASAP7_75t_SL g643 ( 
.A(n_505),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_508),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_508),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_475),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_548),
.B(n_390),
.Y(n_647)
);

OR2x6_ASAP7_75t_L g648 ( 
.A(n_552),
.B(n_447),
.Y(n_648)
);

INVx8_ASAP7_75t_L g649 ( 
.A(n_542),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_485),
.Y(n_650)
);

NAND3xp33_ASAP7_75t_L g651 ( 
.A(n_491),
.B(n_301),
.C(n_293),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_485),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_489),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_478),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_518),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_509),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_509),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_489),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_520),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_520),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_506),
.B(n_452),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_510),
.B(n_452),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_478),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_528),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_490),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_528),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_524),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_478),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_502),
.B(n_456),
.Y(n_669)
);

INVx4_ASAP7_75t_L g670 ( 
.A(n_491),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_542),
.B(n_394),
.Y(n_671)
);

BUFx10_ASAP7_75t_L g672 ( 
.A(n_542),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_529),
.Y(n_673)
);

OAI22xp33_ASAP7_75t_L g674 ( 
.A1(n_552),
.A2(n_342),
.B1(n_331),
.B2(n_308),
.Y(n_674)
);

INVx5_ASAP7_75t_L g675 ( 
.A(n_478),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_515),
.B(n_453),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_529),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_549),
.B(n_453),
.Y(n_678)
);

NAND2xp33_ASAP7_75t_L g679 ( 
.A(n_516),
.B(n_299),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_490),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_493),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_486),
.B(n_299),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_536),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_536),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_535),
.B(n_361),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_493),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_491),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_480),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_514),
.B(n_394),
.Y(n_689)
);

BUFx2_ASAP7_75t_L g690 ( 
.A(n_498),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_514),
.Y(n_691)
);

AOI21x1_ASAP7_75t_L g692 ( 
.A1(n_538),
.A2(n_319),
.B(n_310),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_522),
.Y(n_693)
);

INVxp67_ASAP7_75t_SL g694 ( 
.A(n_541),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_480),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_522),
.Y(n_696)
);

BUFx2_ASAP7_75t_L g697 ( 
.A(n_480),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_492),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_492),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_492),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_503),
.B(n_457),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_530),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_492),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_530),
.B(n_472),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_L g705 ( 
.A1(n_578),
.A2(n_342),
.B1(n_365),
.B2(n_361),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_560),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_606),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_567),
.Y(n_708)
);

NAND3xp33_ASAP7_75t_L g709 ( 
.A(n_579),
.B(n_369),
.C(n_287),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_632),
.B(n_365),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_567),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_632),
.B(n_278),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_694),
.B(n_209),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_592),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_585),
.B(n_216),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_592),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_581),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_628),
.B(n_414),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_581),
.Y(n_719)
);

INVxp67_ASAP7_75t_L g720 ( 
.A(n_669),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_558),
.B(n_246),
.Y(n_721)
);

OAI221xp5_ASAP7_75t_L g722 ( 
.A1(n_590),
.A2(n_334),
.B1(n_306),
.B2(n_313),
.C(n_304),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_572),
.B(n_457),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_SL g724 ( 
.A(n_613),
.B(n_446),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_557),
.B(n_295),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_632),
.B(n_302),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_632),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_SL g728 ( 
.A(n_613),
.B(n_702),
.Y(n_728)
);

INVxp33_ASAP7_75t_L g729 ( 
.A(n_669),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_628),
.B(n_448),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_578),
.A2(n_343),
.B1(n_305),
.B2(n_458),
.Y(n_731)
);

INVxp67_ASAP7_75t_L g732 ( 
.A(n_643),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_629),
.B(n_578),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_629),
.B(n_337),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_578),
.A2(n_343),
.B1(n_305),
.B2(n_458),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_688),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_578),
.B(n_460),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_582),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_555),
.B(n_312),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_655),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_555),
.B(n_318),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_572),
.B(n_460),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_655),
.Y(n_743)
);

NAND2xp33_ASAP7_75t_L g744 ( 
.A(n_578),
.B(n_576),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_578),
.B(n_461),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_637),
.B(n_461),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_704),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_583),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_637),
.B(n_462),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_555),
.B(n_324),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_701),
.B(n_462),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_555),
.B(n_326),
.Y(n_752)
);

NAND3xp33_ASAP7_75t_L g753 ( 
.A(n_571),
.B(n_554),
.C(n_576),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_559),
.B(n_330),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_583),
.Y(n_755)
);

BUFx6f_ASAP7_75t_SL g756 ( 
.A(n_604),
.Y(n_756)
);

INVxp67_ASAP7_75t_L g757 ( 
.A(n_704),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_678),
.B(n_463),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_614),
.B(n_463),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_614),
.A2(n_329),
.B1(n_335),
.B2(n_344),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_569),
.B(n_345),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_622),
.A2(n_347),
.B1(n_353),
.B2(n_358),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_672),
.B(n_363),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_577),
.B(n_346),
.Y(n_764)
);

CKINVDCx14_ASAP7_75t_R g765 ( 
.A(n_574),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_569),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_587),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_622),
.B(n_465),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_620),
.B(n_466),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_615),
.B(n_466),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_615),
.B(n_470),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_564),
.B(n_470),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_688),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_591),
.B(n_471),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_618),
.B(n_348),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_621),
.B(n_349),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_564),
.B(n_405),
.Y(n_777)
);

NAND2xp33_ASAP7_75t_L g778 ( 
.A(n_561),
.B(n_351),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_591),
.B(n_352),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_697),
.B(n_357),
.Y(n_780)
);

INVxp67_ASAP7_75t_L g781 ( 
.A(n_697),
.Y(n_781)
);

INVx4_ASAP7_75t_L g782 ( 
.A(n_649),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_587),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_695),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_605),
.B(n_359),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_605),
.B(n_371),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_672),
.B(n_375),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_616),
.B(n_405),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_589),
.B(n_367),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_695),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_619),
.A2(n_374),
.B(n_376),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_609),
.B(n_189),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_672),
.B(n_343),
.Y(n_793)
);

INVx8_ASAP7_75t_L g794 ( 
.A(n_649),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_617),
.B(n_1),
.Y(n_795)
);

OR2x2_ASAP7_75t_L g796 ( 
.A(n_610),
.B(n_409),
.Y(n_796)
);

HB1xp67_ASAP7_75t_L g797 ( 
.A(n_649),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_604),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_670),
.A2(n_419),
.B1(n_412),
.B2(n_415),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_597),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_609),
.B(n_661),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_619),
.A2(n_192),
.B1(n_190),
.B2(n_193),
.Y(n_802)
);

AND2x2_ASAP7_75t_SL g803 ( 
.A(n_568),
.B(n_250),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_661),
.B(n_195),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_616),
.B(n_409),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_662),
.B(n_197),
.Y(n_806)
);

INVx1_ASAP7_75t_SL g807 ( 
.A(n_667),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_592),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_662),
.B(n_199),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_676),
.B(n_200),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_676),
.B(n_222),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_556),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_682),
.B(n_2),
.Y(n_813)
);

INVxp67_ASAP7_75t_L g814 ( 
.A(n_599),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_610),
.B(n_412),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_597),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_602),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_602),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_649),
.B(n_4),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_565),
.Y(n_820)
);

INVx8_ASAP7_75t_L g821 ( 
.A(n_596),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_672),
.B(n_230),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_625),
.B(n_233),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_646),
.B(n_238),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_562),
.B(n_239),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_646),
.B(n_650),
.Y(n_826)
);

AND2x6_ASAP7_75t_L g827 ( 
.A(n_650),
.B(n_250),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_612),
.B(n_6),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_604),
.B(n_674),
.Y(n_829)
);

A2O1A1Ixp33_ASAP7_75t_L g830 ( 
.A1(n_652),
.A2(n_416),
.B(n_415),
.C(n_417),
.Y(n_830)
);

INVx8_ASAP7_75t_L g831 ( 
.A(n_596),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_685),
.B(n_244),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_566),
.B(n_245),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_652),
.B(n_249),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_679),
.A2(n_309),
.B1(n_257),
.B2(n_261),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_653),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_670),
.A2(n_421),
.B1(n_419),
.B2(n_417),
.Y(n_837)
);

NAND2x1_ASAP7_75t_L g838 ( 
.A(n_580),
.B(n_594),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_570),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_566),
.B(n_267),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_658),
.B(n_270),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_658),
.B(n_272),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_665),
.B(n_275),
.Y(n_843)
);

A2O1A1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_665),
.A2(n_421),
.B(n_416),
.C(n_282),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_570),
.Y(n_845)
);

AO22x2_ASAP7_75t_L g846 ( 
.A1(n_638),
.A2(n_532),
.B1(n_8),
.B2(n_9),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_680),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_680),
.B(n_281),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_681),
.B(n_292),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_600),
.B(n_6),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_681),
.B(n_8),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_686),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_686),
.B(n_13),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_R g854 ( 
.A(n_603),
.B(n_296),
.Y(n_854)
);

BUFx2_ASAP7_75t_L g855 ( 
.A(n_596),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_691),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_575),
.Y(n_857)
);

OR2x2_ASAP7_75t_L g858 ( 
.A(n_563),
.B(n_15),
.Y(n_858)
);

INVxp67_ASAP7_75t_SL g859 ( 
.A(n_607),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_691),
.B(n_300),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_740),
.Y(n_861)
);

NAND2xp33_ASAP7_75t_R g862 ( 
.A(n_812),
.B(n_690),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_765),
.Y(n_863)
);

BUFx2_ASAP7_75t_L g864 ( 
.A(n_718),
.Y(n_864)
);

NAND2x1p5_ASAP7_75t_L g865 ( 
.A(n_782),
.B(n_607),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_715),
.B(n_693),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_725),
.B(n_693),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_706),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_743),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_720),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_725),
.B(n_696),
.Y(n_871)
);

INVx4_ASAP7_75t_L g872 ( 
.A(n_794),
.Y(n_872)
);

NOR3xp33_ASAP7_75t_SL g873 ( 
.A(n_753),
.B(n_696),
.C(n_647),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_757),
.B(n_596),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_814),
.B(n_608),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_803),
.A2(n_772),
.B1(n_846),
.B2(n_690),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_708),
.Y(n_877)
);

NOR3xp33_ASAP7_75t_SL g878 ( 
.A(n_739),
.B(n_726),
.C(n_712),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_757),
.B(n_596),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_820),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_803),
.A2(n_846),
.B1(n_777),
.B2(n_735),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_711),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_846),
.A2(n_648),
.B1(n_588),
.B2(n_638),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_717),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_782),
.B(n_727),
.Y(n_885)
);

BUFx2_ASAP7_75t_SL g886 ( 
.A(n_756),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_744),
.A2(n_648),
.B1(n_573),
.B2(n_588),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_719),
.Y(n_888)
);

O2A1O1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_858),
.A2(n_584),
.B(n_689),
.C(n_630),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_738),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_781),
.B(n_648),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_807),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_733),
.B(n_627),
.Y(n_893)
);

AOI22xp5_ASAP7_75t_SL g894 ( 
.A1(n_720),
.A2(n_532),
.B1(n_648),
.B2(n_556),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_748),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_755),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_814),
.B(n_624),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_731),
.A2(n_648),
.B1(n_588),
.B2(n_670),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_741),
.A2(n_573),
.B1(n_633),
.B2(n_631),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_756),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_758),
.B(n_671),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_732),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_730),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_781),
.B(n_670),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_767),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_783),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_729),
.B(n_664),
.Y(n_907)
);

INVxp67_ASAP7_75t_L g908 ( 
.A(n_747),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_731),
.A2(n_687),
.B1(n_651),
.B2(n_683),
.Y(n_909)
);

BUFx2_ASAP7_75t_L g910 ( 
.A(n_732),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_800),
.Y(n_911)
);

A2O1A1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_813),
.A2(n_651),
.B(n_631),
.C(n_627),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_788),
.B(n_664),
.Y(n_913)
);

AO22x1_ASAP7_75t_L g914 ( 
.A1(n_828),
.A2(n_687),
.B1(n_336),
.B2(n_320),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_741),
.A2(n_631),
.B1(n_627),
.B2(n_687),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_727),
.B(n_592),
.Y(n_916)
);

INVxp67_ASAP7_75t_L g917 ( 
.A(n_737),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_839),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_845),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_707),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_R g921 ( 
.A(n_728),
.B(n_692),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_816),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_817),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_818),
.Y(n_924)
);

INVx4_ASAP7_75t_L g925 ( 
.A(n_794),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_794),
.Y(n_926)
);

OR2x6_ASAP7_75t_L g927 ( 
.A(n_821),
.B(n_687),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_713),
.B(n_666),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_836),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_847),
.Y(n_930)
);

OR2x6_ASAP7_75t_L g931 ( 
.A(n_821),
.B(n_666),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_L g932 ( 
.A1(n_852),
.A2(n_580),
.B1(n_594),
.B2(n_626),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_801),
.B(n_594),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_797),
.B(n_611),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_735),
.A2(n_805),
.B1(n_815),
.B2(n_723),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_750),
.B(n_673),
.Y(n_936)
);

AOI22xp5_ASAP7_75t_L g937 ( 
.A1(n_750),
.A2(n_626),
.B1(n_611),
.B2(n_623),
.Y(n_937)
);

NOR3xp33_ASAP7_75t_SL g938 ( 
.A(n_752),
.B(n_307),
.C(n_311),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_856),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_797),
.B(n_592),
.Y(n_940)
);

INVx8_ASAP7_75t_L g941 ( 
.A(n_821),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_752),
.B(n_673),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_826),
.Y(n_943)
);

OR2x6_ASAP7_75t_SL g944 ( 
.A(n_724),
.B(n_327),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_721),
.B(n_723),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_826),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_855),
.B(n_623),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_742),
.Y(n_948)
);

AO22x1_ASAP7_75t_L g949 ( 
.A1(n_828),
.A2(n_372),
.B1(n_373),
.B2(n_370),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_742),
.B(n_769),
.Y(n_950)
);

CKINVDCx11_ASAP7_75t_R g951 ( 
.A(n_831),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_R g952 ( 
.A(n_766),
.B(n_692),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_796),
.B(n_677),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_770),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_785),
.B(n_677),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_819),
.B(n_705),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_831),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_854),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_819),
.B(n_593),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_786),
.B(n_684),
.Y(n_960)
);

NAND3xp33_ASAP7_75t_SL g961 ( 
.A(n_854),
.B(n_350),
.C(n_354),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_831),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_754),
.B(n_575),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_771),
.Y(n_964)
);

INVx1_ASAP7_75t_SL g965 ( 
.A(n_774),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_754),
.B(n_586),
.Y(n_966)
);

INVxp67_ASAP7_75t_L g967 ( 
.A(n_745),
.Y(n_967)
);

NAND3xp33_ASAP7_75t_L g968 ( 
.A(n_813),
.B(n_700),
.C(n_586),
.Y(n_968)
);

OAI21x1_ASAP7_75t_L g969 ( 
.A1(n_857),
.A2(n_654),
.B(n_598),
.Y(n_969)
);

AO22x1_ASAP7_75t_L g970 ( 
.A1(n_795),
.A2(n_355),
.B1(n_601),
.B2(n_598),
.Y(n_970)
);

AND2x2_ASAP7_75t_SL g971 ( 
.A(n_851),
.B(n_284),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_795),
.A2(n_601),
.B1(n_593),
.B2(n_595),
.Y(n_972)
);

AOI22xp33_ASAP7_75t_L g973 ( 
.A1(n_799),
.A2(n_642),
.B1(n_644),
.B2(n_645),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_736),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_764),
.B(n_654),
.Y(n_975)
);

O2A1O1Ixp5_ASAP7_75t_L g976 ( 
.A1(n_851),
.A2(n_654),
.B(n_700),
.C(n_699),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_746),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_764),
.B(n_634),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_714),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_714),
.B(n_593),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_714),
.B(n_595),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_716),
.B(n_595),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_759),
.B(n_768),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_SL g984 ( 
.A(n_798),
.B(n_634),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_773),
.Y(n_985)
);

INVx1_ASAP7_75t_SL g986 ( 
.A(n_779),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_749),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_776),
.B(n_635),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_L g989 ( 
.A1(n_799),
.A2(n_642),
.B1(n_644),
.B2(n_635),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_751),
.B(n_639),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_716),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_734),
.B(n_595),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_784),
.Y(n_993)
);

INVx1_ASAP7_75t_SL g994 ( 
.A(n_780),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_790),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_716),
.Y(n_996)
);

INVx5_ASAP7_75t_L g997 ( 
.A(n_716),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_789),
.B(n_804),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_789),
.B(n_639),
.Y(n_999)
);

AOI22xp33_ASAP7_75t_L g1000 ( 
.A1(n_837),
.A2(n_656),
.B1(n_640),
.B2(n_641),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_806),
.B(n_640),
.Y(n_1001)
);

INVx2_ASAP7_75t_SL g1002 ( 
.A(n_829),
.Y(n_1002)
);

AOI22xp33_ASAP7_75t_SL g1003 ( 
.A1(n_775),
.A2(n_284),
.B1(n_297),
.B2(n_321),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_809),
.B(n_641),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_810),
.B(n_645),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_811),
.B(n_656),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_830),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_859),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_761),
.B(n_657),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_853),
.Y(n_1010)
);

INVxp67_ASAP7_75t_SL g1011 ( 
.A(n_859),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_853),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_850),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_838),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_792),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_837),
.B(n_657),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_850),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_787),
.B(n_659),
.Y(n_1018)
);

INVx6_ASAP7_75t_L g1019 ( 
.A(n_808),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_824),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_760),
.B(n_659),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_762),
.B(n_660),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_808),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_775),
.B(n_660),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_776),
.B(n_703),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_832),
.Y(n_1026)
);

INVx2_ASAP7_75t_SL g1027 ( 
.A(n_793),
.Y(n_1027)
);

OAI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_722),
.A2(n_703),
.B1(n_699),
.B2(n_698),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_834),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_860),
.Y(n_1030)
);

AOI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_763),
.A2(n_698),
.B1(n_668),
.B2(n_663),
.Y(n_1031)
);

INVx2_ASAP7_75t_SL g1032 ( 
.A(n_833),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_763),
.B(n_668),
.Y(n_1033)
);

OR2x6_ASAP7_75t_L g1034 ( 
.A(n_825),
.B(n_636),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_SL g1035 ( 
.A(n_827),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_709),
.B(n_823),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_920),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_867),
.A2(n_822),
.B(n_849),
.Y(n_1038)
);

NAND2x1_ASAP7_75t_L g1039 ( 
.A(n_872),
.B(n_636),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_1015),
.B(n_710),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_1010),
.A2(n_848),
.B1(n_843),
.B2(n_842),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_R g1042 ( 
.A(n_863),
.B(n_778),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_1012),
.A2(n_841),
.B1(n_791),
.B2(n_844),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_965),
.B(n_802),
.Y(n_1044)
);

NOR3xp33_ASAP7_75t_SL g1045 ( 
.A(n_958),
.B(n_840),
.C(n_18),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_994),
.B(n_835),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_1013),
.A2(n_636),
.B1(n_663),
.B2(n_668),
.Y(n_1047)
);

AND2x2_ASAP7_75t_SL g1048 ( 
.A(n_881),
.B(n_284),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_953),
.B(n_827),
.Y(n_1049)
);

AND2x4_ASAP7_75t_SL g1050 ( 
.A(n_926),
.B(n_636),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_868),
.Y(n_1051)
);

HB1xp67_ASAP7_75t_L g1052 ( 
.A(n_910),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_986),
.B(n_636),
.Y(n_1053)
);

OR2x6_ASAP7_75t_SL g1054 ( 
.A(n_900),
.B(n_902),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_1017),
.A2(n_16),
.B(n_19),
.C(n_20),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_983),
.A2(n_663),
.B1(n_668),
.B2(n_675),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_945),
.B(n_663),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_SL g1058 ( 
.A1(n_933),
.A2(n_675),
.B(n_827),
.C(n_25),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_941),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_1011),
.A2(n_668),
.B(n_663),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_998),
.B(n_874),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_1011),
.A2(n_675),
.B(n_284),
.Y(n_1062)
);

NOR2x1_ASAP7_75t_SL g1063 ( 
.A(n_927),
.B(n_675),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_866),
.A2(n_675),
.B(n_521),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_913),
.B(n_827),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_874),
.B(n_19),
.Y(n_1066)
);

INVx1_ASAP7_75t_SL g1067 ( 
.A(n_892),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_950),
.B(n_827),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_SL g1069 ( 
.A1(n_876),
.A2(n_21),
.B1(n_26),
.B2(n_28),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_935),
.B(n_675),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_935),
.B(n_32),
.Y(n_1071)
);

NAND2xp33_ASAP7_75t_SL g1072 ( 
.A(n_872),
.B(n_33),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_SL g1073 ( 
.A1(n_876),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_957),
.B(n_38),
.Y(n_1074)
);

OAI22x1_ASAP7_75t_L g1075 ( 
.A1(n_879),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_1075)
);

INVx1_ASAP7_75t_SL g1076 ( 
.A(n_864),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_SL g1077 ( 
.A(n_971),
.B(n_321),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_969),
.A2(n_297),
.B(n_321),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_903),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_879),
.B(n_41),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_861),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_1017),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_926),
.B(n_521),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_870),
.B(n_51),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_877),
.Y(n_1085)
);

BUFx2_ASAP7_75t_R g1086 ( 
.A(n_944),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_956),
.A2(n_51),
.B(n_52),
.C(n_54),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_948),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_870),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_882),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_1020),
.B(n_55),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_SL g1092 ( 
.A1(n_894),
.A2(n_321),
.B1(n_297),
.B2(n_55),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_1029),
.B(n_57),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_1030),
.B(n_57),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_956),
.A2(n_891),
.B1(n_971),
.B2(n_862),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_884),
.Y(n_1096)
);

OAI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_976),
.A2(n_321),
.B(n_297),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_977),
.B(n_321),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_948),
.B(n_521),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_987),
.B(n_297),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_875),
.B(n_297),
.Y(n_1101)
);

OA22x2_ASAP7_75t_L g1102 ( 
.A1(n_908),
.A2(n_69),
.B1(n_70),
.B2(n_74),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_891),
.B(n_521),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_908),
.B(n_1002),
.Y(n_1104)
);

AOI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_862),
.A2(n_521),
.B1(n_500),
.B2(n_95),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_926),
.B(n_500),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_869),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_975),
.A2(n_500),
.B(n_91),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_881),
.A2(n_500),
.B1(n_102),
.B2(n_117),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_888),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_941),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_936),
.A2(n_79),
.B(n_124),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_942),
.A2(n_125),
.B(n_126),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_897),
.B(n_141),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_890),
.Y(n_1115)
);

OAI21xp33_ASAP7_75t_L g1116 ( 
.A1(n_904),
.A2(n_142),
.B(n_149),
.Y(n_1116)
);

BUFx3_ASAP7_75t_L g1117 ( 
.A(n_951),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_1036),
.A2(n_152),
.B(n_163),
.C(n_174),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_895),
.Y(n_1119)
);

AOI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1036),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_963),
.A2(n_966),
.B(n_978),
.Y(n_1121)
);

BUFx4f_ASAP7_75t_L g1122 ( 
.A(n_941),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_1025),
.A2(n_904),
.B(n_933),
.C(n_955),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_880),
.Y(n_1124)
);

OAI21xp33_ASAP7_75t_L g1125 ( 
.A1(n_938),
.A2(n_946),
.B(n_943),
.Y(n_1125)
);

OR2x6_ASAP7_75t_L g1126 ( 
.A(n_931),
.B(n_927),
.Y(n_1126)
);

NAND2xp33_ASAP7_75t_L g1127 ( 
.A(n_926),
.B(n_1008),
.Y(n_1127)
);

INVx5_ASAP7_75t_L g1128 ( 
.A(n_927),
.Y(n_1128)
);

AO32x2_ASAP7_75t_L g1129 ( 
.A1(n_932),
.A2(n_1027),
.A3(n_1026),
.B1(n_1032),
.B2(n_883),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_1025),
.A2(n_960),
.B(n_964),
.C(n_954),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_925),
.B(n_934),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_896),
.A2(n_939),
.B1(n_922),
.B2(n_911),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_925),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_918),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1008),
.B(n_907),
.Y(n_1135)
);

NOR2xp67_ASAP7_75t_L g1136 ( 
.A(n_961),
.B(n_905),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_906),
.Y(n_1137)
);

INVx3_ASAP7_75t_L g1138 ( 
.A(n_1019),
.Y(n_1138)
);

AOI22x1_ASAP7_75t_L g1139 ( 
.A1(n_923),
.A2(n_929),
.B1(n_924),
.B2(n_930),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_901),
.B(n_988),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_919),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_917),
.B(n_967),
.Y(n_1142)
);

OAI21xp33_ASAP7_75t_SL g1143 ( 
.A1(n_915),
.A2(n_899),
.B(n_959),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_SL g1144 ( 
.A(n_931),
.B(n_997),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_976),
.A2(n_912),
.B(n_1007),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_980),
.A2(n_982),
.B(n_981),
.Y(n_1146)
);

OR2x6_ASAP7_75t_L g1147 ( 
.A(n_931),
.B(n_886),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_974),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_928),
.B(n_949),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_993),
.Y(n_1150)
);

CKINVDCx11_ASAP7_75t_R g1151 ( 
.A(n_979),
.Y(n_1151)
);

AOI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_883),
.A2(n_1003),
.B1(n_898),
.B2(n_985),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_947),
.B(n_878),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_1019),
.Y(n_1154)
);

OAI22x1_ASAP7_75t_L g1155 ( 
.A1(n_887),
.A2(n_1018),
.B1(n_1009),
.B2(n_947),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_SL g1156 ( 
.A1(n_996),
.A2(n_984),
.B(n_937),
.C(n_1023),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_934),
.B(n_889),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_995),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_878),
.B(n_938),
.Y(n_1159)
);

INVx6_ASAP7_75t_L g1160 ( 
.A(n_997),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_898),
.B(n_999),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_R g1162 ( 
.A(n_997),
.B(n_1019),
.Y(n_1162)
);

A2O1A1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_1003),
.A2(n_968),
.B(n_873),
.C(n_959),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_1014),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_980),
.A2(n_981),
.B(n_982),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1021),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_970),
.B(n_1004),
.Y(n_1167)
);

NAND2x1p5_ASAP7_75t_L g1168 ( 
.A(n_996),
.B(n_991),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1024),
.B(n_1018),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1009),
.B(n_1006),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1022),
.Y(n_1171)
);

NOR3xp33_ASAP7_75t_SL g1172 ( 
.A(n_1028),
.B(n_916),
.C(n_885),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_873),
.A2(n_909),
.B1(n_1016),
.B2(n_1001),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_909),
.A2(n_1005),
.B1(n_1028),
.B2(n_972),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_990),
.B(n_991),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_940),
.A2(n_893),
.B(n_992),
.C(n_1033),
.Y(n_1176)
);

AND2x2_ASAP7_75t_SL g1177 ( 
.A(n_979),
.B(n_991),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_921),
.Y(n_1178)
);

O2A1O1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1034),
.A2(n_865),
.B(n_973),
.C(n_1000),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_921),
.B(n_973),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_979),
.B(n_952),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1031),
.A2(n_989),
.B(n_1000),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_989),
.B(n_952),
.Y(n_1183)
);

AO31x2_ASAP7_75t_L g1184 ( 
.A1(n_1121),
.A2(n_1035),
.A3(n_1174),
.B(n_1173),
.Y(n_1184)
);

AO21x2_ASAP7_75t_L g1185 ( 
.A1(n_1097),
.A2(n_1161),
.B(n_1145),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1123),
.A2(n_1047),
.B(n_1056),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1037),
.Y(n_1187)
);

O2A1O1Ixp5_ASAP7_75t_SL g1188 ( 
.A1(n_1097),
.A2(n_1082),
.B(n_1109),
.C(n_1041),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1078),
.A2(n_1165),
.B(n_1146),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1061),
.B(n_1140),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1051),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1089),
.B(n_1088),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_SL g1193 ( 
.A1(n_1092),
.A2(n_1082),
.B(n_1080),
.Y(n_1193)
);

OAI21xp33_ASAP7_75t_SL g1194 ( 
.A1(n_1048),
.A2(n_1102),
.B(n_1066),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1077),
.A2(n_1095),
.B(n_1093),
.C(n_1094),
.Y(n_1195)
);

CKINVDCx8_ASAP7_75t_R g1196 ( 
.A(n_1079),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1166),
.B(n_1171),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1169),
.B(n_1130),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_SL g1199 ( 
.A1(n_1109),
.A2(n_1179),
.B(n_1102),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1047),
.A2(n_1056),
.B(n_1077),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1145),
.A2(n_1060),
.B(n_1108),
.Y(n_1201)
);

NOR2x1_ASAP7_75t_L g1202 ( 
.A(n_1081),
.B(n_1117),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1176),
.A2(n_1062),
.B(n_1064),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_1107),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_1046),
.B(n_1149),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_SL g1206 ( 
.A1(n_1055),
.A2(n_1084),
.B(n_1087),
.Y(n_1206)
);

AO31x2_ASAP7_75t_L g1207 ( 
.A1(n_1174),
.A2(n_1173),
.A3(n_1155),
.B(n_1163),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1040),
.B(n_1044),
.Y(n_1208)
);

AO31x2_ASAP7_75t_L g1209 ( 
.A1(n_1182),
.A2(n_1041),
.A3(n_1043),
.B(n_1167),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1038),
.A2(n_1116),
.B(n_1127),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1181),
.A2(n_1112),
.B(n_1113),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1170),
.B(n_1180),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1135),
.B(n_1076),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1052),
.B(n_1104),
.Y(n_1214)
);

INVx1_ASAP7_75t_SL g1215 ( 
.A(n_1067),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_SL g1216 ( 
.A(n_1162),
.B(n_1157),
.Y(n_1216)
);

O2A1O1Ixp5_ASAP7_75t_SL g1217 ( 
.A1(n_1043),
.A2(n_1132),
.B(n_1150),
.C(n_1158),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1076),
.B(n_1142),
.Y(n_1218)
);

INVxp67_ASAP7_75t_SL g1219 ( 
.A(n_1053),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1091),
.A2(n_1071),
.B(n_1136),
.C(n_1143),
.Y(n_1220)
);

INVx5_ASAP7_75t_L g1221 ( 
.A(n_1126),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_1067),
.B(n_1122),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_SL g1223 ( 
.A1(n_1114),
.A2(n_1183),
.B(n_1175),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1069),
.A2(n_1073),
.B1(n_1139),
.B2(n_1132),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1122),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1070),
.A2(n_1098),
.B(n_1100),
.Y(n_1226)
);

BUFx10_ASAP7_75t_L g1227 ( 
.A(n_1074),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1159),
.A2(n_1152),
.B1(n_1119),
.B2(n_1137),
.Y(n_1228)
);

NAND3xp33_ASAP7_75t_SL g1229 ( 
.A(n_1045),
.B(n_1042),
.C(n_1072),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_1177),
.B(n_1178),
.Y(n_1230)
);

INVx1_ASAP7_75t_SL g1231 ( 
.A(n_1151),
.Y(n_1231)
);

NAND3xp33_ASAP7_75t_L g1232 ( 
.A(n_1125),
.B(n_1172),
.C(n_1120),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_1164),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1059),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1059),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1085),
.B(n_1096),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1153),
.B(n_1115),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1156),
.A2(n_1103),
.B(n_1144),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1090),
.A2(n_1110),
.B1(n_1105),
.B2(n_1126),
.Y(n_1239)
);

A2O1A1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1057),
.A2(n_1068),
.B(n_1101),
.C(n_1118),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_1160),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1168),
.A2(n_1039),
.B(n_1083),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1144),
.A2(n_1058),
.B(n_1131),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1106),
.A2(n_1126),
.B(n_1063),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1065),
.A2(n_1050),
.B(n_1049),
.Y(n_1245)
);

BUFx12f_ASAP7_75t_L g1246 ( 
.A(n_1059),
.Y(n_1246)
);

A2O1A1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_1099),
.A2(n_1138),
.B(n_1154),
.C(n_1141),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1138),
.A2(n_1154),
.B(n_1134),
.C(n_1148),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1133),
.A2(n_1128),
.B(n_1147),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1133),
.A2(n_1124),
.B(n_1128),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1129),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1111),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1128),
.A2(n_1086),
.B1(n_1160),
.B2(n_1111),
.Y(n_1253)
);

AO31x2_ASAP7_75t_L g1254 ( 
.A1(n_1075),
.A2(n_1121),
.A3(n_1174),
.B(n_1173),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1129),
.Y(n_1255)
);

AOI21xp33_ASAP7_75t_L g1256 ( 
.A1(n_1128),
.A2(n_1048),
.B(n_1077),
.Y(n_1256)
);

INVx5_ASAP7_75t_L g1257 ( 
.A(n_1129),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1061),
.B(n_1140),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1061),
.B(n_1140),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1061),
.B(n_965),
.Y(n_1260)
);

AO31x2_ASAP7_75t_L g1261 ( 
.A1(n_1121),
.A2(n_1174),
.A3(n_1173),
.B(n_1109),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1061),
.B(n_1140),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1089),
.B(n_720),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1046),
.B(n_613),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1126),
.B(n_962),
.Y(n_1265)
);

OAI21xp33_ASAP7_75t_L g1266 ( 
.A1(n_1066),
.A2(n_725),
.B(n_613),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1061),
.B(n_965),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1121),
.A2(n_871),
.B(n_867),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1121),
.A2(n_871),
.B(n_867),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1061),
.B(n_965),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1061),
.B(n_1140),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1123),
.A2(n_1145),
.B(n_976),
.Y(n_1272)
);

NAND3xp33_ASAP7_75t_L g1273 ( 
.A(n_1066),
.B(n_725),
.C(n_545),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_1117),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1048),
.A2(n_1010),
.B1(n_1012),
.B2(n_935),
.Y(n_1275)
);

AND2x2_ASAP7_75t_SL g1276 ( 
.A(n_1048),
.B(n_881),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1046),
.B(n_613),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1061),
.B(n_965),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1117),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1051),
.Y(n_1280)
);

AND2x6_ASAP7_75t_SL g1281 ( 
.A(n_1046),
.B(n_552),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1061),
.B(n_965),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_1042),
.Y(n_1283)
);

OAI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1123),
.A2(n_1145),
.B(n_976),
.Y(n_1284)
);

AO21x1_ASAP7_75t_L g1285 ( 
.A1(n_1077),
.A2(n_1109),
.B(n_956),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1078),
.A2(n_969),
.B(n_1146),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1121),
.A2(n_871),
.B(n_867),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1117),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_1151),
.Y(n_1289)
);

NAND3xp33_ASAP7_75t_SL g1290 ( 
.A(n_1092),
.B(n_576),
.C(n_512),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1061),
.B(n_965),
.Y(n_1291)
);

NAND3xp33_ASAP7_75t_L g1292 ( 
.A(n_1066),
.B(n_725),
.C(n_545),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1061),
.B(n_965),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1061),
.B(n_965),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1123),
.A2(n_1145),
.B(n_976),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1117),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1061),
.B(n_1140),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1051),
.Y(n_1298)
);

AO31x2_ASAP7_75t_L g1299 ( 
.A1(n_1121),
.A2(n_1174),
.A3(n_1173),
.B(n_1109),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1126),
.B(n_962),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1061),
.B(n_1140),
.Y(n_1301)
);

AO31x2_ASAP7_75t_L g1302 ( 
.A1(n_1121),
.A2(n_1174),
.A3(n_1173),
.B(n_1109),
.Y(n_1302)
);

AOI221x1_ASAP7_75t_L g1303 ( 
.A1(n_1109),
.A2(n_1069),
.B1(n_1073),
.B2(n_1075),
.C(n_1163),
.Y(n_1303)
);

BUFx2_ASAP7_75t_SL g1304 ( 
.A(n_1117),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1042),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1051),
.Y(n_1306)
);

OAI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1123),
.A2(n_1145),
.B(n_976),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1046),
.B(n_613),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1061),
.B(n_1140),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1046),
.B(n_613),
.Y(n_1310)
);

AO31x2_ASAP7_75t_L g1311 ( 
.A1(n_1121),
.A2(n_1174),
.A3(n_1173),
.B(n_1109),
.Y(n_1311)
);

INVx1_ASAP7_75t_SL g1312 ( 
.A(n_1079),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1061),
.B(n_1140),
.Y(n_1313)
);

AOI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1046),
.A2(n_576),
.B1(n_724),
.B2(n_628),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1061),
.B(n_1140),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1061),
.B(n_1140),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1122),
.Y(n_1317)
);

OAI22x1_ASAP7_75t_L g1318 ( 
.A1(n_1095),
.A2(n_610),
.B1(n_616),
.B2(n_564),
.Y(n_1318)
);

AO31x2_ASAP7_75t_L g1319 ( 
.A1(n_1121),
.A2(n_1174),
.A3(n_1173),
.B(n_1109),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_1122),
.Y(n_1320)
);

OAI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1123),
.A2(n_1145),
.B(n_976),
.Y(n_1321)
);

O2A1O1Ixp5_ASAP7_75t_L g1322 ( 
.A1(n_1145),
.A2(n_914),
.B(n_956),
.C(n_949),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1121),
.A2(n_871),
.B(n_867),
.Y(n_1323)
);

INVxp67_ASAP7_75t_L g1324 ( 
.A(n_1079),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1151),
.Y(n_1325)
);

BUFx2_ASAP7_75t_R g1326 ( 
.A(n_1054),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1190),
.B(n_1258),
.Y(n_1327)
);

NOR2x1_ASAP7_75t_L g1328 ( 
.A(n_1229),
.B(n_1222),
.Y(n_1328)
);

NAND2x1p5_ASAP7_75t_L g1329 ( 
.A(n_1221),
.B(n_1216),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1221),
.B(n_1265),
.Y(n_1330)
);

OA21x2_ASAP7_75t_L g1331 ( 
.A1(n_1201),
.A2(n_1186),
.B(n_1189),
.Y(n_1331)
);

AOI21xp33_ASAP7_75t_SL g1332 ( 
.A1(n_1264),
.A2(n_1308),
.B(n_1277),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1273),
.A2(n_1292),
.B(n_1188),
.Y(n_1333)
);

OA21x2_ASAP7_75t_L g1334 ( 
.A1(n_1272),
.A2(n_1295),
.B(n_1284),
.Y(n_1334)
);

OA21x2_ASAP7_75t_L g1335 ( 
.A1(n_1272),
.A2(n_1295),
.B(n_1284),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1193),
.A2(n_1276),
.B1(n_1275),
.B2(n_1199),
.Y(n_1336)
);

OR2x6_ASAP7_75t_L g1337 ( 
.A(n_1253),
.B(n_1249),
.Y(n_1337)
);

BUFx12f_ASAP7_75t_L g1338 ( 
.A(n_1305),
.Y(n_1338)
);

A2O1A1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1194),
.A2(n_1193),
.B(n_1200),
.C(n_1195),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1191),
.Y(n_1340)
);

AO31x2_ASAP7_75t_L g1341 ( 
.A1(n_1285),
.A2(n_1251),
.A3(n_1240),
.B(n_1303),
.Y(n_1341)
);

AOI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1310),
.A2(n_1266),
.B1(n_1314),
.B2(n_1224),
.Y(n_1342)
);

INVx6_ASAP7_75t_L g1343 ( 
.A(n_1246),
.Y(n_1343)
);

OA21x2_ASAP7_75t_L g1344 ( 
.A1(n_1307),
.A2(n_1321),
.B(n_1286),
.Y(n_1344)
);

INVx2_ASAP7_75t_SL g1345 ( 
.A(n_1233),
.Y(n_1345)
);

AO21x2_ASAP7_75t_L g1346 ( 
.A1(n_1256),
.A2(n_1223),
.B(n_1238),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1211),
.A2(n_1226),
.B(n_1210),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1192),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_SL g1349 ( 
.A(n_1256),
.B(n_1275),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1190),
.B(n_1258),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1217),
.A2(n_1287),
.B(n_1323),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1221),
.B(n_1265),
.Y(n_1352)
);

INVx3_ASAP7_75t_L g1353 ( 
.A(n_1225),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1245),
.A2(n_1307),
.B(n_1321),
.Y(n_1354)
);

OA21x2_ASAP7_75t_L g1355 ( 
.A1(n_1322),
.A2(n_1220),
.B(n_1198),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1318),
.A2(n_1224),
.B1(n_1228),
.B2(n_1290),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1250),
.A2(n_1243),
.B(n_1242),
.Y(n_1357)
);

AO31x2_ASAP7_75t_L g1358 ( 
.A1(n_1255),
.A2(n_1228),
.A3(n_1239),
.B(n_1198),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1221),
.B(n_1300),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1232),
.A2(n_1206),
.B(n_1297),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1206),
.A2(n_1297),
.B(n_1301),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1244),
.A2(n_1239),
.B(n_1197),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1259),
.B(n_1262),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1197),
.A2(n_1298),
.B(n_1306),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1185),
.A2(n_1271),
.B(n_1259),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1185),
.A2(n_1301),
.B(n_1262),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1271),
.A2(n_1316),
.B(n_1309),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1280),
.A2(n_1230),
.B(n_1237),
.Y(n_1368)
);

OA21x2_ASAP7_75t_L g1369 ( 
.A1(n_1247),
.A2(n_1248),
.B(n_1212),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1253),
.A2(n_1205),
.B(n_1219),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1309),
.B(n_1313),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1213),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1218),
.Y(n_1373)
);

CKINVDCx11_ASAP7_75t_R g1374 ( 
.A(n_1196),
.Y(n_1374)
);

OA21x2_ASAP7_75t_L g1375 ( 
.A1(n_1313),
.A2(n_1316),
.B(n_1315),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1315),
.A2(n_1208),
.B1(n_1293),
.B2(n_1291),
.Y(n_1376)
);

NAND3xp33_ASAP7_75t_L g1377 ( 
.A(n_1260),
.B(n_1270),
.C(n_1267),
.Y(n_1377)
);

AOI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1278),
.A2(n_1282),
.B(n_1294),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1209),
.B(n_1207),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1209),
.Y(n_1380)
);

INVxp67_ASAP7_75t_SL g1381 ( 
.A(n_1263),
.Y(n_1381)
);

AO32x2_ASAP7_75t_L g1382 ( 
.A1(n_1257),
.A2(n_1209),
.A3(n_1207),
.B1(n_1311),
.B2(n_1319),
.Y(n_1382)
);

NAND2x1p5_ASAP7_75t_L g1383 ( 
.A(n_1215),
.B(n_1312),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1317),
.A2(n_1320),
.B(n_1241),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1312),
.A2(n_1324),
.B1(n_1214),
.B2(n_1257),
.Y(n_1385)
);

OAI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1252),
.A2(n_1261),
.B(n_1299),
.Y(n_1386)
);

NOR2x1_ASAP7_75t_SL g1387 ( 
.A(n_1289),
.B(n_1325),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_SL g1388 ( 
.A1(n_1202),
.A2(n_1288),
.B(n_1326),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1257),
.A2(n_1299),
.B(n_1302),
.Y(n_1389)
);

O2A1O1Ixp33_ASAP7_75t_SL g1390 ( 
.A1(n_1231),
.A2(n_1319),
.B(n_1311),
.C(n_1302),
.Y(n_1390)
);

NAND2x1p5_ASAP7_75t_L g1391 ( 
.A(n_1289),
.B(n_1325),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1254),
.B(n_1302),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1235),
.B(n_1234),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1254),
.B(n_1319),
.Y(n_1394)
);

OA21x2_ASAP7_75t_L g1395 ( 
.A1(n_1184),
.A2(n_1281),
.B(n_1227),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1234),
.A2(n_1304),
.B(n_1204),
.Y(n_1396)
);

NAND2x1p5_ASAP7_75t_L g1397 ( 
.A(n_1325),
.B(n_1274),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1279),
.A2(n_1200),
.B(n_1268),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1296),
.A2(n_1203),
.B(n_1189),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1318),
.A2(n_803),
.B1(n_1048),
.B2(n_1276),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1203),
.A2(n_1189),
.B(n_1201),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1190),
.B(n_1258),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1193),
.A2(n_1048),
.B1(n_1292),
.B2(n_1273),
.Y(n_1403)
);

OA21x2_ASAP7_75t_L g1404 ( 
.A1(n_1201),
.A2(n_1186),
.B(n_1189),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1203),
.A2(n_1189),
.B(n_1201),
.Y(n_1405)
);

INVx3_ASAP7_75t_L g1406 ( 
.A(n_1225),
.Y(n_1406)
);

AOI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1193),
.A2(n_1264),
.B1(n_1308),
.B2(n_1277),
.Y(n_1407)
);

AO21x1_ASAP7_75t_L g1408 ( 
.A1(n_1224),
.A2(n_1193),
.B(n_1275),
.Y(n_1408)
);

INVx4_ASAP7_75t_SL g1409 ( 
.A(n_1207),
.Y(n_1409)
);

AO21x2_ASAP7_75t_L g1410 ( 
.A1(n_1200),
.A2(n_1285),
.B(n_1199),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1236),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1236),
.Y(n_1412)
);

BUFx3_ASAP7_75t_L g1413 ( 
.A(n_1233),
.Y(n_1413)
);

NAND3xp33_ASAP7_75t_L g1414 ( 
.A(n_1273),
.B(n_1292),
.C(n_1266),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1283),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1193),
.A2(n_1048),
.B1(n_1292),
.B2(n_1273),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1236),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1236),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1236),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1221),
.B(n_1265),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1209),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1273),
.A2(n_1292),
.B(n_1188),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1187),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1236),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1193),
.A2(n_1048),
.B1(n_1292),
.B2(n_1273),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_L g1426 ( 
.A(n_1266),
.B(n_1273),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1212),
.B(n_1213),
.Y(n_1427)
);

AOI21xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1264),
.A2(n_576),
.B(n_613),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1283),
.Y(n_1429)
);

AND2x2_ASAP7_75t_SL g1430 ( 
.A(n_1276),
.B(n_1048),
.Y(n_1430)
);

INVx6_ASAP7_75t_L g1431 ( 
.A(n_1246),
.Y(n_1431)
);

OA21x2_ASAP7_75t_L g1432 ( 
.A1(n_1201),
.A2(n_1186),
.B(n_1189),
.Y(n_1432)
);

OR2x6_ASAP7_75t_L g1433 ( 
.A(n_1199),
.B(n_1126),
.Y(n_1433)
);

AO31x2_ASAP7_75t_L g1434 ( 
.A1(n_1285),
.A2(n_1109),
.A3(n_1251),
.B(n_1174),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1318),
.A2(n_803),
.B1(n_1048),
.B2(n_1276),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1221),
.B(n_1265),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1203),
.A2(n_1189),
.B(n_1201),
.Y(n_1437)
);

NAND3xp33_ASAP7_75t_L g1438 ( 
.A(n_1273),
.B(n_1292),
.C(n_1266),
.Y(n_1438)
);

NOR2xp67_ASAP7_75t_SL g1439 ( 
.A(n_1289),
.B(n_1325),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1193),
.A2(n_1048),
.B1(n_1292),
.B2(n_1273),
.Y(n_1440)
);

CKINVDCx11_ASAP7_75t_R g1441 ( 
.A(n_1196),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1187),
.Y(n_1442)
);

O2A1O1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1266),
.A2(n_1193),
.B(n_1292),
.C(n_1273),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1200),
.A2(n_1269),
.B(n_1268),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1209),
.Y(n_1445)
);

NAND3xp33_ASAP7_75t_SL g1446 ( 
.A(n_1266),
.B(n_1292),
.C(n_1273),
.Y(n_1446)
);

OR2x6_ASAP7_75t_L g1447 ( 
.A(n_1199),
.B(n_1126),
.Y(n_1447)
);

BUFx6f_ASAP7_75t_L g1448 ( 
.A(n_1246),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1221),
.B(n_1265),
.Y(n_1449)
);

OR2x6_ASAP7_75t_L g1450 ( 
.A(n_1199),
.B(n_1126),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1212),
.B(n_1213),
.Y(n_1451)
);

A2O1A1Ixp33_ASAP7_75t_L g1452 ( 
.A1(n_1194),
.A2(n_1193),
.B(n_1200),
.C(n_1195),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1342),
.A2(n_1407),
.B1(n_1425),
.B2(n_1440),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1381),
.B(n_1348),
.Y(n_1454)
);

INVx3_ASAP7_75t_L g1455 ( 
.A(n_1396),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_1413),
.Y(n_1456)
);

O2A1O1Ixp33_ASAP7_75t_L g1457 ( 
.A1(n_1403),
.A2(n_1416),
.B(n_1440),
.C(n_1425),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1330),
.B(n_1352),
.Y(n_1458)
);

O2A1O1Ixp33_ASAP7_75t_L g1459 ( 
.A1(n_1403),
.A2(n_1416),
.B(n_1443),
.C(n_1446),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1365),
.B(n_1366),
.Y(n_1460)
);

OR2x6_ASAP7_75t_L g1461 ( 
.A(n_1337),
.B(n_1433),
.Y(n_1461)
);

O2A1O1Ixp5_ASAP7_75t_L g1462 ( 
.A1(n_1408),
.A2(n_1452),
.B(n_1339),
.C(n_1336),
.Y(n_1462)
);

O2A1O1Ixp5_ASAP7_75t_L g1463 ( 
.A1(n_1339),
.A2(n_1452),
.B(n_1336),
.C(n_1360),
.Y(n_1463)
);

BUFx3_ASAP7_75t_L g1464 ( 
.A(n_1397),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1365),
.B(n_1366),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1360),
.A2(n_1356),
.B1(n_1430),
.B2(n_1361),
.Y(n_1466)
);

NOR2xp67_ASAP7_75t_L g1467 ( 
.A(n_1377),
.B(n_1376),
.Y(n_1467)
);

OA21x2_ASAP7_75t_L g1468 ( 
.A1(n_1351),
.A2(n_1347),
.B(n_1444),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1375),
.B(n_1376),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1375),
.B(n_1327),
.Y(n_1470)
);

O2A1O1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1443),
.A2(n_1446),
.B(n_1332),
.C(n_1426),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1327),
.B(n_1350),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1427),
.B(n_1451),
.Y(n_1473)
);

O2A1O1Ixp5_ASAP7_75t_L g1474 ( 
.A1(n_1333),
.A2(n_1422),
.B(n_1426),
.C(n_1398),
.Y(n_1474)
);

OA21x2_ASAP7_75t_L g1475 ( 
.A1(n_1401),
.A2(n_1437),
.B(n_1405),
.Y(n_1475)
);

OAI31xp33_ASAP7_75t_L g1476 ( 
.A1(n_1356),
.A2(n_1414),
.A3(n_1438),
.B(n_1400),
.Y(n_1476)
);

O2A1O1Ixp33_ASAP7_75t_L g1477 ( 
.A1(n_1333),
.A2(n_1422),
.B(n_1428),
.C(n_1390),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1368),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1340),
.Y(n_1479)
);

O2A1O1Ixp33_ASAP7_75t_L g1480 ( 
.A1(n_1390),
.A2(n_1367),
.B(n_1371),
.C(n_1350),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1363),
.B(n_1371),
.Y(n_1481)
);

BUFx6f_ASAP7_75t_L g1482 ( 
.A(n_1448),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1364),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1363),
.B(n_1402),
.Y(n_1484)
);

AOI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1410),
.A2(n_1430),
.B(n_1334),
.Y(n_1485)
);

O2A1O1Ixp5_ASAP7_75t_L g1486 ( 
.A1(n_1386),
.A2(n_1385),
.B(n_1394),
.C(n_1392),
.Y(n_1486)
);

NOR2xp67_ASAP7_75t_L g1487 ( 
.A(n_1345),
.B(n_1378),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1373),
.B(n_1372),
.Y(n_1489)
);

OAI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1400),
.A2(n_1435),
.B1(n_1334),
.B2(n_1335),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1417),
.B(n_1418),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1419),
.B(n_1424),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1435),
.A2(n_1335),
.B1(n_1447),
.B2(n_1433),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1359),
.B(n_1420),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1358),
.B(n_1362),
.Y(n_1495)
);

A2O1A1Ixp33_ASAP7_75t_L g1496 ( 
.A1(n_1349),
.A2(n_1389),
.B(n_1370),
.C(n_1385),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1393),
.B(n_1391),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1421),
.A2(n_1445),
.B(n_1389),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1358),
.B(n_1355),
.Y(n_1499)
);

A2O1A1Ixp33_ASAP7_75t_L g1500 ( 
.A1(n_1349),
.A2(n_1379),
.B(n_1328),
.C(n_1354),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1447),
.A2(n_1450),
.B1(n_1397),
.B2(n_1406),
.Y(n_1501)
);

INVxp67_ASAP7_75t_L g1502 ( 
.A(n_1448),
.Y(n_1502)
);

OA21x2_ASAP7_75t_L g1503 ( 
.A1(n_1386),
.A2(n_1399),
.B(n_1380),
.Y(n_1503)
);

AOI31xp33_ASAP7_75t_L g1504 ( 
.A1(n_1329),
.A2(n_1449),
.A3(n_1436),
.B(n_1421),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1395),
.B(n_1387),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1395),
.B(n_1450),
.Y(n_1506)
);

AOI21xp5_ASAP7_75t_SL g1507 ( 
.A1(n_1337),
.A2(n_1369),
.B(n_1346),
.Y(n_1507)
);

BUFx3_ASAP7_75t_L g1508 ( 
.A(n_1338),
.Y(n_1508)
);

O2A1O1Ixp33_ASAP7_75t_L g1509 ( 
.A1(n_1388),
.A2(n_1406),
.B(n_1353),
.C(n_1445),
.Y(n_1509)
);

A2O1A1Ixp33_ASAP7_75t_L g1510 ( 
.A1(n_1434),
.A2(n_1384),
.B(n_1357),
.C(n_1439),
.Y(n_1510)
);

O2A1O1Ixp5_ASAP7_75t_L g1511 ( 
.A1(n_1341),
.A2(n_1434),
.B(n_1442),
.C(n_1423),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1343),
.A2(n_1431),
.B1(n_1337),
.B2(n_1344),
.Y(n_1512)
);

OAI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1343),
.A2(n_1431),
.B1(n_1344),
.B2(n_1329),
.Y(n_1513)
);

O2A1O1Ixp33_ASAP7_75t_L g1514 ( 
.A1(n_1346),
.A2(n_1369),
.B(n_1331),
.C(n_1432),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_L g1515 ( 
.A(n_1374),
.Y(n_1515)
);

CKINVDCx20_ASAP7_75t_R g1516 ( 
.A(n_1374),
.Y(n_1516)
);

OAI211xp5_ASAP7_75t_L g1517 ( 
.A1(n_1441),
.A2(n_1404),
.B(n_1415),
.C(n_1429),
.Y(n_1517)
);

CKINVDCx20_ASAP7_75t_R g1518 ( 
.A(n_1441),
.Y(n_1518)
);

INVxp67_ASAP7_75t_L g1519 ( 
.A(n_1343),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1382),
.B(n_1409),
.Y(n_1520)
);

AOI21x1_ASAP7_75t_SL g1521 ( 
.A1(n_1431),
.A2(n_1434),
.B(n_1382),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1434),
.B(n_1409),
.Y(n_1522)
);

AOI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1382),
.A2(n_1200),
.B(n_1444),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1375),
.B(n_1376),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1342),
.A2(n_1407),
.B1(n_1193),
.B2(n_1403),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1375),
.B(n_1376),
.Y(n_1526)
);

CKINVDCx20_ASAP7_75t_R g1527 ( 
.A(n_1374),
.Y(n_1527)
);

BUFx3_ASAP7_75t_L g1528 ( 
.A(n_1413),
.Y(n_1528)
);

O2A1O1Ixp5_ASAP7_75t_L g1529 ( 
.A1(n_1408),
.A2(n_1452),
.B(n_1339),
.C(n_1416),
.Y(n_1529)
);

A2O1A1Ixp33_ASAP7_75t_L g1530 ( 
.A1(n_1339),
.A2(n_1266),
.B(n_1194),
.C(n_1193),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1381),
.B(n_1348),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1381),
.B(n_1348),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1381),
.B(n_1330),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1342),
.A2(n_1407),
.B1(n_1193),
.B2(n_1403),
.Y(n_1534)
);

OA21x2_ASAP7_75t_L g1535 ( 
.A1(n_1351),
.A2(n_1347),
.B(n_1444),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1381),
.B(n_1348),
.Y(n_1536)
);

INVxp67_ASAP7_75t_SL g1537 ( 
.A(n_1421),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1342),
.A2(n_1407),
.B1(n_1193),
.B2(n_1403),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1381),
.B(n_1348),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1340),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_1415),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1365),
.B(n_1366),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1365),
.B(n_1366),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1383),
.Y(n_1544)
);

AOI21xp5_ASAP7_75t_L g1545 ( 
.A1(n_1444),
.A2(n_1200),
.B(n_1199),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_1415),
.Y(n_1546)
);

AOI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1444),
.A2(n_1200),
.B(n_1199),
.Y(n_1547)
);

O2A1O1Ixp33_ASAP7_75t_L g1548 ( 
.A1(n_1403),
.A2(n_1266),
.B(n_1425),
.C(n_1416),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1340),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1444),
.A2(n_1200),
.B(n_1199),
.Y(n_1550)
);

A2O1A1Ixp33_ASAP7_75t_L g1551 ( 
.A1(n_1339),
.A2(n_1266),
.B(n_1194),
.C(n_1193),
.Y(n_1551)
);

OA21x2_ASAP7_75t_L g1552 ( 
.A1(n_1351),
.A2(n_1347),
.B(n_1444),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1342),
.A2(n_1407),
.B1(n_1193),
.B2(n_1403),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1511),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1479),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1456),
.B(n_1528),
.Y(n_1556)
);

AOI21xp5_ASAP7_75t_SL g1557 ( 
.A1(n_1530),
.A2(n_1551),
.B(n_1457),
.Y(n_1557)
);

BUFx6f_ASAP7_75t_L g1558 ( 
.A(n_1503),
.Y(n_1558)
);

INVxp67_ASAP7_75t_SL g1559 ( 
.A(n_1495),
.Y(n_1559)
);

BUFx3_ASAP7_75t_L g1560 ( 
.A(n_1533),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1529),
.A2(n_1462),
.B(n_1463),
.Y(n_1561)
);

OA21x2_ASAP7_75t_L g1562 ( 
.A1(n_1460),
.A2(n_1542),
.B(n_1465),
.Y(n_1562)
);

AO21x2_ASAP7_75t_L g1563 ( 
.A1(n_1460),
.A2(n_1542),
.B(n_1465),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1483),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1540),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1549),
.Y(n_1566)
);

AO21x2_ASAP7_75t_L g1567 ( 
.A1(n_1543),
.A2(n_1523),
.B(n_1550),
.Y(n_1567)
);

INVx2_ASAP7_75t_SL g1568 ( 
.A(n_1455),
.Y(n_1568)
);

AOI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1467),
.A2(n_1487),
.B(n_1512),
.Y(n_1569)
);

OR2x6_ASAP7_75t_L g1570 ( 
.A(n_1507),
.B(n_1461),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1470),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1469),
.B(n_1524),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1454),
.B(n_1531),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1526),
.Y(n_1574)
);

AO21x2_ASAP7_75t_L g1575 ( 
.A1(n_1545),
.A2(n_1547),
.B(n_1499),
.Y(n_1575)
);

INVx3_ASAP7_75t_L g1576 ( 
.A(n_1475),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1536),
.B(n_1539),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1478),
.Y(n_1578)
);

OA21x2_ASAP7_75t_L g1579 ( 
.A1(n_1474),
.A2(n_1498),
.B(n_1495),
.Y(n_1579)
);

OAI21x1_ASAP7_75t_L g1580 ( 
.A1(n_1514),
.A2(n_1521),
.B(n_1552),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1488),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1532),
.Y(n_1582)
);

AOI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1525),
.A2(n_1553),
.B1(n_1538),
.B2(n_1534),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1491),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_1541),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1520),
.B(n_1468),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1480),
.B(n_1472),
.Y(n_1587)
);

AOI21xp5_ASAP7_75t_SL g1588 ( 
.A1(n_1459),
.A2(n_1548),
.B(n_1553),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1468),
.B(n_1535),
.Y(n_1589)
);

OAI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1525),
.A2(n_1534),
.B(n_1538),
.Y(n_1590)
);

OA21x2_ASAP7_75t_L g1591 ( 
.A1(n_1486),
.A2(n_1485),
.B(n_1496),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1535),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1492),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1537),
.Y(n_1594)
);

AO21x2_ASAP7_75t_L g1595 ( 
.A1(n_1522),
.A2(n_1490),
.B(n_1510),
.Y(n_1595)
);

AO21x2_ASAP7_75t_L g1596 ( 
.A1(n_1490),
.A2(n_1500),
.B(n_1453),
.Y(n_1596)
);

AOI21x1_ASAP7_75t_L g1597 ( 
.A1(n_1512),
.A2(n_1513),
.B(n_1453),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1473),
.B(n_1484),
.Y(n_1598)
);

AO21x2_ASAP7_75t_L g1599 ( 
.A1(n_1493),
.A2(n_1466),
.B(n_1513),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1481),
.B(n_1466),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1519),
.B(n_1546),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1544),
.B(n_1489),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1590),
.A2(n_1583),
.B1(n_1476),
.B2(n_1596),
.Y(n_1603)
);

A2O1A1Ixp33_ASAP7_75t_L g1604 ( 
.A1(n_1590),
.A2(n_1476),
.B(n_1471),
.C(n_1477),
.Y(n_1604)
);

INVx1_ASAP7_75t_SL g1605 ( 
.A(n_1602),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1586),
.B(n_1493),
.Y(n_1606)
);

INVxp33_ASAP7_75t_L g1607 ( 
.A(n_1556),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1572),
.B(n_1504),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1583),
.A2(n_1501),
.B1(n_1515),
.B2(n_1505),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1564),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1564),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1559),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1572),
.B(n_1504),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1596),
.A2(n_1501),
.B1(n_1515),
.B2(n_1506),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1574),
.B(n_1509),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1562),
.B(n_1563),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1562),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1562),
.B(n_1517),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1562),
.B(n_1497),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1563),
.B(n_1458),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1576),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1557),
.A2(n_1518),
.B1(n_1516),
.B2(n_1527),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1576),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1567),
.B(n_1494),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1555),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_1585),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1555),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1619),
.B(n_1573),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1603),
.A2(n_1596),
.B1(n_1599),
.B2(n_1595),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1603),
.A2(n_1596),
.B1(n_1599),
.B2(n_1595),
.Y(n_1630)
);

OAI31xp33_ASAP7_75t_L g1631 ( 
.A1(n_1604),
.A2(n_1600),
.A3(n_1557),
.B(n_1588),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1624),
.B(n_1620),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1610),
.Y(n_1633)
);

INVxp67_ASAP7_75t_SL g1634 ( 
.A(n_1615),
.Y(n_1634)
);

NAND3xp33_ASAP7_75t_L g1635 ( 
.A(n_1604),
.B(n_1588),
.C(n_1561),
.Y(n_1635)
);

BUFx2_ASAP7_75t_L g1636 ( 
.A(n_1610),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_L g1637 ( 
.A(n_1607),
.B(n_1515),
.Y(n_1637)
);

OAI31xp33_ASAP7_75t_L g1638 ( 
.A1(n_1618),
.A2(n_1600),
.A3(n_1587),
.B(n_1571),
.Y(n_1638)
);

AOI211xp5_ASAP7_75t_SL g1639 ( 
.A1(n_1622),
.A2(n_1587),
.B(n_1578),
.C(n_1594),
.Y(n_1639)
);

NAND3xp33_ASAP7_75t_L g1640 ( 
.A(n_1616),
.B(n_1591),
.C(n_1579),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1625),
.Y(n_1641)
);

INVxp67_ASAP7_75t_SL g1642 ( 
.A(n_1615),
.Y(n_1642)
);

BUFx2_ASAP7_75t_L g1643 ( 
.A(n_1611),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_R g1644 ( 
.A(n_1626),
.B(n_1508),
.Y(n_1644)
);

AOI211xp5_ASAP7_75t_L g1645 ( 
.A1(n_1622),
.A2(n_1580),
.B(n_1554),
.C(n_1558),
.Y(n_1645)
);

OAI332xp33_ASAP7_75t_L g1646 ( 
.A1(n_1617),
.A2(n_1581),
.A3(n_1584),
.B1(n_1571),
.B2(n_1554),
.B3(n_1593),
.C1(n_1566),
.C2(n_1565),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1619),
.B(n_1573),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1606),
.A2(n_1599),
.B1(n_1595),
.B2(n_1614),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1605),
.B(n_1582),
.Y(n_1649)
);

OA21x2_ASAP7_75t_L g1650 ( 
.A1(n_1617),
.A2(n_1589),
.B(n_1592),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1606),
.A2(n_1599),
.B1(n_1595),
.B2(n_1614),
.Y(n_1651)
);

OAI221xp5_ASAP7_75t_L g1652 ( 
.A1(n_1618),
.A2(n_1597),
.B1(n_1591),
.B2(n_1569),
.C(n_1584),
.Y(n_1652)
);

INVx1_ASAP7_75t_SL g1653 ( 
.A(n_1626),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1619),
.B(n_1577),
.Y(n_1654)
);

NOR3xp33_ASAP7_75t_L g1655 ( 
.A(n_1618),
.B(n_1578),
.C(n_1568),
.Y(n_1655)
);

AOI22xp5_ASAP7_75t_L g1656 ( 
.A1(n_1609),
.A2(n_1591),
.B1(n_1575),
.B2(n_1567),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1612),
.B(n_1598),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1624),
.B(n_1560),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1624),
.B(n_1620),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1627),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1650),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1635),
.B(n_1607),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1650),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1650),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1641),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1650),
.Y(n_1666)
);

BUFx2_ASAP7_75t_L g1667 ( 
.A(n_1640),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1631),
.B(n_1638),
.Y(n_1668)
);

INVx4_ASAP7_75t_SL g1669 ( 
.A(n_1658),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1633),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1635),
.B(n_1634),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1641),
.Y(n_1672)
);

INVx3_ASAP7_75t_L g1673 ( 
.A(n_1632),
.Y(n_1673)
);

OAI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1631),
.A2(n_1591),
.B(n_1616),
.Y(n_1674)
);

INVx2_ASAP7_75t_SL g1675 ( 
.A(n_1658),
.Y(n_1675)
);

BUFx2_ASAP7_75t_L g1676 ( 
.A(n_1636),
.Y(n_1676)
);

INVx3_ASAP7_75t_SL g1677 ( 
.A(n_1659),
.Y(n_1677)
);

OA21x2_ASAP7_75t_L g1678 ( 
.A1(n_1629),
.A2(n_1617),
.B(n_1621),
.Y(n_1678)
);

BUFx3_ASAP7_75t_L g1679 ( 
.A(n_1656),
.Y(n_1679)
);

BUFx6f_ASAP7_75t_L g1680 ( 
.A(n_1659),
.Y(n_1680)
);

BUFx2_ASAP7_75t_L g1681 ( 
.A(n_1636),
.Y(n_1681)
);

BUFx2_ASAP7_75t_L g1682 ( 
.A(n_1643),
.Y(n_1682)
);

OA21x2_ASAP7_75t_L g1683 ( 
.A1(n_1630),
.A2(n_1621),
.B(n_1623),
.Y(n_1683)
);

OR2x6_ASAP7_75t_L g1684 ( 
.A(n_1679),
.B(n_1570),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1667),
.B(n_1642),
.Y(n_1685)
);

AND2x4_ASAP7_75t_L g1686 ( 
.A(n_1669),
.B(n_1659),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1667),
.B(n_1659),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1667),
.B(n_1646),
.Y(n_1688)
);

NAND3xp33_ASAP7_75t_L g1689 ( 
.A(n_1671),
.B(n_1645),
.C(n_1639),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1661),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1661),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1671),
.B(n_1668),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1662),
.B(n_1653),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1679),
.A2(n_1668),
.B1(n_1648),
.B2(n_1651),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1677),
.B(n_1628),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1677),
.B(n_1647),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1665),
.Y(n_1697)
);

NOR2xp67_ASAP7_75t_L g1698 ( 
.A(n_1674),
.B(n_1652),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1679),
.B(n_1657),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1665),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1669),
.B(n_1658),
.Y(n_1701)
);

CKINVDCx16_ASAP7_75t_R g1702 ( 
.A(n_1662),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1661),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1661),
.Y(n_1704)
);

BUFx2_ASAP7_75t_L g1705 ( 
.A(n_1676),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1669),
.B(n_1654),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1661),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1679),
.B(n_1657),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1669),
.B(n_1645),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1679),
.B(n_1637),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1670),
.B(n_1660),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1666),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1670),
.B(n_1660),
.Y(n_1713)
);

OAI21xp33_ASAP7_75t_L g1714 ( 
.A1(n_1674),
.A2(n_1656),
.B(n_1655),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1674),
.B(n_1649),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1676),
.B(n_1643),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1669),
.B(n_1624),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1665),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1672),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1676),
.B(n_1612),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1683),
.A2(n_1613),
.B1(n_1608),
.B2(n_1567),
.Y(n_1721)
);

HB1xp67_ASAP7_75t_L g1722 ( 
.A(n_1681),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1666),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1697),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1692),
.B(n_1681),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1697),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1705),
.Y(n_1727)
);

INVx2_ASAP7_75t_SL g1728 ( 
.A(n_1686),
.Y(n_1728)
);

INVx2_ASAP7_75t_SL g1729 ( 
.A(n_1686),
.Y(n_1729)
);

NOR4xp25_ASAP7_75t_L g1730 ( 
.A(n_1692),
.B(n_1666),
.C(n_1664),
.D(n_1663),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1702),
.B(n_1681),
.Y(n_1731)
);

INVxp67_ASAP7_75t_SL g1732 ( 
.A(n_1693),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1700),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1686),
.B(n_1669),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1700),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1718),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1718),
.Y(n_1737)
);

INVx1_ASAP7_75t_SL g1738 ( 
.A(n_1702),
.Y(n_1738)
);

INVx3_ASAP7_75t_L g1739 ( 
.A(n_1686),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1686),
.B(n_1669),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1719),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1689),
.A2(n_1673),
.B1(n_1675),
.B2(n_1680),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1719),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1722),
.Y(n_1744)
);

INVxp67_ASAP7_75t_L g1745 ( 
.A(n_1710),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1687),
.B(n_1669),
.Y(n_1746)
);

NOR2x2_ASAP7_75t_L g1747 ( 
.A(n_1684),
.B(n_1644),
.Y(n_1747)
);

INVxp67_ASAP7_75t_L g1748 ( 
.A(n_1705),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1711),
.Y(n_1749)
);

OR2x6_ASAP7_75t_L g1750 ( 
.A(n_1689),
.B(n_1482),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1690),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1711),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1687),
.B(n_1673),
.Y(n_1753)
);

OR2x6_ASAP7_75t_L g1754 ( 
.A(n_1698),
.B(n_1502),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1699),
.B(n_1649),
.Y(n_1755)
);

OR2x6_ASAP7_75t_L g1756 ( 
.A(n_1698),
.B(n_1464),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1687),
.B(n_1673),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1688),
.B(n_1682),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1699),
.B(n_1708),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1713),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1738),
.B(n_1688),
.Y(n_1761)
);

BUFx2_ASAP7_75t_L g1762 ( 
.A(n_1750),
.Y(n_1762)
);

NAND2x1p5_ASAP7_75t_L g1763 ( 
.A(n_1739),
.B(n_1709),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1732),
.B(n_1714),
.Y(n_1764)
);

OA21x2_ASAP7_75t_L g1765 ( 
.A1(n_1758),
.A2(n_1694),
.B(n_1714),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1745),
.B(n_1685),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1746),
.B(n_1701),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1746),
.B(n_1701),
.Y(n_1768)
);

INVx1_ASAP7_75t_SL g1769 ( 
.A(n_1747),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1753),
.Y(n_1770)
);

NOR2x1_ASAP7_75t_L g1771 ( 
.A(n_1750),
.B(n_1685),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1727),
.Y(n_1772)
);

INVxp67_ASAP7_75t_L g1773 ( 
.A(n_1731),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1727),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1739),
.B(n_1701),
.Y(n_1775)
);

INVxp67_ASAP7_75t_L g1776 ( 
.A(n_1725),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_SL g1777 ( 
.A1(n_1750),
.A2(n_1709),
.B1(n_1715),
.B2(n_1683),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1739),
.B(n_1701),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1744),
.B(n_1708),
.Y(n_1779)
);

INVxp67_ASAP7_75t_L g1780 ( 
.A(n_1759),
.Y(n_1780)
);

AOI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1750),
.A2(n_1721),
.B1(n_1683),
.B2(n_1678),
.Y(n_1781)
);

OR2x6_ASAP7_75t_L g1782 ( 
.A(n_1756),
.B(n_1684),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1748),
.B(n_1682),
.Y(n_1783)
);

HB1xp67_ASAP7_75t_L g1784 ( 
.A(n_1755),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1724),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1728),
.B(n_1729),
.Y(n_1786)
);

AOI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1754),
.A2(n_1683),
.B1(n_1678),
.B2(n_1684),
.Y(n_1787)
);

NAND2x1p5_ASAP7_75t_L g1788 ( 
.A(n_1771),
.B(n_1728),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1765),
.B(n_1730),
.Y(n_1789)
);

OAI221xp5_ASAP7_75t_L g1790 ( 
.A1(n_1777),
.A2(n_1754),
.B1(n_1756),
.B2(n_1715),
.C(n_1683),
.Y(n_1790)
);

A2O1A1Ixp33_ASAP7_75t_L g1791 ( 
.A1(n_1781),
.A2(n_1666),
.B(n_1664),
.C(n_1663),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1765),
.A2(n_1764),
.B1(n_1787),
.B2(n_1761),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1774),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1763),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1774),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1772),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1784),
.B(n_1749),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_SL g1798 ( 
.A1(n_1765),
.A2(n_1754),
.B1(n_1742),
.B2(n_1756),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_L g1799 ( 
.A(n_1769),
.B(n_1729),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1776),
.B(n_1752),
.Y(n_1800)
);

INVxp67_ASAP7_75t_L g1801 ( 
.A(n_1762),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1779),
.B(n_1760),
.Y(n_1802)
);

OAI21xp5_ASAP7_75t_SL g1803 ( 
.A1(n_1763),
.A2(n_1740),
.B(n_1734),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1780),
.B(n_1726),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1785),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1767),
.B(n_1734),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1766),
.Y(n_1807)
);

AOI321xp33_ASAP7_75t_L g1808 ( 
.A1(n_1770),
.A2(n_1751),
.A3(n_1690),
.B1(n_1691),
.B2(n_1703),
.C(n_1704),
.Y(n_1808)
);

INVx3_ASAP7_75t_L g1809 ( 
.A(n_1763),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1788),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1801),
.Y(n_1811)
);

NOR2xp33_ASAP7_75t_L g1812 ( 
.A(n_1789),
.B(n_1773),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1806),
.B(n_1767),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1799),
.B(n_1768),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1789),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1797),
.B(n_1762),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1807),
.B(n_1768),
.Y(n_1817)
);

INVxp67_ASAP7_75t_L g1818 ( 
.A(n_1809),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1809),
.B(n_1786),
.Y(n_1819)
);

NOR2xp33_ASAP7_75t_L g1820 ( 
.A(n_1793),
.B(n_1786),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1817),
.B(n_1820),
.Y(n_1821)
);

NAND3xp33_ASAP7_75t_L g1822 ( 
.A(n_1812),
.B(n_1792),
.C(n_1808),
.Y(n_1822)
);

AOI221xp5_ASAP7_75t_L g1823 ( 
.A1(n_1812),
.A2(n_1790),
.B1(n_1791),
.B2(n_1798),
.C(n_1800),
.Y(n_1823)
);

NAND4xp25_ASAP7_75t_L g1824 ( 
.A(n_1816),
.B(n_1804),
.C(n_1796),
.D(n_1794),
.Y(n_1824)
);

AOI22xp5_ASAP7_75t_L g1825 ( 
.A1(n_1815),
.A2(n_1782),
.B1(n_1803),
.B2(n_1788),
.Y(n_1825)
);

NAND3xp33_ASAP7_75t_SL g1826 ( 
.A(n_1816),
.B(n_1804),
.C(n_1802),
.Y(n_1826)
);

NAND4xp25_ASAP7_75t_L g1827 ( 
.A(n_1820),
.B(n_1795),
.C(n_1805),
.D(n_1783),
.Y(n_1827)
);

AOI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1814),
.A2(n_1782),
.B1(n_1770),
.B2(n_1751),
.Y(n_1828)
);

HAxp5_ASAP7_75t_SL g1829 ( 
.A(n_1811),
.B(n_1747),
.CON(n_1829),
.SN(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1813),
.B(n_1753),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1826),
.B(n_1830),
.Y(n_1831)
);

AOI221xp5_ASAP7_75t_L g1832 ( 
.A1(n_1822),
.A2(n_1823),
.B1(n_1824),
.B2(n_1827),
.C(n_1810),
.Y(n_1832)
);

OAI222xp33_ASAP7_75t_L g1833 ( 
.A1(n_1825),
.A2(n_1828),
.B1(n_1810),
.B2(n_1782),
.C1(n_1821),
.C2(n_1818),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1829),
.Y(n_1834)
);

INVxp67_ASAP7_75t_L g1835 ( 
.A(n_1821),
.Y(n_1835)
);

AOI211xp5_ASAP7_75t_SL g1836 ( 
.A1(n_1826),
.A2(n_1819),
.B(n_1778),
.C(n_1775),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1834),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1835),
.Y(n_1838)
);

NOR2x1_ASAP7_75t_L g1839 ( 
.A(n_1831),
.B(n_1775),
.Y(n_1839)
);

INVxp67_ASAP7_75t_L g1840 ( 
.A(n_1836),
.Y(n_1840)
);

OAI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1832),
.A2(n_1735),
.B(n_1733),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1833),
.B(n_1778),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1839),
.B(n_1757),
.Y(n_1843)
);

NOR2x1_ASAP7_75t_SL g1844 ( 
.A(n_1842),
.B(n_1782),
.Y(n_1844)
);

INVxp33_ASAP7_75t_SL g1845 ( 
.A(n_1837),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1838),
.Y(n_1846)
);

AOI322xp5_ASAP7_75t_L g1847 ( 
.A1(n_1840),
.A2(n_1691),
.A3(n_1707),
.B1(n_1704),
.B2(n_1703),
.C1(n_1690),
.C2(n_1712),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1844),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1843),
.Y(n_1849)
);

AOI22xp5_ASAP7_75t_SL g1850 ( 
.A1(n_1845),
.A2(n_1841),
.B1(n_1740),
.B2(n_1757),
.Y(n_1850)
);

NOR3xp33_ASAP7_75t_L g1851 ( 
.A(n_1848),
.B(n_1846),
.C(n_1841),
.Y(n_1851)
);

AOI322xp5_ASAP7_75t_L g1852 ( 
.A1(n_1851),
.A2(n_1849),
.A3(n_1850),
.B1(n_1847),
.B2(n_1691),
.C1(n_1707),
.C2(n_1712),
.Y(n_1852)
);

NAND3xp33_ASAP7_75t_L g1853 ( 
.A(n_1852),
.B(n_1704),
.C(n_1703),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1852),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1854),
.Y(n_1855)
);

XOR2x1_ASAP7_75t_L g1856 ( 
.A(n_1853),
.B(n_1701),
.Y(n_1856)
);

OA22x2_ASAP7_75t_L g1857 ( 
.A1(n_1855),
.A2(n_1743),
.B1(n_1741),
.B2(n_1737),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1856),
.A2(n_1736),
.B1(n_1723),
.B2(n_1707),
.Y(n_1858)
);

OR3x1_ASAP7_75t_L g1859 ( 
.A(n_1857),
.B(n_1601),
.C(n_1672),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1859),
.A2(n_1858),
.B1(n_1723),
.B2(n_1712),
.Y(n_1860)
);

OA21x2_ASAP7_75t_L g1861 ( 
.A1(n_1860),
.A2(n_1716),
.B(n_1720),
.Y(n_1861)
);

AOI22x1_ASAP7_75t_L g1862 ( 
.A1(n_1861),
.A2(n_1682),
.B1(n_1723),
.B2(n_1706),
.Y(n_1862)
);

AO22x2_ASAP7_75t_L g1863 ( 
.A1(n_1862),
.A2(n_1716),
.B1(n_1720),
.B2(n_1713),
.Y(n_1863)
);

AOI211xp5_ASAP7_75t_L g1864 ( 
.A1(n_1863),
.A2(n_1717),
.B(n_1695),
.C(n_1696),
.Y(n_1864)
);


endmodule