module real_jpeg_32410_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_131;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_0),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_1),
.B(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_1),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_1),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_2),
.B(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_2),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_3),
.B(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_3),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_3),
.B(n_82),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_3),
.Y(n_123)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_4),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_5),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_8),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_8),
.B(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_9),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_10),
.B(n_44),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_28),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_11),
.B(n_86),
.Y(n_85)
);

AND2x4_ASAP7_75t_SL g118 ( 
.A(n_11),
.B(n_119),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_104),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_69),
.B(n_103),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_36),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_16),
.B(n_36),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_27),
.C(n_31),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_17),
.A2(n_18),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.Y(n_18)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_22),
.B(n_26),
.Y(n_47)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_27),
.B(n_31),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_30),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_35),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_50),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_38),
.B(n_49),
.C(n_50),
.Y(n_106)
);

AO22x1_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_38)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_43),
.B(n_45),
.Y(n_127)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_56),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_51),
.B(n_63),
.C(n_68),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_63),
.B1(n_64),
.B2(n_68),
.Y(n_56)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OA21x2_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_96),
.B(n_102),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_90),
.B(n_95),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_80),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_84),
.B1(n_85),
.B2(n_89),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_84),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_99),
.Y(n_102)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_141),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

NOR2xp67_ASAP7_75t_SL g142 ( 
.A(n_106),
.B(n_107),
.Y(n_142)
);

XNOR2x1_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_126),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_121),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_117),
.B2(n_118),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_SL g121 ( 
.A(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2x2_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_137),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_129)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);


endmodule