module fake_jpeg_17063_n_132 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_8),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_0),
.B(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_24),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_0),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_17),
.A2(n_1),
.B(n_2),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_18),
.B1(n_13),
.B2(n_24),
.Y(n_30)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_9),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_19),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_37),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_18),
.B1(n_21),
.B2(n_11),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_33),
.A2(n_18),
.B1(n_12),
.B2(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_29),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_44),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_26),
.C(n_25),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_42),
.B(n_17),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_50),
.Y(n_62)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_45),
.B(n_37),
.Y(n_60)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_48),
.Y(n_70)
);

AND2x4_ASAP7_75t_SL g47 ( 
.A(n_32),
.B(n_22),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_12),
.B(n_17),
.Y(n_69)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_55),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_54),
.A2(n_14),
.B1(n_21),
.B2(n_16),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_11),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_59),
.A2(n_20),
.B1(n_23),
.B2(n_3),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_60),
.B(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_32),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_31),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_67),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_17),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_71),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_14),
.B(n_10),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_28),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_23),
.Y(n_90)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_16),
.Y(n_73)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_66),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_76),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_42),
.B(n_41),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_81),
.B(n_86),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_80),
.B(n_61),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_SL g81 ( 
.A1(n_69),
.A2(n_47),
.B(n_54),
.C(n_28),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_68),
.A2(n_27),
.B1(n_46),
.B2(n_49),
.Y(n_84)
);

AOI221xp5_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_89),
.B1(n_59),
.B2(n_73),
.C(n_62),
.Y(n_91)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_87),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_90),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_91),
.A2(n_87),
.B1(n_76),
.B2(n_63),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_67),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_79),
.B(n_60),
.Y(n_95)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_62),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_97),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_65),
.C(n_70),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_25),
.C(n_63),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_102),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_83),
.B1(n_90),
.B2(n_81),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_104),
.A2(n_108),
.B(n_105),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_81),
.B(n_86),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_107),
.A2(n_101),
.B(n_100),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_81),
.B1(n_84),
.B2(n_88),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_93),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_98),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_99),
.Y(n_114)
);

BUFx24_ASAP7_75t_SL g112 ( 
.A(n_106),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_115),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_108),
.B(n_104),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_114),
.A2(n_116),
.B(n_117),
.Y(n_119)
);

OA21x2_ASAP7_75t_SL g117 ( 
.A1(n_103),
.A2(n_96),
.B(n_77),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_109),
.C(n_103),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_123),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_120),
.A2(n_122),
.B(n_121),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_116),
.A2(n_109),
.B(n_56),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_40),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_119),
.A2(n_1),
.B(n_2),
.Y(n_124)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_125),
.B(n_5),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_127),
.A2(n_7),
.B(n_8),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_SL g129 ( 
.A1(n_128),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_130),
.B1(n_7),
.B2(n_8),
.Y(n_131)
);

BUFx24_ASAP7_75t_SL g132 ( 
.A(n_131),
.Y(n_132)
);


endmodule