module real_jpeg_21930_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_35;
wire n_38;
wire n_33;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_40;
wire n_39;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx14_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_0),
.B(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_1),
.B(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_2),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g8 ( 
.A(n_3),
.B(n_9),
.Y(n_8)
);

OR2x2_ASAP7_75t_SL g23 ( 
.A(n_3),
.B(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

AO21x1_ASAP7_75t_SL g25 ( 
.A1(n_5),
.A2(n_14),
.B(n_17),
.Y(n_25)
);

OAI211xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_10),
.B(n_19),
.C(n_35),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_8),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_8),
.B(n_18),
.Y(n_27)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_9),
.B(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_11),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_18),
.Y(n_11)
);

AOI221xp5_ASAP7_75t_L g35 ( 
.A1(n_12),
.A2(n_15),
.B1(n_36),
.B2(n_38),
.C(n_40),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_SL g12 ( 
.A1(n_13),
.A2(n_14),
.B(n_17),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_13),
.B(n_18),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_16),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_16),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_22),
.Y(n_39)
);

AOI221xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.C(n_28),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);


endmodule