module fake_jpeg_19497_n_346 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_346);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_346;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_23),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_59),
.B(n_28),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_26),
.B1(n_24),
.B2(n_27),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_62),
.B1(n_48),
.B2(n_44),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_26),
.B1(n_24),
.B2(n_27),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_43),
.B1(n_39),
.B2(n_42),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_63),
.A2(n_44),
.B1(n_47),
.B2(n_46),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_25),
.Y(n_65)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_75),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_59),
.B(n_23),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_96),
.Y(n_124)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_48),
.B1(n_45),
.B2(n_39),
.Y(n_73)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_73),
.A2(n_74),
.B1(n_53),
.B2(n_52),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_33),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

BUFx2_ASAP7_75t_SL g77 ( 
.A(n_51),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_38),
.B1(n_43),
.B2(n_39),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_82),
.A2(n_88),
.B1(n_94),
.B2(n_97),
.Y(n_118)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

BUFx10_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

AO22x1_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_48),
.B1(n_49),
.B2(n_47),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_67),
.B(n_66),
.C(n_58),
.Y(n_107)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_66),
.B1(n_64),
.B2(n_61),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_90),
.Y(n_126)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

AND2x4_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_48),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_53),
.B(n_58),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_64),
.A2(n_45),
.B1(n_44),
.B2(n_46),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_34),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_25),
.Y(n_113)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_53),
.A2(n_44),
.B1(n_19),
.B2(n_28),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_100),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_67),
.B1(n_58),
.B2(n_60),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_104),
.A2(n_115),
.B(n_125),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_107),
.Y(n_159)
);

INVx2_ASAP7_75t_R g110 ( 
.A(n_93),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_110),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_114),
.Y(n_143)
);

AOI32xp33_ASAP7_75t_L g114 ( 
.A1(n_78),
.A2(n_93),
.A3(n_89),
.B1(n_74),
.B2(n_79),
.Y(n_114)
);

BUFx24_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_121),
.A2(n_127),
.B1(n_21),
.B2(n_17),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_78),
.A2(n_86),
.B(n_62),
.C(n_97),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_34),
.B1(n_33),
.B2(n_19),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_82),
.B(n_30),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_18),
.C(n_21),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_83),
.B(n_30),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_87),
.B(n_19),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_133),
.B(n_99),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_134),
.A2(n_102),
.B1(n_109),
.B2(n_112),
.Y(n_162)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_119),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_145),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_138),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_129),
.B(n_110),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_81),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_148),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_94),
.B1(n_100),
.B2(n_69),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_142),
.A2(n_158),
.B1(n_47),
.B2(n_46),
.Y(n_186)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_125),
.A2(n_73),
.B(n_17),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_146),
.A2(n_18),
.B(n_22),
.Y(n_187)
);

MAJx2_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_73),
.C(n_92),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_147),
.A2(n_157),
.B(n_122),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_80),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_124),
.B(n_69),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_122),
.Y(n_176)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_138),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_122),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_161),
.Y(n_182)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_109),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

MAJx2_ASAP7_75t_L g157 ( 
.A(n_104),
.B(n_118),
.C(n_126),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_104),
.A2(n_85),
.B1(n_49),
.B2(n_47),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_130),
.A2(n_35),
.B1(n_31),
.B2(n_18),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_160),
.A2(n_132),
.B1(n_31),
.B2(n_35),
.Y(n_178)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_103),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_162),
.A2(n_163),
.B1(n_168),
.B2(n_188),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_159),
.A2(n_106),
.B1(n_112),
.B2(n_105),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_167),
.B(n_179),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_146),
.A2(n_111),
.B1(n_108),
.B2(n_105),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_111),
.C(n_123),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_171),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_123),
.C(n_108),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_173),
.A2(n_183),
.B(n_187),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_132),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_176),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_178),
.A2(n_186),
.B1(n_154),
.B2(n_153),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_49),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_184),
.Y(n_212)
);

AOI22x1_ASAP7_75t_SL g183 ( 
.A1(n_141),
.A2(n_31),
.B1(n_35),
.B2(n_18),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_139),
.B(n_49),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_145),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_157),
.A2(n_46),
.B1(n_41),
.B2(n_40),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_190),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_135),
.B(n_41),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_155),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_156),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_157),
.A2(n_41),
.B1(n_40),
.B2(n_37),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_192),
.A2(n_40),
.B1(n_37),
.B2(n_32),
.Y(n_224)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_193),
.Y(n_244)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_194),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_165),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_196),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_140),
.B(n_154),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_197),
.A2(n_202),
.B1(n_221),
.B2(n_163),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_165),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_203),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_174),
.A2(n_134),
.B1(n_147),
.B2(n_152),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_182),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_174),
.A2(n_147),
.B(n_136),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_206),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_192),
.A2(n_144),
.B1(n_150),
.B2(n_161),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_205),
.A2(n_224),
.B1(n_181),
.B2(n_184),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_180),
.Y(n_206)
);

NOR2x1p5_ASAP7_75t_SL g208 ( 
.A(n_188),
.B(n_151),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_208),
.Y(n_227)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_209),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_169),
.Y(n_235)
);

OAI21xp33_ASAP7_75t_L g211 ( 
.A1(n_183),
.A2(n_11),
.B(n_16),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_SL g246 ( 
.A1(n_211),
.A2(n_9),
.B(n_16),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_172),
.B(n_156),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_217),
.Y(n_242)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_216),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_175),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_218),
.Y(n_243)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_176),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_219),
.A2(n_220),
.B1(n_222),
.B2(n_223),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_186),
.A2(n_41),
.B1(n_40),
.B2(n_37),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_166),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_166),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_185),
.C(n_171),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_208),
.C(n_196),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_228),
.A2(n_229),
.B1(n_233),
.B2(n_250),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_200),
.A2(n_172),
.B1(n_170),
.B2(n_187),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_230),
.A2(n_234),
.B1(n_238),
.B2(n_224),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_200),
.A2(n_162),
.B1(n_191),
.B2(n_164),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_202),
.A2(n_164),
.B1(n_169),
.B2(n_180),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_235),
.B(n_239),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_213),
.A2(n_180),
.B1(n_22),
.B2(n_32),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_237),
.A2(n_246),
.B1(n_249),
.B2(n_206),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_197),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_22),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_201),
.B(n_214),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_247),
.B(n_248),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_22),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_213),
.A2(n_32),
.B1(n_9),
.B2(n_10),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_215),
.A2(n_32),
.B1(n_1),
.B2(n_2),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_252),
.B(n_264),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_240),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_253),
.B(n_255),
.Y(n_284)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_242),
.Y(n_254)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_244),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_209),
.Y(n_256)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_256),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_193),
.Y(n_257)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_257),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_236),
.B(n_194),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_258),
.B(n_267),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_199),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_259),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_219),
.C(n_218),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_248),
.C(n_234),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_204),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_261),
.B(n_228),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_212),
.Y(n_262)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_262),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_263),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_226),
.A2(n_207),
.B(n_244),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_265),
.A2(n_266),
.B1(n_238),
.B2(n_230),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_232),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_231),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_250),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_270),
.A2(n_271),
.B1(n_254),
.B2(n_266),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_243),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_261),
.B(n_247),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_273),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_269),
.B(n_235),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_275),
.C(n_290),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_229),
.C(n_233),
.Y(n_275)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_280),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_269),
.B(n_227),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_289),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_287),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_252),
.B(n_268),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_207),
.C(n_223),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_267),
.C(n_251),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_293),
.B(n_295),
.C(n_299),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_284),
.Y(n_294)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_294),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_251),
.C(n_262),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_276),
.A2(n_264),
.B(n_259),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_297),
.A2(n_10),
.B1(n_13),
.B2(n_16),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_263),
.C(n_259),
.Y(n_299)
);

OAI21x1_ASAP7_75t_L g300 ( 
.A1(n_277),
.A2(n_227),
.B(n_232),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_285),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_212),
.C(n_205),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_0),
.C(n_3),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_278),
.A2(n_206),
.B1(n_221),
.B2(n_11),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_303),
.A2(n_306),
.B1(n_302),
.B2(n_279),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_272),
.B(n_8),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_281),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_288),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_305),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_283),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_290),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_310),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_308),
.B(n_316),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_312),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_273),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_313),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_299),
.A2(n_279),
.B1(n_289),
.B2(n_4),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_291),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_318),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_314),
.B(n_295),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_320),
.B(n_316),
.Y(n_330)
);

FAx1_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_298),
.CI(n_296),
.CON(n_322),
.SN(n_322)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_324),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_301),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_315),
.A2(n_312),
.B(n_293),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_304),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_315),
.C(n_326),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g337 ( 
.A(n_328),
.B(n_332),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_326),
.B(n_298),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_333),
.C(n_323),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_330),
.B(n_334),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_296),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_325),
.B(n_305),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_335),
.A2(n_336),
.B1(n_329),
.B2(n_333),
.Y(n_339)
);

INVxp33_ASAP7_75t_L g336 ( 
.A(n_331),
.Y(n_336)
);

A2O1A1Ixp33_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_337),
.B(n_322),
.C(n_338),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_319),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_322),
.B1(n_10),
.B2(n_13),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_3),
.B(n_5),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_343),
.B(n_6),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_7),
.Y(n_345)
);

MAJx2_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_7),
.C(n_343),
.Y(n_346)
);


endmodule