module fake_jpeg_12563_n_69 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_69);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_69;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_43;
wire n_50;
wire n_29;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

BUFx16f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx2_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx10_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_0),
.B(n_4),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_24),
.Y(n_32)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_13),
.B(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_11),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_20),
.A2(n_10),
.B1(n_11),
.B2(n_14),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_23),
.B(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_12),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_35),
.B(n_15),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_38),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_L g38 ( 
.A1(n_26),
.A2(n_13),
.B(n_15),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_41),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_46),
.B(n_47),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_5),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_43),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_28),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_37),
.B(n_36),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_36),
.B1(n_30),
.B2(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_29),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_49),
.B(n_39),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_56),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_25),
.C(n_9),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_52),
.C(n_51),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_59),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_55),
.A2(n_52),
.B1(n_53),
.B2(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_60),
.B(n_6),
.Y(n_62)
);

OA21x2_ASAP7_75t_SL g64 ( 
.A1(n_62),
.A2(n_7),
.B(n_9),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_60),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_64),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_63),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_9),
.B(n_16),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_19),
.Y(n_69)
);


endmodule