module real_aes_8932_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_478;
wire n_356;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_552;
wire n_402;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g246 ( .A(n_0), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g84 ( .A1(n_1), .A2(n_34), .B1(n_85), .B2(n_102), .Y(n_84) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_2), .A2(n_58), .B1(n_195), .B2(n_196), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_2), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g301 ( .A1(n_2), .A2(n_32), .B1(n_236), .B2(n_283), .Y(n_301) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_3), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_4), .B(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g209 ( .A(n_5), .Y(n_209) );
AND2x6_ASAP7_75t_L g251 ( .A(n_5), .B(n_207), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_5), .B(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_6), .B(n_255), .Y(n_263) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_7), .A2(n_186), .B1(n_187), .B2(n_193), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_7), .Y(n_186) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_8), .A2(n_28), .B1(n_91), .B2(n_96), .Y(n_99) );
INVx1_ASAP7_75t_L g227 ( .A(n_9), .Y(n_227) );
INVx1_ASAP7_75t_L g230 ( .A(n_10), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_11), .B(n_232), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_12), .B(n_223), .Y(n_329) );
AO32x2_ASAP7_75t_L g299 ( .A1(n_13), .A2(n_222), .A3(n_255), .B1(n_274), .B2(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g296 ( .A(n_14), .B(n_236), .Y(n_296) );
AO22x2_ASAP7_75t_L g101 ( .A1(n_15), .A2(n_30), .B1(n_91), .B2(n_92), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_16), .B(n_223), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_17), .A2(n_42), .B1(n_236), .B2(n_283), .Y(n_302) );
AOI22xp33_ASAP7_75t_SL g285 ( .A1(n_18), .A2(n_64), .B1(n_232), .B2(n_236), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_19), .B(n_236), .Y(n_315) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_20), .Y(n_147) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_21), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_22), .B(n_276), .Y(n_275) );
CKINVDCx20_ASAP7_75t_R g143 ( .A(n_23), .Y(n_143) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_24), .A2(n_33), .B1(n_189), .B2(n_190), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_24), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_25), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_26), .B(n_276), .Y(n_317) );
INVx2_ASAP7_75t_L g234 ( .A(n_27), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_29), .A2(n_188), .B1(n_191), .B2(n_192), .Y(n_187) );
INVx1_ASAP7_75t_L g191 ( .A(n_29), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_29), .B(n_236), .Y(n_267) );
OAI221xp5_ASAP7_75t_L g200 ( .A1(n_30), .A2(n_46), .B1(n_56), .B2(n_201), .C(n_202), .Y(n_200) );
INVxp67_ASAP7_75t_L g203 ( .A(n_30), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_31), .B(n_276), .Y(n_298) );
INVx1_ASAP7_75t_L g190 ( .A(n_33), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_35), .B(n_236), .Y(n_258) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_36), .Y(n_178) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_37), .A2(n_72), .B1(n_283), .B2(n_284), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_38), .B(n_236), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_39), .B(n_236), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_40), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_41), .B(n_244), .Y(n_262) );
AOI22xp33_ASAP7_75t_SL g327 ( .A1(n_43), .A2(n_47), .B1(n_232), .B2(n_236), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_44), .B(n_236), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_45), .B(n_236), .Y(n_291) );
AO22x2_ASAP7_75t_L g90 ( .A1(n_46), .A2(n_68), .B1(n_91), .B2(n_92), .Y(n_90) );
INVxp67_ASAP7_75t_L g204 ( .A(n_46), .Y(n_204) );
INVx1_ASAP7_75t_L g207 ( .A(n_48), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_49), .A2(n_81), .B1(n_183), .B2(n_548), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_49), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_50), .B(n_236), .Y(n_247) );
INVx1_ASAP7_75t_L g226 ( .A(n_51), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_52), .Y(n_201) );
AO32x2_ASAP7_75t_L g280 ( .A1(n_53), .A2(n_255), .A3(n_274), .B1(n_281), .B2(n_286), .Y(n_280) );
INVx1_ASAP7_75t_L g270 ( .A(n_54), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g107 ( .A1(n_55), .A2(n_65), .B1(n_108), .B2(n_115), .Y(n_107) );
AO22x2_ASAP7_75t_L g95 ( .A1(n_56), .A2(n_74), .B1(n_91), .B2(n_96), .Y(n_95) );
INVx1_ASAP7_75t_L g312 ( .A(n_57), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_57), .A2(n_81), .B1(n_183), .B2(n_312), .Y(n_538) );
CKINVDCx14_ASAP7_75t_R g196 ( .A(n_58), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_59), .B(n_232), .Y(n_313) );
INVx1_ASAP7_75t_L g546 ( .A(n_59), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_60), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_61), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_62), .Y(n_131) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_63), .A2(n_81), .B1(n_182), .B2(n_183), .Y(n_80) );
CKINVDCx16_ASAP7_75t_R g182 ( .A(n_63), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_66), .B(n_283), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g316 ( .A(n_67), .B(n_232), .Y(n_316) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_69), .Y(n_160) );
INVx2_ASAP7_75t_L g224 ( .A(n_70), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_71), .B(n_232), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_73), .A2(n_77), .B1(n_232), .B2(n_233), .Y(n_326) );
INVx1_ASAP7_75t_L g91 ( .A(n_75), .Y(n_91) );
INVx1_ASAP7_75t_L g93 ( .A(n_75), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_76), .B(n_232), .Y(n_268) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_197), .B1(n_210), .B2(n_531), .C(n_537), .Y(n_78) );
XNOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_184), .Y(n_79) );
INVx1_ASAP7_75t_L g183 ( .A(n_81), .Y(n_183) );
AND2x2_ASAP7_75t_SL g81 ( .A(n_82), .B(n_141), .Y(n_81) );
NOR3xp33_ASAP7_75t_L g82 ( .A(n_83), .B(n_120), .C(n_130), .Y(n_82) );
NAND2xp5_ASAP7_75t_L g83 ( .A(n_84), .B(n_107), .Y(n_83) );
BUFx3_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_97), .Y(n_87) );
AND2x6_ASAP7_75t_L g104 ( .A(n_88), .B(n_105), .Y(n_104) );
AND2x4_ASAP7_75t_L g125 ( .A(n_88), .B(n_114), .Y(n_125) );
AND2x6_ASAP7_75t_L g159 ( .A(n_88), .B(n_152), .Y(n_159) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_94), .Y(n_88) );
AND2x2_ASAP7_75t_L g135 ( .A(n_89), .B(n_95), .Y(n_135) );
INVx2_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
AND2x2_ASAP7_75t_L g112 ( .A(n_90), .B(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_90), .B(n_95), .Y(n_119) );
AND2x2_ASAP7_75t_L g145 ( .A(n_90), .B(n_99), .Y(n_145) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g96 ( .A(n_93), .Y(n_96) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx1_ASAP7_75t_L g113 ( .A(n_95), .Y(n_113) );
INVx1_ASAP7_75t_L g166 ( .A(n_95), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_97), .B(n_112), .Y(n_129) );
AND2x4_ASAP7_75t_L g134 ( .A(n_97), .B(n_135), .Y(n_134) );
AND2x4_ASAP7_75t_L g139 ( .A(n_97), .B(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g97 ( .A(n_98), .B(n_100), .Y(n_97) );
OR2x2_ASAP7_75t_L g106 ( .A(n_98), .B(n_101), .Y(n_106) );
AND2x2_ASAP7_75t_L g114 ( .A(n_98), .B(n_101), .Y(n_114) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x2_ASAP7_75t_L g152 ( .A(n_99), .B(n_101), .Y(n_152) );
INVx1_ASAP7_75t_L g146 ( .A(n_100), .Y(n_146) );
AND2x2_ASAP7_75t_L g165 ( .A(n_100), .B(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g118 ( .A(n_101), .Y(n_118) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx11_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OR2x2_ASAP7_75t_L g176 ( .A(n_106), .B(n_177), .Y(n_176) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx8_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_114), .Y(n_111) );
INVx1_ASAP7_75t_L g154 ( .A(n_113), .Y(n_154) );
NAND2x1p5_ASAP7_75t_L g181 ( .A(n_114), .B(n_135), .Y(n_181) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx6_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
OR2x6_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
INVx1_ASAP7_75t_L g140 ( .A(n_119), .Y(n_140) );
OAI22xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_122), .B1(n_126), .B2(n_127), .Y(n_120) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx6_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OAI22xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_132), .B1(n_136), .B2(n_137), .Y(n_130) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g177 ( .A(n_135), .Y(n_177) );
INVxp67_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NOR3xp33_ASAP7_75t_SL g141 ( .A(n_142), .B(n_155), .C(n_173), .Y(n_141) );
OAI22xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_144), .B1(n_147), .B2(n_148), .Y(n_142) );
NAND2x1p5_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AND2x4_ASAP7_75t_L g164 ( .A(n_145), .B(n_165), .Y(n_164) );
AND2x4_ASAP7_75t_L g171 ( .A(n_145), .B(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
CKINVDCx16_ASAP7_75t_R g149 ( .A(n_150), .Y(n_149) );
OR2x6_ASAP7_75t_L g150 ( .A(n_151), .B(n_153), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
OAI221xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_160), .B1(n_161), .B2(n_167), .C(n_168), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx4_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx4_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_SL g161 ( .A(n_162), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g172 ( .A(n_166), .Y(n_172) );
BUFx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OAI22xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B1(n_178), .B2(n_179), .Y(n_173) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
XNOR2xp5_ASAP7_75t_L g184 ( .A(n_185), .B(n_194), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g193 ( .A(n_187), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_188), .Y(n_192) );
CKINVDCx16_ASAP7_75t_R g197 ( .A(n_198), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_199), .Y(n_198) );
AND3x1_ASAP7_75t_SL g199 ( .A(n_200), .B(n_205), .C(n_208), .Y(n_199) );
INVxp67_ASAP7_75t_L g542 ( .A(n_200), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
OAI21xp5_ASAP7_75t_L g544 ( .A1(n_205), .A2(n_533), .B(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g552 ( .A(n_205), .Y(n_552) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
OAI322xp33_ASAP7_75t_L g537 ( .A1(n_206), .A2(n_538), .A3(n_539), .B1(n_543), .B2(n_546), .C1(n_547), .C2(n_549), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_206), .B(n_209), .Y(n_545) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
OR2x2_ASAP7_75t_SL g551 ( .A(n_208), .B(n_552), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_SL g211 ( .A(n_212), .B(n_497), .Y(n_211) );
NOR3xp33_ASAP7_75t_L g212 ( .A(n_213), .B(n_401), .C(n_485), .Y(n_212) );
NAND4xp25_ASAP7_75t_L g213 ( .A(n_214), .B(n_344), .C(n_366), .D(n_382), .Y(n_213) );
AOI221xp5_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_277), .B1(n_303), .B2(n_322), .C(n_330), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_253), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g356 ( .A(n_217), .B(n_322), .Y(n_356) );
NAND4xp25_ASAP7_75t_L g396 ( .A(n_217), .B(n_384), .C(n_397), .D(n_399), .Y(n_396) );
INVxp67_ASAP7_75t_L g513 ( .A(n_217), .Y(n_513) );
INVx3_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
OR2x2_ASAP7_75t_L g395 ( .A(n_218), .B(n_333), .Y(n_395) );
AND2x2_ASAP7_75t_L g419 ( .A(n_218), .B(n_253), .Y(n_419) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g386 ( .A(n_219), .B(n_321), .Y(n_386) );
AND2x2_ASAP7_75t_L g426 ( .A(n_219), .B(n_407), .Y(n_426) );
AND2x2_ASAP7_75t_L g443 ( .A(n_219), .B(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_219), .B(n_254), .Y(n_467) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g320 ( .A(n_220), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g338 ( .A(n_220), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g350 ( .A(n_220), .B(n_254), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_220), .B(n_264), .Y(n_372) );
OA21x2_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_228), .B(n_252), .Y(n_220) );
OA21x2_ASAP7_75t_L g264 ( .A1(n_221), .A2(n_265), .B(n_275), .Y(n_264) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_223), .Y(n_255) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
AND2x2_ASAP7_75t_SL g276 ( .A(n_224), .B(n_225), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
OAI21xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_242), .B(n_251), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_235), .C(n_238), .Y(n_229) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx3_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g237 ( .A(n_234), .Y(n_237) );
INVx1_ASAP7_75t_L g245 ( .A(n_234), .Y(n_245) );
INVx3_ASAP7_75t_L g311 ( .A(n_236), .Y(n_311) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g283 ( .A(n_237), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_237), .Y(n_284) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_239), .A2(n_315), .B(n_316), .Y(n_314) );
INVx4_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g536 ( .A(n_240), .Y(n_536) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx3_ASAP7_75t_L g250 ( .A(n_241), .Y(n_250) );
BUFx6f_ASAP7_75t_L g273 ( .A(n_241), .Y(n_273) );
INVx1_ASAP7_75t_L g294 ( .A(n_241), .Y(n_294) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_246), .B(n_247), .C(n_248), .Y(n_242) );
O2A1O1Ixp5_ASAP7_75t_L g269 ( .A1(n_243), .A2(n_270), .B(n_271), .C(n_272), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_243), .B(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_248), .A2(n_261), .B(n_262), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_248), .A2(n_273), .B1(n_301), .B2(n_302), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_248), .A2(n_273), .B1(n_326), .B2(n_327), .Y(n_325) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_249), .A2(n_258), .B(n_259), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_249), .A2(n_267), .B(n_268), .Y(n_266) );
O2A1O1Ixp5_ASAP7_75t_SL g310 ( .A1(n_249), .A2(n_311), .B(n_312), .C(n_313), .Y(n_310) );
INVx5_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
OAI22xp5_ASAP7_75t_SL g281 ( .A1(n_250), .A2(n_273), .B1(n_282), .B2(n_285), .Y(n_281) );
OAI21xp5_ASAP7_75t_L g256 ( .A1(n_251), .A2(n_257), .B(n_260), .Y(n_256) );
BUFx3_ASAP7_75t_L g274 ( .A(n_251), .Y(n_274) );
OAI21xp5_ASAP7_75t_L g289 ( .A1(n_251), .A2(n_290), .B(n_295), .Y(n_289) );
OAI21xp5_ASAP7_75t_L g309 ( .A1(n_251), .A2(n_310), .B(n_314), .Y(n_309) );
AND2x2_ASAP7_75t_L g353 ( .A(n_253), .B(n_354), .Y(n_353) );
AOI221xp5_ASAP7_75t_L g402 ( .A1(n_253), .A2(n_403), .B1(n_406), .B2(n_408), .C(n_412), .Y(n_402) );
AND2x2_ASAP7_75t_L g461 ( .A(n_253), .B(n_426), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_253), .B(n_443), .Y(n_495) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_264), .Y(n_253) );
INVx3_ASAP7_75t_L g321 ( .A(n_254), .Y(n_321) );
AND2x2_ASAP7_75t_L g370 ( .A(n_254), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g424 ( .A(n_254), .B(n_339), .Y(n_424) );
AND2x2_ASAP7_75t_L g482 ( .A(n_254), .B(n_483), .Y(n_482) );
OA21x2_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_256), .B(n_263), .Y(n_254) );
INVx4_ASAP7_75t_L g324 ( .A(n_255), .Y(n_324) );
AND2x2_ASAP7_75t_L g322 ( .A(n_264), .B(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g339 ( .A(n_264), .Y(n_339) );
INVx1_ASAP7_75t_L g394 ( .A(n_264), .Y(n_394) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_264), .Y(n_400) );
AND2x2_ASAP7_75t_L g445 ( .A(n_264), .B(n_321), .Y(n_445) );
OR2x2_ASAP7_75t_L g484 ( .A(n_264), .B(n_323), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_269), .B(n_274), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_272), .A2(n_296), .B(n_297), .Y(n_295) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND3xp33_ASAP7_75t_L g343 ( .A(n_274), .B(n_324), .C(n_325), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_274), .B(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g286 ( .A(n_276), .Y(n_286) );
OA21x2_ASAP7_75t_L g288 ( .A1(n_276), .A2(n_289), .B(n_298), .Y(n_288) );
OA21x2_ASAP7_75t_L g308 ( .A1(n_276), .A2(n_309), .B(n_317), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_277), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_287), .Y(n_277) );
AND2x2_ASAP7_75t_L g480 ( .A(n_278), .B(n_477), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_278), .B(n_462), .Y(n_512) );
BUFx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g411 ( .A(n_279), .B(n_335), .Y(n_411) );
AND2x2_ASAP7_75t_L g460 ( .A(n_279), .B(n_306), .Y(n_460) );
INVx1_ASAP7_75t_L g506 ( .A(n_279), .Y(n_506) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_280), .Y(n_319) );
AND2x2_ASAP7_75t_L g361 ( .A(n_280), .B(n_335), .Y(n_361) );
INVx1_ASAP7_75t_L g378 ( .A(n_280), .Y(n_378) );
AND2x2_ASAP7_75t_L g384 ( .A(n_280), .B(n_299), .Y(n_384) );
AND2x2_ASAP7_75t_L g452 ( .A(n_287), .B(n_360), .Y(n_452) );
INVx2_ASAP7_75t_L g517 ( .A(n_287), .Y(n_517) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_299), .Y(n_287) );
AND2x2_ASAP7_75t_L g334 ( .A(n_288), .B(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g347 ( .A(n_288), .B(n_307), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_288), .B(n_306), .Y(n_375) );
INVx1_ASAP7_75t_L g381 ( .A(n_288), .Y(n_381) );
INVx1_ASAP7_75t_L g398 ( .A(n_288), .Y(n_398) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_288), .Y(n_410) );
INVx2_ASAP7_75t_L g478 ( .A(n_288), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_292), .B(n_293), .Y(n_290) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g335 ( .A(n_299), .Y(n_335) );
BUFx2_ASAP7_75t_L g432 ( .A(n_299), .Y(n_432) );
AND2x2_ASAP7_75t_L g477 ( .A(n_299), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_318), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_305), .B(n_414), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_305), .A2(n_476), .B(n_490), .Y(n_500) );
AND2x2_ASAP7_75t_L g525 ( .A(n_305), .B(n_411), .Y(n_525) );
BUFx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g447 ( .A(n_307), .Y(n_447) );
AND2x2_ASAP7_75t_L g476 ( .A(n_307), .B(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_308), .Y(n_360) );
INVx2_ASAP7_75t_L g379 ( .A(n_308), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_308), .B(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx2_ASAP7_75t_L g333 ( .A(n_319), .Y(n_333) );
OR2x2_ASAP7_75t_L g346 ( .A(n_319), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g414 ( .A(n_319), .B(n_410), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_319), .B(n_510), .Y(n_509) );
OR2x2_ASAP7_75t_L g515 ( .A(n_319), .B(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_319), .B(n_452), .Y(n_527) );
AND2x2_ASAP7_75t_L g406 ( .A(n_320), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g429 ( .A(n_320), .B(n_322), .Y(n_429) );
INVx2_ASAP7_75t_L g341 ( .A(n_321), .Y(n_341) );
AND2x2_ASAP7_75t_L g369 ( .A(n_321), .B(n_342), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_321), .B(n_394), .Y(n_450) );
AND2x2_ASAP7_75t_L g364 ( .A(n_322), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g511 ( .A(n_322), .Y(n_511) );
AND2x2_ASAP7_75t_L g523 ( .A(n_322), .B(n_386), .Y(n_523) );
AND2x2_ASAP7_75t_L g349 ( .A(n_323), .B(n_339), .Y(n_349) );
INVx1_ASAP7_75t_L g444 ( .A(n_323), .Y(n_444) );
AO21x1_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_325), .B(n_328), .Y(n_323) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x4_ASAP7_75t_L g342 ( .A(n_329), .B(n_343), .Y(n_342) );
INVxp67_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_336), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_333), .B(n_380), .Y(n_389) );
OR2x2_ASAP7_75t_L g521 ( .A(n_333), .B(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g438 ( .A(n_334), .B(n_379), .Y(n_438) );
AND2x2_ASAP7_75t_L g446 ( .A(n_334), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g505 ( .A(n_334), .B(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g529 ( .A(n_334), .B(n_376), .Y(n_529) );
NOR2xp67_ASAP7_75t_L g487 ( .A(n_335), .B(n_488), .Y(n_487) );
OR2x2_ASAP7_75t_L g516 ( .A(n_335), .B(n_379), .Y(n_516) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2x1p5_ASAP7_75t_L g337 ( .A(n_338), .B(n_340), .Y(n_337) );
AND2x2_ASAP7_75t_L g368 ( .A(n_338), .B(n_369), .Y(n_368) );
INVxp67_ASAP7_75t_L g530 ( .A(n_338), .Y(n_530) );
NOR2x1_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g365 ( .A(n_341), .Y(n_365) );
AND2x2_ASAP7_75t_L g416 ( .A(n_341), .B(n_349), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_341), .B(n_484), .Y(n_510) );
INVx2_ASAP7_75t_L g355 ( .A(n_342), .Y(n_355) );
INVx3_ASAP7_75t_L g407 ( .A(n_342), .Y(n_407) );
OR2x2_ASAP7_75t_L g435 ( .A(n_342), .B(n_436), .Y(n_435) );
AOI311xp33_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_348), .A3(n_350), .B(n_351), .C(n_362), .Y(n_344) );
O2A1O1Ixp33_ASAP7_75t_L g382 ( .A1(n_345), .A2(n_383), .B(n_385), .C(n_387), .Y(n_382) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_SL g367 ( .A(n_347), .Y(n_367) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g385 ( .A(n_349), .B(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_349), .B(n_365), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_349), .B(n_350), .Y(n_518) );
AND2x2_ASAP7_75t_L g440 ( .A(n_350), .B(n_354), .Y(n_440) );
AOI21xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_356), .B(n_357), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g498 ( .A(n_354), .B(n_386), .Y(n_498) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_355), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g392 ( .A(n_355), .Y(n_392) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_361), .Y(n_358) );
AND2x2_ASAP7_75t_L g383 ( .A(n_359), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g428 ( .A(n_361), .Y(n_428) );
AND2x4_ASAP7_75t_L g490 ( .A(n_361), .B(n_459), .Y(n_490) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AOI222xp33_ASAP7_75t_L g441 ( .A1(n_364), .A2(n_430), .B1(n_442), .B2(n_446), .C1(n_448), .C2(n_452), .Y(n_441) );
A2O1A1Ixp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B(n_370), .C(n_373), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_367), .B(n_411), .Y(n_434) );
INVx1_ASAP7_75t_L g456 ( .A(n_369), .Y(n_456) );
INVx1_ASAP7_75t_L g390 ( .A(n_371), .Y(n_390) );
OR2x2_ASAP7_75t_L g455 ( .A(n_372), .B(n_456), .Y(n_455) );
OAI21xp33_ASAP7_75t_SL g373 ( .A1(n_374), .A2(n_376), .B(n_380), .Y(n_373) );
NAND3xp33_ASAP7_75t_L g391 ( .A(n_374), .B(n_392), .C(n_393), .Y(n_391) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_374), .A2(n_411), .B(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_378), .Y(n_431) );
AND2x2_ASAP7_75t_SL g397 ( .A(n_379), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g488 ( .A(n_379), .Y(n_488) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_379), .Y(n_504) );
INVx2_ASAP7_75t_L g462 ( .A(n_380), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_384), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g436 ( .A(n_386), .Y(n_436) );
OAI221xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_390), .B1(n_391), .B2(n_395), .C(n_396), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_390), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_SL g524 ( .A(n_390), .Y(n_524) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g405 ( .A(n_397), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_397), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g463 ( .A(n_397), .B(n_411), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_397), .B(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g496 ( .A(n_397), .B(n_431), .Y(n_496) );
BUFx3_ASAP7_75t_L g459 ( .A(n_398), .Y(n_459) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NAND5xp2_ASAP7_75t_L g401 ( .A(n_402), .B(n_420), .C(n_441), .D(n_453), .E(n_468), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AOI32xp33_ASAP7_75t_L g493 ( .A1(n_405), .A2(n_432), .A3(n_448), .B1(n_494), .B2(n_496), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_407), .B(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_411), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g417 ( .A(n_411), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_415), .B1(n_417), .B2(n_418), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_427), .B1(n_429), .B2(n_430), .C(n_433), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_425), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g492 ( .A(n_424), .B(n_443), .Y(n_492) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g507 ( .A1(n_429), .A2(n_490), .B1(n_508), .B2(n_513), .C(n_514), .Y(n_507) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx2_ASAP7_75t_L g473 ( .A(n_432), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B1(n_437), .B2(n_439), .Y(n_433) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_445), .Y(n_442) );
INVx1_ASAP7_75t_L g451 ( .A(n_443), .Y(n_451) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
AOI222xp33_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_457), .B1(n_461), .B2(n_462), .C1(n_463), .C2(n_464), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_460), .Y(n_457) );
INVxp67_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OAI22xp33_ASAP7_75t_L g508 ( .A1(n_462), .A2(n_509), .B1(n_511), .B2(n_512), .Y(n_508) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_471), .B(n_474), .Y(n_468) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AOI21xp33_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_479), .B(n_481), .Y(n_474) );
INVx2_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g522 ( .A(n_477), .Y(n_522) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
A2O1A1Ixp33_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_489), .B(n_491), .C(n_493), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AOI211xp5_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_499), .B(n_501), .C(n_526), .Y(n_497) );
CKINVDCx16_ASAP7_75t_R g502 ( .A(n_498), .Y(n_502) );
INVxp67_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OAI211xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_503), .B(n_507), .C(n_519), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
AOI21xp33_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_517), .B(n_518), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_523), .B1(n_524), .B2(n_525), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AOI21xp33_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_528), .B(n_530), .Y(n_526) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_532), .Y(n_531) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
CKINVDCx14_ASAP7_75t_R g539 ( .A(n_540), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_541), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_544), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_550), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_551), .Y(n_550) );
endmodule