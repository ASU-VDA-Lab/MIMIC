module fake_jpeg_3490_n_206 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_206);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_19),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_5),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_24),
.B(n_15),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_9),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_28),
.B(n_20),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_30),
.Y(n_73)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_60),
.Y(n_75)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_78),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_66),
.Y(n_93)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_68),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_23),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_81),
.B(n_64),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_59),
.B1(n_58),
.B2(n_72),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_82),
.A2(n_90),
.B1(n_75),
.B2(n_74),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_84),
.B(n_88),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_65),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_91),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_93),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_79),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_67),
.B1(n_56),
.B2(n_52),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_58),
.Y(n_91)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_92),
.Y(n_95)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_90),
.A2(n_76),
.B1(n_52),
.B2(n_62),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_62),
.B1(n_67),
.B2(n_77),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_76),
.B1(n_78),
.B2(n_55),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_97),
.A2(n_102),
.B1(n_109),
.B2(n_77),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_69),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_103),
.B(n_104),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_69),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_65),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_107),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_81),
.B(n_59),
.C(n_73),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_106),
.A2(n_110),
.B(n_83),
.C(n_61),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_94),
.B(n_63),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_73),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_71),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_78),
.B1(n_74),
.B2(n_56),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_51),
.B(n_53),
.C(n_57),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_112),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_86),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_116),
.B1(n_118),
.B2(n_126),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_99),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_115),
.B(n_117),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_71),
.B1(n_63),
.B2(n_83),
.Y(n_118)
);

NOR3xp33_ASAP7_75t_SL g151 ( 
.A(n_120),
.B(n_119),
.C(n_132),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_70),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_122),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_0),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_124),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_26),
.C(n_50),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_112),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_127),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_89),
.B1(n_2),
.B2(n_3),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_1),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_95),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_130),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_89),
.B1(n_27),
.B2(n_31),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_129),
.A2(n_132),
.B1(n_7),
.B2(n_8),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_89),
.B1(n_4),
.B2(n_5),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_101),
.A2(n_1),
.B1(n_4),
.B2(n_6),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_110),
.B(n_101),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_125),
.A2(n_6),
.B(n_7),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_138),
.A2(n_136),
.B(n_139),
.Y(n_159)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_140),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_143),
.Y(n_166)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_130),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_146),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_8),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_145),
.B(n_149),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_36),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_10),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_152),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_10),
.Y(n_152)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_37),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_11),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_49),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_163),
.C(n_165),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_158),
.B(n_170),
.Y(n_184)
);

AOI221xp5_ASAP7_75t_L g178 ( 
.A1(n_159),
.A2(n_151),
.B1(n_147),
.B2(n_140),
.C(n_148),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_153),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_162),
.A2(n_147),
.B1(n_155),
.B2(n_134),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_146),
.Y(n_163)
);

OA21x2_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_35),
.B(n_47),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_164),
.A2(n_138),
.B(n_144),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_34),
.C(n_46),
.Y(n_165)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_137),
.Y(n_174)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_183),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_48),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_181),
.C(n_182),
.Y(n_190)
);

OAI322xp33_ASAP7_75t_L g180 ( 
.A1(n_160),
.A2(n_45),
.A3(n_44),
.B1(n_43),
.B2(n_39),
.C1(n_38),
.C2(n_21),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_165),
.C(n_156),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_22),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_12),
.C(n_13),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_181),
.A2(n_159),
.B(n_166),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_191),
.C(n_175),
.Y(n_197)
);

OAI321xp33_ASAP7_75t_L g186 ( 
.A1(n_184),
.A2(n_164),
.A3(n_171),
.B1(n_173),
.B2(n_169),
.C(n_162),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_186),
.B(n_187),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_176),
.A2(n_172),
.B(n_167),
.Y(n_191)
);

AO21x1_ASAP7_75t_L g192 ( 
.A1(n_179),
.A2(n_158),
.B(n_161),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_192),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_182),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_196),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_192),
.Y(n_196)
);

AOI31xp67_ASAP7_75t_L g198 ( 
.A1(n_197),
.A2(n_175),
.A3(n_190),
.B(n_21),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_199),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_16),
.C(n_17),
.Y(n_199)
);

AOI21x1_ASAP7_75t_L g202 ( 
.A1(n_201),
.A2(n_200),
.B(n_193),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_193),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_203),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_22),
.Y(n_205)
);

BUFx24_ASAP7_75t_SL g206 ( 
.A(n_205),
.Y(n_206)
);


endmodule