module fake_jpeg_27209_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_6),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_19),
.Y(n_25)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_18),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_8),
.B(n_16),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_22),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

AO21x1_ASAP7_75t_L g30 ( 
.A1(n_24),
.A2(n_13),
.B(n_21),
.Y(n_30)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_34),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_24),
.A2(n_15),
.B(n_14),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_31),
.A2(n_32),
.B(n_36),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_23),
.A2(n_17),
.B1(n_15),
.B2(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_37),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_25),
.A2(n_20),
.B1(n_18),
.B2(n_11),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_10),
.B1(n_12),
.B2(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_12),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_27),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_41),
.C(n_32),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_27),
.C(n_10),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2x1_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_26),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_46),
.B1(n_47),
.B2(n_44),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_10),
.C(n_3),
.Y(n_47)
);

INVxp67_ASAP7_75t_SL g49 ( 
.A(n_48),
.Y(n_49)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_R g51 ( 
.A1(n_45),
.A2(n_44),
.B(n_40),
.C(n_43),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_53),
.A2(n_51),
.B(n_38),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_55),
.B1(n_53),
.B2(n_52),
.Y(n_56)
);

OAI321xp33_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_41),
.A3(n_49),
.B1(n_42),
.B2(n_7),
.C(n_4),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_52),
.C(n_3),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_52),
.Y(n_59)
);


endmodule