module fake_netlist_6_772_n_20591 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_135, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_20591);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_135;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_20591;

wire n_5643;
wire n_18652;
wire n_2817;
wire n_18318;
wire n_2576;
wire n_1674;
wire n_16664;
wire n_19057;
wire n_11926;
wire n_6441;
wire n_8668;
wire n_1212;
wire n_208;
wire n_4251;
wire n_11111;
wire n_7933;
wire n_578;
wire n_4395;
wire n_19613;
wire n_1061;
wire n_16335;
wire n_5653;
wire n_4978;
wire n_13125;
wire n_3088;
wire n_8186;
wire n_6725;
wire n_6126;
wire n_4699;
wire n_17647;
wire n_8899;
wire n_5345;
wire n_17634;
wire n_10053;
wire n_1930;
wire n_19785;
wire n_8534;
wire n_3376;
wire n_4868;
wire n_10020;
wire n_19715;
wire n_17991;
wire n_15665;
wire n_19382;
wire n_1555;
wire n_17735;
wire n_20091;
wire n_19161;
wire n_7161;
wire n_19232;
wire n_830;
wire n_7868;
wire n_15764;
wire n_5725;
wire n_447;
wire n_5229;
wire n_3427;
wire n_18903;
wire n_18105;
wire n_5101;
wire n_3071;
wire n_8561;
wire n_14998;
wire n_14944;
wire n_11954;
wire n_19220;
wire n_14341;
wire n_10392;
wire n_15074;
wire n_5545;
wire n_2321;
wire n_15253;
wire n_4501;
wire n_9626;
wire n_5598;
wire n_20377;
wire n_19097;
wire n_15898;
wire n_18013;
wire n_7389;
wire n_10719;
wire n_20151;
wire n_5259;
wire n_6913;
wire n_10015;
wire n_6948;
wire n_3929;
wire n_3048;
wire n_9362;
wire n_7401;
wire n_7516;
wire n_12767;
wire n_16095;
wire n_18502;
wire n_5930;
wire n_9658;
wire n_1971;
wire n_5354;
wire n_8426;
wire n_5908;
wire n_953;
wire n_19755;
wire n_3664;
wire n_13681;
wire n_5420;
wire n_17209;
wire n_6243;
wire n_4414;
wire n_6585;
wire n_16553;
wire n_18122;
wire n_2625;
wire n_11543;
wire n_4646;
wire n_7651;
wire n_2843;
wire n_3760;
wire n_14662;
wire n_13247;
wire n_16286;
wire n_7956;
wire n_20321;
wire n_7369;
wire n_16549;
wire n_15421;
wire n_5136;
wire n_20011;
wire n_15964;
wire n_5638;
wire n_9100;
wire n_6784;
wire n_18310;
wire n_10868;
wire n_9067;
wire n_6323;
wire n_17847;
wire n_14431;
wire n_17478;
wire n_13515;
wire n_6110;
wire n_1967;
wire n_11684;
wire n_16324;
wire n_14410;
wire n_15800;
wire n_9400;
wire n_1911;
wire n_13139;
wire n_7774;
wire n_15600;
wire n_16267;
wire n_20471;
wire n_6951;
wire n_15899;
wire n_19991;
wire n_279;
wire n_18317;
wire n_2735;
wire n_13729;
wire n_4671;
wire n_18709;
wire n_14813;
wire n_4314;
wire n_18002;
wire n_19810;
wire n_323;
wire n_14628;
wire n_8421;
wire n_1381;
wire n_331;
wire n_2093;
wire n_18863;
wire n_17854;
wire n_10114;
wire n_10357;
wire n_15762;
wire n_2770;
wire n_16351;
wire n_15883;
wire n_17706;
wire n_8389;
wire n_2917;
wire n_13711;
wire n_16721;
wire n_12742;
wire n_3923;
wire n_11768;
wire n_9267;
wire n_939;
wire n_19401;
wire n_9652;
wire n_5493;
wire n_8849;
wire n_9059;
wire n_15332;
wire n_5346;
wire n_5252;
wire n_3446;
wire n_18445;
wire n_5309;
wire n_1895;
wire n_4698;
wire n_16254;
wire n_7564;
wire n_3859;
wire n_14989;
wire n_17564;
wire n_10204;
wire n_6383;
wire n_3397;
wire n_18669;
wire n_11637;
wire n_3575;
wire n_8151;
wire n_2469;
wire n_9038;
wire n_16004;
wire n_8748;
wire n_20487;
wire n_13984;
wire n_5452;
wire n_6794;
wire n_18608;
wire n_8718;
wire n_2764;
wire n_9935;
wire n_6990;
wire n_14288;
wire n_14824;
wire n_18699;
wire n_8223;
wire n_4856;
wire n_3492;
wire n_9135;
wire n_16800;
wire n_13771;
wire n_18644;
wire n_11295;
wire n_4291;
wire n_13960;
wire n_5532;
wire n_5897;
wire n_2434;
wire n_9070;
wire n_11708;
wire n_15629;
wire n_14401;
wire n_10827;
wire n_3247;
wire n_5922;
wire n_14922;
wire n_7569;
wire n_7823;
wire n_9477;
wire n_7062;
wire n_12158;
wire n_14769;
wire n_355;
wire n_14961;
wire n_8577;
wire n_20559;
wire n_8594;
wire n_8428;
wire n_9829;
wire n_13341;
wire n_20345;
wire n_2254;
wire n_5058;
wire n_10685;
wire n_1926;
wire n_17139;
wire n_15185;
wire n_12083;
wire n_12014;
wire n_14803;
wire n_19270;
wire n_19816;
wire n_1747;
wire n_16035;
wire n_10607;
wire n_15490;
wire n_18033;
wire n_5042;
wire n_19569;
wire n_8164;
wire n_20485;
wire n_4072;
wire n_835;
wire n_928;
wire n_15100;
wire n_10368;
wire n_19137;
wire n_9088;
wire n_10183;
wire n_17161;
wire n_6952;
wire n_11464;
wire n_19421;
wire n_3997;
wire n_14878;
wire n_15046;
wire n_2468;
wire n_5144;
wire n_10383;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_3434;
wire n_4510;
wire n_6776;
wire n_13550;
wire n_17601;
wire n_13348;
wire n_2812;
wire n_10724;
wire n_16398;
wire n_19396;
wire n_9988;
wire n_7009;
wire n_2136;
wire n_2409;
wire n_3834;
wire n_12795;
wire n_11553;
wire n_2075;
wire n_10876;
wire n_18780;
wire n_9137;
wire n_11180;
wire n_14043;
wire n_18820;
wire n_3192;
wire n_8995;
wire n_1546;
wire n_4394;
wire n_6010;
wire n_20006;
wire n_3352;
wire n_8711;
wire n_12505;
wire n_18602;
wire n_2150;
wire n_4082;
wire n_1420;
wire n_13721;
wire n_18430;
wire n_20018;
wire n_10820;
wire n_13514;
wire n_8306;
wire n_7488;
wire n_2558;
wire n_13194;
wire n_8887;
wire n_18677;
wire n_16183;
wire n_4289;
wire n_11866;
wire n_13575;
wire n_11450;
wire n_12522;
wire n_15659;
wire n_1487;
wire n_9578;
wire n_13109;
wire n_7438;
wire n_20003;
wire n_20224;
wire n_16631;
wire n_14355;
wire n_7337;
wire n_9489;
wire n_14123;
wire n_5957;
wire n_10728;
wire n_6357;
wire n_925;
wire n_6800;
wire n_18962;
wire n_4322;
wire n_10655;
wire n_9797;
wire n_1249;
wire n_2693;
wire n_8332;
wire n_9478;
wire n_2767;
wire n_11379;
wire n_16627;
wire n_19571;
wire n_19659;
wire n_19944;
wire n_10670;
wire n_5929;
wire n_5787;
wire n_11981;
wire n_19181;
wire n_9351;
wire n_5445;
wire n_14556;
wire n_6839;
wire n_532;
wire n_173;
wire n_9189;
wire n_413;
wire n_18888;
wire n_16528;
wire n_2170;
wire n_4156;
wire n_14701;
wire n_7098;
wire n_16587;
wire n_19933;
wire n_18936;
wire n_3158;
wire n_1788;
wire n_20502;
wire n_8921;
wire n_20404;
wire n_9356;
wire n_15880;
wire n_16499;
wire n_1835;
wire n_5076;
wire n_18328;
wire n_5870;
wire n_9175;
wire n_6508;
wire n_12013;
wire n_11835;
wire n_4995;
wire n_10959;
wire n_6809;
wire n_11233;
wire n_4310;
wire n_7782;
wire n_5212;
wire n_13385;
wire n_2689;
wire n_1473;
wire n_6636;
wire n_5286;
wire n_16339;
wire n_1246;
wire n_4528;
wire n_899;
wire n_13992;
wire n_17429;
wire n_19103;
wire n_13790;
wire n_4914;
wire n_499;
wire n_3418;
wire n_705;
wire n_1004;
wire n_10624;
wire n_13304;
wire n_14633;
wire n_15699;
wire n_11900;
wire n_2297;
wire n_5901;
wire n_6538;
wire n_5599;
wire n_12883;
wire n_5324;
wire n_2103;
wire n_8983;
wire n_10422;
wire n_3770;
wire n_9818;
wire n_4402;
wire n_927;
wire n_16503;
wire n_18974;
wire n_12367;
wire n_17360;
wire n_5009;
wire n_13526;
wire n_12563;
wire n_7243;
wire n_13321;
wire n_15042;
wire n_15519;
wire n_14722;
wire n_13427;
wire n_4627;
wire n_4079;
wire n_9909;
wire n_19607;
wire n_8620;
wire n_19204;
wire n_15264;
wire n_13270;
wire n_10052;
wire n_10109;
wire n_18151;
wire n_3390;
wire n_19582;
wire n_10448;
wire n_11196;
wire n_16239;
wire n_11963;
wire n_16334;
wire n_9571;
wire n_8424;
wire n_2137;
wire n_16003;
wire n_4798;
wire n_2532;
wire n_12655;
wire n_7941;
wire n_16096;
wire n_18628;
wire n_11483;
wire n_15067;
wire n_19591;
wire n_19345;
wire n_5089;
wire n_13356;
wire n_2849;
wire n_14912;
wire n_1398;
wire n_884;
wire n_19177;
wire n_731;
wire n_8907;
wire n_11080;
wire n_958;
wire n_5137;
wire n_20447;
wire n_17557;
wire n_14079;
wire n_15168;
wire n_9894;
wire n_8324;
wire n_15411;
wire n_9441;
wire n_6380;
wire n_10906;
wire n_7913;
wire n_15144;
wire n_5288;
wire n_3606;
wire n_819;
wire n_14224;
wire n_2788;
wire n_10380;
wire n_6449;
wire n_18687;
wire n_6461;
wire n_3892;
wire n_18273;
wire n_4069;
wire n_14682;
wire n_2748;
wire n_5194;
wire n_1834;
wire n_9033;
wire n_2331;
wire n_15031;
wire n_12933;
wire n_15718;
wire n_9537;
wire n_11297;
wire n_14635;
wire n_17076;
wire n_13893;
wire n_5947;
wire n_1877;
wire n_2030;
wire n_11946;
wire n_9443;
wire n_9996;
wire n_14950;
wire n_20205;
wire n_7800;
wire n_13795;
wire n_3026;
wire n_17501;
wire n_14547;
wire n_15416;
wire n_221;
wire n_20562;
wire n_3847;
wire n_2552;
wire n_17942;
wire n_18735;
wire n_9938;
wire n_7261;
wire n_9023;
wire n_14415;
wire n_11818;
wire n_16298;
wire n_18739;
wire n_6773;
wire n_13569;
wire n_7455;
wire n_18042;
wire n_19105;
wire n_2160;
wire n_9201;
wire n_6531;
wire n_10952;
wire n_2131;
wire n_13628;
wire n_18958;
wire n_9559;
wire n_11803;
wire n_15738;
wire n_16301;
wire n_8015;
wire n_18507;
wire n_1933;
wire n_19102;
wire n_15613;
wire n_14786;
wire n_4411;
wire n_9184;
wire n_13585;
wire n_18418;
wire n_18472;
wire n_8024;
wire n_12562;
wire n_18396;
wire n_4180;
wire n_16531;
wire n_20243;
wire n_3354;
wire n_11090;
wire n_19035;
wire n_5740;
wire n_5820;
wire n_13266;
wire n_13957;
wire n_9403;
wire n_9875;
wire n_5180;
wire n_2049;
wire n_5182;
wire n_11561;
wire n_19956;
wire n_5534;
wire n_8003;
wire n_8785;
wire n_3566;
wire n_17826;
wire n_2829;
wire n_8692;
wire n_6889;
wire n_16142;
wire n_9183;
wire n_3804;
wire n_4207;
wire n_14326;
wire n_5196;
wire n_16381;
wire n_10852;
wire n_4470;
wire n_9529;
wire n_3901;
wire n_465;
wire n_11425;
wire n_4704;
wire n_2142;
wire n_4596;
wire n_6478;
wire n_820;
wire n_6100;
wire n_6516;
wire n_17845;
wire n_6977;
wire n_16854;
wire n_17542;
wire n_7660;
wire n_2263;
wire n_6911;
wire n_6599;
wire n_6522;
wire n_17189;
wire n_5660;
wire n_2756;
wire n_5334;
wire n_9347;
wire n_807;
wire n_4761;
wire n_18879;
wire n_16395;
wire n_13603;
wire n_6207;
wire n_6931;
wire n_7948;
wire n_238;
wire n_9082;
wire n_1595;
wire n_8685;
wire n_6963;
wire n_16252;
wire n_4932;
wire n_19358;
wire n_5456;
wire n_10618;
wire n_9594;
wire n_7837;
wire n_19531;
wire n_9445;
wire n_7627;
wire n_9803;
wire n_20572;
wire n_16698;
wire n_17041;
wire n_7601;
wire n_3195;
wire n_6346;
wire n_19833;
wire n_4274;
wire n_15729;
wire n_17519;
wire n_5386;
wire n_14737;
wire n_11676;
wire n_12266;
wire n_2595;
wire n_16949;
wire n_12287;
wire n_19713;
wire n_13485;
wire n_12991;
wire n_11134;
wire n_13735;
wire n_8886;
wire n_7211;
wire n_10933;
wire n_5618;
wire n_8506;
wire n_2264;
wire n_6494;
wire n_16365;
wire n_13041;
wire n_11548;
wire n_17037;
wire n_13154;
wire n_7822;
wire n_6453;
wire n_9307;
wire n_10762;
wire n_11342;
wire n_7785;
wire n_1891;
wire n_1213;
wire n_2235;
wire n_11266;
wire n_19706;
wire n_5082;
wire n_5338;
wire n_12479;
wire n_8352;
wire n_18941;
wire n_10360;
wire n_9450;
wire n_2298;
wire n_490;
wire n_3594;
wire n_5689;
wire n_16777;
wire n_4165;
wire n_12454;
wire n_8143;
wire n_10480;
wire n_4626;
wire n_4144;
wire n_12537;
wire n_17183;
wire n_9693;
wire n_17582;
wire n_12921;
wire n_2169;
wire n_13567;
wire n_11957;
wire n_10633;
wire n_13686;
wire n_13645;
wire n_16753;
wire n_12215;
wire n_18473;
wire n_9880;
wire n_12467;
wire n_6329;
wire n_11607;
wire n_11546;
wire n_15259;
wire n_16946;
wire n_15460;
wire n_330;
wire n_7158;
wire n_20546;
wire n_1406;
wire n_13400;
wire n_9905;
wire n_18717;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_13331;
wire n_9456;
wire n_20285;
wire n_7044;
wire n_9710;
wire n_8623;
wire n_11113;
wire n_18593;
wire n_2518;
wire n_17769;
wire n_19193;
wire n_13812;
wire n_14970;
wire n_7838;
wire n_4842;
wire n_204;
wire n_482;
wire n_4135;
wire n_16969;
wire n_1845;
wire n_12731;
wire n_7518;
wire n_2798;
wire n_6147;
wire n_9199;
wire n_13544;
wire n_7791;
wire n_2753;
wire n_2007;
wire n_2039;
wire n_18172;
wire n_12616;
wire n_1544;
wire n_18333;
wire n_3437;
wire n_4111;
wire n_14375;
wire n_12653;
wire n_533;
wire n_7146;
wire n_18081;
wire n_16580;
wire n_18498;
wire n_4859;
wire n_9363;
wire n_12047;
wire n_12587;
wire n_10747;
wire n_13110;
wire n_16628;
wire n_2973;
wire n_9422;
wire n_18344;
wire n_5218;
wire n_12348;
wire n_3665;
wire n_16929;
wire n_273;
wire n_16099;
wire n_15590;
wire n_10843;
wire n_7888;
wire n_11823;
wire n_5358;
wire n_6397;
wire n_16869;
wire n_3174;
wire n_10997;
wire n_1948;
wire n_19855;
wire n_9010;
wire n_13707;
wire n_15241;
wire n_19640;
wire n_6073;
wire n_19157;
wire n_6331;
wire n_13498;
wire n_2283;
wire n_9341;
wire n_7848;
wire n_6939;
wire n_18289;
wire n_11408;
wire n_4196;
wire n_2056;
wire n_13183;
wire n_12519;
wire n_17184;
wire n_4902;
wire n_6405;
wire n_7580;
wire n_14077;
wire n_13007;
wire n_2680;
wire n_10112;
wire n_7304;
wire n_3713;
wire n_1931;
wire n_502;
wire n_1257;
wire n_20065;
wire n_3197;
wire n_7223;
wire n_7833;
wire n_14868;
wire n_5512;
wire n_9297;
wire n_2398;
wire n_6206;
wire n_9068;
wire n_8136;
wire n_5033;
wire n_9808;
wire n_18534;
wire n_2695;
wire n_4035;
wire n_7445;
wire n_11086;
wire n_6529;
wire n_1949;
wire n_3759;
wire n_4516;
wire n_1804;
wire n_11710;
wire n_251;
wire n_6290;
wire n_10253;
wire n_6025;
wire n_1337;
wire n_6455;
wire n_15277;
wire n_18435;
wire n_13804;
wire n_12455;
wire n_13099;
wire n_4492;
wire n_19524;
wire n_18516;
wire n_5607;
wire n_7695;
wire n_7179;
wire n_7122;
wire n_12157;
wire n_5999;
wire n_19676;
wire n_6203;
wire n_15806;
wire n_13064;
wire n_7630;
wire n_16246;
wire n_20013;
wire n_8643;
wire n_15660;
wire n_15357;
wire n_8565;
wire n_10821;
wire n_19784;
wire n_13648;
wire n_4542;
wire n_6892;
wire n_4462;
wire n_15722;
wire n_14181;
wire n_15278;
wire n_18054;
wire n_13338;
wire n_6685;
wire n_11639;
wire n_4931;
wire n_14213;
wire n_17320;
wire n_17885;
wire n_7051;
wire n_8477;
wire n_19766;
wire n_9793;
wire n_11692;
wire n_15054;
wire n_14842;
wire n_13115;
wire n_1291;
wire n_11759;
wire n_20195;
wire n_8230;
wire n_12549;
wire n_20388;
wire n_5911;
wire n_11601;
wire n_11971;
wire n_2122;
wire n_12314;
wire n_3503;
wire n_1065;
wire n_11116;
wire n_12604;
wire n_13305;
wire n_1255;
wire n_8876;
wire n_5124;
wire n_19017;
wire n_3951;
wire n_9359;
wire n_14189;
wire n_3874;
wire n_15761;
wire n_5123;
wire n_8060;
wire n_3027;
wire n_4083;
wire n_11124;
wire n_6392;
wire n_182;
wire n_17470;
wire n_15301;
wire n_7351;
wire n_9352;
wire n_2746;
wire n_389;
wire n_7608;
wire n_17053;
wire n_15567;
wire n_6832;
wire n_7394;
wire n_13202;
wire n_15350;
wire n_13638;
wire n_4171;
wire n_17948;
wire n_14392;
wire n_19953;
wire n_19347;
wire n_7027;
wire n_1105;
wire n_7992;
wire n_6912;
wire n_10330;
wire n_1461;
wire n_8276;
wire n_2076;
wire n_3567;
wire n_11465;
wire n_8027;
wire n_4705;
wire n_3807;
wire n_17808;
wire n_11265;
wire n_11125;
wire n_1114;
wire n_17244;
wire n_20348;
wire n_7783;
wire n_13220;
wire n_10276;
wire n_191;
wire n_10594;
wire n_8978;
wire n_8245;
wire n_15072;
wire n_12910;
wire n_18725;
wire n_18215;
wire n_8454;
wire n_2881;
wire n_1116;
wire n_8891;
wire n_1219;
wire n_11690;
wire n_18719;
wire n_19142;
wire n_16194;
wire n_3897;
wire n_5591;
wire n_11373;
wire n_3372;
wire n_6403;
wire n_7947;
wire n_1221;
wire n_16826;
wire n_20370;
wire n_6491;
wire n_19519;
wire n_16321;
wire n_14072;
wire n_17120;
wire n_11412;
wire n_13039;
wire n_13130;
wire n_10441;
wire n_19500;
wire n_17237;
wire n_5518;
wire n_15671;
wire n_9124;
wire n_6661;
wire n_13719;
wire n_8847;
wire n_14548;
wire n_19099;
wire n_4068;
wire n_10841;
wire n_16076;
wire n_12313;
wire n_18071;
wire n_2743;
wire n_4766;
wire n_20266;
wire n_14661;
wire n_8356;
wire n_6136;
wire n_16384;
wire n_16416;
wire n_3378;
wire n_15305;
wire n_15588;
wire n_3745;
wire n_8888;
wire n_11810;
wire n_14267;
wire n_5357;
wire n_3523;
wire n_2222;
wire n_13062;
wire n_7857;
wire n_3176;
wire n_7481;
wire n_14130;
wire n_14930;
wire n_5541;
wire n_10576;
wire n_16596;
wire n_334;
wire n_6668;
wire n_2999;
wire n_15548;
wire n_1239;
wire n_3697;
wire n_16714;
wire n_19168;
wire n_2408;
wire n_6859;
wire n_18752;
wire n_13752;
wire n_10237;
wire n_19484;
wire n_13596;
wire n_12889;
wire n_18092;
wire n_12050;
wire n_12922;
wire n_12250;
wire n_9515;
wire n_6971;
wire n_17957;
wire n_9642;
wire n_393;
wire n_20470;
wire n_14231;
wire n_12385;
wire n_13219;
wire n_17449;
wire n_5443;
wire n_5673;
wire n_6351;
wire n_9382;
wire n_16392;
wire n_6212;
wire n_7668;
wire n_9775;
wire n_19207;
wire n_13295;
wire n_3936;
wire n_1349;
wire n_16906;
wire n_18194;
wire n_17693;
wire n_6829;
wire n_2723;
wire n_17981;
wire n_3496;
wire n_13160;
wire n_15249;
wire n_11071;
wire n_5473;
wire n_17337;
wire n_10072;
wire n_10708;
wire n_13818;
wire n_15024;
wire n_8803;
wire n_3239;
wire n_3902;
wire n_4062;
wire n_18478;
wire n_4396;
wire n_19898;
wire n_9706;
wire n_3101;
wire n_15174;
wire n_17904;
wire n_3374;
wire n_10387;
wire n_13764;
wire n_20258;
wire n_19408;
wire n_1552;
wire n_11224;
wire n_8790;
wire n_15569;
wire n_4293;
wire n_10219;
wire n_1031;
wire n_11924;
wire n_15193;
wire n_9591;
wire n_6137;
wire n_14833;
wire n_10364;
wire n_11422;
wire n_8338;
wire n_4412;
wire n_14480;
wire n_12489;
wire n_8491;
wire n_2217;
wire n_4781;
wire n_16610;
wire n_9283;
wire n_19299;
wire n_12030;
wire n_206;
wire n_20330;
wire n_633;
wire n_12565;
wire n_15236;
wire n_1040;
wire n_3059;
wire n_9468;
wire n_14098;
wire n_14482;
wire n_17174;
wire n_14223;
wire n_15962;
wire n_5424;
wire n_12415;
wire n_3017;
wire n_1805;
wire n_17332;
wire n_10559;
wire n_13173;
wire n_15355;
wire n_15945;
wire n_14848;
wire n_18548;
wire n_7154;
wire n_16232;
wire n_8304;
wire n_19644;
wire n_19012;
wire n_11418;
wire n_6655;
wire n_19694;
wire n_19187;
wire n_3274;
wire n_9958;
wire n_14544;
wire n_4457;
wire n_7320;
wire n_4928;
wire n_5769;
wire n_16122;
wire n_722;
wire n_5613;
wire n_18852;
wire n_14604;
wire n_14735;
wire n_2223;
wire n_1621;
wire n_19572;
wire n_19688;
wire n_13101;
wire n_6786;
wire n_8315;
wire n_16446;
wire n_15885;
wire n_17528;
wire n_18964;
wire n_11040;
wire n_11754;
wire n_14916;
wire n_9756;
wire n_4762;
wire n_192;
wire n_13748;
wire n_11672;
wire n_3113;
wire n_10353;
wire n_10847;
wire n_10451;
wire n_1458;
wire n_15801;
wire n_17778;
wire n_5303;
wire n_12240;
wire n_12003;
wire n_7496;
wire n_223;
wire n_4154;
wire n_12165;
wire n_19894;
wire n_10866;
wire n_18127;
wire n_9940;
wire n_6200;
wire n_4504;
wire n_14600;
wire n_3844;
wire n_1237;
wire n_11763;
wire n_15010;
wire n_8465;
wire n_6670;
wire n_3741;
wire n_18730;
wire n_10653;
wire n_8535;
wire n_11587;
wire n_6373;
wire n_12280;
wire n_13461;
wire n_20253;
wire n_12492;
wire n_19535;
wire n_16282;
wire n_17011;
wire n_2243;
wire n_4898;
wire n_5601;
wire n_13188;
wire n_4819;
wire n_17639;
wire n_7131;
wire n_20271;
wire n_20416;
wire n_9586;
wire n_8909;
wire n_3332;
wire n_18977;
wire n_16356;
wire n_11843;
wire n_2570;
wire n_14614;
wire n_4645;
wire n_11629;
wire n_15147;
wire n_9554;
wire n_18246;
wire n_5635;
wire n_17180;
wire n_5091;
wire n_6546;
wire n_4302;
wire n_15927;
wire n_3395;
wire n_7060;
wire n_19439;
wire n_13217;
wire n_5363;
wire n_4178;
wire n_5165;
wire n_16332;
wire n_1711;
wire n_20489;
wire n_14397;
wire n_17971;
wire n_10853;
wire n_13802;
wire n_18559;
wire n_7761;
wire n_20055;
wire n_10338;
wire n_12978;
wire n_1422;
wire n_15668;
wire n_15137;
wire n_8496;
wire n_1842;
wire n_12476;
wire n_8568;
wire n_516;
wire n_8852;
wire n_18423;
wire n_12023;
wire n_20560;
wire n_17655;
wire n_8637;
wire n_2703;
wire n_6168;
wire n_16225;
wire n_16677;
wire n_4606;
wire n_13413;
wire n_6450;
wire n_15153;
wire n_13203;
wire n_2058;
wire n_2660;
wire n_19128;
wire n_14462;
wire n_8456;
wire n_4962;
wire n_4563;
wire n_7137;
wire n_14933;
wire n_5056;
wire n_9920;
wire n_12598;
wire n_9039;
wire n_11854;
wire n_8573;
wire n_2124;
wire n_19070;
wire n_5336;
wire n_18623;
wire n_5447;
wire n_17389;
wire n_13230;
wire n_7743;
wire n_6179;
wire n_19230;
wire n_9125;
wire n_20244;
wire n_9139;
wire n_20080;
wire n_17941;
wire n_5747;
wire n_12733;
wire n_13750;
wire n_8775;
wire n_14104;
wire n_808;
wire n_20228;
wire n_18695;
wire n_14684;
wire n_5753;
wire n_12245;
wire n_15713;
wire n_1193;
wire n_18124;
wire n_14572;
wire n_9972;
wire n_6083;
wire n_12909;
wire n_6434;
wire n_551;
wire n_9157;
wire n_16417;
wire n_3884;
wire n_17880;
wire n_9324;
wire n_5808;
wire n_8807;
wire n_6933;
wire n_8521;
wire n_6547;
wire n_5193;
wire n_9442;
wire n_20145;
wire n_1481;
wire n_19374;
wire n_6984;
wire n_18394;
wire n_17392;
wire n_10763;
wire n_9957;
wire n_12759;
wire n_11793;
wire n_7106;
wire n_7213;
wire n_17586;
wire n_5961;
wire n_18757;
wire n_6507;
wire n_9313;
wire n_6687;
wire n_9173;
wire n_6690;
wire n_7412;
wire n_12144;
wire n_9160;
wire n_219;
wire n_9974;
wire n_19365;
wire n_12129;
wire n_14753;
wire n_13658;
wire n_5533;
wire n_20222;
wire n_14671;
wire n_4257;
wire n_16454;
wire n_17977;
wire n_18441;
wire n_13572;
wire n_15547;
wire n_12032;
wire n_4720;
wire n_14674;
wire n_3857;
wire n_243;
wire n_1873;
wire n_19496;
wire n_3630;
wire n_6524;
wire n_3518;
wire n_12835;
wire n_10129;
wire n_16089;
wire n_1330;
wire n_7523;
wire n_8654;
wire n_2876;
wire n_15060;
wire n_14229;
wire n_11241;
wire n_15520;
wire n_5953;
wire n_14188;
wire n_11508;
wire n_7141;
wire n_5198;
wire n_16139;
wire n_5718;
wire n_6505;
wire n_1663;
wire n_12636;
wire n_4172;
wire n_3403;
wire n_11227;
wire n_1107;
wire n_20221;
wire n_3294;
wire n_6001;
wire n_11218;
wire n_4502;
wire n_318;
wire n_10195;
wire n_13722;
wire n_3490;
wire n_4849;
wire n_277;
wire n_4319;
wire n_7327;
wire n_3369;
wire n_12938;
wire n_13057;
wire n_8367;
wire n_7367;
wire n_3581;
wire n_16439;
wire n_6023;
wire n_14897;
wire n_19251;
wire n_12173;
wire n_6905;
wire n_17520;
wire n_15925;
wire n_18255;
wire n_19275;
wire n_7368;
wire n_429;
wire n_5553;
wire n_8011;
wire n_4066;
wire n_10263;
wire n_4340;
wire n_5790;
wire n_15141;
wire n_12411;
wire n_10280;
wire n_20484;
wire n_4004;
wire n_5404;
wire n_18634;
wire n_4292;
wire n_8570;
wire n_6163;
wire n_7628;
wire n_9074;
wire n_5549;
wire n_9408;
wire n_267;
wire n_6553;
wire n_1124;
wire n_1624;
wire n_19190;
wire n_12568;
wire n_3280;
wire n_16163;
wire n_13478;
wire n_18256;
wire n_12970;
wire n_1515;
wire n_8902;
wire n_14295;
wire n_7557;
wire n_20022;
wire n_593;
wire n_7128;
wire n_14367;
wire n_637;
wire n_13915;
wire n_7594;
wire n_15057;
wire n_19479;
wire n_16300;
wire n_19236;
wire n_18288;
wire n_10504;
wire n_2525;
wire n_7788;
wire n_13783;
wire n_5154;
wire n_10658;
wire n_11590;
wire n_11238;
wire n_3889;
wire n_2687;
wire n_2887;
wire n_2194;
wire n_5637;
wire n_1987;
wire n_7586;
wire n_968;
wire n_7767;
wire n_8294;
wire n_12279;
wire n_9419;
wire n_16402;
wire n_13705;
wire n_17986;
wire n_17771;
wire n_9277;
wire n_9257;
wire n_17773;
wire n_2391;
wire n_2431;
wire n_17070;
wire n_5843;
wire n_8170;
wire n_18515;
wire n_11558;
wire n_9159;
wire n_7744;
wire n_10595;
wire n_7748;
wire n_6827;
wire n_20167;
wire n_19958;
wire n_18914;
wire n_11073;
wire n_1208;
wire n_20308;
wire n_1072;
wire n_815;
wire n_7485;
wire n_18867;
wire n_11974;
wire n_12881;
wire n_15736;
wire n_14986;
wire n_14920;
wire n_8671;
wire n_19196;
wire n_15313;
wire n_284;
wire n_3436;
wire n_9671;
wire n_1026;
wire n_289;
wire n_14994;
wire n_10080;
wire n_16505;
wire n_12228;
wire n_10570;
wire n_16120;
wire n_20119;
wire n_12929;
wire n_16065;
wire n_685;
wire n_3240;
wire n_15075;
wire n_12261;
wire n_18007;
wire n_12106;
wire n_5333;
wire n_5594;
wire n_12291;
wire n_14510;
wire n_12124;
wire n_11755;
wire n_9510;
wire n_18055;
wire n_13497;
wire n_15406;
wire n_19529;
wire n_14396;
wire n_2517;
wire n_2713;
wire n_11918;
wire n_11748;
wire n_12433;
wire n_5000;
wire n_5551;
wire n_8701;
wire n_16810;
wire n_6499;
wire n_19678;
wire n_18158;
wire n_12217;
wire n_15922;
wire n_12097;
wire n_5257;
wire n_8097;
wire n_13851;
wire n_9679;
wire n_8645;
wire n_13272;
wire n_18954;
wire n_4688;
wire n_4058;
wire n_3082;
wire n_4848;
wire n_16411;
wire n_19507;
wire n_156;
wire n_16717;
wire n_8824;
wire n_11673;
wire n_2407;
wire n_3799;
wire n_7712;
wire n_2574;
wire n_4475;
wire n_6276;
wire n_10499;
wire n_8340;
wire n_5854;
wire n_11387;
wire n_19975;
wire n_11333;
wire n_2667;
wire n_18425;
wire n_1571;
wire n_2948;
wire n_8455;
wire n_7208;
wire n_13613;
wire n_947;
wire n_12185;
wire n_9770;
wire n_1992;
wire n_8681;
wire n_11417;
wire n_7406;
wire n_16044;
wire n_18656;
wire n_3140;
wire n_4749;
wire n_9592;
wire n_5155;
wire n_17507;
wire n_9180;
wire n_10922;
wire n_926;
wire n_19013;
wire n_10718;
wire n_1698;
wire n_4100;
wire n_13821;
wire n_19198;
wire n_13712;
wire n_9625;
wire n_777;
wire n_15041;
wire n_4085;
wire n_15393;
wire n_4464;
wire n_14144;
wire n_6851;
wire n_6460;
wire n_19429;
wire n_4659;
wire n_5217;
wire n_6650;
wire n_8221;
wire n_11682;
wire n_20583;
wire n_15595;
wire n_8255;
wire n_15081;
wire n_8461;
wire n_6368;
wire n_1857;
wire n_16474;
wire n_20184;
wire n_6583;
wire n_4866;
wire n_4889;
wire n_3638;
wire n_16940;
wire n_4816;
wire n_17419;
wire n_20295;
wire n_12520;
wire n_2110;
wire n_1659;
wire n_3393;
wire n_17134;
wire n_3451;
wire n_11459;
wire n_4937;
wire n_10904;
wire n_11317;
wire n_5277;
wire n_8792;
wire n_12436;
wire n_16344;
wire n_2053;
wire n_12808;
wire n_4222;
wire n_18275;
wire n_2710;
wire n_6064;
wire n_1966;
wire n_13801;
wire n_5793;
wire n_19286;
wire n_19920;
wire n_8523;
wire n_12143;
wire n_4976;
wire n_13879;
wire n_5578;
wire n_18064;
wire n_231;
wire n_1457;
wire n_20084;
wire n_1993;
wire n_11806;
wire n_2617;
wire n_19682;
wire n_1466;
wire n_11050;
wire n_5207;
wire n_17714;
wire n_5676;
wire n_1893;
wire n_4665;
wire n_11484;
wire n_2387;
wire n_19483;
wire n_2846;
wire n_19183;
wire n_10295;
wire n_1980;
wire n_5464;
wire n_2237;
wire n_20418;
wire n_10336;
wire n_4362;
wire n_7716;
wire n_17903;
wire n_20256;
wire n_8954;
wire n_12212;
wire n_20277;
wire n_7540;
wire n_775;
wire n_13231;
wire n_12624;
wire n_1531;
wire n_453;
wire n_8552;
wire n_17412;
wire n_7558;
wire n_4261;
wire n_8373;
wire n_13165;
wire n_426;
wire n_3986;
wire n_12151;
wire n_17407;
wire n_15204;
wire n_2556;
wire n_4747;
wire n_5251;
wire n_18284;
wire n_20188;
wire n_9970;
wire n_11365;
wire n_18138;
wire n_3175;
wire n_17016;
wire n_16081;
wire n_5475;
wire n_15341;
wire n_4448;
wire n_1096;
wire n_15477;
wire n_6233;
wire n_6377;
wire n_12402;
wire n_17959;
wire n_18782;
wire n_19942;
wire n_688;
wire n_1077;
wire n_4132;
wire n_10361;
wire n_1437;
wire n_7143;
wire n_10424;
wire n_8965;
wire n_4355;
wire n_18454;
wire n_2276;
wire n_13476;
wire n_2803;
wire n_379;
wire n_18399;
wire n_12162;
wire n_3202;
wire n_602;
wire n_17087;
wire n_7497;
wire n_4655;
wire n_11829;
wire n_11517;
wire n_7793;
wire n_16102;
wire n_587;
wire n_16274;
wire n_3554;
wire n_6991;
wire n_10556;
wire n_13776;
wire n_7248;
wire n_7204;
wire n_15835;
wire n_12852;
wire n_10567;
wire n_7578;
wire n_3462;
wire n_13343;
wire n_7654;
wire n_5132;
wire n_17339;
wire n_10230;
wire n_12675;
wire n_5627;
wire n_5774;
wire n_13907;
wire n_4846;
wire n_2984;
wire n_5187;
wire n_12821;
wire n_14782;
wire n_4024;
wire n_18756;
wire n_7120;
wire n_6335;
wire n_12837;
wire n_8728;
wire n_8386;
wire n_14070;
wire n_14330;
wire n_13491;
wire n_4860;
wire n_18654;
wire n_15748;
wire n_3414;
wire n_17995;
wire n_14235;
wire n_6173;
wire n_14851;
wire n_18012;
wire n_10058;
wire n_16471;
wire n_2563;
wire n_19434;
wire n_4989;
wire n_7757;
wire n_1683;
wire n_17539;
wire n_280;
wire n_6630;
wire n_1187;
wire n_4558;
wire n_16560;
wire n_8396;
wire n_6612;
wire n_13450;
wire n_6606;
wire n_3550;
wire n_19533;
wire n_14178;
wire n_5508;
wire n_20314;
wire n_12907;
wire n_15500;
wire n_14891;
wire n_17051;
wire n_9318;
wire n_6158;
wire n_11917;
wire n_9028;
wire n_17217;
wire n_4328;
wire n_8020;
wire n_1057;
wire n_9374;
wire n_20386;
wire n_2785;
wire n_2636;
wire n_13634;
wire n_18027;
wire n_10413;
wire n_3399;
wire n_19268;
wire n_1611;
wire n_19948;
wire n_2740;
wire n_17786;
wire n_4808;
wire n_5767;
wire n_1589;
wire n_12708;
wire n_4712;
wire n_10369;
wire n_2309;
wire n_6821;
wire n_5462;
wire n_9983;
wire n_6688;
wire n_8580;
wire n_9993;
wire n_3533;
wire n_13622;
wire n_4725;
wire n_11207;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3132;
wire n_16951;
wire n_6798;
wire n_10838;
wire n_10530;
wire n_14794;
wire n_17684;
wire n_9237;
wire n_13931;
wire n_14404;
wire n_6557;
wire n_18302;
wire n_6753;
wire n_18164;
wire n_17151;
wire n_7341;
wire n_4908;
wire n_12088;
wire n_15423;
wire n_14377;
wire n_6639;
wire n_12508;
wire n_12096;
wire n_5150;
wire n_8832;
wire n_3819;
wire n_20059;
wire n_2050;
wire n_19412;
wire n_19399;
wire n_2164;
wire n_11098;
wire n_15815;
wire n_20537;
wire n_5179;
wire n_7957;
wire n_10938;
wire n_6627;
wire n_17147;
wire n_3544;
wire n_2904;
wire n_18019;
wire n_10927;
wire n_4616;
wire n_4982;
wire n_370;
wire n_8592;
wire n_11204;
wire n_6190;
wire n_1979;
wire n_2738;
wire n_16920;
wire n_12701;
wire n_20187;
wire n_10578;
wire n_4323;
wire n_16199;
wire n_19113;
wire n_6615;
wire n_17331;
wire n_2342;
wire n_2167;
wire n_7294;
wire n_4017;
wire n_11811;
wire n_13745;
wire n_10569;
wire n_2541;
wire n_8622;
wire n_2940;
wire n_4739;
wire n_15367;
wire n_19095;
wire n_8104;
wire n_2768;
wire n_18511;
wire n_17428;
wire n_4298;
wire n_2314;
wire n_10746;
wire n_9188;
wire n_16407;
wire n_18009;
wire n_4644;
wire n_19002;
wire n_8779;
wire n_5503;
wire n_5945;
wire n_10697;
wire n_11714;
wire n_16179;
wire n_2390;
wire n_15070;
wire n_1343;
wire n_20040;
wire n_2734;
wire n_7250;
wire n_8762;
wire n_17503;
wire n_18365;
wire n_17358;
wire n_1900;
wire n_3381;
wire n_13419;
wire n_9207;
wire n_11860;
wire n_17057;
wire n_10926;
wire n_8897;
wire n_11503;
wire n_17104;
wire n_4672;
wire n_8376;
wire n_18271;
wire n_2939;
wire n_18998;
wire n_5749;
wire n_1672;
wire n_15640;
wire n_6271;
wire n_15683;
wire n_16202;
wire n_4598;
wire n_8599;
wire n_13460;
wire n_15451;
wire n_5993;
wire n_15233;
wire n_6716;
wire n_9637;
wire n_11636;
wire n_9418;
wire n_8616;
wire n_13105;
wire n_14467;
wire n_20154;
wire n_14789;
wire n_13076;
wire n_15526;
wire n_12950;
wire n_8628;
wire n_19867;
wire n_15150;
wire n_13028;
wire n_8547;
wire n_4424;
wire n_7113;
wire n_1751;
wire n_20510;
wire n_10433;
wire n_285;
wire n_9116;
wire n_14096;
wire n_11983;
wire n_10839;
wire n_11813;
wire n_3506;
wire n_1928;
wire n_14583;
wire n_4317;
wire n_14893;
wire n_20148;
wire n_20504;
wire n_8275;
wire n_6198;
wire n_5418;
wire n_18270;
wire n_6762;
wire n_4088;
wire n_3711;
wire n_19826;
wire n_9035;
wire n_729;
wire n_16960;
wire n_3642;
wire n_14915;
wire n_4650;
wire n_17780;
wire n_438;
wire n_17075;
wire n_2874;
wire n_1200;
wire n_4967;
wire n_9678;
wire n_8247;
wire n_6577;
wire n_12956;
wire n_17373;
wire n_14856;
wire n_15235;
wire n_4912;
wire n_9284;
wire n_5086;
wire n_4735;
wire n_187;
wire n_20039;
wire n_3300;
wire n_2978;
wire n_15711;
wire n_1050;
wire n_5170;
wire n_7604;
wire n_3515;
wire n_1150;
wire n_9606;
wire n_17018;
wire n_13459;
wire n_1023;
wire n_1118;
wire n_14268;
wire n_194;
wire n_2949;
wire n_10297;
wire n_12553;
wire n_19928;
wire n_5028;
wire n_5839;
wire n_1814;
wire n_1631;
wire n_14127;
wire n_440;
wire n_3806;
wire n_8827;
wire n_2931;
wire n_19884;
wire n_3866;
wire n_17937;
wire n_9549;
wire n_14894;
wire n_12866;
wire n_17801;
wire n_4157;
wire n_6845;
wire n_9482;
wire n_3629;
wire n_969;
wire n_8877;
wire n_9412;
wire n_15561;
wire n_6321;
wire n_6819;
wire n_10136;
wire n_15148;
wire n_16457;
wire n_19560;
wire n_11356;
wire n_1379;
wire n_15955;
wire n_214;
wire n_8688;
wire n_4910;
wire n_20250;
wire n_3083;
wire n_10692;
wire n_14826;
wire n_16421;
wire n_15776;
wire n_11280;
wire n_14987;
wire n_8686;
wire n_12239;
wire n_17641;
wire n_19823;
wire n_3830;
wire n_8403;
wire n_11493;
wire n_17742;
wire n_3117;
wire n_8588;
wire n_15229;
wire n_11339;
wire n_15804;
wire n_5623;
wire n_15269;
wire n_20394;
wire n_10471;
wire n_2385;
wire n_4112;
wire n_3739;
wire n_14946;
wire n_18727;
wire n_15674;
wire n_4352;
wire n_17933;
wire n_8780;
wire n_17384;
wire n_7958;
wire n_18037;
wire n_4980;
wire n_11885;
wire n_1924;
wire n_15855;
wire n_3363;
wire n_10777;
wire n_3721;
wire n_16490;
wire n_7760;
wire n_13306;
wire n_9753;
wire n_8722;
wire n_16489;
wire n_19580;
wire n_8589;
wire n_3969;
wire n_20130;
wire n_7573;
wire n_6281;
wire n_7364;
wire n_5647;
wire n_13133;
wire n_4256;
wire n_4938;
wire n_8608;
wire n_12874;
wire n_11480;
wire n_11194;
wire n_10469;
wire n_445;
wire n_18650;
wire n_930;
wire n_9342;
wire n_18062;
wire n_2620;
wire n_9329;
wire n_1945;
wire n_5426;
wire n_19257;
wire n_17119;
wire n_9868;
wire n_1414;
wire n_7048;
wire n_944;
wire n_16491;
wire n_2744;
wire n_1011;
wire n_1566;
wire n_8145;
wire n_8928;
wire n_17638;
wire n_7682;
wire n_990;
wire n_18584;
wire n_6231;
wire n_12509;
wire n_14902;
wire n_6932;
wire n_13527;
wire n_7901;
wire n_870;
wire n_366;
wire n_5709;
wire n_7658;
wire n_10055;
wire n_10979;
wire n_19753;
wire n_19765;
wire n_3802;
wire n_6996;
wire n_15935;
wire n_17674;
wire n_376;
wire n_2111;
wire n_10408;
wire n_16180;
wire n_8572;
wire n_17182;
wire n_6337;
wire n_18212;
wire n_3643;
wire n_2425;
wire n_8227;
wire n_12936;
wire n_18424;
wire n_19947;
wire n_3060;
wire n_10482;
wire n_4105;
wire n_7405;
wire n_14151;
wire n_4926;
wire n_1518;
wire n_20538;
wire n_9386;
wire n_15120;
wire n_8314;
wire n_11121;
wire n_3038;
wire n_11270;
wire n_6310;
wire n_11689;
wire n_10003;
wire n_15601;
wire n_15936;
wire n_20426;
wire n_10321;
wire n_5310;
wire n_9661;
wire n_20452;
wire n_14284;
wire n_3863;
wire n_5722;
wire n_4640;
wire n_13232;
wire n_13001;
wire n_17377;
wire n_9901;
wire n_17334;
wire n_2805;
wire n_5593;
wire n_4769;
wire n_8934;
wire n_13059;
wire n_6365;
wire n_4628;
wire n_8407;
wire n_15455;
wire n_8567;
wire n_11288;
wire n_12772;
wire n_5237;
wire n_409;
wire n_11042;
wire n_10726;
wire n_16534;
wire n_19304;
wire n_4460;
wire n_4108;
wire n_14681;
wire n_11272;
wire n_14230;
wire n_5853;
wire n_8283;
wire n_5011;
wire n_14546;
wire n_20361;
wire n_9882;
wire n_16484;
wire n_10637;
wire n_9205;
wire n_17464;
wire n_7972;
wire n_1675;
wire n_13512;
wire n_7916;
wire n_9368;
wire n_13069;
wire n_12362;
wire n_19038;
wire n_6167;
wire n_13233;
wire n_18495;
wire n_8008;
wire n_18833;
wire n_13297;
wire n_20551;
wire n_2553;
wire n_6307;
wire n_149;
wire n_632;
wire n_2038;
wire n_7483;
wire n_14873;
wire n_19891;
wire n_9504;
wire n_14840;
wire n_16556;
wire n_6267;
wire n_5998;
wire n_17861;
wire n_6568;
wire n_19083;
wire n_7507;
wire n_7159;
wire n_18038;
wire n_6028;
wire n_1417;
wire n_16072;
wire n_14083;
wire n_681;
wire n_10189;
wire n_8697;
wire n_6813;
wire n_6669;
wire n_422;
wire n_8420;
wire n_8297;
wire n_3079;
wire n_10881;
wire n_13519;
wire n_16583;
wire n_20425;
wire n_15641;
wire n_16007;
wire n_17129;
wire n_19869;
wire n_4853;
wire n_8639;
wire n_16796;
wire n_16510;
wire n_531;
wire n_15892;
wire n_4272;
wire n_14049;
wire n_1025;
wire n_7562;
wire n_3111;
wire n_336;
wire n_12019;
wire n_8176;
wire n_14529;
wire n_17624;
wire n_16106;
wire n_10891;
wire n_9026;
wire n_10803;
wire n_13190;
wire n_6188;
wire n_5262;
wire n_4670;
wire n_4882;
wire n_11695;
wire n_17595;
wire n_4738;
wire n_8113;
wire n_18922;
wire n_15877;
wire n_1307;
wire n_11453;
wire n_19233;
wire n_17896;
wire n_19088;
wire n_5713;
wire n_16445;
wire n_168;
wire n_6318;
wire n_2353;
wire n_16997;
wire n_4099;
wire n_14690;
wire n_19252;
wire n_17356;
wire n_1738;
wire n_10290;
wire n_19705;
wire n_11862;
wire n_14839;
wire n_15409;
wire n_16207;
wire n_9433;
wire n_18568;
wire n_11660;
wire n_14249;
wire n_14241;
wire n_6604;
wire n_2386;
wire n_5373;
wire n_1724;
wire n_16101;
wire n_3708;
wire n_6391;
wire n_10284;
wire n_14446;
wire n_14719;
wire n_15575;
wire n_19896;
wire n_8522;
wire n_12971;
wire n_7942;
wire n_16599;
wire n_6473;
wire n_18620;
wire n_15696;
wire n_14558;
wire n_19695;
wire n_11318;
wire n_17198;
wire n_7725;
wire n_16950;
wire n_20517;
wire n_20131;
wire n_8626;
wire n_1393;
wire n_1867;
wire n_1603;
wire n_19277;
wire n_5466;
wire n_19475;
wire n_15095;
wire n_5955;
wire n_658;
wire n_1874;
wire n_11487;
wire n_2825;
wire n_8441;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_7778;
wire n_758;
wire n_2256;
wire n_4060;
wire n_8397;
wire n_5796;
wire n_17916;
wire n_8726;
wire n_17250;
wire n_770;
wire n_6958;
wire n_15417;
wire n_16615;
wire n_14667;
wire n_6523;
wire n_14713;
wire n_4687;
wire n_7531;
wire n_18686;
wire n_1404;
wire n_13214;
wire n_8615;
wire n_15975;
wire n_11062;
wire n_14202;
wire n_15859;
wire n_11933;
wire n_14554;
wire n_9887;
wire n_4600;
wire n_20380;
wire n_13211;
wire n_8316;
wire n_5829;
wire n_19654;
wire n_8057;
wire n_5191;
wire n_1231;
wire n_14874;
wire n_20566;
wire n_18198;
wire n_2370;
wire n_18550;
wire n_4253;
wire n_407;
wire n_913;
wire n_16824;
wire n_15098;
wire n_867;
wire n_16832;
wire n_13336;
wire n_1333;
wire n_2496;
wire n_16074;
wire n_3189;
wire n_19487;
wire n_18664;
wire n_13102;
wire n_4691;
wire n_12894;
wire n_10492;
wire n_15769;
wire n_4297;
wire n_17340;
wire n_9247;
wire n_8378;
wire n_2907;
wire n_577;
wire n_10526;
wire n_5575;
wire n_8725;
wire n_9570;
wire n_5675;
wire n_12356;
wire n_2778;
wire n_19454;
wire n_11077;
wire n_1909;
wire n_5020;
wire n_9846;
wire n_13262;
wire n_1123;
wire n_10764;
wire n_18005;
wire n_18429;
wire n_9677;
wire n_3934;
wire n_4033;
wire n_6804;
wire n_6603;
wire n_17812;
wire n_3193;
wire n_7534;
wire n_8201;
wire n_4354;
wire n_16485;
wire n_9348;
wire n_14262;
wire n_1530;
wire n_8696;
wire n_938;
wire n_6396;
wire n_20072;
wire n_12630;
wire n_6890;
wire n_549;
wire n_4377;
wire n_12022;
wire n_19929;
wire n_905;
wire n_10741;
wire n_6109;
wire n_14727;
wire n_12425;
wire n_14762;
wire n_322;
wire n_689;
wire n_13507;
wire n_10915;
wire n_18290;
wire n_558;
wire n_3036;
wire n_7943;
wire n_11743;
wire n_8892;
wire n_12199;
wire n_17133;
wire n_17729;
wire n_15410;
wire n_4511;
wire n_2908;
wire n_9707;
wire n_16002;
wire n_16258;
wire n_13594;
wire n_20096;
wire n_10680;
wire n_3599;
wire n_5543;
wire n_5885;
wire n_14228;
wire n_5356;
wire n_3772;
wire n_5458;
wire n_16131;
wire n_11473;
wire n_5038;
wire n_1760;
wire n_19856;
wire n_4585;
wire n_2664;
wire n_1722;
wire n_11726;
wire n_15944;
wire n_12574;
wire n_20407;
wire n_8833;
wire n_10142;
wire n_7828;
wire n_9918;
wire n_18643;
wire n_15932;
wire n_16345;
wire n_4427;
wire n_9390;
wire n_19997;
wire n_10069;
wire n_17325;
wire n_3549;
wire n_5714;
wire n_8541;
wire n_2804;
wire n_2453;
wire n_18233;
wire n_5510;
wire n_5555;
wire n_13678;
wire n_12458;
wire n_19291;
wire n_6066;
wire n_14582;
wire n_6897;
wire n_13523;
wire n_9619;
wire n_11171;
wire n_15117;
wire n_19868;
wire n_4886;
wire n_9187;
wire n_2733;
wire n_16621;
wire n_13819;
wire n_15777;
wire n_14424;
wire n_18398;
wire n_14523;
wire n_11063;
wire n_18846;
wire n_20435;
wire n_9989;
wire n_8319;
wire n_4200;
wire n_3460;
wire n_12853;
wire n_12942;
wire n_9259;
wire n_3519;
wire n_12397;
wire n_16555;
wire n_15336;
wire n_14161;
wire n_6573;
wire n_16760;
wire n_7634;
wire n_5078;
wire n_13290;
wire n_13500;
wire n_11440;
wire n_16844;
wire n_10483;
wire n_17758;
wire n_4737;
wire n_4116;
wire n_20158;
wire n_7285;
wire n_11337;
wire n_12005;
wire n_11243;
wire n_8929;
wire n_9360;
wire n_18610;
wire n_9824;
wire n_342;
wire n_15089;
wire n_2658;
wire n_2665;
wire n_20088;
wire n_8233;
wire n_6130;
wire n_7273;
wire n_14750;
wire n_17939;
wire n_5976;
wire n_14074;
wire n_20325;
wire n_840;
wire n_2913;
wire n_12800;
wire n_2230;
wire n_1969;
wire n_1565;
wire n_16574;
wire n_15145;
wire n_17516;
wire n_8187;
wire n_9399;
wire n_15838;
wire n_15297;
wire n_13979;
wire n_9740;
wire n_615;
wire n_12947;
wire n_5371;
wire n_20297;
wire n_20327;
wire n_4651;
wire n_17178;
wire n_20576;
wire n_9764;
wire n_4854;
wire n_20349;
wire n_15160;
wire n_3789;
wire n_605;
wire n_12354;
wire n_12666;
wire n_14297;
wire n_7597;
wire n_17388;
wire n_16368;
wire n_12631;
wire n_1646;
wire n_19154;
wire n_14969;
wire n_14820;
wire n_10133;
wire n_18426;
wire n_18073;
wire n_19995;
wire n_6921;
wire n_14675;
wire n_18905;
wire n_9826;
wire n_3171;
wire n_3608;
wire n_11942;
wire n_15998;
wire n_3459;
wire n_19138;
wire n_6624;
wire n_6956;
wire n_12966;
wire n_15851;
wire n_15884;
wire n_5656;
wire n_5125;
wire n_7329;
wire n_14502;
wire n_14533;
wire n_5652;
wire n_17935;
wire n_10752;
wire n_18630;
wire n_10067;
wire n_18021;
wire n_19841;
wire n_10399;
wire n_12498;
wire n_656;
wire n_11010;
wire n_9590;
wire n_16017;
wire n_2717;
wire n_11588;
wire n_16346;
wire n_738;
wire n_13956;
wire n_3497;
wire n_7418;
wire n_6880;
wire n_19305;
wire n_3580;
wire n_12387;
wire n_19783;
wire n_9497;
wire n_13255;
wire n_15911;
wire n_2307;
wire n_3704;
wire n_684;
wire n_9219;
wire n_17376;
wire n_8028;
wire n_4280;
wire n_8914;
wire n_1181;
wire n_15276;
wire n_8391;
wire n_16343;
wire n_13749;
wire n_15552;
wire n_17722;
wire n_19370;
wire n_16228;
wire n_803;
wire n_1817;
wire n_12862;
wire n_13621;
wire n_8216;
wire n_2868;
wire n_16953;
wire n_2231;
wire n_3609;
wire n_9982;
wire n_7804;
wire n_18948;
wire n_12656;
wire n_8313;
wire n_14828;
wire n_7656;
wire n_19150;
wire n_19971;
wire n_8263;
wire n_6438;
wire n_11936;
wire n_19132;
wire n_10374;
wire n_7332;
wire n_10382;
wire n_18247;
wire n_4455;
wire n_8374;
wire n_13223;
wire n_13451;
wire n_4514;
wire n_13939;
wire n_18909;
wire n_13728;
wire n_4806;
wire n_7386;
wire n_17824;
wire n_11018;
wire n_10981;
wire n_16014;
wire n_2682;
wire n_13379;
wire n_13781;
wire n_19311;
wire n_5098;
wire n_17513;
wire n_10344;
wire n_5707;
wire n_14613;
wire n_19451;
wire n_11515;
wire n_17466;
wire n_3505;
wire n_15881;
wire n_7637;
wire n_16577;
wire n_10318;
wire n_4796;
wire n_4442;
wire n_18422;
wire n_2581;
wire n_18091;
wire n_12890;
wire n_20067;
wire n_3590;
wire n_13994;
wire n_954;
wire n_5344;
wire n_4419;
wire n_17060;
wire n_11972;
wire n_13484;
wire n_17298;
wire n_8460;
wire n_3327;
wire n_20462;
wire n_17468;
wire n_14593;
wire n_2701;
wire n_16013;
wire n_1080;
wire n_7409;
wire n_19266;
wire n_10735;
wire n_17153;
wire n_13807;
wire n_9825;
wire n_2784;
wire n_5494;
wire n_7444;
wire n_16942;
wire n_2421;
wire n_17569;
wire n_4387;
wire n_2618;
wire n_2464;
wire n_5128;
wire n_18661;
wire n_14033;
wire n_2224;
wire n_10393;
wire n_1092;
wire n_15221;
wire n_5467;
wire n_16090;
wire n_18467;
wire n_4890;
wire n_1784;
wire n_9045;
wire n_12281;
wire n_9373;
wire n_14337;
wire n_2929;
wire n_11809;
wire n_17994;
wire n_9967;
wire n_13553;
wire n_20291;
wire n_4236;
wire n_7187;
wire n_19039;
wire n_17063;
wire n_19692;
wire n_1831;
wire n_9182;
wire n_5079;
wire n_9365;
wire n_18960;
wire n_10909;
wire n_6336;
wire n_10083;
wire n_18891;
wire n_9224;
wire n_10347;
wire n_6541;
wire n_12410;
wire n_4706;
wire n_16327;
wire n_19238;
wire n_14707;
wire n_16043;
wire n_19677;
wire n_4622;
wire n_14612;
wire n_12294;
wire n_7603;
wire n_10667;
wire n_2732;
wire n_17688;
wire n_4206;
wire n_2249;
wire n_18794;
wire n_5835;
wire n_7979;
wire n_13382;
wire n_11675;
wire n_20094;
wire n_15543;
wire n_15906;
wire n_8657;
wire n_8006;
wire n_8296;
wire n_2955;
wire n_11083;
wire n_17418;
wire n_2158;
wire n_7866;
wire n_3367;
wire n_7205;
wire n_18283;
wire n_2202;
wire n_736;
wire n_11728;
wire n_2993;
wire n_4754;
wire n_11698;
wire n_4647;
wire n_9556;
wire n_8590;
wire n_16682;
wire n_4030;
wire n_1995;
wire n_17038;
wire n_15798;
wire n_4760;
wire n_11326;
wire n_6421;
wire n_19743;
wire n_11870;
wire n_7407;
wire n_20193;
wire n_6328;
wire n_11283;
wire n_6236;
wire n_11834;
wire n_13361;
wire n_17286;
wire n_4509;
wire n_15061;
wire n_2875;
wire n_1103;
wire n_6144;
wire n_11506;
wire n_10135;
wire n_13161;
wire n_144;
wire n_2219;
wire n_14010;
wire n_16413;
wire n_999;
wire n_4897;
wire n_19796;
wire n_15030;
wire n_18205;
wire n_9152;
wire n_3539;
wire n_16451;
wire n_19965;
wire n_19590;
wire n_8364;
wire n_3276;
wire n_15228;
wire n_15832;
wire n_10720;
wire n_10535;
wire n_19349;
wire n_17629;
wire n_17536;
wire n_3886;
wire n_6708;
wire n_11236;
wire n_18793;
wire n_4420;
wire n_892;
wire n_19987;
wire n_18529;
wire n_6242;
wire n_12379;
wire n_1468;
wire n_2855;
wire n_2156;
wire n_18222;
wire n_12932;
wire n_14078;
wire n_3548;
wire n_18985;
wire n_8548;
wire n_19793;
wire n_10672;
wire n_7645;
wire n_14222;
wire n_16990;
wire n_20155;
wire n_3141;
wire n_5096;
wire n_1841;
wire n_12114;
wire n_10308;
wire n_11608;
wire n_14430;
wire n_1015;
wire n_10623;
wire n_4797;
wire n_6285;
wire n_4270;
wire n_16545;
wire n_19339;
wire n_13709;
wire n_4945;
wire n_17713;
wire n_5677;
wire n_9454;
wire n_10586;
wire n_8742;
wire n_12626;
wire n_11967;
wire n_9253;
wire n_15084;
wire n_13559;
wire n_20332;
wire n_8874;
wire n_5927;
wire n_15071;
wire n_11996;
wire n_9566;
wire n_11338;
wire n_13426;
wire n_1356;
wire n_4333;
wire n_18826;
wire n_7666;
wire n_11250;
wire n_15328;
wire n_1452;
wire n_2854;
wire n_7963;
wire n_6398;
wire n_8329;
wire n_302;
wire n_9503;
wire n_8270;
wire n_16051;
wire n_11738;
wire n_18196;
wire n_3217;
wire n_1983;
wire n_11522;
wire n_7737;
wire n_16569;
wire n_8614;
wire n_18459;
wire n_9568;
wire n_15621;
wire n_18411;
wire n_20170;
wire n_8816;
wire n_9119;
wire n_19337;
wire n_13529;
wire n_6224;
wire n_3279;
wire n_18293;
wire n_2402;
wire n_20455;
wire n_1081;
wire n_19616;
wire n_1084;
wire n_6614;
wire n_5912;
wire n_18395;
wire n_20379;
wire n_3501;
wire n_374;
wire n_12554;
wire n_8035;
wire n_12722;
wire n_6735;
wire n_17445;
wire n_20581;
wire n_10491;
wire n_921;
wire n_12037;
wire n_15371;
wire n_17572;
wire n_13453;
wire n_15080;
wire n_20178;
wire n_5265;
wire n_2257;
wire n_9943;
wire n_12391;
wire n_14242;
wire n_15622;
wire n_7152;
wire n_2200;
wire n_9575;
wire n_10409;
wire n_4548;
wire n_11822;
wire n_10521;
wire n_9610;
wire n_16483;
wire n_14016;
wire n_12323;
wire n_15566;
wire n_20298;
wire n_10527;
wire n_3115;
wire n_7570;
wire n_2084;
wire n_4875;
wire n_7817;
wire n_5682;
wire n_5387;
wire n_654;
wire n_11394;
wire n_2458;
wire n_3050;
wire n_9928;
wire n_11820;
wire n_13897;
wire n_2527;
wire n_14792;
wire n_16290;
wire n_14248;
wire n_8370;
wire n_164;
wire n_13300;
wire n_16296;
wire n_5681;
wire n_20521;
wire n_7566;
wire n_11940;
wire n_1271;
wire n_4901;
wire n_9217;
wire n_12901;
wire n_4040;
wire n_10518;
wire n_20480;
wire n_2406;
wire n_7617;
wire n_15170;
wire n_16936;
wire n_19262;
wire n_9771;
wire n_15774;
wire n_5316;
wire n_7718;
wire n_244;
wire n_13844;
wire n_19246;
wire n_7396;
wire n_282;
wire n_18543;
wire n_5703;
wire n_18930;
wire n_833;
wire n_523;
wire n_7998;
wire n_12432;
wire n_7561;
wire n_18349;
wire n_6810;
wire n_2196;
wire n_17010;
wire n_17040;
wire n_16130;
wire n_12879;
wire n_5564;
wire n_13746;
wire n_12559;
wire n_13508;
wire n_14660;
wire n_4530;
wire n_9899;
wire n_19930;
wire n_13004;
wire n_5406;
wire n_13479;
wire n_8277;
wire n_652;
wire n_18014;
wire n_1906;
wire n_14437;
wire n_4841;
wire n_1758;
wire n_13759;
wire n_5806;
wire n_4338;
wire n_10486;
wire n_306;
wire n_16613;
wire n_8724;
wire n_5738;
wire n_15938;
wire n_17216;
wire n_3151;
wire n_15146;
wire n_3779;
wire n_2388;
wire n_3984;
wire n_9995;
wire n_5710;
wire n_9076;
wire n_12351;
wire n_16360;
wire n_19146;
wire n_19878;
wire n_13359;
wire n_10372;
wire n_3558;
wire n_14867;
wire n_1984;
wire n_2236;
wire n_6044;
wire n_8867;
wire n_9491;
wire n_4326;
wire n_12702;
wire n_17811;
wire n_15188;
wire n_2834;
wire n_12439;
wire n_19478;
wire n_11008;
wire n_6125;
wire n_7314;
wire n_786;
wire n_14186;
wire n_7526;
wire n_17816;
wire n_5040;
wire n_14023;
wire n_19758;
wire n_17890;
wire n_10736;
wire n_19550;
wire n_11575;
wire n_7004;
wire n_14418;
wire n_8308;
wire n_18897;
wire n_151;
wire n_8165;
wire n_14283;
wire n_4788;
wire n_8400;
wire n_18177;
wire n_5977;
wire n_10446;
wire n_7879;
wire n_16372;
wire n_1908;
wire n_15958;
wire n_18853;
wire n_7696;
wire n_11570;
wire n_16567;
wire n_12952;
wire n_19096;
wire n_2045;
wire n_14795;
wire n_3687;
wire n_2216;
wire n_19318;
wire n_3621;
wire n_19886;
wire n_16425;
wire n_16769;
wire n_8217;
wire n_12004;
wire n_6962;
wire n_10603;
wire n_12830;
wire n_8858;
wire n_7246;
wire n_10255;
wire n_20172;
wire n_20420;
wire n_2719;
wire n_11490;
wire n_8689;
wire n_10113;
wire n_15086;
wire n_680;
wire n_3339;
wire n_6853;
wire n_10188;
wire n_10686;
wire n_9841;
wire n_19916;
wire n_8743;
wire n_7087;
wire n_8753;
wire n_6191;
wire n_4741;
wire n_16838;
wire n_10974;
wire n_11067;
wire n_8627;
wire n_20294;
wire n_13659;
wire n_12034;
wire n_16586;
wire n_1399;
wire n_16056;
wire n_13303;
wire n_6894;
wire n_13346;
wire n_13702;
wire n_9179;
wire n_2358;
wire n_15894;
wire n_8752;
wire n_2186;
wire n_18237;
wire n_3034;
wire n_4408;
wire n_18367;
wire n_10937;
wire n_643;
wire n_12134;
wire n_400;
wire n_12449;
wire n_2814;
wire n_16399;
wire n_789;
wire n_327;
wire n_6284;
wire n_10167;
wire n_12524;
wire n_18113;
wire n_6883;
wire n_12963;
wire n_10428;
wire n_16860;
wire n_17869;
wire n_20140;
wire n_19199;
wire n_18682;
wire n_12366;
wire n_747;
wire n_14951;
wire n_11068;
wire n_11035;
wire n_5495;
wire n_535;
wire n_19148;
wire n_12729;
wire n_13292;
wire n_12198;
wire n_9420;
wire n_3851;
wire n_16995;
wire n_14336;
wire n_7825;
wire n_10079;
wire n_7212;
wire n_19436;
wire n_6966;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_6035;
wire n_1652;
wire n_15435;
wire n_8634;
wire n_9531;
wire n_12605;
wire n_20202;
wire n_1258;
wire n_2438;
wire n_6253;
wire n_2914;
wire n_12828;
wire n_10258;
wire n_5786;
wire n_14960;
wire n_19109;
wire n_8532;
wire n_12661;
wire n_10588;
wire n_8991;
wire n_8065;
wire n_3100;
wire n_11140;
wire n_3573;
wire n_17882;
wire n_17677;
wire n_8518;
wire n_19845;
wire n_197;
wire n_18226;
wire n_13017;
wire n_1083;
wire n_16884;
wire n_15199;
wire n_18153;
wire n_1721;
wire n_9812;
wire n_1737;
wire n_15419;
wire n_752;
wire n_7361;
wire n_9949;
wire n_20200;
wire n_1028;
wire n_14889;
wire n_7228;
wire n_9576;
wire n_5872;
wire n_1973;
wire n_3181;
wire n_6338;
wire n_15267;
wire n_19366;
wire n_1500;
wire n_3699;
wire n_854;
wire n_4913;
wire n_6266;
wire n_14796;
wire n_2242;
wire n_19125;
wire n_11364;
wire n_12790;
wire n_4266;
wire n_8632;
wire n_2466;
wire n_19069;
wire n_17397;
wire n_19952;
wire n_5873;
wire n_7018;
wire n_7975;
wire n_10009;
wire n_9279;
wire n_11902;
wire n_924;
wire n_16782;
wire n_11993;
wire n_2318;
wire n_10443;
wire n_3170;
wire n_17317;
wire n_12813;
wire n_13534;
wire n_3304;
wire n_4968;
wire n_10384;
wire n_5085;
wire n_5736;
wire n_2433;
wire n_829;
wire n_7978;
wire n_10293;
wire n_17422;
wire n_20036;
wire n_12312;
wire n_10074;
wire n_13097;
wire n_17850;
wire n_15786;
wire n_4208;
wire n_9632;
wire n_20542;
wire n_12256;
wire n_11812;
wire n_9711;
wire n_9431;
wire n_4779;
wire n_14650;
wire n_18068;
wire n_481;
wire n_14610;
wire n_997;
wire n_11505;
wire n_4437;
wire n_7316;
wire n_17938;
wire n_1306;
wire n_3264;
wire n_18955;
wire n_7103;
wire n_14601;
wire n_436;
wire n_11363;
wire n_15794;
wire n_20164;
wire n_17066;
wire n_2426;
wire n_2478;
wire n_14645;
wire n_1133;
wire n_4642;
wire n_11151;
wire n_15825;
wire n_10716;
wire n_10664;
wire n_2578;
wire n_19819;
wire n_20392;
wire n_3709;
wire n_11434;
wire n_3738;
wire n_6873;
wire n_4186;
wire n_8494;
wire n_20056;
wire n_5812;
wire n_12468;
wire n_9429;
wire n_8544;
wire n_19536;
wire n_4998;
wire n_10749;
wire n_3330;
wire n_8788;
wire n_10992;
wire n_19380;
wire n_1629;
wire n_10160;
wire n_10560;
wire n_7404;
wire n_12857;
wire n_13171;
wire n_18615;
wire n_1260;
wire n_309;
wire n_9854;
wire n_14854;
wire n_812;
wire n_15266;
wire n_1006;
wire n_7271;
wire n_9713;
wire n_16501;
wire n_257;
wire n_19264;
wire n_1311;
wire n_10300;
wire n_9588;
wire n_14218;
wire n_15107;
wire n_6842;
wire n_13876;
wire n_4803;
wire n_18935;
wire n_6030;
wire n_1242;
wire n_2086;
wire n_14487;
wire n_9127;
wire n_5996;
wire n_20019;
wire n_16767;
wire n_9869;
wire n_315;
wire n_14449;
wire n_17094;
wire n_12885;
wire n_2579;
wire n_15539;
wire n_2105;
wire n_9715;
wire n_17112;
wire n_8618;
wire n_18916;
wire n_3387;
wire n_12108;
wire n_7535;
wire n_20469;
wire n_11531;
wire n_19450;
wire n_9407;
wire n_2912;
wire n_14476;
wire n_3409;
wire n_15244;
wire n_2320;
wire n_19574;
wire n_11824;
wire n_1259;
wire n_20201;
wire n_6957;
wire n_9361;
wire n_13976;
wire n_16578;
wire n_18949;
wire n_13579;
wire n_11566;
wire n_17452;
wire n_16650;
wire n_14639;
wire n_8990;
wire n_17067;
wire n_6444;
wire n_19170;
wire n_226;
wire n_7944;
wire n_19235;
wire n_11374;
wire n_8647;
wire n_15857;
wire n_2003;
wire n_7016;
wire n_10782;
wire n_13557;
wire n_3301;
wire n_20162;
wire n_16709;
wire n_6379;
wire n_15589;
wire n_17491;
wire n_2324;
wire n_17757;
wire n_12754;
wire n_245;
wire n_13583;
wire n_2977;
wire n_1739;
wire n_5840;
wire n_17333;
wire n_19043;
wire n_2847;
wire n_17749;
wire n_16658;
wire n_4050;
wire n_13455;
wire n_883;
wire n_19136;
wire n_6232;
wire n_9132;
wire n_1032;
wire n_20339;
wire n_10861;
wire n_17035;
wire n_8879;
wire n_1099;
wire n_19639;
wire n_11203;
wire n_16157;
wire n_11159;
wire n_8052;
wire n_2211;
wire n_6362;
wire n_11956;
wire n_11975;
wire n_12121;
wire n_9332;
wire n_17097;
wire n_369;
wire n_16765;
wire n_11030;
wire n_4179;
wire n_1285;
wire n_6326;
wire n_10073;
wire n_14619;
wire n_1590;
wire n_5072;
wire n_7241;
wire n_10419;
wire n_7172;
wire n_3106;
wire n_15427;
wire n_17364;
wire n_10333;
wire n_12430;
wire n_18330;
wire n_7235;
wire n_6239;
wire n_2340;
wire n_13407;
wire n_5896;
wire n_13676;
wire n_18391;
wire n_16694;
wire n_12557;
wire n_13788;
wire n_6974;
wire n_16537;
wire n_18227;
wire n_18666;
wire n_8939;
wire n_13584;
wire n_428;
wire n_15471;
wire n_12139;
wire n_9030;
wire n_7657;
wire n_822;
wire n_20075;
wire n_2791;
wire n_19433;
wire n_9665;
wire n_5044;
wire n_5134;
wire n_7096;
wire n_3063;
wire n_13327;
wire n_1550;
wire n_19098;
wire n_11197;
wire n_491;
wire n_7442;
wire n_1591;
wire n_3632;
wire n_10093;
wire n_20351;
wire n_15428;
wire n_15014;
wire n_1344;
wire n_6174;
wire n_2730;
wire n_7999;
wire n_10675;
wire n_6087;
wire n_16311;
wire n_538;
wire n_4164;
wire n_10107;
wire n_3225;
wire n_15536;
wire n_20061;
wire n_13224;
wire n_11469;
wire n_5022;
wire n_14046;
wire n_7041;
wire n_10742;
wire n_10829;
wire n_19115;
wire n_12389;
wire n_9309;
wire n_19632;
wire n_10620;
wire n_13971;
wire n_16750;
wire n_7672;
wire n_2551;
wire n_5047;
wire n_7318;
wire n_20368;
wire n_19325;
wire n_12995;
wire n_18261;
wire n_14406;
wire n_13209;
wire n_11883;
wire n_14959;
wire n_19979;
wire n_3269;
wire n_15387;
wire n_11901;
wire n_6352;
wire n_15973;
wire n_8542;
wire n_19747;
wire n_10859;
wire n_18446;
wire n_8576;
wire n_14807;
wire n_8038;
wire n_11572;
wire n_5141;
wire n_3603;
wire n_14493;
wire n_18306;
wire n_13113;
wire n_13387;
wire n_8716;
wire n_3822;
wire n_5535;
wire n_19411;
wire n_3812;
wire n_16807;
wire n_18538;
wire n_2696;
wire n_17576;
wire n_4080;
wire n_6002;
wire n_541;
wire n_18665;
wire n_15538;
wire n_2073;
wire n_2273;
wire n_4941;
wire n_5506;
wire n_11399;
wire n_17578;
wire n_8768;
wire n_10884;
wire n_1162;
wire n_15870;
wire n_12035;
wire n_13006;
wire n_12791;
wire n_7600;
wire n_14742;
wire n_2831;
wire n_4158;
wire n_6644;
wire n_17878;
wire n_4795;
wire n_19528;
wire n_12810;
wire n_16930;
wire n_3824;
wire n_13947;
wire n_11322;
wire n_17562;
wire n_4544;
wire n_5841;
wire n_12241;
wire n_9343;
wire n_15895;
wire n_16554;
wire n_17779;
wire n_5108;
wire n_7347;
wire n_11057;
wire n_2355;
wire n_10969;
wire n_14474;
wire n_7383;
wire n_2751;
wire n_6805;
wire n_8863;
wire n_18501;
wire n_7759;
wire n_11551;
wire n_18049;
wire n_7479;
wire n_2866;
wire n_10598;
wire n_8947;
wire n_15494;
wire n_10717;
wire n_11118;
wire n_18579;
wire n_3649;
wire n_2821;
wire n_6067;
wire n_12674;
wire n_17727;
wire n_17839;
wire n_8510;
wire n_11410;
wire n_12230;
wire n_19282;
wire n_1563;
wire n_9942;
wire n_11712;
wire n_9703;
wire n_17122;
wire n_1359;
wire n_5367;
wire n_16778;
wire n_3794;
wire n_12220;
wire n_6868;
wire n_1335;
wire n_5970;
wire n_16133;
wire n_12283;
wire n_7174;
wire n_9421;
wire n_5202;
wire n_19055;
wire n_13383;
wire n_18787;
wire n_17079;
wire n_8021;
wire n_3346;
wire n_15124;
wire n_7803;
wire n_12595;
wire n_11429;
wire n_15802;
wire n_15163;
wire n_13983;
wire n_9416;
wire n_6225;
wire n_5502;
wire n_3428;
wire n_4552;
wire n_6218;
wire n_17489;
wire n_9929;
wire n_12920;
wire n_13317;
wire n_2519;
wire n_9953;
wire n_1063;
wire n_6648;
wire n_15578;
wire n_10955;
wire n_7927;
wire n_11011;
wire n_9998;
wire n_11795;
wire n_5521;
wire n_4837;
wire n_9850;
wire n_12141;
wire n_20553;
wire n_9346;
wire n_7920;
wire n_437;
wire n_12774;
wire n_4169;
wire n_14687;
wire n_20283;
wire n_11904;
wire n_8480;
wire n_697;
wire n_17399;
wire n_388;
wire n_7025;
wire n_15886;
wire n_17022;
wire n_15856;
wire n_1757;
wire n_8484;
wire n_9472;
wire n_14304;
wire n_14357;
wire n_13044;
wire n_13228;
wire n_13518;
wire n_4070;
wire n_19763;
wire n_3885;
wire n_1369;
wire n_14008;
wire n_17069;
wire n_12746;
wire n_4031;
wire n_16162;
wire n_10970;
wire n_16285;
wire n_14927;
wire n_13881;
wire n_3209;
wire n_17205;
wire n_5547;
wire n_13747;
wire n_1391;
wire n_12532;
wire n_10238;
wire n_8931;
wire n_5596;
wire n_4653;
wire n_4435;
wire n_8334;
wire n_4019;
wire n_1071;
wire n_11681;
wire n_10890;
wire n_11202;
wire n_19513;
wire n_10552;
wire n_5815;
wire n_15254;
wire n_6595;
wire n_8539;
wire n_10205;
wire n_16947;
wire n_15747;
wire n_3727;
wire n_13899;
wire n_6306;
wire n_19386;
wire n_1714;
wire n_16235;
wire n_11663;
wire n_542;
wire n_11331;
wire n_305;
wire n_19472;
wire n_9528;
wire n_14348;
wire n_12201;
wire n_7583;
wire n_14086;
wire n_12499;
wire n_19334;
wire n_19173;
wire n_12448;
wire n_10610;
wire n_11187;
wire n_12761;
wire n_16455;
wire n_15004;
wire n_16625;
wire n_16025;
wire n_5520;
wire n_2638;
wire n_14552;
wire n_7353;
wire n_9490;
wire n_19767;
wire n_5669;
wire n_14575;
wire n_9574;
wire n_9024;
wire n_11694;
wire n_5772;
wire n_7571;
wire n_145;
wire n_4775;
wire n_16249;
wire n_16435;
wire n_4674;
wire n_16723;
wire n_11446;
wire n_10910;
wire n_294;
wire n_8242;
wire n_20132;
wire n_11540;
wire n_13248;
wire n_17296;
wire n_19237;
wire n_9819;
wire n_15338;
wire n_8184;
wire n_425;
wire n_20254;
wire n_6525;
wire n_4286;
wire n_13119;
wire n_2958;
wire n_12642;
wire n_3731;
wire n_1822;
wire n_12484;
wire n_6128;
wire n_13549;
wire n_2489;
wire n_17361;
wire n_16080;
wire n_4525;
wire n_9992;
wire n_15180;
wire n_15692;
wire n_19976;
wire n_5712;
wire n_12669;
wire n_14296;
wire n_6702;
wire n_19490;
wire n_11179;
wire n_17074;
wire n_2520;
wire n_446;
wire n_7749;
wire n_10078;
wire n_11321;
wire n_14313;
wire n_9500;
wire n_18496;
wire n_8705;
wire n_19107;
wire n_11779;
wire n_7508;
wire n_2501;
wire n_3203;
wire n_5694;
wire n_14211;
wire n_7574;
wire n_4306;
wire n_13516;
wire n_14273;
wire n_20063;
wire n_12462;
wire n_4453;
wire n_16462;
wire n_18648;
wire n_4005;
wire n_6169;
wire n_18775;
wire n_15230;
wire n_3546;
wire n_3661;
wire n_12735;
wire n_10709;
wire n_12646;
wire n_19849;
wire n_15875;
wire n_7352;
wire n_10244;
wire n_755;
wire n_20128;
wire n_18512;
wire n_12999;
wire n_12682;
wire n_14802;
wire n_6848;
wire n_17415;
wire n_3509;
wire n_10043;
wire n_14834;
wire n_5919;
wire n_8159;
wire n_14346;
wire n_16955;
wire n_7439;
wire n_17653;
wire n_2504;
wire n_14506;
wire n_2623;
wire n_18822;
wire n_16018;
wire n_14615;
wire n_15222;
wire n_6850;
wire n_18991;
wire n_15285;
wire n_5005;
wire n_13294;
wire n_6098;
wire n_20446;
wire n_7112;
wire n_11307;
wire n_19021;
wire n_17860;
wire n_18274;
wire n_9545;
wire n_596;
wire n_9629;
wire n_9603;
wire n_18003;
wire n_12719;
wire n_10342;
wire n_15361;
wire n_3322;
wire n_19037;
wire n_16244;
wire n_17862;
wire n_4654;
wire n_13438;
wire n_3640;
wire n_1159;
wire n_995;
wire n_15850;
wire n_9930;
wire n_14371;
wire n_12925;
wire n_5775;
wire n_14988;
wire n_9659;
wire n_3226;
wire n_2780;
wire n_16293;
wire n_9897;
wire n_9241;
wire n_14590;
wire n_14603;
wire n_8185;
wire n_11466;
wire n_5061;
wire n_15265;
wire n_15040;
wire n_6775;
wire n_9291;
wire n_4063;
wire n_11982;
wire n_2601;
wire n_773;
wire n_11873;
wire n_15821;
wire n_920;
wire n_10185;
wire n_11182;
wire n_20037;
wire n_3212;
wire n_16250;
wire n_15768;
wire n_8220;
wire n_18807;
wire n_4721;
wire n_14145;
wire n_11991;
wire n_848;
wire n_12875;
wire n_15064;
wire n_11807;
wire n_9262;
wire n_7426;
wire n_4247;
wire n_13918;
wire n_13775;
wire n_9851;
wire n_11799;
wire n_8009;
wire n_7852;
wire n_1881;
wire n_10983;
wire n_9987;
wire n_7984;
wire n_18307;
wire n_2720;
wire n_19860;
wire n_18110;
wire n_14973;
wire n_16751;
wire n_7220;
wire n_18015;
wire n_20300;
wire n_1323;
wire n_2627;
wire n_18242;
wire n_6550;
wire n_3004;
wire n_8841;
wire n_12196;
wire n_5483;
wire n_3625;
wire n_15136;
wire n_1764;
wire n_10354;
wire n_7465;
wire n_13177;
wire n_4546;
wire n_12724;
wire n_14958;
wire n_6672;
wire n_16744;
wire n_17876;
wire n_1551;
wire n_15992;
wire n_7738;
wire n_17406;
wire n_19079;
wire n_8395;
wire n_6634;
wire n_14758;
wire n_18392;
wire n_8961;
wire n_10849;
wire n_7462;
wire n_4635;
wire n_16802;
wire n_17909;
wire n_18439;
wire n_5735;
wire n_19022;
wire n_13311;
wire n_19700;
wire n_2278;
wire n_20587;
wire n_16020;
wire n_11513;
wire n_7464;
wire n_8937;
wire n_7115;
wire n_2924;
wire n_12087;
wire n_13675;
wire n_15022;
wire n_18693;
wire n_3595;
wire n_6104;
wire n_10537;
wire n_421;
wire n_6082;
wire n_18305;
wire n_1270;
wire n_10426;
wire n_1852;
wire n_9167;
wire n_12082;
wire n_9655;
wire n_20448;
wire n_11436;
wire n_11729;
wire n_3230;
wire n_19276;
wire n_1499;
wire n_12989;
wire n_504;
wire n_5877;
wire n_8845;
wire n_15198;
wire n_6018;
wire n_17902;
wire n_13620;
wire n_1503;
wire n_7702;
wire n_6676;
wire n_2819;
wire n_9976;
wire n_2423;
wire n_8042;
wire n_17144;
wire n_12464;
wire n_9560;
wire n_18362;
wire n_18886;
wire n_20264;
wire n_1182;
wire n_15007;
wire n_15197;
wire n_167;
wire n_8519;
wire n_5582;
wire n_5886;
wire n_1216;
wire n_6032;
wire n_18982;
wire n_9319;
wire n_5446;
wire n_3010;
wire n_12450;
wire n_5224;
wire n_19776;
wire n_14648;
wire n_11767;
wire n_2486;
wire n_3560;
wire n_10985;
wire n_9401;
wire n_11586;
wire n_12149;
wire n_12002;
wire n_12836;
wire n_19506;
wire n_17084;
wire n_13548;
wire n_15710;
wire n_2232;
wire n_11195;
wire n_4038;
wire n_16240;
wire n_2790;
wire n_9747;
wire n_5414;
wire n_14526;
wire n_13487;
wire n_17190;
wire n_3784;
wire n_17973;
wire n_220;
wire n_8586;
wire n_9058;
wire n_18707;
wire n_1472;
wire n_18547;
wire n_16700;
wire n_5454;
wire n_800;
wire n_10780;
wire n_17940;
wire n_8756;
wire n_1840;
wire n_4434;
wire n_13406;
wire n_16371;
wire n_7923;
wire n_14040;
wire n_8602;
wire n_14054;
wire n_1346;
wire n_13469;
wire n_10411;
wire n_13249;
wire n_12984;
wire n_18840;
wire n_13587;
wire n_5913;
wire n_10090;
wire n_14872;
wire n_1102;
wire n_8112;
wire n_18959;
wire n_258;
wire n_11567;
wire n_2766;
wire n_19428;
wire n_9292;
wire n_18771;
wire n_12197;
wire n_356;
wire n_17753;
wire n_19134;
wire n_4833;
wire n_11580;
wire n_13326;
wire n_6474;
wire n_13082;
wire n_5230;
wire n_5944;
wire n_6226;
wire n_152;
wire n_18518;
wire n_10856;
wire n_12403;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_2782;
wire n_9584;
wire n_13692;
wire n_8194;
wire n_8055;
wire n_8579;
wire n_10914;
wire n_8360;
wire n_4279;
wire n_20340;
wire n_6425;
wire n_1456;
wire n_6493;
wire n_14382;
wire n_13396;
wire n_10071;
wire n_8755;
wire n_2099;
wire n_11565;
wire n_3388;
wire n_14911;
wire n_15405;
wire n_5810;
wire n_4461;
wire n_3245;
wire n_4007;
wire n_15643;
wire n_15420;
wire n_13052;
wire n_11013;
wire n_5991;
wire n_1676;
wire n_20486;
wire n_1319;
wire n_16634;
wire n_16762;
wire n_10035;
wire n_5702;
wire n_18094;
wire n_20247;
wire n_18673;
wire n_18980;
wire n_14962;
wire n_1633;
wire n_17435;
wire n_8108;
wire n_2820;
wire n_17065;
wire n_12068;
wire n_5250;
wire n_3074;
wire n_17285;
wire n_10041;
wire n_15499;
wire n_5590;
wire n_14514;
wire n_17612;
wire n_8498;
wire n_14256;
wire n_17073;
wire n_16773;
wire n_2727;
wire n_2533;
wire n_5349;
wire n_19320;
wire n_2759;
wire n_2361;
wire n_2266;
wire n_14082;
wire n_20160;
wire n_7280;
wire n_5833;
wire n_7886;
wire n_15728;
wire n_6884;
wire n_7664;
wire n_18292;
wire n_7012;
wire n_299;
wire n_1248;
wire n_17354;
wire n_12486;
wire n_902;
wire n_2189;
wire n_7376;
wire n_5816;
wire n_15347;
wire n_10137;
wire n_12084;
wire n_16517;
wire n_706;
wire n_1794;
wire n_20032;
wire n_1236;
wire n_11863;
wire n_17868;
wire n_17033;
wire n_17234;
wire n_430;
wire n_16174;
wire n_18059;
wire n_19015;
wire n_10794;
wire n_14703;
wire n_13533;
wire n_6274;
wire n_16283;
wire n_12109;
wire n_8838;
wire n_9562;
wire n_3097;
wire n_7007;
wire n_2975;
wire n_16088;
wire n_2856;
wire n_4498;
wire n_12320;
wire n_19245;
wire n_9759;
wire n_6992;
wire n_15226;
wire n_19742;
wire n_646;
wire n_528;
wire n_19859;
wire n_10206;
wire n_1329;
wire n_17736;
wire n_6322;
wire n_5167;
wire n_15425;
wire n_5661;
wire n_16878;
wire n_3589;
wire n_262;
wire n_897;
wire n_7616;
wire n_1800;
wire n_18294;
wire n_9733;
wire n_12282;
wire n_8189;
wire n_6498;
wire n_8481;
wire n_13011;
wire n_9981;
wire n_18514;
wire n_5558;
wire n_5687;
wire n_16513;
wire n_6378;
wire n_14495;
wire n_1759;
wire n_16879;
wire n_12269;
wire n_853;
wire n_13486;
wire n_11463;
wire n_3585;
wire n_17541;
wire n_5954;
wire n_5025;
wire n_933;
wire n_17394;
wire n_7587;
wire n_3135;
wire n_17496;
wire n_6930;
wire n_17472;
wire n_19121;
wire n_12802;
wire n_11569;
wire n_10064;
wire n_7197;
wire n_9676;
wire n_7393;
wire n_11332;
wire n_13629;
wire n_13207;
wire n_310;
wire n_5766;
wire n_18025;
wire n_7358;
wire n_2796;
wire n_9950;
wire n_18088;
wire n_13589;
wire n_15730;
wire n_18089;
wire n_4534;
wire n_17967;
wire n_19731;
wire n_6929;
wire n_16706;
wire n_11309;
wire n_955;
wire n_8045;
wire n_16032;
wire n_19740;
wire n_19741;
wire n_18910;
wire n_2969;
wire n_2395;
wire n_16959;
wire n_8209;
wire n_14477;
wire n_9213;
wire n_7291;
wire n_14522;
wire n_669;
wire n_16971;
wire n_2290;
wire n_19998;
wire n_20526;
wire n_2005;
wire n_13561;
wire n_14720;
wire n_7437;
wire n_16873;
wire n_1408;
wire n_7618;
wire n_8575;
wire n_5733;
wire n_6620;
wire n_6597;
wire n_11105;
wire n_13698;
wire n_13894;
wire n_452;
wire n_6586;
wire n_10474;
wire n_12689;
wire n_18939;
wire n_8789;
wire n_7953;
wire n_19775;
wire n_13540;
wire n_6428;
wire n_5328;
wire n_14642;
wire n_12042;
wire n_14827;
wire n_15481;
wire n_5657;
wire n_174;
wire n_1173;
wire n_13465;
wire n_11130;
wire n_16149;
wire n_11664;
wire n_18705;
wire n_17430;
wire n_15388;
wire n_19242;
wire n_10652;
wire n_13733;
wire n_13098;
wire n_3334;
wire n_20029;
wire n_9388;
wire n_12654;
wire n_4985;
wire n_10869;
wire n_3823;
wire n_18708;
wire n_19112;
wire n_11783;
wire n_2255;
wire n_17837;
wire n_4678;
wire n_2649;
wire n_9911;
wire n_19603;
wire n_5579;
wire n_414;
wire n_16317;
wire n_1922;
wire n_15187;
wire n_10346;
wire n_12419;
wire n_13763;
wire n_17897;
wire n_4363;
wire n_10473;
wire n_15712;
wire n_5107;
wire n_16985;
wire n_5095;
wire n_19941;
wire n_8493;
wire n_10957;
wire n_13517;
wire n_20049;
wire n_11188;
wire n_3404;
wire n_10442;
wire n_1509;
wire n_3290;
wire n_13973;
wire n_7150;
wire n_8252;
wire n_11774;
wire n_3671;
wire n_7015;
wire n_2015;
wire n_3982;
wire n_13206;
wire n_7249;
wire n_1161;
wire n_15939;
wire n_3840;
wire n_3461;
wire n_7985;
wire n_13637;
wire n_3513;
wire n_16705;
wire n_18163;
wire n_8893;
wire n_6372;
wire n_3995;
wire n_4076;
wire n_15904;
wire n_592;
wire n_12768;
wire n_1156;
wire n_18369;
wire n_16047;
wire n_3508;
wire n_10165;
wire n_8156;
wire n_868;
wire n_19674;
wire n_14923;
wire n_13031;
wire n_19029;
wire n_19316;
wire n_17912;
wire n_13155;
wire n_469;
wire n_1218;
wire n_13410;
wire n_19581;
wire n_7814;
wire n_8660;
wire n_985;
wire n_2440;
wire n_13124;
wire n_6054;
wire n_11095;
wire n_19546;
wire n_561;
wire n_8606;
wire n_9663;
wire n_16584;
wire n_18340;
wire n_1244;
wire n_9743;
wire n_19048;
wire n_11584;
wire n_2285;
wire n_5280;
wire n_14169;
wire n_7700;
wire n_4451;
wire n_10158;
wire n_10582;
wire n_16151;
wire n_10427;
wire n_11816;
wire n_18808;
wire n_3563;
wire n_16420;
wire n_201;
wire n_11693;
wire n_3495;
wire n_15429;
wire n_9248;
wire n_6138;
wire n_5369;
wire n_10835;
wire n_975;
wire n_11411;
wire n_5576;
wire n_19681;
wire n_13823;
wire n_11386;
wire n_20159;
wire n_11604;
wire n_13323;
wire n_3359;
wire n_12164;
wire n_16919;
wire n_12824;
wire n_13434;
wire n_16680;
wire n_16938;
wire n_3187;
wire n_10844;
wire n_17793;
wire n_14153;
wire n_6802;
wire n_10654;
wire n_6909;
wire n_13445;
wire n_17177;
wire n_19074;
wire n_18182;
wire n_4336;
wire n_15760;
wire n_16712;
wire n_14746;
wire n_11097;
wire n_4981;
wire n_14606;
wire n_12052;
wire n_9746;
wire n_8073;
wire n_1166;
wire n_5440;
wire n_2891;
wire n_8821;
wire n_19922;
wire n_9440;
wire n_3955;
wire n_17253;
wire n_2280;
wire n_20457;
wire n_203;
wire n_20212;
wire n_20142;
wire n_1868;
wire n_17264;
wire n_2079;
wire n_15475;
wire n_8663;
wire n_20114;
wire n_2185;
wire n_5861;
wire n_1836;
wire n_10553;
wire n_19770;
wire n_8309;
wire n_1486;
wire n_5258;
wire n_8945;
wire n_15121;
wire n_10988;
wire n_19209;
wire n_784;
wire n_20175;
wire n_6112;
wire n_16192;
wire n_18030;
wire n_9041;
wire n_862;
wire n_8166;
wire n_2098;
wire n_5606;
wire n_1935;
wire n_10108;
wire n_13865;
wire n_5920;
wire n_10307;
wire n_1449;
wire n_361;
wire n_8215;
wire n_19538;
wire n_17497;
wire n_6180;
wire n_8809;
wire n_12382;
wire n_5527;
wire n_6476;
wire n_14428;
wire n_6566;
wire n_5172;
wire n_11173;
wire n_16218;
wire n_6872;
wire n_13998;
wire n_5254;
wire n_17825;
wire n_10587;
wire n_8713;
wire n_15450;
wire n_7111;
wire n_13522;
wire n_7967;
wire n_15609;
wire n_16423;
wire n_9002;
wire n_14670;
wire n_9130;
wire n_19016;
wire n_7180;
wire n_13530;
wire n_8604;
wire n_16362;
wire n_7263;
wire n_1342;
wire n_4829;
wire n_5393;
wire n_677;
wire n_14318;
wire n_4686;
wire n_17673;
wire n_17004;
wire n_11802;
wire n_20215;
wire n_3706;
wire n_8005;
wire n_2179;
wire n_13942;
wire n_18230;
wire n_1547;
wire n_12570;
wire n_11905;
wire n_19326;
wire n_893;
wire n_20007;
wire n_3801;
wire n_5267;
wire n_10202;
wire n_3564;
wire n_15295;
wire n_9104;
wire n_17050;
wire n_17408;
wire n_15445;
wire n_8272;
wire n_13997;
wire n_14402;
wire n_14882;
wire n_11051;
wire n_11214;
wire n_2628;
wire n_7000;
wire n_7398;
wire n_18335;
wire n_1078;
wire n_14232;
wire n_12882;
wire n_19300;
wire n_18057;
wire n_12617;
wire n_8236;
wire n_13137;
wire n_3345;
wire n_19612;
wire n_15933;
wire n_17188;
wire n_6325;
wire n_4724;
wire n_9840;
wire n_10348;
wire n_12495;
wire n_9581;
wire n_8070;
wire n_4696;
wire n_18468;
wire n_16786;
wire n_7802;
wire n_17118;
wire n_3877;
wire n_15353;
wire n_19623;
wire n_1455;
wire n_15993;
wire n_6629;
wire n_5279;
wire n_5894;
wire n_17699;
wire n_19605;
wire n_8175;
wire n_567;
wire n_8953;
wire n_17546;
wire n_17279;
wire n_19111;
wire n_4814;
wire n_10373;
wire n_3979;
wire n_3077;
wire n_9525;
wire n_10816;
wire n_9725;
wire n_19511;
wire n_6914;
wire n_14121;
wire n_10381;
wire n_713;
wire n_1400;
wire n_20163;
wire n_10947;
wire n_16984;
wire n_6015;
wire n_11261;
wire n_16012;
wire n_1560;
wire n_734;
wire n_13929;
wire n_17739;
wire n_10767;
wire n_19684;
wire n_14646;
wire n_14095;
wire n_15069;
wire n_14520;
wire n_14780;
wire n_4950;
wire n_19828;
wire n_19966;
wire n_4729;
wire n_4268;
wire n_11447;
wire n_12652;
wire n_15507;
wire n_8142;
wire n_11627;
wire n_6404;
wire n_12209;
wire n_5680;
wire n_6674;
wire n_17883;
wire n_13606;
wire n_11659;
wire n_13501;
wire n_4102;
wire n_9106;
wire n_4662;
wire n_8869;
wire n_3959;
wire n_2268;
wire n_8381;
wire n_1367;
wire n_5504;
wire n_1336;
wire n_17149;
wire n_9520;
wire n_2080;
wire n_14931;
wire n_18774;
wire n_7770;
wire n_6968;
wire n_16268;
wire n_12371;
wire n_4507;
wire n_20027;
wire n_11497;
wire n_14900;
wire n_792;
wire n_15846;
wire n_13454;
wire n_5306;
wire n_16662;
wire n_9042;
wire n_17329;
wire n_3488;
wire n_8987;
wire n_11805;
wire n_1910;
wire n_14935;
wire n_2998;
wire n_237;
wire n_6282;
wire n_12770;
wire n_4294;
wire n_19551;
wire n_11635;
wire n_15434;
wire n_16530;
wire n_12951;
wire n_9453;
wire n_8118;
wire n_12393;
wire n_16442;
wire n_9718;
wire n_10281;
wire n_3927;
wire n_3888;
wire n_764;
wire n_12831;
wire n_2895;
wire n_6431;
wire n_733;
wire n_19620;
wire n_19839;
wire n_15767;
wire n_1290;
wire n_12427;
wire n_1354;
wire n_7533;
wire n_7221;
wire n_16026;
wire n_15159;
wire n_1701;
wire n_10656;
wire n_6575;
wire n_6055;
wire n_8246;
wire n_8952;
wire n_3875;
wire n_5609;
wire n_4717;
wire n_871;
wire n_15154;
wire n_9680;
wire n_12172;
wire n_5658;
wire n_4731;
wire n_12923;
wire n_12147;
wire n_3052;
wire n_19624;
wire n_20204;
wire n_13227;
wire n_19683;
wire n_8848;
wire n_12825;
wire n_5667;
wire n_8259;
wire n_2624;
wire n_5865;
wire n_15182;
wire n_8349;
wire n_6836;
wire n_11998;
wire n_19900;
wire n_8776;
wire n_19391;
wire n_7753;
wire n_6771;
wire n_14732;
wire n_9947;
wire n_16659;
wire n_1750;
wire n_1462;
wire n_10138;
wire n_12117;
wire n_10375;
wire n_14535;
wire n_6795;
wire n_5314;
wire n_12960;
wire n_18972;
wire n_14094;
wire n_13033;
wire n_15703;
wire n_19353;
wire n_7648;
wire n_515;
wire n_4418;
wire n_12131;
wire n_12851;
wire n_19854;
wire n_7452;
wire n_5226;
wire n_9269;
wire n_10320;
wire n_514;
wire n_15518;
wire n_14217;
wire n_10903;
wire n_17596;
wire n_15574;
wire n_14062;
wire n_8453;
wire n_12740;
wire n_2393;
wire n_2921;
wire n_3237;
wire n_8949;
wire n_10831;
wire n_9131;
wire n_17580;
wire n_10517;
wire n_16889;
wire n_10323;
wire n_10842;
wire n_17620;
wire n_3542;
wire n_16465;
wire n_2763;
wire n_2762;
wire n_20519;
wire n_11146;
wire n_10883;
wire n_17785;
wire n_1296;
wire n_19249;
wire n_3073;
wire n_5343;
wire n_20493;
wire n_1294;
wire n_3696;
wire n_20106;
wire n_12278;
wire n_18918;
wire n_19018;
wire n_1779;
wire n_524;
wire n_17672;
wire n_4329;
wire n_18036;
wire n_5135;
wire n_17414;
wire n_10123;
wire n_10651;
wire n_4697;
wire n_3763;
wire n_17483;
wire n_17689;
wire n_18975;
wire n_14785;
wire n_8500;
wire n_17857;
wire n_2145;
wire n_4964;
wire n_12804;
wire n_20458;
wire n_12116;
wire n_17438;
wire n_1932;
wire n_13755;
wire n_1101;
wire n_10468;
wire n_4636;
wire n_14105;
wire n_14126;
wire n_8285;
wire n_8483;
wire n_4946;
wire n_4767;
wire n_4287;
wire n_19145;
wire n_17696;
wire n_1451;
wire n_639;
wire n_11370;
wire n_16731;
wire n_4576;
wire n_9020;
wire n_4615;
wire n_1018;
wire n_9895;
wire n_16452;
wire n_11585;
wire n_13140;
wire n_13962;
wire n_4389;
wire n_13753;
wire n_1376;
wire n_15365;
wire n_17141;
wire n_948;
wire n_12560;
wire n_19295;
wire n_18171;
wire n_977;
wire n_13610;
wire n_536;
wire n_8851;
wire n_13332;
wire n_15293;
wire n_19405;
wire n_6097;
wire n_19214;
wire n_19779;
wire n_7093;
wire n_4098;
wire n_5026;
wire n_4476;
wire n_432;
wire n_3700;
wire n_3104;
wire n_2239;
wire n_7840;
wire n_18797;
wire n_10024;
wire n_16386;
wire n_17101;
wire n_15695;
wire n_7080;
wire n_17984;
wire n_2191;
wire n_14156;
wire n_10711;
wire n_7624;
wire n_1426;
wire n_19915;
wire n_16185;
wire n_10818;
wire n_9186;
wire n_1529;
wire n_4634;
wire n_2069;
wire n_18851;
wire n_2362;
wire n_4096;
wire n_15178;
wire n_2698;
wire n_11951;
wire n_12222;
wire n_7003;
wire n_13604;
wire n_5427;
wire n_10788;
wire n_17163;
wire n_10563;
wire n_8810;
wire n_20427;
wire n_3631;
wire n_2772;
wire n_14518;
wire n_16310;
wire n_16477;
wire n_13397;
wire n_10178;
wire n_5052;
wire n_4541;
wire n_17731;
wire n_15360;
wire n_929;
wire n_4551;
wire n_2857;
wire n_13132;
wire n_6609;
wire n_10115;
wire n_17157;
wire n_5326;
wire n_16927;
wire n_12793;
wire n_11778;
wire n_1183;
wire n_2494;
wire n_12406;
wire n_998;
wire n_717;
wire n_1383;
wire n_7484;
wire n_16639;
wire n_6414;
wire n_1000;
wire n_9470;
wire n_3810;
wire n_552;
wire n_15516;
wire n_3006;
wire n_216;
wire n_13792;
wire n_5010;
wire n_1201;
wire n_4592;
wire n_18229;
wire n_9405;
wire n_1395;
wire n_6264;
wire n_2199;
wire n_17426;
wire n_13480;
wire n_1955;
wire n_20233;
wire n_19583;
wire n_312;
wire n_13571;
wire n_10984;
wire n_5104;
wire n_19723;
wire n_20249;
wire n_18742;
wire n_20255;
wire n_12001;
wire n_7883;
wire n_589;
wire n_1310;
wire n_13715;
wire n_3591;
wire n_16675;
wire n_2797;
wire n_7458;
wire n_4746;
wire n_15186;
wire n_16935;
wire n_18576;
wire n_13810;
wire n_14403;
wire n_7435;
wire n_6997;
wire n_10509;
wire n_5952;
wire n_3964;
wire n_19292;
wire n_13473;
wire n_18267;
wire n_5985;
wire n_556;
wire n_15963;
wire n_14353;
wire n_16589;
wire n_1602;
wire n_19213;
wire n_11742;
wire n_6891;
wire n_10031;
wire n_276;
wire n_19163;
wire n_12235;
wire n_5232;
wire n_7663;
wire n_12204;
wire n_10898;
wire n_5116;
wire n_14386;
wire n_18784;
wire n_16472;
wire n_17830;
wire n_12098;
wire n_4428;
wire n_1533;
wire n_7917;
wire n_12579;
wire n_2274;
wire n_9203;
wire n_15073;
wire n_7532;
wire n_9613;
wire n_5761;
wire n_13982;
wire n_19921;
wire n_18703;
wire n_12611;
wire n_13269;
wire n_7375;
wire n_13369;
wire n_7968;
wire n_6382;
wire n_317;
wire n_18542;
wire n_1679;
wire n_9141;
wire n_15867;
wire n_5760;
wire n_2146;
wire n_11027;
wire n_11852;
wire n_5472;
wire n_8377;
wire n_9913;
wire n_2575;
wire n_19911;
wire n_9286;
wire n_19646;
wire n_7921;
wire n_10044;
wire n_7728;
wire n_4410;
wire n_10819;
wire n_1179;
wire n_324;
wire n_14521;
wire n_20024;
wire n_9704;
wire n_19468;
wire n_19025;
wire n_9046;
wire n_16576;
wire n_6339;
wire n_8814;
wire n_8530;
wire n_9193;
wire n_16882;
wire n_20353;
wire n_7711;
wire n_16181;
wire n_15948;
wire n_8984;
wire n_17123;
wire n_3663;
wire n_3299;
wire n_9290;
wire n_351;
wire n_259;
wire n_14580;
wire n_5745;
wire n_1645;
wire n_14028;
wire n_19131;
wire n_14772;
wire n_956;
wire n_13827;
wire n_14542;
wire n_18632;
wire n_3845;
wire n_664;
wire n_1869;
wire n_7230;
wire n_17552;
wire n_7989;
wire n_9778;
wire n_20511;
wire n_18986;
wire n_2016;
wire n_20109;
wire n_5171;
wire n_18280;
wire n_15003;
wire n_13200;
wire n_1937;
wire n_16783;
wire n_12848;
wire n_18963;
wire n_341;
wire n_1744;
wire n_828;
wire n_10315;
wire n_18321;
wire n_607;
wire n_19104;
wire n_17187;
wire n_4028;
wire n_17031;
wire n_11455;
wire n_12368;
wire n_5255;
wire n_3756;
wire n_17240;
wire n_19795;
wire n_3406;
wire n_13193;
wire n_951;
wire n_19798;
wire n_952;
wire n_8462;
wire n_18953;
wire n_9380;
wire n_19881;
wire n_10062;
wire n_18235;
wire n_20115;
wire n_19476;
wire n_2375;
wire n_1934;
wire n_8429;
wire n_10514;
wire n_1434;
wire n_12785;
wire n_3981;
wire n_15312;
wire n_14155;
wire n_1275;
wire n_1510;
wire n_7620;
wire n_20034;
wire n_5783;
wire n_3120;
wire n_5821;
wire n_15818;
wire n_6079;
wire n_16481;
wire n_16430;
wire n_19313;
wire n_3864;
wire n_16715;
wire n_8492;
wire n_16565;
wire n_248;
wire n_2302;
wire n_8135;
wire n_16620;
wire n_8445;
wire n_1037;
wire n_6427;
wire n_3592;
wire n_468;
wire n_4230;
wire n_14978;
wire n_2637;
wire n_18353;
wire n_12639;
wire n_991;
wire n_8895;
wire n_3817;
wire n_7811;
wire n_340;
wire n_14649;
wire n_15940;
wire n_19955;
wire n_12175;
wire n_5003;
wire n_13536;
wire n_10512;
wire n_14714;
wire n_11384;
wire n_4827;
wire n_8273;
wire n_12353;
wire n_14129;
wire n_6065;
wire n_9761;
wire n_16962;
wire n_4610;
wire n_9087;
wire n_4472;
wire n_17832;
wire n_3081;
wire n_17316;
wire n_15333;
wire n_10434;
wire n_12869;
wire n_8312;
wire n_6781;
wire n_18585;
wire n_13830;
wire n_6133;
wire n_14184;
wire n_11889;
wire n_14183;
wire n_4990;
wire n_6127;
wire n_19172;
wire n_17751;
wire n_2498;
wire n_11362;
wire n_19256;
wire n_8078;
wire n_4515;
wire n_14200;
wire n_6006;
wire n_16558;
wire n_7926;
wire n_19118;
wire n_6598;
wire n_20359;
wire n_172;
wire n_15568;
wire n_12502;
wire n_2392;
wire n_4131;
wire n_16859;
wire n_1043;
wire n_18800;
wire n_16703;
wire n_2305;
wire n_19666;
wire n_13191;
wire n_10131;
wire n_15464;
wire n_17741;
wire n_6867;
wire n_12600;
wire n_14536;
wire n_16338;
wire n_6139;
wire n_12133;
wire n_19939;
wire n_7965;
wire n_12919;
wire n_3356;
wire n_10273;
wire n_11416;
wire n_3210;
wire n_937;
wire n_17485;
wire n_14321;
wire n_1682;
wire n_7474;
wire n_11169;
wire n_8650;
wire n_17843;
wire n_14654;
wire n_10503;
wire n_4905;
wire n_14664;
wire n_13215;
wire n_4601;
wire n_16834;
wire n_962;
wire n_10465;
wire n_16073;
wire n_10590;
wire n_19890;
wire n_3647;
wire n_13782;
wire n_15476;
wire n_8526;
wire n_1186;
wire n_13751;
wire n_19988;
wire n_17150;
wire n_14019;
wire n_19140;
wire n_19418;
wire n_20385;
wire n_6759;
wire n_10786;
wire n_3988;
wire n_19806;
wire n_7028;
wire n_9890;
wire n_11492;
wire n_19653;
wire n_394;
wire n_18904;
wire n_6535;
wire n_18801;
wire n_16644;
wire n_9817;
wire n_1524;
wire n_11160;
wire n_18899;
wire n_9782;
wire n_1920;
wire n_3292;
wire n_1225;
wire n_12319;
wire n_10805;
wire n_17214;
wire n_20356;
wire n_6643;
wire n_17982;
wire n_9471;
wire n_3712;
wire n_4608;
wire n_2506;
wire n_17012;
wire n_14896;
wire n_17440;
wire n_12930;
wire n_17181;
wire n_1567;
wire n_4037;
wire n_8351;
wire n_9069;
wire n_17371;
wire n_3562;
wire n_14030;
wire n_8603;
wire n_17274;
wire n_16660;
wire n_11343;
wire n_3007;
wire n_19143;
wire n_12575;
wire n_11451;
wire n_4571;
wire n_16853;
wire n_20050;
wire n_3698;
wire n_13384;
wire n_3355;
wire n_2114;
wire n_16048;
wire n_16262;
wire n_17127;
wire n_15422;
wire n_9003;
wire n_2154;
wire n_18874;
wire n_12418;
wire n_5290;
wire n_4185;
wire n_14837;
wire n_7312;
wire n_4219;
wire n_11269;
wire n_16849;
wire n_3985;
wire n_1447;
wire n_14103;
wire n_4774;
wire n_6689;
wire n_7632;
wire n_9172;
wire n_14653;
wire n_4232;
wire n_3000;
wire n_19464;
wire n_17275;
wire n_8980;
wire n_5571;
wire n_17573;
wire n_11311;
wire n_6698;
wire n_18553;
wire n_17345;
wire n_17770;
wire n_13242;
wire n_7707;
wire n_13282;
wire n_14436;
wire n_12113;
wire n_14599;
wire n_16087;
wire n_4736;
wire n_1725;
wire n_3743;
wire n_13352;
wire n_17648;
wire n_18116;
wire n_17853;
wire n_14812;
wire n_17871;
wire n_11293;
wire n_14728;
wire n_19184;
wire n_545;
wire n_2671;
wire n_6363;
wire n_2715;
wire n_8619;
wire n_3511;
wire n_19224;
wire n_18217;
wire n_18812;
wire n_15122;
wire n_10134;
wire n_11603;
wire n_1477;
wire n_7277;
wire n_11271;
wire n_14778;
wire n_15714;
wire n_17270;
wire n_12015;
wire n_8146;
wire n_13690;
wire n_2833;
wire n_11562;
wire n_10194;
wire n_17085;
wire n_8910;
wire n_1001;
wire n_6408;
wire n_6150;
wire n_10077;
wire n_4708;
wire n_13619;
wire n_4657;
wire n_18508;
wire n_12031;
wire n_1191;
wire n_9278;
wire n_855;
wire n_10889;
wire n_10010;
wire n_20472;
wire n_14996;
wire n_12126;
wire n_14543;
wire n_8550;
wire n_11094;
wire n_20046;
wire n_14747;
wire n_10599;
wire n_9667;
wire n_6401;
wire n_9739;
wire n_14358;
wire n_4536;
wire n_9480;
wire n_17886;
wire n_1976;
wire n_12195;
wire n_19369;
wire n_6679;
wire n_19294;
wire n_1824;
wire n_13289;
wire n_13182;
wire n_16265;
wire n_16466;
wire n_13324;
wire n_9541;
wire n_11286;
wire n_15215;
wire n_18947;
wire n_17748;
wire n_16379;
wire n_16728;
wire n_823;
wire n_1074;
wire n_7097;
wire n_8140;
wire n_15111;
wire n_1097;
wire n_781;
wire n_18563;
wire n_1810;
wire n_5915;
wire n_8527;
wire n_12899;
wire n_18917;
wire n_1583;
wire n_17621;
wire n_2295;
wire n_1643;
wire n_19570;
wire n_7909;
wire n_6303;
wire n_3652;
wire n_8935;
wire n_15759;
wire n_20556;
wire n_10734;
wire n_16441;
wire n_15383;
wire n_11560;
wire n_10395;
wire n_3617;
wire n_14966;
wire n_11435;
wire n_1598;
wire n_15255;
wire n_6214;
wire n_9370;
wire n_918;
wire n_13136;
wire n_763;
wire n_6692;
wire n_2485;
wire n_14322;
wire n_12331;
wire n_8093;
wire n_6036;
wire n_13349;
wire n_9956;
wire n_17007;
wire n_6552;
wire n_17096;
wire n_8327;
wire n_13096;
wire n_15314;
wire n_10991;
wire n_14173;
wire n_17005;
wire n_1702;
wire n_4947;
wire n_9487;
wire n_16791;
wire n_14608;
wire n_7306;
wire n_16153;
wire n_10118;
wire n_795;
wire n_18791;
wire n_7470;
wire n_13800;
wire n_19593;
wire n_1245;
wire n_7693;
wire n_3215;
wire n_20568;
wire n_4740;
wire n_20498;
wire n_15662;
wire n_20077;
wire n_1112;
wire n_10002;
wire n_2081;
wire n_911;
wire n_11242;
wire n_17974;
wire n_2862;
wire n_472;
wire n_15923;
wire n_20052;
wire n_2474;
wire n_3703;
wire n_13694;
wire n_4863;
wire n_17494;
wire n_2267;
wire n_668;
wire n_1821;
wire n_9660;
wire n_16233;
wire n_20371;
wire n_17344;
wire n_13093;
wire n_9328;
wire n_16511;
wire n_15274;
wire n_16410;
wire n_7653;
wire n_8354;
wire n_14276;
wire n_6959;
wire n_8353;
wire n_6388;
wire n_5045;
wire n_13185;
wire n_11053;
wire n_18635;
wire n_12159;
wire n_9434;
wire n_18450;
wire n_13855;
wire n_10902;
wire n_19596;
wire n_8348;
wire n_7032;
wire n_19086;
wire n_18806;
wire n_8211;
wire n_1816;
wire n_11304;
wire n_9681;
wire n_5848;
wire n_10485;
wire n_7475;
wire n_18448;
wire n_4612;
wire n_6435;
wire n_10536;
wire n_2531;
wire n_9079;
wire n_15544;
wire n_18738;
wire n_19564;
wire n_16145;
wire n_19424;
wire n_17512;
wire n_18931;
wire n_18988;
wire n_714;
wire n_8653;
wire n_8920;
wire n_17521;
wire n_10950;
wire n_5485;
wire n_17477;
wire n_6682;
wire n_6823;
wire n_14550;
wire n_9089;
wire n_4390;
wire n_15346;
wire n_13477;
wire n_18200;
wire n_2095;
wire n_8942;
wire n_10978;
wire n_8222;
wire n_13808;
wire n_6822;
wire n_3295;
wire n_8553;
wire n_1998;
wire n_240;
wire n_19608;
wire n_17068;
wire n_10187;
wire n_11014;
wire n_17508;
wire n_15033;
wire n_2640;
wire n_3288;
wire n_583;
wire n_17789;
wire n_3876;
wire n_9564;
wire n_7391;
wire n_9230;
wire n_19301;
wire n_941;
wire n_19297;
wire n_10768;
wire n_14067;
wire n_6389;
wire n_15903;
wire n_2471;
wire n_6983;
wire n_10494;
wire n_8398;
wire n_13970;
wire n_19866;
wire n_15247;
wire n_16656;
wire n_4580;
wire n_1055;
wire n_2197;
wire n_10065;
wire n_8700;
wire n_4148;
wire n_2461;
wire n_271;
wire n_13408;
wire n_17585;
wire n_15248;
wire n_13727;
wire n_17500;
wire n_13025;
wire n_10268;
wire n_18728;
wire n_14801;
wire n_12601;
wire n_15399;
wire n_17549;
wire n_13641;
wire n_2634;
wire n_1761;
wire n_20520;
wire n_19588;
wire n_19493;
wire n_8750;
wire n_17473;
wire n_17746;
wire n_5868;
wire n_10305;
wire n_2308;
wire n_16862;
wire n_3001;
wire n_12807;
wire n_15669;
wire n_18018;
wire n_3795;
wire n_7321;
wire n_5289;
wire n_8200;
wire n_4138;
wire n_16055;
wire n_19053;
wire n_18179;
wire n_18564;
wire n_3815;
wire n_12981;
wire n_19950;
wire n_6254;
wire n_1862;
wire n_5989;
wire n_339;
wire n_434;
wire n_13542;
wire n_288;
wire n_8212;
wire n_5612;
wire n_20293;
wire n_20047;
wire n_9016;
wire n_14426;
wire n_15456;
wire n_11545;
wire n_8846;
wire n_4834;
wire n_12665;
wire n_19469;
wire n_16526;
wire n_16397;
wire n_11850;
wire n_9194;
wire n_8760;
wire n_12592;
wire n_17467;
wire n_9029;
wire n_6837;
wire n_3813;
wire n_18860;
wire n_1613;
wire n_11043;
wire n_9414;
wire n_18539;
wire n_7023;
wire n_9615;
wire n_14205;
wire n_1189;
wire n_18532;
wire n_5034;
wire n_726;
wire n_10779;
wire n_11061;
wire n_16495;
wire n_17922;
wire n_5375;
wire n_15742;
wire n_16686;
wire n_16347;
wire n_5370;
wire n_9811;
wire n_5784;
wire n_3443;
wire n_7899;
wire n_8631;
wire n_16385;
wire n_19141;
wire n_1708;
wire n_805;
wire n_14723;
wire n_2051;
wire n_5112;
wire n_19205;
wire n_1402;
wire n_1691;
wire n_10520;
wire n_17437;
wire n_13531;
wire n_7797;
wire n_3668;
wire n_18641;
wire n_13880;
wire n_7687;
wire n_2491;
wire n_19992;
wire n_1264;
wire n_18251;
wire n_4087;
wire n_7582;
wire n_10541;
wire n_14587;
wire n_8959;
wire n_17326;
wire n_10614;
wire n_18834;
wire n_7809;
wire n_461;
wire n_16877;
wire n_18169;
wire n_8425;
wire n_11257;
wire n_15176;
wire n_9910;
wire n_16790;
wire n_10217;
wire n_17255;
wire n_2513;
wire n_10743;
wire n_2247;
wire n_13424;
wire n_14658;
wire n_15066;
wire n_1579;
wire n_20481;
wire n_9651;
wire n_3275;
wire n_836;
wire n_15474;
wire n_15316;
wire n_10270;
wire n_11115;
wire n_8001;
wire n_2094;
wire n_1511;
wire n_17417;
wire n_20260;
wire n_7529;
wire n_14233;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_1313;
wire n_3607;
wire n_3316;
wire n_2418;
wire n_6881;
wire n_3371;
wire n_19269;
wire n_9544;
wire n_3261;
wire n_17324;
wire n_666;
wire n_7520;
wire n_9831;
wire n_4187;
wire n_940;
wire n_18245;
wire n_9697;
wire n_18878;
wire n_5317;
wire n_18414;
wire n_494;
wire n_8362;
wire n_2394;
wire n_5540;
wire n_6300;
wire n_8256;
wire n_5716;
wire n_9310;
wire n_10132;
wire n_3948;
wire n_12091;
wire n_8704;
wire n_17589;
wire n_6132;
wire n_5211;
wire n_17493;
wire n_9294;
wire n_11747;
wire n_6395;
wire n_976;
wire n_7054;
wire n_2686;
wire n_5327;
wire n_4392;
wire n_11858;
wire n_14027;
wire n_7433;
wire n_16316;
wire n_10075;
wire n_10423;
wire n_17762;
wire n_4334;
wire n_3351;
wire n_6171;
wire n_17291;
wire n_17895;
wire n_5519;
wire n_11895;
wire n_13458;
wire n_4047;
wire n_7092;
wire n_6980;
wire n_11213;
wire n_10886;
wire n_18720;
wire n_13091;
wire n_3791;
wire n_13003;
wire n_6387;
wire n_10192;
wire n_9465;
wire n_13811;
wire n_5139;
wire n_757;
wire n_19459;
wire n_14011;
wire n_166;
wire n_10436;
wire n_19026;
wire n_12794;
wire n_15496;
wire n_6342;
wire n_17744;
wire n_15260;
wire n_15104;
wire n_12483;
wire n_20086;
wire n_16374;
wire n_18173;
wire n_17251;
wire n_3883;
wire n_18945;
wire n_261;
wire n_5866;
wire n_3728;
wire n_2925;
wire n_5822;
wire n_17381;
wire n_9959;
wire n_15055;
wire n_3949;
wire n_11015;
wire n_18712;
wire n_5364;
wire n_3315;
wire n_9631;
wire n_14751;
wire n_6194;
wire n_20226;
wire n_4893;
wire n_18313;
wire n_12815;
wire n_15913;
wire n_10431;
wire n_9945;
wire n_1413;
wire n_2228;
wire n_17694;
wire n_5039;
wire n_16314;
wire n_2455;
wire n_4772;
wire n_15115;
wire n_8746;
wire n_20319;
wire n_11183;
wire n_10019;
wire n_8531;
wire n_12093;
wire n_19296;
wire n_11581;
wire n_4468;
wire n_4161;
wire n_6459;
wire n_8379;
wire n_13100;
wire n_4961;
wire n_4454;
wire n_16154;
wire n_12334;
wire n_18397;
wire n_9209;
wire n_7311;
wire n_3686;
wire n_18234;
wire n_7669;
wire n_8793;
wire n_12355;
wire n_19340;
wire n_15052;
wire n_9838;
wire n_9767;
wire n_1713;
wire n_4277;
wire n_9300;
wire n_11500;
wire n_12943;
wire n_17598;
wire n_530;
wire n_17956;
wire n_618;
wire n_11021;
wire n_8543;
wire n_16502;
wire n_3069;
wire n_7189;
wire n_13067;
wire n_6258;
wire n_16688;
wire n_10243;
wire n_9700;
wire n_18114;
wire n_18802;
wire n_3725;
wire n_8533;
wire n_15483;
wire n_9118;
wire n_11122;
wire n_6657;
wire n_5554;
wire n_1175;
wire n_10596;
wire n_20512;
wire n_19671;
wire n_903;
wire n_12140;
wire n_1802;
wire n_286;
wire n_254;
wire n_8063;
wire n_3961;
wire n_12599;
wire n_2347;
wire n_19419;
wire n_816;
wire n_8032;
wire n_7427;
wire n_2967;
wire n_13250;
wire n_11190;
wire n_11794;
wire n_10519;
wire n_2467;
wire n_17630;
wire n_10163;
wire n_17409;
wire n_3983;
wire n_3538;
wire n_20186;
wire n_16544;
wire n_2824;
wire n_17529;
wire n_18979;
wire n_12330;
wire n_950;
wire n_15871;
wire n_14819;
wire n_14890;
wire n_8129;
wire n_13906;
wire n_3009;
wire n_5824;
wire n_6760;
wire n_14265;
wire n_13664;
wire n_13566;
wire n_12591;
wire n_12466;
wire n_9509;
wire n_3526;
wire n_20089;
wire n_4367;
wire n_10874;
wire n_6825;
wire n_19558;
wire n_11831;
wire n_16213;
wire n_14399;
wire n_9628;
wire n_18940;
wire n_19348;
wire n_2583;
wire n_18279;
wire n_19655;
wire n_10250;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_18658;
wire n_14063;
wire n_16657;
wire n_2078;
wire n_2932;
wire n_3431;
wire n_3450;
wire n_17584;
wire n_12041;
wire n_449;
wire n_16734;
wire n_17783;
wire n_2728;
wire n_15157;
wire n_13074;
wire n_3183;
wire n_1067;
wire n_14716;
wire n_255;
wire n_1952;
wire n_12876;
wire n_15286;
wire n_14698;
wire n_19152;
wire n_18633;
wire n_6468;
wire n_3937;
wire n_3159;
wire n_14323;
wire n_18565;
wire n_13071;
wire n_6857;
wire n_3576;
wire n_1863;
wire n_12536;
wire n_10795;
wire n_16333;
wire n_872;
wire n_15116;
wire n_8049;
wire n_7762;
wire n_9467;
wire n_7186;
wire n_13739;
wire n_11157;
wire n_19809;
wire n_9097;
wire n_1513;
wire n_14364;
wire n_15472;
wire n_837;
wire n_5087;
wire n_13234;
wire n_9314;
wire n_7017;
wire n_16718;
wire n_2060;
wire n_7830;
wire n_5131;
wire n_19217;
wire n_17380;
wire n_8084;
wire n_14113;
wire n_8289;
wire n_11178;
wire n_20492;
wire n_5887;
wire n_16428;
wire n_19010;
wire n_14938;
wire n_14784;
wire n_2816;
wire n_11432;
wire n_14179;
wire n_17755;
wire n_7191;
wire n_14979;
wire n_10412;
wire n_12650;
wire n_19935;
wire n_4443;
wire n_14324;
wire n_614;
wire n_5460;
wire n_1615;
wire n_4114;
wire n_12859;
wire n_2119;
wire n_17763;
wire n_7961;
wire n_5899;
wire n_17176;
wire n_10617;
wire n_3185;
wire n_2605;
wire n_16524;
wire n_10544;
wire n_13030;
wire n_2848;
wire n_919;
wire n_17819;
wire n_18475;
wire n_15094;
wire n_16880;
wire n_20287;
wire n_20153;
wire n_11952;
wire n_6422;
wire n_1299;
wire n_13896;
wire n_5339;
wire n_3837;
wire n_16473;
wire n_1436;
wire n_9873;
wire n_13299;
wire n_13042;
wire n_4818;
wire n_15658;
wire n_10095;
wire n_15873;
wire n_8268;
wire n_6160;
wire n_19749;
wire n_7066;
wire n_18128;
wire n_796;
wire n_7789;
wire n_184;
wire n_6192;
wire n_10056;
wire n_16597;
wire n_17627;
wire n_18815;
wire n_6039;
wire n_2144;
wire n_20296;
wire n_11919;
wire n_1142;
wire n_11414;
wire n_17705;
wire n_5719;
wire n_17728;
wire n_19457;
wire n_17618;
wire n_7344;
wire n_9888;
wire n_10037;
wire n_2259;
wire n_18029;
wire n_6707;
wire n_12744;
wire n_19601;
wire n_11136;
wire n_19790;
wire n_3142;
wire n_19527;
wire n_19672;
wire n_6787;
wire n_11620;
wire n_15480;
wire n_10179;
wire n_4709;
wire n_2132;
wire n_14038;
wire n_18726;
wire n_11215;
wire n_2860;
wire n_2330;
wire n_11890;
wire n_9366;
wire n_14253;
wire n_7915;
wire n_5893;
wire n_9077;
wire n_2281;
wire n_8406;
wire n_15919;
wire n_16652;
wire n_12443;
wire n_6463;
wire n_11683;
wire n_20135;
wire n_8554;
wire n_386;
wire n_6051;
wire n_2301;
wire n_7538;
wire n_12934;
wire n_3270;
wire n_19547;
wire n_18981;
wire n_970;
wire n_6799;
wire n_19368;
wire n_444;
wire n_3913;
wire n_3311;
wire n_6487;
wire n_8818;
wire n_16648;
wire n_4348;
wire n_16724;
wire n_10466;
wire n_11953;
wire n_4404;
wire n_439;
wire n_6563;
wire n_20415;
wire n_2828;
wire n_7554;
wire n_2384;
wire n_4204;
wire n_19005;
wire n_759;
wire n_18881;
wire n_2724;
wire n_15926;
wire n_20210;
wire n_4513;
wire n_16943;
wire n_11089;
wire n_6341;
wire n_13422;
wire n_7421;
wire n_10166;
wire n_7489;
wire n_1647;
wire n_14702;
wire n_13179;
wire n_15844;
wire n_2306;
wire n_11839;
wire n_18039;
wire n_3683;
wire n_4801;
wire n_19874;
wire n_13834;
wire n_401;
wire n_18277;
wire n_2550;
wire n_8341;
wire n_11193;
wire n_17800;
wire n_17613;
wire n_7188;
wire n_3736;
wire n_11217;
wire n_15651;
wire n_17759;
wire n_20014;
wire n_6923;
wire n_9287;
wire n_7991;
wire n_10877;
wire n_16737;
wire n_14686;
wire n_3284;
wire n_12214;
wire n_427;
wire n_16259;
wire n_8926;
wire n_2995;
wire n_10766;
wire n_4438;
wire n_4844;
wire n_10086;
wire n_4836;
wire n_5439;
wire n_13924;
wire n_4149;
wire n_9608;
wire n_501;
wire n_19539;
wire n_20313;
wire n_20251;
wire n_8817;
wire n_8190;
wire n_1668;
wire n_2777;
wire n_11488;
wire n_13671;
wire n_14876;
wire n_18571;
wire n_1129;
wire n_6987;
wire n_18265;
wire n_11037;
wire n_16925;
wire n_18740;
wire n_14319;
wire n_2911;
wire n_1429;
wire n_5706;
wire n_16763;
wire n_3429;
wire n_17462;
wire n_1593;
wire n_15287;
wire n_1202;
wire n_7671;
wire n_13150;
wire n_5431;
wire n_15103;
wire n_12541;
wire n_8649;
wire n_19757;
wire n_14818;
wire n_19508;
wire n_20422;
wire n_8303;
wire n_6153;
wire n_16512;
wire n_13809;
wire n_8059;
wire n_18364;
wire n_11665;
wire n_6579;
wire n_13590;
wire n_16747;
wire n_11138;
wire n_5798;
wire n_575;
wire n_11731;
wire n_5875;
wire n_16257;
wire n_5621;
wire n_16200;
wire n_16023;
wire n_732;
wire n_2983;
wire n_16041;
wire n_6789;
wire n_12100;
wire n_1042;
wire n_15327;
wire n_17718;
wire n_1728;
wire n_13471;
wire n_17615;
wire n_845;
wire n_19063;
wire n_140;
wire n_8862;
wire n_16161;
wire n_10580;
wire n_17287;
wire n_4870;
wire n_6164;
wire n_13261;
wire n_768;
wire n_9675;
wire n_7786;
wire n_16923;
wire n_11454;
wire n_7609;
wire n_3449;
wire n_2598;
wire n_8900;
wire n_597;
wire n_12523;
wire n_6934;
wire n_1403;
wire n_6737;
wire n_18388;
wire n_4488;
wire n_3767;
wire n_8478;
wire n_16988;
wire n_6695;
wire n_12395;
wire n_4211;
wire n_5867;
wire n_17475;
wire n_17363;
wire n_4656;
wire n_3839;
wire n_10770;
wire n_8497;
wire n_6410;
wire n_17873;
wire n_4915;
wire n_15592;
wire n_16064;
wire n_18524;
wire n_15319;
wire n_235;
wire n_5662;
wire n_3730;
wire n_14452;
wire n_17894;
wire n_13464;
wire n_12670;
wire n_16817;
wire n_18336;
wire n_7667;
wire n_10203;
wire n_10980;
wire n_9174;
wire n_17835;
wire n_2737;
wire n_17459;
wire n_10082;
wire n_7182;
wire n_7365;
wire n_10467;
wire n_9849;
wire n_1622;
wire n_17476;
wire n_9856;
wire n_18449;
wire n_17591;
wire n_18672;
wire n_18848;
wire n_11668;
wire n_7885;
wire n_15684;
wire n_2171;
wire n_16720;
wire n_9349;
wire n_17423;
wire n_3136;
wire n_11091;
wire n_4192;
wire n_10940;
wire n_16463;
wire n_15976;
wire n_2808;
wire n_18100;
wire n_17723;
wire n_8839;
wire n_4174;
wire n_12891;
wire n_11615;
wire n_1171;
wire n_11059;
wire n_16403;
wire n_1827;
wire n_14616;
wire n_16799;
wire n_2187;
wire n_6058;
wire n_17965;
wire n_7745;
wire n_12941;
wire n_20219;
wire n_2872;
wire n_14258;
wire n_12200;
wire n_14024;
wire n_2046;
wire n_17212;
wire n_8684;
wire n_13682;
wire n_6249;
wire n_11060;
wire n_5480;
wire n_18943;
wire n_4831;
wire n_11461;
wire n_10714;
wire n_6969;
wire n_7459;
wire n_6161;
wire n_2970;
wire n_8206;
wire n_18070;
wire n_2882;
wire n_4260;
wire n_18338;
wire n_19908;
wire n_6607;
wire n_9335;
wire n_1974;
wire n_4122;
wire n_9452;
wire n_11427;
wire n_19293;
wire n_934;
wire n_5284;
wire n_12673;
wire n_14694;
wire n_8513;
wire n_10120;
wire n_9474;
wire n_19818;
wire n_19208;
wire n_9427;
wire n_17817;
wire n_6294;
wire n_543;
wire n_9611;
wire n_18371;
wire n_9021;
wire n_16269;
wire n_9250;
wire n_11212;
wire n_13145;
wire n_804;
wire n_9550;
wire n_16591;
wire n_11263;
wire n_10641;
wire n_959;
wire n_4312;
wire n_18805;
wire n_16566;
wire n_13195;
wire n_8694;
wire n_13965;
wire n_5048;
wire n_11994;
wire n_13358;
wire n_2195;
wire n_3208;
wire n_18759;
wire n_16693;
wire n_14519;
wire n_6123;
wire n_11000;
wire n_16125;
wire n_20430;
wire n_4935;
wire n_19403;
wire n_8191;
wire n_10325;
wire n_16354;
wire n_10298;
wire n_6922;
wire n_16701;
wire n_7698;
wire n_12854;
wire n_16427;
wire n_16336;
wire n_8431;
wire n_19631;
wire n_2945;
wire n_3061;
wire n_16248;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_10400;
wire n_19081;
wire n_9177;
wire n_9060;
wire n_11947;
wire n_14496;
wire n_9096;
wire n_13952;
wire n_11697;
wire n_16963;
wire n_18074;
wire n_7891;
wire n_14413;
wire n_8517;
wire n_3008;
wire n_4776;
wire n_4153;
wire n_10901;
wire n_11034;
wire n_10549;
wire n_12115;
wire n_1962;
wire n_11499;
wire n_10825;
wire n_4723;
wire n_17292;
wire n_4269;
wire n_18023;
wire n_14777;
wire n_14057;
wire n_5459;
wire n_17788;
wire n_4143;
wire n_876;
wire n_16406;
wire n_12558;
wire n_11984;
wire n_11948;
wire n_4719;
wire n_7477;
wire n_17028;
wire n_15654;
wire n_1904;
wire n_17289;
wire n_2588;
wire n_11402;
wire n_1353;
wire n_11401;
wire n_17828;
wire n_19679;
wire n_17820;
wire n_2366;
wire n_10581;
wire n_14949;
wire n_17487;
wire n_4423;
wire n_2210;
wire n_3602;
wire n_18372;
wire n_12086;
wire n_1411;
wire n_16952;
wire n_566;
wire n_16449;
wire n_2951;
wire n_11589;
wire n_11246;
wire n_1807;
wire n_18266;
wire n_16606;
wire n_14460;
wire n_13216;
wire n_209;
wire n_12849;
wire n_11312;
wire n_13786;
wire n_5909;
wire n_9344;
wire n_671;
wire n_19719;
wire n_10865;
wire n_740;
wire n_10738;
wire n_7378;
wire n_9798;
wire n_15491;
wire n_14925;
wire n_11612;
wire n_4229;
wire n_12447;
wire n_13417;
wire n_12296;
wire n_13414;
wire n_3865;
wire n_4073;
wire n_5400;
wire n_7498;
wire n_3846;
wire n_11916;
wire n_180;
wire n_3512;
wire n_7501;
wire n_5201;
wire n_10421;
wire n_10976;
wire n_6465;
wire n_9447;
wire n_12764;
wire n_15325;
wire n_1326;
wire n_4783;
wire n_18987;
wire n_20268;
wire n_19091;
wire n_14238;
wire n_16918;
wire n_12409;
wire n_11625;
wire n_1130;
wire n_17054;
wire n_20053;
wire n_6592;
wire n_9712;
wire n_6626;
wire n_8585;
wire n_19877;
wire n_14042;
wire n_9220;
wire n_17312;
wire n_12763;
wire n_378;
wire n_18460;
wire n_17272;
wire n_16394;
wire n_18869;
wire n_20136;
wire n_15310;
wire n_17989;
wire n_1283;
wire n_4917;
wire n_8698;
wire n_12584;
wire n_14435;
wire n_4432;
wire n_10376;
wire n_15510;
wire n_7515;
wire n_17567;
wire n_344;
wire n_9994;
wire n_14226;
wire n_7309;
wire n_15811;
wire n_5114;
wire n_1392;
wire n_8559;
wire n_20123;
wire n_5693;
wire n_17670;
wire n_15618;
wire n_2463;
wire n_10224;
wire n_15849;
wire n_611;
wire n_18758;
wire n_3062;
wire n_2679;
wire n_20545;
wire n_19951;
wire n_9391;
wire n_16105;
wire n_8514;
wire n_14515;
wire n_14159;
wire n_9134;
wire n_12268;
wire n_18990;
wire n_12077;
wire n_15321;
wire n_14757;
wire n_1017;
wire n_5396;
wire n_12534;
wire n_6846;
wire n_13271;
wire n_11481;
wire n_10175;
wire n_15812;
wire n_16292;
wire n_18458;
wire n_6886;
wire n_17019;
wire n_5365;
wire n_8405;
wire n_15223;
wire n_11350;
wire n_626;
wire n_11925;
wire n_16033;
wire n_8672;
wire n_1104;
wire n_4920;
wire n_1253;
wire n_6446;
wire n_3256;
wire n_9430;
wire n_19279;
wire n_7218;
wire n_11407;
wire n_2118;
wire n_19548;
wire n_12710;
wire n_19331;
wire n_2188;
wire n_8440;
wire n_7005;
wire n_9776;
wire n_16736;
wire n_6777;
wire n_18156;
wire n_11987;
wire n_18208;
wire n_19206;
wire n_8475;
wire n_8029;
wire n_18845;
wire n_18527;
wire n_4861;
wire n_4064;
wire n_1829;
wire n_13089;
wire n_15459;
wire n_15192;
wire n_5266;
wire n_4828;
wire n_1638;
wire n_18360;
wire n_16836;
wire n_13167;
wire n_12329;
wire n_519;
wire n_15013;
wire n_6953;
wire n_3669;
wire n_16710;
wire n_14945;
wire n_4316;
wire n_5122;
wire n_5390;
wire n_18660;
wire n_18348;
wire n_19658;
wire n_18487;
wire n_9834;
wire n_16353;
wire n_2047;
wire n_12318;
wire n_5385;
wire n_13278;
wire n_13597;
wire n_5322;
wire n_3989;
wire n_7089;
wire n_2490;
wire n_18232;
wire n_3841;
wire n_20317;
wire n_1996;
wire n_6332;
wire n_1442;
wire n_20206;
wire n_7403;
wire n_7338;
wire n_5917;
wire n_7129;
wire n_4909;
wire n_13938;
wire n_13251;
wire n_8566;
wire n_7343;
wire n_12766;
wire n_18913;
wire n_8317;
wire n_12229;
wire n_269;
wire n_6116;
wire n_7492;
wire n_13319;
wire n_9071;
wire n_10415;
wire n_7694;
wire n_11711;
wire n_18637;
wire n_15666;
wire n_20509;
wire n_11931;
wire n_8109;
wire n_2055;
wire n_18971;
wire n_12780;
wire n_14017;
wire n_13267;
wire n_7987;
wire n_9133;
wire n_16054;
wire n_12664;
wire n_14942;
wire n_7434;
wire n_9009;
wire n_6155;
wire n_20449;
wire n_7269;
wire n_9777;
wire n_15359;
wire n_9063;
wire n_7787;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_5304;
wire n_15035;
wire n_18500;
wire n_19085;
wire n_18536;
wire n_6261;
wire n_4281;
wire n_19893;
wire n_4648;
wire n_10096;
wire n_13617;
wire n_10025;
wire n_412;
wire n_18779;
wire n_6299;
wire n_20573;
wire n_11753;
wire n_7425;
wire n_19061;
wire n_1059;
wire n_11150;
wire n_18199;
wire n_4360;
wire n_16111;
wire n_3263;
wire n_6316;
wire n_6292;
wire n_9726;
wire n_1748;
wire n_13884;
wire n_17125;
wire n_7719;
wire n_5615;
wire n_6220;
wire n_12783;
wire n_1885;
wire n_1240;
wire n_17671;
wire n_1234;
wire n_14195;
wire n_18363;
wire n_3254;
wire n_3684;
wire n_20479;
wire n_7938;
wire n_3152;
wire n_7935;
wire n_8458;
wire n_6772;
wire n_16902;
wire n_16646;
wire n_14300;
wire n_6077;
wire n_1003;
wire n_11512;
wire n_17090;
wire n_14678;
wire n_13599;
wire n_17282;
wire n_15008;
wire n_5188;
wire n_13647;
wire n_4490;
wire n_13683;
wire n_1575;
wire n_19094;
wire n_10147;
wire n_17921;
wire n_17197;
wire n_18503;
wire n_20474;
wire n_9298;
wire n_18058;
wire n_16939;
wire n_14497;
wire n_1991;
wire n_5161;
wire n_14280;
wire n_4078;
wire n_13724;
wire n_9301;
wire n_3046;
wire n_5382;
wire n_12054;
wire n_15827;
wire n_5659;
wire n_8099;
wire n_17256;
wire n_11595;
wire n_17806;
wire n_13768;
wire n_1415;
wire n_16707;
wire n_8578;
wire n_1370;
wire n_7222;
wire n_13838;
wire n_10046;
wire n_2291;
wire n_2184;
wire n_10397;
wire n_2982;
wire n_19379;
wire n_10936;
wire n_12442;
wire n_8611;
wire n_1517;
wire n_8819;
wire n_17927;
wire n_2630;
wire n_15123;
wire n_9835;
wire n_15021;
wire n_12839;
wire n_6697;
wire n_7875;
wire n_13153;
wire n_7643;
wire n_13441;
wire n_16082;
wire n_10207;
wire n_13857;
wire n_18872;
wire n_1143;
wire n_10401;
wire n_19352;
wire n_7242;
wire n_17737;
wire n_19240;
wire n_13816;
wire n_18355;
wire n_2013;
wire n_17215;
wire n_19737;
wire n_14736;
wire n_10139;
wire n_13246;
wire n_14061;
wire n_12986;
wire n_11381;
wire n_16378;
wire n_16109;
wire n_7224;
wire n_12441;
wire n_15789;
wire n_16611;
wire n_16172;
wire n_7746;
wire n_3662;
wire n_2981;
wire n_18108;
wire n_16598;
wire n_16277;
wire n_17588;
wire n_12516;
wire n_8414;
wire n_13921;
wire n_6297;
wire n_6653;
wire n_16806;
wire n_15512;
wire n_18836;
wire n_12377;
wire n_638;
wire n_18486;
wire n_5492;
wire n_9965;
wire n_13650;
wire n_16789;
wire n_887;
wire n_15636;
wire n_15946;
wire n_6501;
wire n_18063;
wire n_9990;
wire n_10005;
wire n_12905;
wire n_11426;
wire n_2599;
wire n_15311;
wire n_8505;
wire n_19827;
wire n_3368;
wire n_17667;
wire n_7884;
wire n_11258;
wire n_19879;
wire n_15498;
wire n_20477;
wire n_7417;
wire n_18097;
wire n_4881;
wire n_12513;
wire n_5734;
wire n_13395;
wire n_4255;
wire n_4071;
wire n_20016;
wire n_7388;
wire n_3568;
wire n_11657;
wire n_8717;
wire n_5770;
wire n_5705;
wire n_3313;
wire n_9064;
wire n_17420;
wire n_2725;
wire n_14135;
wire n_8571;
wire n_16482;
wire n_4305;
wire n_12514;
wire n_10048;
wire n_16809;
wire n_14194;
wire n_619;
wire n_13825;
wire n_19945;
wire n_18942;
wire n_8243;
wire n_6347;
wire n_9593;
wire n_606;
wire n_13398;
wire n_8449;
wire n_17605;
wire n_630;
wire n_13204;
wire n_4094;
wire n_14331;
wire n_18994;
wire n_4765;
wire n_2522;
wire n_4364;
wire n_9406;
wire n_8967;
wire n_9322;
wire n_15017;
wire n_5959;
wire n_3720;
wire n_8031;
wire n_15591;
wire n_264;
wire n_12188;
wire n_16609;
wire n_4745;
wire n_5642;
wire n_9232;
wire n_15167;
wire n_12299;
wire n_16739;
wire n_15706;
wire n_1680;
wire n_3842;
wire n_993;
wire n_1605;
wire n_11327;
wire n_4979;
wire n_1988;
wire n_15900;
wire n_12000;
wire n_17281;
wire n_19004;
wire n_1233;
wire n_14182;
wire n_241;
wire n_10279;
wire n_15853;
wire n_4520;
wire n_5299;
wire n_3455;
wire n_14352;
wire n_13889;
wire n_17864;
wire n_7081;
wire n_13015;
wire n_20112;
wire n_7319;
wire n_15831;
wire n_7644;
wire n_11176;
wire n_9883;
wire n_11135;
wire n_5668;
wire n_11275;
wire n_268;
wire n_18850;
wire n_5463;
wire n_12700;
wire n_12904;
wire n_5489;
wire n_1165;
wire n_14623;
wire n_4773;
wire n_7910;
wire n_6009;
wire n_3281;
wire n_9034;
wire n_7084;
wire n_5923;
wire n_14073;
wire n_8074;
wire n_13639;
wire n_15989;
wire n_8860;
wire n_2676;
wire n_3940;
wire n_1214;
wire n_15514;
wire n_9266;
wire n_3453;
wire n_3410;
wire n_16210;
wire n_10027;
wire n_12784;
wire n_1813;
wire n_18639;
wire n_825;
wire n_12877;
wire n_14677;
wire n_14261;
wire n_18020;
wire n_10616;
wire n_8587;
wire n_5366;
wire n_16016;
wire n_15550;
wire n_15528;
wire n_6925;
wire n_6878;
wire n_9078;
wire n_16297;
wire n_16896;
wire n_13198;
wire n_15914;
wire n_3289;
wire n_13741;
wire n_12610;
wire n_14416;
wire n_11251;
wire n_12293;
wire n_2036;
wire n_6470;
wire n_11598;
wire n_8368;
wire n_15691;
wire n_17560;
wire n_8322;
wire n_16127;
wire n_6187;
wire n_8300;
wire n_9378;
wire n_678;
wire n_12206;
wire n_18112;
wire n_17488;
wire n_17427;
wire n_11400;
wire n_19532;
wire n_19870;
wire n_6693;
wire n_15848;
wire n_11563;
wire n_362;
wire n_12444;
wire n_18586;
wire n_16409;
wire n_5419;
wire n_14513;
wire n_2943;
wire n_12778;
wire n_12485;
wire n_3253;
wire n_15995;
wire n_14602;
wire n_11468;
wire n_16150;
wire n_4603;
wire n_9683;
wire n_17403;
wire n_15132;
wire n_1527;
wire n_495;
wire n_5732;
wire n_11878;
wire n_15843;
wire n_16666;
wire n_4471;
wire n_15749;
wire n_7449;
wire n_15638;
wire n_16547;
wire n_14289;
wire n_1493;
wire n_16479;
wire n_10751;
wire n_16967;
wire n_10240;
wire n_10691;
wire n_2535;
wire n_9561;
wire n_19351;
wire n_16104;
wire n_20445;
wire n_9773;
wire n_2436;
wire n_3838;
wire n_9745;
wire n_3941;
wire n_15413;
wire n_15628;
wire n_10216;
wire n_17733;
wire n_1514;
wire n_10150;
wire n_12581;
wire n_17395;
wire n_4994;
wire n_6652;
wire n_10971;
wire n_5168;
wire n_4661;
wire n_20116;
wire n_18506;
wire n_7674;
wire n_14516;
wire n_18484;
wire n_12305;
wire n_12170;
wire n_2853;
wire n_9630;
wire n_13927;
wire n_13313;
wire n_15308;
wire n_17025;
wire n_9255;
wire n_10231;
wire n_8310;
wire n_16500;
wire n_9758;
wire n_15175;
wire n_8936;
wire n_7126;
wire n_18413;
wire n_15206;
wire n_9691;
wire n_12997;
wire n_14005;
wire n_14293;
wire n_14334;
wire n_7690;
wire n_15245;
wire n_15225;
wire n_3229;
wire n_11223;
wire n_13562;
wire n_14537;
wire n_6950;
wire n_10038;
wire n_17794;
wire n_15614;
wire n_20234;
wire n_2012;
wire n_5066;
wire n_18101;
wire n_2842;
wire n_19087;
wire n_11221;
wire n_15772;
wire n_14245;
wire n_20322;
wire n_17659;
wire n_11448;
wire n_17321;
wire n_18272;
wire n_1809;
wire n_8328;
wire n_15502;
wire n_15076;
wire n_12576;
wire n_7258;
wire n_10579;
wire n_13345;
wire n_3677;
wire n_8336;
wire n_20376;
wire n_3996;
wire n_17492;
wire n_19324;
wire n_20008;
wire n_4218;
wire n_11445;
wire n_13151;
wire n_3685;
wire n_11552;
wire n_15102;
wire n_14733;
wire n_417;
wire n_14317;
wire n_19807;
wire n_4459;
wire n_16220;
wire n_9852;
wire n_11623;
wire n_3019;
wire n_3471;
wire n_5295;
wire n_2368;
wire n_18599;
wire n_14131;
wire n_8041;
wire n_10676;
wire n_17931;
wire n_4175;
wire n_10540;
wire n_10299;
wire n_16993;
wire n_12845;
wire n_11645;
wire n_10200;
wire n_3259;
wire n_2524;
wire n_13164;
wire n_2460;
wire n_13662;
wire n_3867;
wire n_3593;
wire n_1073;
wire n_16275;
wire n_17062;
wire n_13340;
wire n_17887;
wire n_17192;
wire n_4140;
wire n_2481;
wire n_9939;
wire n_7766;
wire n_19397;
wire n_12797;
wire n_20561;
wire n_6758;
wire n_5160;
wire n_19709;
wire n_9481;
wire n_7955;
wire n_17081;
wire n_1207;
wire n_12012;
wire n_7287;
wire n_10076;
wire n_880;
wire n_6464;
wire n_18675;
wire n_20508;
wire n_3540;
wire n_11554;
wire n_150;
wire n_1478;
wire n_3777;
wire n_4203;
wire n_767;
wire n_1837;
wire n_4533;
wire n_9635;
wire n_19619;
wire n_1410;
wire n_14308;
wire n_5408;
wire n_1736;
wire n_3848;
wire n_319;
wire n_8181;
wire n_2511;
wire n_8254;
wire n_13452;
wire n_8071;
wire n_5271;
wire n_17480;
wire n_562;
wire n_6004;
wire n_5964;
wire n_11628;
wire n_20218;
wire n_1136;
wire n_11549;
wire n_20177;
wire n_17162;
wire n_12286;
wire n_9001;
wire n_19517;
wire n_2329;
wire n_16107;
wire n_14545;
wire n_18031;
wire n_8013;
wire n_146;
wire n_19670;
wire n_193;
wire n_16683;
wire n_17804;
wire n_12347;
wire n_19346;
wire n_17424;
wire n_20262;
wire n_296;
wire n_651;
wire n_3407;
wire n_5992;
wire n_217;
wire n_1185;
wire n_19394;
wire n_215;
wire n_17818;
wire n_20378;
wire n_12698;
wire n_2621;
wire n_6540;
wire n_16086;
wire n_5513;
wire n_5614;
wire n_497;
wire n_17383;
wire n_11871;
wire n_16857;
wire n_1315;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_15326;
wire n_17555;
wire n_18957;
wire n_7722;
wire n_3188;
wire n_1459;
wire n_20329;
wire n_2462;
wire n_4056;
wire n_9240;
wire n_8293;
wire n_14726;
wire n_14180;
wire n_18697;
wire n_10548;
wire n_12957;
wire n_11616;
wire n_8791;
wire n_8288;
wire n_1091;
wire n_1425;
wire n_12786;
wire n_983;
wire n_10678;
wire n_6757;
wire n_17752;
wire n_18045;
wire n_1390;
wire n_2289;
wire n_8323;
wire n_10391;
wire n_13176;
wire n_9784;
wire n_19647;
wire n_7990;
wire n_18368;
wire n_10036;
wire n_17631;
wire n_5278;
wire n_14905;
wire n_15128;
wire n_3688;
wire n_8720;
wire n_12205;
wire n_11989;
wire n_16912;
wire n_16215;
wire n_1905;
wire n_14009;
wire n_3466;
wire n_5704;
wire n_15787;
wire n_19943;
wire n_7148;
wire n_5956;
wire n_9417;
wire n_2139;
wire n_12020;
wire n_18875;
wire n_6835;
wire n_1203;
wire n_11624;
wire n_20275;
wire n_8826;
wire n_15083;
wire n_11352;
wire n_19290;
wire n_5516;
wire n_2841;
wire n_6247;
wire n_11234;
wire n_10919;
wire n_12099;
wire n_12858;
wire n_4399;
wire n_15351;
wire n_2487;
wire n_18170;
wire n_19159;
wire n_7544;
wire n_9336;
wire n_19750;
wire n_3572;
wire n_8854;
wire n_6645;
wire n_16177;
wire n_10727;
wire n_10885;
wire n_443;
wire n_13201;
wire n_14759;
wire n_13274;
wire n_18621;
wire n_9312;
wire n_5174;
wire n_7469;
wire n_5538;
wire n_5017;
wire n_10895;
wire n_198;
wire n_11977;
wire n_15576;
wire n_11696;
wire n_11734;
wire n_9533;
wire n_9494;
wire n_5241;
wire n_11507;
wire n_17290;
wire n_15337;
wire n_17276;
wire n_7082;
wire n_14749;
wire n_18731;
wire n_20000;
wire n_3108;
wire n_19306;
wire n_11320;
wire n_11837;
wire n_19458;
wire n_8260;
wire n_3417;
wire n_13898;
wire n_16507;
wire n_4124;
wire n_16543;
wire n_11938;
wire n_6418;
wire n_17003;
wire n_5153;
wire n_18814;
wire n_609;
wire n_10571;
wire n_19202;
wire n_19664;
wire n_9807;
wire n_9057;
wire n_8706;
wire n_2607;
wire n_7945;
wire n_8894;
wire n_19244;
wire n_2890;
wire n_12053;
wire n_15947;
wire n_17738;
wire n_12619;
wire n_1320;
wire n_20488;
wire n_11289;
wire n_13555;
wire n_2499;
wire n_12582;
wire n_5487;
wire n_18919;
wire n_12423;
wire n_15426;
wire n_14137;
wire n_16905;
wire n_17765;
wire n_14163;
wire n_15523;
wire n_2472;
wire n_7328;
wire n_19298;
wire n_10958;
wire n_15682;
wire n_9479;
wire n_15556;
wire n_3957;
wire n_14041;
wire n_18622;
wire n_9181;
wire n_19338;
wire n_19385;
wire n_6578;
wire n_3040;
wire n_14763;
wire n_19319;
wire n_17686;
wire n_18381;
wire n_10879;
wire n_19481;
wire n_5951;
wire n_6589;
wire n_1864;
wire n_10639;
wire n_16359;
wire n_3475;
wire n_17448;
wire n_18657;
wire n_16037;
wire n_13351;
wire n_9276;
wire n_579;
wire n_5152;
wire n_16805;
wire n_15937;
wire n_20453;
wire n_16141;
wire n_4927;
wire n_5574;
wire n_9821;
wire n_11112;
wire n_4258;
wire n_2699;
wire n_11723;
wire n_650;
wire n_16647;
wire n_1940;
wire n_1405;
wire n_5469;
wire n_14393;
wire n_456;
wire n_12364;
wire n_3878;
wire n_12420;
wire n_6567;
wire n_313;
wire n_20574;
wire n_5895;
wire n_5804;
wire n_9508;
wire n_3134;
wire n_16231;
wire n_896;
wire n_4553;
wire n_3278;
wire n_20423;
wire n_17805;
wire n_20181;
wire n_17318;
wire n_11906;
wire n_20586;
wire n_2673;
wire n_2456;
wire n_14298;
wire n_9741;
wire n_1637;
wire n_3307;
wire n_1407;
wire n_2871;
wire n_420;
wire n_10180;
wire n_4183;
wire n_14112;
wire n_12120;
wire n_10650;
wire n_12021;
wire n_10157;
wire n_7423;
wire n_10402;
wire n_12515;
wire n_17283;
wire n_9166;
wire n_1640;
wire n_12895;
wire n_12045;
wire n_2141;
wire n_6940;
wire n_12726;
wire n_12668;
wire n_7835;
wire n_15437;
wire n_20536;
wire n_6320;
wire n_20570;
wire n_799;
wire n_3044;
wire n_9969;
wire n_11437;
wire n_14068;
wire n_14853;
wire n_16735;
wire n_11869;
wire n_5620;
wire n_20214;
wire n_10836;
wire n_159;
wire n_16375;
wire n_2125;
wire n_8072;
wire n_13117;
wire n_7130;
wire n_2992;
wire n_1241;
wire n_3221;
wire n_11282;
wire n_17720;
wire n_14700;
wire n_16382;
wire n_7491;
wire n_1706;
wire n_18944;
wire n_18474;
wire n_4052;
wire n_20138;
wire n_9636;
wire n_7559;
wire n_13175;
wire n_2441;
wire n_9833;
wire n_9095;
wire n_15757;
wire n_18465;
wire n_5907;
wire n_15979;
wire n_19076;
wire n_1559;
wire n_6731;
wire n_4315;
wire n_2888;
wire n_6154;
wire n_6943;
wire n_4301;
wire n_3744;
wire n_12038;
wire n_8210;
wire n_12644;
wire n_1360;
wire n_11826;
wire n_18241;
wire n_3781;
wire n_10888;
wire n_2484;
wire n_10116;
wire n_16764;
wire n_14808;
wire n_2126;
wire n_18135;
wire n_3843;
wire n_11764;
wire n_6600;
wire n_817;
wire n_14140;
wire n_5402;
wire n_10696;
wire n_7355;
wire n_18688;
wire n_9331;
wire n_10170;
wire n_6031;
wire n_14479;
wire n_20183;
wire n_8331;
wire n_3216;
wire n_332;
wire n_19883;
wire n_1882;
wire n_18109;
wire n_14172;
wire n_7270;
wire n_591;
wire n_18721;
wire n_5417;
wire n_6967;
wire n_19241;
wire n_18117;
wire n_6742;
wire n_13525;
wire n_4923;
wire n_2400;
wire n_5864;
wire n_14997;
wire n_15931;
wire n_6691;
wire n_14799;
wire n_10689;
wire n_13909;
wire n_6172;
wire n_19062;
wire n_12634;
wire n_14774;
wire n_12680;
wire n_11613;
wire n_10233;
wire n_751;
wire n_19721;
wire n_15492;
wire n_18443;
wire n_17343;
wire n_4652;
wire n_10810;
wire n_12176;
wire n_10311;
wire n_9140;
wire n_2163;
wire n_18533;
wire n_2815;
wire n_19427;
wire n_4577;
wire n_4748;
wire n_337;
wire n_5814;
wire n_12094;
wire n_3231;
wire n_9736;
wire n_2979;
wire n_5531;
wire n_12517;
wire n_6517;
wire n_18431;
wire n_15441;
wire n_9225;
wire n_17353;
wire n_2946;
wire n_11923;
wire n_12071;
wire n_13832;
wire n_3430;
wire n_2269;
wire n_8105;
wire n_9031;
wire n_4225;
wire n_19406;
wire n_13087;
wire n_13972;
wire n_15436;
wire n_17920;
wire n_15633;
wire n_19937;
wire n_2565;
wire n_12339;
wire n_10602;
wire n_16630;
wire n_14632;
wire n_5655;
wire n_6393;
wire n_15969;
wire n_8154;
wire n_2175;
wire n_2182;
wire n_13849;
wire n_11131;
wire n_10778;
wire n_17961;
wire n_19912;
wire n_13258;
wire n_1506;
wire n_3473;
wire n_957;
wire n_1994;
wire n_13166;
wire n_9014;
wire n_8509;
wire n_6364;
wire n_16754;
wire n_15482;
wire n_16217;
wire n_19467;
wire n_11003;
wire n_6061;
wire n_18132;
wire n_12723;
wire n_19762;
wire n_14097;
wire n_18741;
wire n_19973;
wire n_2685;
wire n_8372;
wire n_17042;
wire n_10088;
wire n_20552;
wire n_14887;
wire n_7225;
wire n_8077;
wire n_18530;
wire n_20341;
wire n_16948;
wire n_6755;
wire n_18934;
wire n_2265;
wire n_13762;
wire n_13037;
wire n_11573;
wire n_4409;
wire n_7509;
wire n_10145;
wire n_14225;
wire n_11005;
wire n_4629;
wire n_6255;
wire n_18611;
wire n_19903;
wire n_4638;
wire n_6840;
wire n_17675;
wire n_8423;
wire n_9577;
wire n_19149;
wire n_12589;
wire n_14143;
wire n_6488;
wire n_904;
wire n_8337;
wire n_709;
wire n_7164;
wire n_14044;
wire n_17431;
wire n_3868;
wire n_18249;
wire n_18561;
wire n_18134;
wire n_17000;
wire n_12699;
wire n_1085;
wire n_12927;
wire n_2042;
wire n_16588;
wire n_771;
wire n_8199;
wire n_17456;
wire n_1149;
wire n_8656;
wire n_265;
wire n_14909;
wire n_10918;
wire n_13122;
wire n_2592;
wire n_15553;
wire n_2666;
wire n_1585;
wire n_12663;
wire n_1799;
wire n_2564;
wire n_16349;
wire n_17165;
wire n_20125;
wire n_15841;
wire n_17623;
wire n_4259;
wire n_2035;
wire n_11127;
wire n_18083;
wire n_7134;
wire n_4572;
wire n_9547;
wire n_4104;
wire n_16350;
wire n_8346;
wire n_8761;
wire n_15458;
wire n_9085;
wire n_13734;
wire n_8226;
wire n_17532;
wire n_7079;
wire n_9084;
wire n_5928;
wire n_4089;
wire n_5478;
wire n_6016;
wire n_1144;
wire n_3219;
wire n_20365;
wire n_14051;
wire n_20078;
wire n_17680;
wire n_9889;
wire n_12556;
wire n_12375;
wire n_2010;
wire n_1198;
wire n_13723;
wire n_10168;
wire n_2174;
wire n_12156;
wire n_13128;
wire n_13490;
wire n_4727;
wire n_4594;
wire n_17663;
wire n_14913;
wire n_10621;
wire n_9731;
wire n_6572;
wire n_4429;
wire n_9604;
wire n_7962;
wire n_15382;
wire n_4051;
wire n_20466;
wire n_7755;
wire n_16031;
wire n_6080;
wire n_4865;
wire n_8387;
wire n_12076;
wire n_10613;
wire n_6717;
wire n_7473;
wire n_20464;
wire n_11359;
wire n_19404;
wire n_19064;
wire n_15997;
wire n_19562;
wire n_10561;
wire n_19335;
wire n_14695;
wire n_16251;
wire n_13212;
wire n_16978;
wire n_15166;
wire n_18304;
wire n_15138;
wire n_16516;
wire n_18517;
wire n_2879;
wire n_17533;
wire n_14405;
wire n_967;
wire n_7038;
wire n_14081;
wire n_4341;
wire n_1819;
wire n_8177;
wire n_17616;
wire n_12025;
wire n_8962;
wire n_9538;
wire n_14254;
wire n_16137;
wire n_6145;
wire n_6539;
wire n_6926;
wire n_13421;
wire n_1632;
wire n_13495;
wire n_13474;
wire n_14903;
wire n_13949;
wire n_12383;
wire n_11912;
wire n_4973;
wire n_14967;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3950;
wire n_9423;
wire n_16619;
wire n_2927;
wire n_20550;
wire n_4750;
wire n_12962;
wire n_18823;
wire n_16263;
wire n_11666;
wire n_12459;
wire n_2166;
wire n_2899;
wire n_7105;
wire n_14500;
wire n_13568;
wire n_10140;
wire n_12612;
wire n_16369;
wire n_5903;
wire n_17213;
wire n_5986;
wire n_3065;
wire n_6710;
wire n_1423;
wire n_19745;
wire n_18326;
wire n_19402;
wire n_17664;
wire n_4959;
wire n_9056;
wire n_4426;
wire n_12496;
wire n_12814;
wire n_3002;
wire n_649;
wire n_15943;
wire n_18714;
wire n_11921;
wire n_8495;
wire n_14532;
wire n_8783;
wire n_14557;
wire n_19805;
wire n_1199;
wire n_12603;
wire n_15392;
wire n_14340;
wire n_18444;
wire n_14032;
wire n_16944;
wire n_15702;
wire n_7262;
wire n_212;
wire n_3773;
wire n_12967;
wire n_14899;
wire n_12232;
wire n_18115;
wire n_18847;
wire n_11859;
wire n_15773;
wire n_798;
wire n_19771;
wire n_15307;
wire n_14111;
wire n_6719;
wire n_13580;
wire n_7178;
wire n_9553;
wire n_11633;
wire n_7506;
wire n_8551;
wire n_14361;
wire n_12760;
wire n_18291;
wire n_2647;
wire n_19633;
wire n_14943;
wire n_4578;
wire n_4777;
wire n_2672;
wire n_12590;
wire n_2299;
wire n_15605;
wire n_5871;
wire n_18951;
wire n_7142;
wire n_12577;
wire n_17711;
wire n_10182;
wire n_16813;
wire n_13928;
wire n_19342;
wire n_7125;
wire n_1172;
wire n_11655;
wire n_3626;
wire n_2313;
wire n_12069;
wire n_16899;
wire n_15656;
wire n_18455;
wire n_16957;
wire n_10317;
wire n_4029;
wire n_375;
wire n_12270;
wire n_4617;
wire n_16021;
wire n_9196;
wire n_4010;
wire n_1649;
wire n_5882;
wire n_19934;
wire n_5650;
wire n_6057;
wire n_14555;
wire n_10893;
wire n_1572;
wire n_5021;
wire n_9251;
wire n_9973;
wire n_11117;
wire n_8064;
wire n_8468;
wire n_4325;
wire n_3251;
wire n_10201;
wire n_2212;
wire n_12210;
wire n_8778;
wire n_17106;
wire n_14168;
wire n_5249;
wire n_2603;
wire n_2090;
wire n_15342;
wire n_15534;
wire n_10539;
wire n_14080;
wire n_5625;
wire n_11777;
wire n_17402;
wire n_4919;
wire n_3737;
wire n_13975;
wire n_5969;
wire n_10121;
wire n_8198;
wire n_19054;
wire n_6828;
wire n_5158;
wire n_7255;
wire n_12189;
wire n_1211;
wire n_9270;
wire n_14142;
wire n_6041;
wire n_9099;
wire n_7350;
wire n_10814;
wire n_5276;
wire n_16034;
wire n_9627;
wire n_17008;
wire n_16563;
wire n_6664;
wire n_196;
wire n_17575;
wire n_2985;
wire n_13131;
wire n_14941;
wire n_1446;
wire n_3938;
wire n_11154;
wire n_3507;
wire n_11700;
wire n_20428;
wire n_5855;
wire n_3531;
wire n_16128;
wire n_10975;
wire n_1054;
wire n_9460;
wire n_17698;
wire n_11652;
wire n_14320;
wire n_11056;
wire n_19229;
wire n_6238;
wire n_13932;
wire n_2397;
wire n_16804;
wire n_3931;
wire n_15606;
wire n_10459;
wire n_2113;
wire n_1918;
wire n_20501;
wire n_5429;
wire n_6545;
wire n_11583;
wire n_15866;
wire n_9766;
wire n_20041;
wire n_4163;
wire n_10463;
wire n_14764;
wire n_19897;
wire n_645;
wire n_7074;
wire n_8734;
wire n_2633;
wire n_12564;
wire n_19443;
wire n_13433;
wire n_15505;
wire n_10403;
wire n_7037;
wire n_13697;
wire n_11784;
wire n_20549;
wire n_5298;
wire n_9025;
wire n_3396;
wire n_14244;
wire n_7928;
wire n_12886;
wire n_6532;
wire n_821;
wire n_4372;
wire n_7293;
wire n_18638;
wire n_13000;
wire n_14362;
wire n_5640;
wire n_15996;
wire n_408;
wire n_4318;
wire n_6721;
wire n_18825;
wire n_2123;
wire n_3716;
wire n_6108;
wire n_10370;
wire n_8258;
wire n_18537;
wire n_9597;
wire n_11892;
wire n_5744;
wire n_5384;
wire n_3248;
wire n_15731;
wire n_19909;
wire n_8299;
wire n_12473;
wire n_4032;
wire n_1064;
wire n_11421;
wire n_1396;
wire n_18704;
wire n_11966;
wire n_19530;
wire n_17450;
wire n_18011;
wire n_12748;
wire n_4337;
wire n_16829;
wire n_3092;
wire n_9692;
wire n_7395;
wire n_13402;
wire n_3734;
wire n_17305;
wire n_18047;
wire n_7078;
wire n_8188;
wire n_2580;
wire n_13831;
wire n_16792;
wire n_18572;
wire n_11423;
wire n_1875;
wire n_1865;
wire n_5701;
wire n_18378;
wire n_20211;
wire n_9567;
wire n_9061;
wire n_3419;
wire n_1297;
wire n_17154;
wire n_16922;
wire n_8664;
wire n_922;
wire n_16552;
wire n_16867;
wire n_16638;
wire n_14783;
wire n_13268;
wire n_10740;
wire n_10457;
wire n_19042;
wire n_17968;
wire n_1896;
wire n_3058;
wire n_14158;
wire n_9701;
wire n_675;
wire n_19247;
wire n_14236;
wire n_1540;
wire n_18849;
wire n_13510;
wire n_14640;
wire n_6659;
wire n_9709;
wire n_242;
wire n_9295;
wire n_4371;
wire n_2994;
wire n_3689;
wire n_16678;
wire n_10264;
wire n_5850;
wire n_15029;
wire n_14286;
wire n_12528;
wire n_17640;
wire n_6182;
wire n_12717;
wire n_6520;
wire n_12660;
wire n_3918;
wire n_1965;
wire n_2476;
wire n_17651;
wire n_17662;
wire n_598;
wire n_11547;
wire n_19680;
wire n_20273;
wire n_13520;
wire n_19668;
wire n_20028;
wire n_8501;
wire n_10301;
wire n_3271;
wire n_295;
wire n_4248;
wire n_13018;
wire n_18240;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_15139;
wire n_8076;
wire n_6826;
wire n_1792;
wire n_11395;
wire n_9107;
wire n_19630;
wire n_3809;
wire n_11279;
wire n_18370;
wire n_11724;
wire n_20429;
wire n_11789;
wire n_14152;
wire n_3139;
wire n_14869;
wire n_19989;
wire n_19354;
wire n_881;
wire n_8014;
wire n_19030;
wire n_7768;
wire n_8638;
wire n_16294;
wire n_4018;
wire n_14651;
wire n_694;
wire n_7982;
wire n_8804;
wire n_297;
wire n_3337;
wire n_11383;
wire n_1044;
wire n_2165;
wire n_15882;
wire n_17740;
wire n_6879;
wire n_17059;
wire n_7567;
wire n_8433;
wire n_6074;
wire n_4588;
wire n_585;
wire n_10932;
wire n_10619;
wire n_1756;
wire n_5411;
wire n_17263;
wire n_9156;
wire n_16113;
wire n_16848;
wire n_1968;
wire n_4728;
wire n_4385;
wire n_18749;
wire n_20082;
wire n_10248;
wire n_9748;
wire n_3616;
wire n_13365;
wire n_7771;
wire n_11780;
wire n_5695;
wire n_6027;
wire n_2870;
wire n_16289;
wire n_2151;
wire n_7701;
wire n_16342;
wire n_1839;
wire n_17278;
wire n_5235;
wire n_6720;
wire n_11930;
wire n_6888;
wire n_826;
wire n_3747;
wire n_12628;
wire n_8122;
wire n_17095;
wire n_13444;
wire n_16504;
wire n_8432;
wire n_4330;
wire n_7592;
wire n_14209;
wire n_20305;
wire n_19462;
wire n_18651;
wire n_5311;
wire n_6590;
wire n_3522;
wire n_2747;
wire n_18243;
wire n_791;
wire n_11876;
wire n_5572;
wire n_19110;
wire n_7151;
wire n_8950;
wire n_18683;
wire n_10758;
wire n_2861;
wire n_13431;
wire n_3975;
wire n_1838;
wire n_4683;
wire n_12538;
wire n_14025;
wire n_7758;
wire n_13779;
wire n_12446;
wire n_2316;
wire n_15954;
wire n_9355;
wire n_5060;
wire n_15386;
wire n_4986;
wire n_14620;
wire n_5888;
wire n_15349;
wire n_9582;
wire n_2208;
wire n_5884;
wire n_11009;
wire n_9288;
wire n_6308;
wire n_7897;
wire n_17701;
wire n_7118;
wire n_2134;
wire n_8284;
wire n_9702;
wire n_18767;
wire n_15378;
wire n_7422;
wire n_1431;
wire n_17881;
wire n_3835;
wire n_6738;
wire n_12307;
wire n_8703;
wire n_15839;
wire n_16135;
wire n_17661;
wire n_14999;
wire n_2771;
wire n_3020;
wire n_5264;
wire n_19377;
wire n_3557;
wire n_2610;
wire n_3620;
wire n_13720;
wire n_478;
wire n_7339;
wire n_3832;
wire n_13706;
wire n_13903;
wire n_9051;
wire n_3693;
wire n_8545;
wire n_10385;
wire n_10105;
wire n_2372;
wire n_1490;
wire n_15785;
wire n_20530;
wire n_19056;
wire n_3674;
wire n_2959;
wire n_17114;
wire n_10251;
wire n_15234;
wire n_293;
wire n_18796;
wire n_1070;
wire n_2403;
wire n_4700;
wire n_17524;
wire n_9980;
wire n_14394;
wire n_20098;
wire n_4224;
wire n_18679;
wire n_6005;
wire n_17261;
wire n_9555;
wire n_14845;
wire n_19906;
wire n_1358;
wire n_7713;
wire n_4564;
wire n_15372;
wire n_13560;
wire n_15700;
wire n_16182;
wire n_2424;
wire n_3201;
wire n_19239;
wire n_1475;
wire n_10304;
wire n_3103;
wire n_5860;
wire n_6936;
wire n_15934;
wire n_16827;
wire n_16121;
wire n_7487;
wire n_9986;
wire n_527;
wire n_13794;
wire n_3627;
wire n_13537;
wire n_9397;
wire n_18616;
wire n_1137;
wire n_3612;
wire n_17574;
wire n_4695;
wire n_9855;
wire n_10568;
wire n_2966;
wire n_2294;
wire n_13463;
wire n_600;
wire n_9496;
wire n_16241;
wire n_10796;
wire n_10016;
wire n_10030;
wire n_12864;
wire n_9653;
wire n_10272;
wire n_8989;
wire n_9640;
wire n_1339;
wire n_13936;
wire n_13933;
wire n_7815;
wire n_403;
wire n_7934;
wire n_3244;
wire n_11578;
wire n_6865;
wire n_1141;
wire n_7276;
wire n_18595;
wire n_1755;
wire n_5043;
wire n_17078;
wire n_8739;
wire n_6747;
wire n_13714;
wire n_2025;
wire n_12725;
wire n_6640;
wire n_16030;
wire n_2250;
wire n_3033;
wire n_16079;
wire n_11908;
wire n_18166;
wire n_6462;
wire n_17372;
wire n_6034;
wire n_9781;
wire n_13159;
wire n_418;
wire n_14788;
wire n_13287;
wire n_11913;
wire n_7034;
wire n_1618;
wire n_4867;
wire n_13389;
wire n_17726;
wire n_1653;
wire n_9906;
wire n_4237;
wire n_5029;
wire n_12317;
wire n_13302;
wire n_10092;
wire n_6833;
wire n_6793;
wire n_16766;
wire n_17834;
wire n_11815;
wire n_6295;
wire n_3386;
wire n_11231;
wire n_463;
wire n_13740;
wire n_17966;
wire n_19278;
wire n_19926;
wire n_8137;
wire n_12027;
wire n_3205;
wire n_15218;
wire n_17366;
wire n_19114;
wire n_17514;
wire n_17975;
wire n_7014;
wire n_10430;
wire n_16697;
wire n_8305;
wire n_18147;
wire n_1636;
wire n_4001;
wire n_18751;
wire n_6709;
wire n_17525;
wire n_960;
wire n_6712;
wire n_7416;
wire n_778;
wire n_14553;
wire n_5177;
wire n_9657;
wire n_16594;
wire n_16370;
wire n_6743;
wire n_16223;
wire n_1610;
wire n_12412;
wire n_11880;
wire n_5785;
wire n_14528;
wire n_20150;
wire n_4583;
wire n_9485;
wire n_13940;
wire n_2515;
wire n_11249;
wire n_15449;
wire n_4054;
wire n_10119;
wire n_11986;
wire n_14798;
wire n_5966;
wire n_3349;
wire n_17579;
wire n_368;
wire n_12118;
wire n_14409;
wire n_14724;
wire n_18451;
wire n_14291;
wire n_1020;
wire n_8625;
wire n_4214;
wire n_6919;
wire n_13756;
wire n_7805;
wire n_10995;
wire n_19957;
wire n_9192;
wire n_1138;
wire n_5752;
wire n_11618;
wire n_14266;
wire n_12594;
wire n_8179;
wire n_19360;
wire n_11861;
wire n_8511;
wire n_6973;
wire n_12081;
wire n_4413;
wire n_7453;
wire n_10684;
wire n_2381;
wire n_18095;
wire n_2052;
wire n_5081;
wire n_15039;
wire n_17929;
wire n_17027;
wire n_8806;
wire n_17400;
wire n_6619;
wire n_19234;
wire n_16434;
wire n_5189;
wire n_20405;
wire n_13930;
wire n_8149;
wire n_3041;
wire n_603;
wire n_10390;
wire n_1657;
wire n_20073;
wire n_7210;
wire n_5869;
wire n_2439;
wire n_2404;
wire n_6718;
wire n_4238;
wire n_3011;
wire n_15400;
wire n_2061;
wire n_17411;
wire n_16866;
wire n_15485;
wire n_18499;
wire n_18789;
wire n_14841;
wire n_16726;
wire n_13624;
wire n_5632;
wire n_5425;
wire n_18603;
wire n_19480;
wire n_8269;
wire n_13805;
wire n_18786;
wire n_3650;
wire n_8968;
wire n_16243;
wire n_7855;
wire n_14029;
wire n_4590;
wire n_3137;
wire n_14056;
wire n_5678;
wire n_13695;
wire n_6981;
wire n_13288;
wire n_19465;
wire n_16917;
wire n_3238;
wire n_218;
wire n_11519;
wire n_13065;
wire n_11229;
wire n_18655;
wire n_16159;
wire n_17570;
wire n_11397;
wire n_12840;
wire n_5437;
wire n_12846;
wire n_14705;
wire n_17660;
wire n_8401;
wire n_7854;
wire n_10577;
wire n_11324;
wire n_12945;
wire n_5307;
wire n_17385;
wire n_10151;
wire n_6439;
wire n_2446;
wire n_8240;
wire n_12850;
wire n_7714;
wire n_16193;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_9305;
wire n_9999;
wire n_17495;
wire n_1121;
wire n_11361;
wire n_1963;
wire n_6945;
wire n_18617;
wire n_3790;
wire n_7029;
wire n_19009;
wire n_20180;
wire n_10186;
wire n_17236;
wire n_11841;
wire n_6618;
wire n_14453;
wire n_19824;
wire n_19882;
wire n_20389;
wire n_17545;
wire n_13094;
wire n_7317;
wire n_17558;
wire n_3977;
wire n_227;
wire n_9461;
wire n_6816;
wire n_10928;
wire n_5008;
wire n_6502;
wire n_6250;
wire n_6288;
wire n_5974;
wire n_7522;
wire n_4133;
wire n_9618;
wire n_6118;
wire n_18961;
wire n_4561;
wire n_464;
wire n_19772;
wire n_11808;
wire n_17970;
wire n_13257;
wire n_17160;
wire n_18778;
wire n_4239;
wire n_18509;
wire n_4184;
wire n_17636;
wire n_1830;
wire n_13393;
wire n_6251;
wire n_9828;
wire n_3915;
wire n_13922;
wire n_13423;
wire n_18149;
wire n_2835;
wire n_5243;
wire n_1416;
wire n_2293;
wire n_10252;
wire n_16641;
wire n_11555;
wire n_6869;
wire n_3102;
wire n_14625;
wire n_10345;
wire n_2026;
wire n_10059;
wire n_8325;
wire n_7621;
wire n_7359;
wire n_550;
wire n_3321;
wire n_2322;
wire n_12394;
wire n_4782;
wire n_13578;
wire n_19540;
wire n_14204;
wire n_9005;
wire n_4378;
wire n_8274;
wire n_12954;
wire n_4876;
wire n_19703;
wire n_6146;
wire n_8504;
wire n_10464;
wire n_14688;
wire n_10644;
wire n_12801;
wire n_18594;
wire n_13708;
wire n_10365;
wire n_11781;
wire n_20312;
wire n_9648;
wire n_2653;
wire n_12965;
wire n_12788;
wire n_9498;
wire n_15707;
wire n_16328;
wire n_3156;
wire n_20127;
wire n_15396;
wire n_19804;
wire n_15909;
wire n_672;
wire n_3483;
wire n_11884;
wire n_20146;
wire n_19516;
wire n_19734;
wire n_13371;
wire n_4493;
wire n_7971;
wire n_743;
wire n_12264;
wire n_8232;
wire n_9649;
wire n_8904;
wire n_16977;
wire n_19287;
wire n_10629;
wire n_660;
wire n_7070;
wire n_8382;
wire n_4421;
wire n_18950;
wire n_2839;
wire n_4793;
wire n_13856;
wire n_15607;
wire n_15879;
wire n_7259;
wire n_12274;
wire n_14588;
wire n_2944;
wire n_8128;
wire n_15746;
wire n_19985;
wire n_3831;
wire n_15921;
wire n_19545;
wire n_5932;
wire n_5830;
wire n_11345;
wire n_12380;
wire n_13245;
wire n_12586;
wire n_3391;
wire n_8794;
wire n_11760;
wire n_19203;
wire n_1463;
wire n_4505;
wire n_17222;
wire n_1826;
wire n_20505;
wire n_5126;
wire n_8205;
wire n_9907;
wire n_19887;
wire n_13088;
wire n_6976;
wire n_13538;
wire n_11024;
wire n_18437;
wire n_6304;
wire n_5236;
wire n_7640;
wire n_13701;
wire n_10498;
wire n_11424;
wire n_12585;
wire n_5012;
wire n_14021;
wire n_1256;
wire n_10635;
wire n_13626;
wire n_20403;
wire n_19218;
wire n_12832;
wire n_8067;
wire n_12301;
wire n_9643;
wire n_4630;
wire n_18973;
wire n_18402;
wire n_15822;
wire n_11881;
wire n_14980;
wire n_2109;
wire n_7727;
wire n_18968;
wire n_11935;
wire n_17561;
wire n_18766;
wire n_1204;
wire n_18901;
wire n_233;
wire n_8719;
wire n_16140;
wire n_19223;
wire n_18046;
wire n_2787;
wire n_15493;
wire n_12615;
wire n_13357;
wire n_10802;
wire n_17148;
wire n_769;
wire n_4786;
wire n_7565;
wire n_16624;
wire n_20225;
wire n_7631;
wire n_13869;
wire n_16903;
wire n_7387;
wire n_9212;
wire n_12167;
wire n_9473;
wire n_13026;
wire n_10490;
wire n_15019;
wire n_13499;
wire n_17107;
wire n_14843;
wire n_2736;
wire n_10647;
wire n_3493;
wire n_9320;
wire n_10523;
wire n_16781;
wire n_19738;
wire n_12298;
wire n_10081;
wire n_3774;
wire n_12569;
wire n_2910;
wire n_14929;
wire n_18497;
wire n_5148;
wire n_20288;
wire n_2584;
wire n_866;
wire n_12456;
wire n_8655;
wire n_17039;
wire n_10808;
wire n_6333;
wire n_8745;
wire n_5791;
wire n_18504;
wire n_8086;
wire n_15466;
wire n_13943;
wire n_17124;
wire n_7379;
wire n_17530;
wire n_8901;
wire n_11078;
wire n_8695;
wire n_4911;
wire n_8173;
wire n_12072;
wire n_4436;
wire n_10545;
wire n_1174;
wire n_17945;
wire n_16557;
wire n_20093;
wire n_14141;
wire n_5602;
wire n_647;
wire n_9379;
wire n_11992;
wire n_15790;
wire n_844;
wire n_17061;
wire n_14880;
wire n_13142;
wire n_13180;
wire n_3584;
wire n_10453;
wire n_16975;
wire n_3556;
wire n_16716;
wire n_13785;
wire n_5831;
wire n_7742;
wire n_9274;
wire n_3456;
wire n_20395;
wire n_10331;
wire n_11439;
wire n_14655;
wire n_17230;
wire n_12863;
wire n_10352;
wire n_19876;
wire n_19449;
wire n_1122;
wire n_4059;
wire n_16830;
wire n_1109;
wire n_17851;
wire n_8507;
wire n_3309;
wire n_8415;
wire n_2609;
wire n_10713;
wire n_6680;
wire n_10954;
wire n_7432;
wire n_16036;
wire n_13978;
wire n_13941;
wire n_15339;
wire n_13439;
wire n_228;
wire n_16152;
wire n_14133;
wire n_14433;
wire n_13187;
wire n_13162;
wire n_2600;
wire n_7505;
wire n_18521;
wire n_15059;
wire n_8244;
wire n_18380;
wire n_7494;
wire n_4353;
wire n_735;
wire n_17071;
wire n_13661;
wire n_9546;
wire n_7589;
wire n_17764;
wire n_4346;
wire n_4351;
wire n_19969;
wire n_11296;
wire n_13770;
wire n_18636;
wire n_8723;
wire n_13511;
wire n_18016;
wire n_11019;
wire n_980;
wire n_7843;
wire n_1651;
wire n_19544;
wire n_4784;
wire n_19258;
wire n_14569;
wire n_7902;
wire n_1685;
wire n_6496;
wire n_3066;
wire n_15744;
wire n_7756;
wire n_2844;
wire n_15557;
wire n_18244;
wire n_8940;
wire n_8342;
wire n_14154;
wire n_8472;
wire n_4332;
wire n_810;
wire n_10000;
wire n_12812;
wire n_7988;
wire n_14174;
wire n_7500;
wire n_10246;
wire n_3198;
wire n_18236;
wire n_14269;
wire n_9822;
wire n_13991;
wire n_17523;
wire n_14821;
wire n_17330;
wire n_15096;
wire n_5272;
wire n_14992;
wire n_10125;
wire n_9065;
wire n_16637;
wire n_3218;
wire n_18627;
wire n_9086;
wire n_9153;
wire n_10505;
wire n_582;
wire n_861;
wire n_11064;
wire n_6908;
wire n_8237;
wire n_9093;
wire n_19046;
wire n_2968;
wire n_4201;
wire n_7266;
wire n_17928;
wire n_8046;
wire n_5646;
wire n_13284;
wire n_4852;
wire n_4210;
wire n_16521;
wire n_2709;
wire n_9198;
wire n_20580;
wire n_8335;
wire n_9142;
wire n_17697;
wire n_15820;
wire n_18239;
wire n_5214;
wire n_15486;
wire n_9493;
wire n_19371;
wire n_11330;
wire n_12720;
wire n_7794;
wire n_19139;
wire n_20431;
wire n_13318;
wire n_15917;
wire n_1274;
wire n_3333;
wire n_6605;
wire n_19748;
wire n_12687;
wire n_18278;
wire n_17510;
wire n_19106;
wire n_13208;
wire n_13867;
wire n_15594;
wire n_17807;
wire n_17841;
wire n_5380;
wire n_5776;
wire n_11796;
wire n_18339;
wire n_16881;
wire n_12789;
wire n_2677;
wire n_12127;
wire n_17232;
wire n_3283;
wire n_16976;
wire n_8037;
wire n_14119;
wire n_13673;
wire n_1742;
wire n_16775;
wire n_12573;
wire n_2542;
wire n_1671;
wire n_19400;
wire n_15214;
wire n_13045;
wire n_741;
wire n_1351;
wire n_19913;
wire n_17347;
wire n_18684;
wire n_6806;
wire n_13146;
wire n_13235;
wire n_15125;
wire n_5019;
wire n_2332;
wire n_5138;
wire n_4388;
wire n_6960;
wire n_3089;
wire n_8169;
wire n_12265;
wire n_783;
wire n_5409;
wire n_5301;
wire n_17777;
wire n_188;
wire n_1854;
wire n_3222;
wire n_7504;
wire n_15971;
wire n_442;
wire n_11678;
wire n_19814;
wire n_8023;
wire n_12251;
wire n_1975;
wire n_16307;
wire n_8130;
wire n_16911;
wire n_15294;
wire n_5055;
wire n_18676;
wire n_16288;
wire n_7116;
wire n_4249;
wire n_17992;
wire n_6999;
wire n_14741;
wire n_20436;
wire n_11046;
wire n_11079;
wire n_5548;
wire n_15581;
wire n_11065;
wire n_8339;
wire n_19058;
wire n_14215;
wire n_20290;
wire n_17368;
wire n_852;
wire n_544;
wire n_5900;
wire n_4273;
wire n_18104;
wire n_8499;
wire n_15356;
wire n_18525;
wire n_6882;
wire n_10775;
wire n_2129;
wire n_9526;
wire n_17511;
wire n_18762;
wire n_15571;
wire n_7983;
wire n_10863;
wire n_4997;
wire n_2399;
wire n_4843;
wire n_1232;
wire n_17138;
wire n_17700;
wire n_13993;
wire n_10986;
wire n_8366;
wire n_8102;
wire n_19126;
wire n_18087;
wire n_8022;
wire n_17226;
wire n_19212;
wire n_10262;
wire n_5239;
wire n_1781;
wire n_10239;
wire n_14577;
wire n_5332;
wire n_14984;
wire n_20514;
wire n_2004;
wire n_1106;
wire n_18183;
wire n_8913;
wire n_155;
wire n_4956;
wire n_16772;
wire n_14699;
wire n_454;
wire n_20074;
wire n_10335;
wire n_15362;
wire n_5129;
wire n_11301;
wire n_15101;
wire n_5070;
wire n_18154;
wire n_11703;
wire n_6374;
wire n_17013;
wire n_6628;
wire n_13483;
wire n_18923;
wire n_4262;
wire n_16551;
wire n_17803;
wire n_1894;
wire n_6570;
wire n_20358;
wire n_8556;
wire n_8040;
wire n_11821;
wire n_13121;
wire n_13989;
wire n_10755;
wire n_16998;
wire n_15200;
wire n_17349;
wire n_10682;
wire n_3928;
wire n_6371;
wire n_8079;
wire n_2613;
wire n_3535;
wire n_8595;
wire n_2708;
wire n_1648;
wire n_2011;
wire n_5684;
wire n_15887;
wire n_10022;
wire n_5729;
wire n_13803;
wire n_14066;
wire n_7856;
wire n_564;
wire n_6148;
wire n_7625;
wire n_686;
wire n_1641;
wire n_3871;
wire n_12775;
wire n_6989;
wire n_7863;
wire n_8958;
wire n_12833;
wire n_5099;
wire n_12090;
wire n_6896;
wire n_13687;
wire n_19852;
wire n_7623;
wire n_7217;
wire n_1699;
wire n_14540;
wire n_16784;
wire n_8115;
wire n_608;
wire n_2101;
wire n_9398;
wire n_15320;
wire n_3484;
wire n_4677;
wire n_12915;
wire n_6196;
wire n_13149;
wire n_18748;
wire n_2616;
wire n_5275;
wire n_14091;
wire n_15755;
wire n_8412;
wire n_2811;
wire n_6485;
wire n_14478;
wire n_17848;
wire n_10177;
wire n_6107;
wire n_16689;
wire n_11944;
wire n_1075;
wire n_7796;
wire n_6994;
wire n_15986;
wire n_14570;
wire n_16068;
wire n_13797;
wire n_13013;
wire n_13238;
wire n_4810;
wire n_175;
wire n_9446;
wire n_11129;
wire n_7234;
wire n_3914;
wire n_10296;
wire n_8119;
wire n_8641;
wire n_12988;
wire n_17136;
wire n_20524;
wire n_13344;
wire n_11139;
wire n_17766;
wire n_8436;
wire n_12685;
wire n_14239;
wire n_8659;
wire n_14045;
wire n_19575;
wire n_4369;
wire n_7849;
wire n_12667;
wire n_18747;
wire n_15635;
wire n_4331;
wire n_7297;
wire n_10018;
wire n_15183;
wire n_4972;
wire n_4993;
wire n_7298;
wire n_15118;
wire n_5536;
wire n_10141;
wire n_9129;
wire n_14162;
wire n_8224;
wire n_20522;
wire n_2678;
wire n_15679;
wire n_4613;
wire n_13014;
wire n_19744;
wire n_1167;
wire n_2428;
wire n_10897;
wire n_210;
wire n_10449;
wire n_7861;
wire n_14303;
wire n_7039;
wire n_11349;
wire n_5046;
wire n_2749;
wire n_3273;
wire n_7077;
wire n_12540;
wire n_19160;
wire n_5305;
wire n_4681;
wire n_13239;
wire n_15942;
wire n_17583;
wire n_4752;
wire n_18552;
wire n_9143;
wire n_8287;
wire n_2092;
wire n_19967;
wire n_7950;
wire n_8607;
wire n_2514;
wire n_604;
wire n_17032;
wire n_6248;
wire n_16768;
wire n_16134;
wire n_20149;
wire n_10452;
wire n_7806;
wire n_3942;
wire n_15928;
wire n_16092;
wire n_7595;
wire n_8066;
wire n_5795;
wire n_12349;
wire n_14282;
wire n_5552;
wire n_6715;
wire n_6714;
wire n_11308;
wire n_890;
wire n_16266;
wire n_8416;
wire n_4518;
wire n_20070;
wire n_14167;
wire n_9113;
wire n_7149;
wire n_5291;
wire n_10363;
wire n_2252;
wire n_13623;
wire n_11511;
wire n_15833;
wire n_16046;
wire n_760;
wire n_9393;
wire n_15974;
wire n_13845;
wire n_12709;
wire n_13432;
wire n_12771;
wire n_17760;
wire n_20523;
wire n_1858;
wire n_14787;
wire n_19502;
wire n_7303;
wire n_3021;
wire n_6616;
wire n_17100;
wire n_10781;
wire n_7315;
wire n_9886;
wire n_1164;
wire n_13244;
wire n_4288;
wire n_18969;
wire n_6185;
wire n_5529;
wire n_3733;
wire n_10943;
wire n_12344;
wire n_6042;
wire n_13843;
wire n_17191;
wire n_13404;
wire n_3614;
wire n_874;
wire n_382;
wire n_5183;
wire n_18689;
wire n_7268;
wire n_4228;
wire n_3423;
wire n_10094;
wire n_16295;
wire n_10084;
wire n_19259;
wire n_13870;
wire n_13791;
wire n_3644;
wire n_6955;
wire n_2706;
wire n_1127;
wire n_1512;
wire n_9932;
wire n_16745;
wire n_320;
wire n_13900;
wire n_16224;
wire n_14652;
wire n_1139;
wire n_3179;
wire n_8741;
wire n_4000;
wire n_2897;
wire n_3970;
wire n_7232;
wire n_7377;
wire n_19461;
wire n_996;
wire n_16132;
wire n_19425;
wire n_6646;
wire n_19789;
wire n_15149;
wire n_14844;
wire n_16907;
wire n_14391;
wire n_6033;
wire n_11541;
wire n_15495;
wire n_4873;
wire n_9801;
wire n_19312;
wire n_3782;
wire n_8773;
wire n_6369;
wire n_19837;
wire n_8394;
wire n_3470;
wire n_11155;
wire n_581;
wire n_7542;
wire n_5636;
wire n_13213;
wire n_12231;
wire n_989;
wire n_17643;
wire n_8410;
wire n_14756;
wire n_18144;
wire n_7739;
wire n_4939;
wire n_19474;
wire n_14384;
wire n_15905;
wire n_5530;
wire n_2473;
wire n_12552;
wire n_11069;
wire n_2539;
wire n_4123;
wire n_9941;
wire n_16795;
wire n_5595;
wire n_20282;
wire n_17131;
wire n_3119;
wire n_3735;
wire n_11369;
wire n_4379;
wire n_14210;
wire n_486;
wire n_5388;
wire n_4718;
wire n_15788;
wire n_13362;
wire n_5962;
wire n_7010;
wire n_648;
wire n_9728;
wire n_16690;
wire n_20111;
wire n_2057;
wire n_7219;
wire n_9662;
wire n_12896;
wire n_15694;
wire n_8774;
wire n_18690;
wire n_19494;
wire n_7299;
wire n_4872;
wire n_9936;
wire n_6195;
wire n_9530;
wire n_14692;
wire n_7471;
wire n_15488;
wire n_10455;
wire n_5300;
wire n_11393;
wire n_7741;
wire n_5035;
wire n_9466;
wire n_16525;
wire n_7790;
wire n_16315;
wire n_19283;
wire n_6149;
wire n_17918;
wire n_7002;
wire n_12428;
wire n_3025;
wire n_1626;
wire n_15814;
wire n_1388;
wire n_10265;
wire n_16676;
wire n_18736;
wire n_15756;
wire n_19495;
wire n_2296;
wire n_3633;
wire n_5352;
wire n_11995;
wire n_14378;
wire n_18299;
wire n_11371;
wire n_5394;
wire n_14191;
wire n_19267;
wire n_16546;
wire n_18252;
wire n_17454;
wire n_16144;
wire n_16669;
wire n_474;
wire n_6902;
wire n_3331;
wire n_10100;
wire n_18607;
wire n_5741;
wire n_15743;
wire n_2773;
wire n_7478;
wire n_19587;
wire n_19130;
wire n_5405;
wire n_7456;
wire n_13600;
wire n_964;
wire n_8503;
wire n_4756;
wire n_8196;
wire n_16062;
wire n_17712;
wire n_9787;
wire n_10846;
wire n_13363;
wire n_19648;
wire n_4970;
wire n_211;
wire n_9786;
wire n_18681;
wire n_14908;
wire n_2292;
wire n_12908;
wire n_18692;
wire n_3441;
wire n_17168;
wire n_2416;
wire n_311;
wire n_14201;
wire n_8923;
wire n_13315;
wire n_18900;
wire n_6736;
wire n_19231;
wire n_1769;
wire n_14597;
wire n_15663;
wire n_3605;
wire n_4633;
wire n_3306;
wire n_9115;
wire n_4584;
wire n_3090;
wire n_11833;
wire n_3724;
wire n_4276;
wire n_11897;
wire n_2990;
wire n_19675;
wire n_1773;
wire n_5001;
wire n_5176;
wire n_7443;
wire n_11285;
wire n_3323;
wire n_9977;
wire n_8051;
wire n_16719;
wire n_518;
wire n_9242;
wire n_4618;
wire n_4679;
wire n_914;
wire n_11262;
wire n_4496;
wire n_12880;
wire n_4805;
wire n_8651;
wire n_13959;
wire n_3454;
wire n_10732;
wire n_6885;
wire n_10851;
wire n_10221;
wire n_3547;
wire n_9299;
wire n_11162;
wire n_13685;
wire n_3816;
wire n_14693;
wire n_8842;
wire n_3214;
wire n_19780;
wire n_16915;
wire n_1917;
wire n_14486;
wire n_1580;
wire n_7730;
wire n_11592;
wire n_15090;
wire n_8467;
wire n_17043;
wire n_15385;
wire n_3109;
wire n_16094;
wire n_2863;
wire n_6417;
wire n_13281;
wire n_1731;
wire n_5648;
wire n_15627;
wire n_2135;
wire n_4707;
wire n_1832;
wire n_10996;
wire n_858;
wire n_8676;
wire n_9853;
wire n_13192;
wire n_7448;
wire n_17170;
wire n_19045;
wire n_410;
wire n_17351;
wire n_18060;
wire n_1594;
wire n_15048;
wire n_16393;
wire n_17135;
wire n_20292;
wire n_6199;
wire n_9823;
wire n_15739;
wire n_12937;
wire n_10698;
wire n_16891;
wire n_18118;
wire n_14665;
wire n_6726;
wire n_580;
wire n_7011;
wire n_5261;
wire n_10870;
wire n_11066;
wire n_17327;
wire n_4252;
wire n_13886;
wire n_16887;
wire n_6576;
wire n_2448;
wire n_8906;
wire n_17117;
wire n_8482;
wire n_7952;
wire n_16242;
wire n_14489;
wire n_13774;
wire n_13847;
wire n_6915;
wire n_19645;
wire n_12529;
wire n_20414;
wire n_12103;
wire n_7834;
wire n_17072;
wire n_5185;
wire n_8409;
wire n_17889;
wire n_974;
wire n_14053;
wire n_5023;
wire n_2656;
wire n_4952;
wire n_19321;
wire n_5906;
wire n_8930;
wire n_16564;
wire n_14581;
wire n_628;
wire n_18811;
wire n_1573;
wire n_7890;
wire n_3973;
wire n_11950;
wire n_6024;
wire n_12461;
wire n_485;
wire n_11415;
wire n_7265;
wire n_7986;
wire n_17809;
wire n_2024;
wire n_17900;
wire n_202;
wire n_9879;
wire n_1749;
wire n_18744;
wire n_3474;
wire n_11390;
wire n_20021;
wire n_17238;
wire n_11669;
wire n_1669;
wire n_1024;
wire n_14712;
wire n_15717;
wire n_5556;
wire n_8250;
wire n_10601;
wire n_9158;
wire n_18591;
wire n_1667;
wire n_16945;
wire n_7717;
wire n_9518;
wire n_18187;
wire n_18462;
wire n_18260;
wire n_5143;
wire n_11739;
wire n_10497;
wire n_14561;
wire n_18405;
wire n_1639;
wire n_13301;
wire n_8298;
wire n_466;
wire n_5215;
wire n_7860;
wire n_14212;
wire n_2548;
wire n_7335;
wire n_4189;
wire n_9815;
wire n_13158;
wire n_1108;
wire n_11044;
wire n_15967;
wire n_15530;
wire n_1601;
wire n_11679;
wire n_8450;
wire n_17665;
wire n_3648;
wire n_17799;
wire n_7499;
wire n_3042;
wire n_19718;
wire n_7292;
wire n_12398;
wire n_17089;
wire n_5433;
wire n_9043;
wire n_6075;
wire n_7397;
wire n_10789;
wire n_17020;
wire n_12705;
wire n_1430;
wire n_1316;
wire n_7977;
wire n_12847;
wire n_13047;
wire n_6861;
wire n_14470;
wire n_15497;
wire n_7847;
wire n_15952;
wire n_13178;
wire n_19777;
wire n_3723;
wire n_18609;
wire n_1190;
wire n_12404;
wire n_397;
wire n_11606;
wire n_19817;
wire n_5978;
wire n_11452;
wire n_15734;
wire n_6217;
wire n_20152;
wire n_5031;
wire n_10797;
wire n_7289;
wire n_17656;
wire n_14110;
wire n_14806;
wire n_1673;
wire n_7354;
wire n_18312;
wire n_13824;
wire n_3424;
wire n_239;
wire n_7960;
wire n_15620;
wire n_2326;
wire n_18053;
wire n_12912;
wire n_12211;
wire n_6115;
wire n_13377;
wire n_2120;
wire n_16493;
wire n_6048;
wire n_6416;
wire n_2964;
wire n_352;
wire n_6838;
wire n_10068;
wire n_11988;
wire n_19927;
wire n_3485;
wire n_4077;
wire n_1361;
wire n_19034;
wire n_6256;
wire n_15645;
wire n_6613;
wire n_11438;
wire n_15965;
wire n_5221;
wire n_5641;
wire n_18877;
wire n_6361;
wire n_14981;
wire n_11348;
wire n_9685;
wire n_11685;
wire n_5731;
wire n_6678;
wire n_8662;
wire n_15058;
wire n_16539;
wire n_14971;
wire n_19801;
wire n_12429;
wire n_14734;
wire n_20265;
wire n_14494;
wire n_14956;
wire n_4623;
wire n_7325;
wire n_14866;
wire n_19123;
wire n_5007;
wire n_3320;
wire n_6370;
wire n_9923;
wire n_13743;
wire n_7166;
wire n_7356;
wire n_13378;
wire n_11319;
wire n_3476;
wire n_16981;
wire n_5629;
wire n_3439;
wire n_7873;
wire n_2688;
wire n_1489;
wire n_16418;
wire n_20189;
wire n_19363;
wire n_17795;
wire n_12640;
wire n_10063;
wire n_13092;
wire n_2852;
wire n_14292;
wire n_20289;
wire n_8419;
wire n_1496;
wire n_19497;
wire n_9862;
wire n_11385;
wire n_1485;
wire n_11355;
wire n_18659;
wire n_11674;
wire n_1846;
wire n_12535;
wire n_19031;
wire n_12327;
wire n_879;
wire n_2310;
wire n_10091;
wire n_11638;
wire n_6157;
wire n_8430;
wire n_15719;
wire n_12058;
wire n_14879;
wire n_16143;
wire n_18387;
wire n_5852;
wire n_15164;
wire n_7052;
wire n_16755;
wire n_10496;
wire n_5960;
wire n_14149;
wire n_2454;
wire n_18225;
wire n_5321;
wire n_9960;
wire n_157;
wire n_4215;
wire n_10998;
wire n_19180;
wire n_7502;
wire n_1484;
wire n_14216;
wire n_16380;
wire n_3752;
wire n_7919;
wire n_20554;
wire n_10800;
wire n_17962;
wire n_7085;
wire n_1373;
wire n_12065;
wire n_3958;
wire n_13950;
wire n_18952;
wire n_5210;
wire n_13732;
wire n_16422;
wire n_14968;
wire n_10993;
wire n_15542;
wire n_14985;
wire n_15910;
wire n_20267;
wire n_17734;
wire n_14443;
wire n_1047;
wire n_3899;
wire n_16136;
wire n_14285;
wire n_1385;
wire n_9734;
wire n_7288;
wire n_16325;
wire n_16842;
wire n_17355;
wire n_20281;
wire n_4987;
wire n_10495;
wire n_9004;
wire n_834;
wire n_19981;
wire n_3818;
wire n_6610;
wire n_3124;
wire n_10612;
wire n_1741;
wire n_10260;
wire n_12285;
wire n_6750;
wire n_9150;
wire n_14508;
wire n_15092;
wire n_20259;
wire n_12683;
wire n_18535;
wire n_2614;
wire n_19691;
wire n_18457;
wire n_3694;
wire n_14566;
wire n_2937;
wire n_7869;
wire n_7165;
wire n_13386;
wire n_13846;
wire n_4376;
wire n_7683;
wire n_16437;
wire n_9587;
wire n_1076;
wire n_10671;
wire n_10193;
wire n_1377;
wire n_11718;
wire n_19333;
wire n_695;
wire n_14383;
wire n_16695;
wire n_4081;
wire n_11680;
wire n_14683;
wire n_18685;
wire n_17052;
wire n_7322;
wire n_17378;
wire n_11658;
wire n_12226;
wire n_13492;
wire n_14001;
wire n_5562;
wire n_15397;
wire n_978;
wire n_15840;
wire n_7880;
wire n_20567;
wire n_4382;
wire n_749;
wire n_16855;
wire n_19120;
wire n_16937;
wire n_2140;
wire n_9919;
wire n_12135;
wire n_19485;
wire n_5577;
wire n_568;
wire n_17092;
wire n_8829;
wire n_19308;
wire n_13381;
wire n_739;
wire n_5413;
wire n_8971;
wire n_18076;
wire n_16667;
wire n_1338;
wire n_16897;
wire n_10558;
wire n_9579;
wire n_9475;
wire n_17603;
wire n_20366;
wire n_15273;
wire n_573;
wire n_9049;
wire n_13718;
wire n_18701;
wire n_4480;
wire n_14775;
wire n_18809;
wire n_11045;
wire n_16756;
wire n_222;
wire n_11340;
wire n_16965;
wire n_7675;
wire n_11903;
wire n_13279;
wire n_20410;
wire n_19704;
wire n_13644;
wire n_20242;
wire n_13291;
wire n_742;
wire n_691;
wire n_10174;
wire n_20324;
wire n_377;
wire n_7524;
wire n_2935;
wire n_15897;
wire n_4046;
wire n_11564;
wire n_14015;
wire n_8925;
wire n_12946;
wire n_16729;
wire n_18406;
wire n_13513;
wire n_4027;
wire n_12916;
wire n_1227;
wire n_3520;
wire n_8471;
wire n_12521;
wire n_18925;
wire n_9800;
wire n_11382;
wire n_19578;
wire n_10098;
wire n_11745;
wire n_1570;
wire n_15240;
wire n_1780;
wire n_15564;
wire n_1347;
wire n_17002;
wire n_14350;
wire n_7733;
wire n_17405;
wire n_18711;
wire n_4631;
wire n_19090;
wire n_1561;
wire n_13773;
wire n_14109;
wire n_6982;
wire n_20117;
wire n_2168;
wire n_5847;
wire n_7345;
wire n_17526;
wire n_14136;
wire n_7385;
wire n_10923;
wire n_5159;
wire n_2615;
wire n_20528;
wire n_14176;
wire n_4625;
wire n_11149;
wire n_19889;
wire n_12635;
wire n_3962;
wire n_8488;
wire n_9543;
wire n_11443;
wire n_15765;
wire n_6855;
wire n_18176;
wire n_3362;
wire n_10665;
wire n_4744;
wire n_12906;
wire n_4188;
wire n_13467;
wire n_3667;
wire n_712;
wire n_18374;
wire n_18700;
wire n_7907;
wire n_5568;
wire n_6312;
wire n_11532;
wire n_2505;
wire n_9415;
wire n_4115;
wire n_14343;
wire n_18619;
wire n_9147;
wire n_470;
wire n_11209;
wire n_3680;
wire n_15918;
wire n_5723;
wire n_5918;
wire n_16212;
wire n_11790;
wire n_1972;
wire n_19189;
wire n_4491;
wire n_19444;
wire n_363;
wire n_18148;
wire n_16313;
wire n_10420;
wire n_17058;
wire n_18309;
wire n_16363;
wire n_503;
wire n_6131;
wire n_15232;
wire n_20491;
wire n_12105;
wire n_14329;
wire n_19392;
wire n_15721;
wire n_5163;
wire n_307;
wire n_10444;
wire n_3361;
wire n_11377;
wire n_3478;
wire n_8018;
wire n_18557;
wire n_7937;
wire n_9176;
wire n_20103;
wire n_7819;
wire n_10631;
wire n_7305;
wire n_6334;
wire n_16780;
wire n_3096;
wire n_2651;
wire n_8884;
wire n_5537;
wire n_19222;
wire n_1574;
wire n_20171;
wire n_253;
wire n_2918;
wire n_8751;
wire n_4307;
wire n_11864;
wire n_11006;
wire n_15018;
wire n_6617;
wire n_3552;
wire n_7511;
wire n_6533;
wire n_849;
wire n_4091;
wire n_14108;
wire n_1753;
wire n_19829;
wire n_3095;
wire n_15439;
wire n_16049;
wire n_19875;
wire n_2807;
wire n_8178;
wire n_14000;
wire n_14372;
wire n_3618;
wire n_4758;
wire n_17911;
wire n_12046;
wire n_10212;
wire n_18566;
wire n_5335;
wire n_9425;
wire n_12917;
wire n_14629;
wire n_11172;
wire n_10089;
wire n_14947;
wire n_5505;
wire n_8560;
wire n_14748;
wire n_18895;
wire n_20068;
wire n_19722;
wire n_18466;
wire n_10004;
wire n_12488;
wire n_3852;
wire n_1365;
wire n_11110;
wire n_17338;
wire n_16211;
wire n_15001;
wire n_3896;
wire n_8674;
wire n_5274;
wire n_5401;
wire n_12977;
wire n_7584;
wire n_13328;
wire n_4093;
wire n_10892;
wire n_18556;
wire n_10493;
wire n_19195;
wire n_10405;
wire n_15037;
wire n_4794;
wire n_17386;
wire n_7964;
wire n_17091;
wire n_629;
wire n_14349;
wire n_6278;
wire n_7022;
wire n_12691;
wire n_11033;
wire n_19760;
wire n_19072;
wire n_18203;
wire n_14356;
wire n_19028;
wire n_5581;
wire n_16926;
wire n_16006;
wire n_992;
wire n_12651;
wire n_19194;
wire n_16476;
wire n_7486;
wire n_6756;
wire n_16373;
wire n_18792;
wire n_14190;
wire n_8563;
wire n_17223;
wire n_15546;
wire n_14157;
wire n_11534;
wire n_14344;
wire n_9221;
wire n_509;
wire n_1209;
wire n_7906;
wire n_5248;
wire n_6411;
wire n_350;
wire n_10285;
wire n_4370;
wire n_14488;
wire n_11032;
wire n_2359;
wire n_13582;
wire n_142;
wire n_17950;
wire n_7302;
wire n_18162;
wire n_19725;
wire n_11174;
wire n_18574;
wire n_6381;
wire n_7030;
wire n_6656;
wire n_9730;
wire n_18544;
wire n_10294;
wire n_4359;
wire n_10106;
wire n_17865;
wire n_9934;
wire n_3487;
wire n_287;
wire n_9234;
wire n_10674;
wire n_6534;
wire n_3340;
wire n_230;
wire n_5227;
wire n_16011;
wire n_6265;
wire n_2989;
wire n_5778;
wire n_18185;
wire n_8087;
wire n_7607;
wire n_14458;
wire n_17540;
wire n_12073;
wire n_13655;
wire n_6898;
wire n_6596;
wire n_20543;
wire n_13565;
wire n_14643;
wire n_10249;
wire n_8361;
wire n_10705;
wire n_8007;
wire n_9246;
wire n_522;
wire n_18965;
wire n_3440;
wire n_13784;
wire n_13468;
wire n_2356;
wire n_12363;
wire n_18201;
wire n_7553;
wire n_1772;
wire n_1119;
wire n_6824;
wire n_19625;
wire n_5788;
wire n_11788;
wire n_2739;
wire n_12544;
wire n_20240;
wire n_13036;
wire n_20496;
wire n_14146;
wire n_13199;
wire n_20248;
wire n_6903;
wire n_2864;
wire n_13009;
wire n_1180;
wire n_10908;
wire n_10339;
wire n_9908;
wire n_9486;
wire n_13002;
wire n_13868;
wire n_7903;
wire n_18596;
wire n_11877;
wire n_8864;
wire n_7384;
wire n_18674;
wire n_13285;
wire n_20476;
wire n_8610;
wire n_19075;
wire n_7894;
wire n_11750;
wire n_3532;
wire n_7055;
wire n_18722;
wire n_8520;
wire n_16458;
wire n_13374;
wire n_12055;
wire n_381;
wire n_7639;
wire n_16520;
wire n_4327;
wire n_3765;
wire n_4125;
wire n_20231;
wire n_12811;
wire n_12186;
wire n_13032;
wire n_3067;
wire n_2155;
wire n_11001;
wire n_9512;
wire n_14199;
wire n_17858;
wire n_13684;
wire n_2364;
wire n_9170;
wire n_15108;
wire n_9616;
wire n_3803;
wire n_2085;
wire n_917;
wire n_16898;
wire n_3639;
wire n_9073;
wire n_12897;
wire n_5192;
wire n_18325;
wire n_12272;
wire n_9302;
wire n_19068;
wire n_13948;
wire n_11798;
wire n_9062;
wire n_3413;
wire n_9171;
wire n_3412;
wire n_8279;
wire n_12191;
wire n_17432;
wire n_9580;
wire n_8019;
wire n_13963;
wire n_17707;
wire n_4575;
wire n_699;
wire n_4320;
wire n_18842;
wire n_7832;
wire n_9540;
wire n_17242;
wire n_11137;
wire n_451;
wire n_8390;
wire n_8898;
wire n_14316;
wire n_5231;
wire n_2190;
wire n_8613;
wire n_3438;
wire n_18300;
wire n_8464;
wire n_15701;
wire n_6423;
wire n_1441;
wire n_15612;
wire n_3373;
wire n_18804;
wire n_7441;
wire n_513;
wire n_12112;
wire n_13060;
wire n_16187;
wire n_9449;
wire n_19787;
wire n_14817;
wire n_9050;
wire n_433;
wire n_6121;
wire n_5726;
wire n_14087;
wire n_2792;
wire n_15980;
wire n_3798;
wire n_788;
wire n_20066;
wire n_329;
wire n_14438;
wire n_2674;
wire n_4641;
wire n_16253;
wire n_7133;
wire n_12202;
wire n_13836;
wire n_1866;
wire n_8661;
wire n_2130;
wire n_7424;
wire n_3714;
wire n_19774;
wire n_16671;
wire n_12870;
wire n_11156;
wire n_10611;
wire n_10715;
wire n_12333;
wire n_8609;
wire n_17666;
wire n_17219;
wire n_13576;
wire n_7626;
wire n_2714;
wire n_2245;
wire n_7310;
wire n_17451;
wire n_12119;
wire n_12618;
wire n_16093;
wire n_1265;
wire n_17266;
wire n_20213;
wire n_15129;
wire n_17146;
wire n_16209;
wire n_14306;
wire n_8873;
wire n_11891;
wire n_16276;
wire n_199;
wire n_18427;
wire n_12401;
wire n_13055;
wire n_7323;
wire n_7301;
wire n_3715;
wire n_18600;
wire n_612;
wire n_17633;
wire n_13829;
wire n_16533;
wire n_8089;
wire n_9218;
wire n_6704;
wire n_14657;
wire n_3933;
wire n_20577;
wire n_17815;
wire n_7244;
wire n_10745;
wire n_2311;
wire n_1012;
wire n_3691;
wire n_7633;
wire n_18760;
wire n_13937;
wire n_4146;
wire n_5711;
wire n_9437;
wire n_18724;
wire n_14359;
wire n_8640;
wire n_4855;
wire n_6186;
wire n_16933;
wire n_6803;
wire n_8437;
wire n_8427;
wire n_1188;
wire n_10605;
wire n_14013;
wire n_14419;
wire n_9933;
wire n_11449;
wire n_2916;
wire n_15251;
wire n_9892;
wire n_18976;
wire n_16727;
wire n_9462;
wire n_5972;
wire n_19447;
wire n_15854;
wire n_3145;
wire n_19438;
wire n_5444;
wire n_12501;
wire n_961;
wire n_4356;
wire n_17518;
wire n_8843;
wire n_9891;
wire n_15810;
wire n_2377;
wire n_701;
wire n_10643;
wire n_16974;
wire n_3719;
wire n_4361;
wire n_10872;
wire n_13987;
wire n_15626;
wire n_1630;
wire n_4136;
wire n_13416;
wire n_12798;
wire n_14885;
wire n_2619;
wire n_5329;
wire n_9925;
wire n_16066;
wire n_9757;
wire n_10008;
wire n_13726;
wire n_507;
wire n_14412;
wire n_17587;
wire n_2271;
wire n_12243;
wire n_8562;
wire n_19714;
wire n_12614;
wire n_11378;
wire n_2606;
wire n_14631;
wire n_5728;
wire n_10032;
wire n_462;
wire n_304;
wire n_13425;
wire n_9806;
wire n_17105;
wire n_17233;
wire n_7021;
wire n_13591;
wire n_18296;
wire n_11713;
wire n_16972;
wire n_15586;
wire n_6355;
wire n_2954;
wire n_17821;
wire n_12931;
wire n_15525;
wire n_7215;
wire n_17790;
wire n_2493;
wire n_4802;
wire n_17566;
wire n_2705;
wire n_5523;
wire n_14332;
wire n_18379;
wire n_3405;
wire n_8016;
wire n_5423;
wire n_10645;
wire n_11096;
wire n_10604;
wire n_5074;
wire n_17398;
wire n_4044;
wire n_6564;
wire n_11161;
wire n_8709;
wire n_2631;
wire n_12491;
wire n_11216;
wire n_14368;
wire n_1293;
wire n_18390;
wire n_4701;
wire n_10966;
wire n_794;
wire n_727;
wire n_19310;
wire n_19871;
wire n_20110;
wire n_3385;
wire n_19650;
wire n_4851;
wire n_6442;
wire n_18359;
wire n_3293;
wire n_5204;
wire n_7925;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_15126;
wire n_4991;
wire n_19289;
wire n_20097;
wire n_5422;
wire n_6871;
wire n_16846;
wire n_9389;
wire n_1913;
wire n_12074;
wire n_8357;
wire n_6904;
wire n_10912;
wire n_5292;
wire n_19665;
wire n_12745;
wire n_9752;
wire n_14473;
wire n_12887;
wire n_18997;
wire n_10341;
wire n_19521;
wire n_4011;
wire n_15816;
wire n_18314;
wire n_7138;
wire n_17341;
wire n_4753;
wire n_8712;
wire n_631;
wire n_2262;
wire n_3611;
wire n_19254;
wire n_20363;
wire n_5059;
wire n_8837;
wire n_843;
wire n_17652;
wire n_2604;
wire n_14641;
wire n_16506;
wire n_17543;
wire n_15433;
wire n_15953;
wire n_5219;
wire n_9721;
wire n_11344;
wire n_3537;
wire n_12658;
wire n_1022;
wire n_9197;
wire n_19167;
wire n_1474;
wire n_14740;
wire n_9210;
wire n_6893;
wire n_5686;
wire n_8905;
wire n_13008;
wire n_18832;
wire n_18691;
wire n_7807;
wire n_18126;
wire n_14198;
wire n_14846;
wire n_3654;
wire n_1849;
wire n_9917;
wire n_12056;
wire n_14539;
wire n_8106;
wire n_20381;
wire n_4264;
wire n_12238;
wire n_5937;
wire n_19226;
wire n_12976;
wire n_14420;
wire n_18562;
wire n_6040;
wire n_11888;
wire n_13243;
wire n_14314;
wire n_16642;
wire n_14227;
wire n_10309;
wire n_11099;
wire n_5465;
wire n_8974;
wire n_4339;
wire n_14164;
wire n_3324;
wire n_9871;
wire n_10050;
wire n_19652;
wire n_19996;
wire n_1195;
wire n_10306;
wire n_7606;
wire n_1811;
wire n_7193;
wire n_3987;
wire n_1519;
wire n_18180;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_5721;
wire n_1048;
wire n_18142;
wire n_13632;
wire n_13020;
wire n_6012;
wire n_13148;
wire n_1418;
wire n_10429;
wire n_292;
wire n_11470;
wire n_3072;
wire n_13871;
wire n_4874;
wire n_4401;
wire n_889;
wire n_20387;
wire n_9903;
wire n_17208;
wire n_11102;
wire n_1110;
wire n_9228;
wire n_11539;
wire n_7710;
wire n_17792;
wire n_16166;
wire n_11899;
wire n_7892;
wire n_13168;
wire n_9522;
wire n_15617;
wire n_15463;
wire n_4658;
wire n_11076;
wire n_14339;
wire n_505;
wire n_1787;
wire n_16005;
wire n_6769;
wire n_9148;
wire n_11054;
wire n_2776;
wire n_10754;
wire n_5742;
wire n_3909;
wire n_9275;
wire n_10223;
wire n_1220;
wire n_8896;
wire n_19727;
wire n_7206;
wire n_5539;
wire n_6895;
wire n_13598;
wire n_2488;
wire n_17979;
wire n_10228;
wire n_1252;
wire n_511;
wire n_8758;
wire n_6026;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_8617;
wire n_17953;
wire n_13966;
wire n_12530;
wire n_1597;
wire n_9463;
wire n_4839;
wire n_2596;
wire n_1153;
wire n_13077;
wire n_16309;
wire n_10425;
wire n_8069;
wire n_6481;
wire n_19144;
wire n_4006;
wire n_15201;
wire n_9997;
wire n_6384;
wire n_13828;
wire n_7541;
wire n_6906;
wire n_14562;
wire n_9844;
wire n_12826;
wire n_8318;
wire n_10366;
wire n_15015;
wire n_19122;
wire n_7334;
wire n_5807;
wire n_20280;
wire n_16376;
wire n_2227;
wire n_5216;
wire n_14991;
wire n_10225;
wire n_4869;
wire n_6257;
wire n_4386;
wire n_20490;
wire n_20360;
wire n_8383;
wire n_12621;
wire n_4955;
wire n_11290;
wire n_17080;
wire n_12518;
wire n_19033;
wire n_3234;
wire n_14047;
wire n_9052;
wire n_856;
wire n_17447;
wire n_2830;
wire n_17678;
wire n_6587;
wire n_7781;
wire n_7360;
wire n_14568;
wire n_2181;
wire n_11702;
wire n_19395;
wire n_16970;
wire n_11372;
wire n_20424;
wire n_2826;
wire n_10817;
wire n_15324;
wire n_326;
wire n_8355;
wire n_19501;
wire n_17098;
wire n_12741;
wire n_18041;
wire n_7101;
wire n_1635;
wire n_7530;
wire n_15006;
wire n_20113;
wire n_15619;
wire n_19914;
wire n_20460;
wire n_18911;
wire n_9860;
wire n_12510;
wire n_11756;
wire n_2851;
wire n_8369;
wire n_9022;
wire n_160;
wire n_9103;
wire n_17142;
wire n_8831;
wire n_1508;
wire n_5608;
wire n_2240;
wire n_392;
wire n_12233;
wire n_8853;
wire n_4582;
wire n_6252;
wire n_18403;
wire n_6211;
wire n_15716;
wire n_5844;
wire n_17499;
wire n_1549;
wire n_17898;
wire n_17172;
wire n_8081;
wire n_16608;
wire n_17310;
wire n_13442;
wire n_1916;
wire n_14444;
wire n_18531;
wire n_10484;
wire n_11744;
wire n_17247;
wire n_10288;
wire n_18838;
wire n_10388;
wire n_6189;
wire n_20209;
wire n_15299;
wire n_4016;
wire n_11072;
wire n_621;
wire n_750;
wire n_19836;
wire n_2823;
wire n_5597;
wire n_13944;
wire n_9492;
wire n_6413;
wire n_7419;
wire n_6506;
wire n_18476;
wire n_1997;
wire n_710;
wire n_1818;
wire n_17086;
wire n_6935;
wire n_9727;
wire n_13019;
wire n_12703;
wire n_13079;
wire n_4397;
wire n_18343;
wire n_5050;
wire n_746;
wire n_3416;
wire n_3498;
wire n_15369;
wire n_15134;
wire n_16110;
wire n_2957;
wire n_1740;
wire n_19420;
wire n_9375;
wire n_17715;
wire n_5980;
wire n_8770;
wire n_3672;
wire n_15453;
wire n_5318;
wire n_6105;
wire n_6022;
wire n_10964;
wire n_3382;
wire n_19739;
wire n_12493;
wire n_13135;
wire n_8075;
wire n_5053;
wire n_7841;
wire n_9458;
wire n_20335;
wire n_8466;
wire n_6527;
wire n_15275;
wire n_19092;
wire n_8094;
wire n_4824;
wire n_2037;
wire n_4567;
wire n_6430;
wire n_782;
wire n_18268;
wire n_809;
wire n_10987;
wire n_4778;
wire n_5477;
wire n_12684;
wire n_1797;
wire n_4595;
wire n_402;
wire n_1870;
wire n_20473;
wire n_11965;
wire n_4904;
wire n_1152;
wire n_14696;
wire n_5988;
wire n_5585;
wire n_15093;
wire n_12324;
wire n_711;
wire n_3105;
wire n_14006;
wire n_6666;
wire n_3692;
wire n_8321;
wire n_20126;
wire n_19116;
wire n_9954;
wire n_8735;
wire n_1695;
wire n_11722;
wire n_2272;
wire n_2760;
wire n_972;
wire n_12310;
wire n_5348;
wire n_6594;
wire n_624;
wire n_19471;
wire n_20197;
wire n_7095;
wire n_3045;
wire n_16672;
wire n_11701;
wire n_885;
wire n_3666;
wire n_4916;
wire n_18010;
wire n_13917;
wire n_7184;
wire n_9617;
wire n_13546;
wire n_14595;
wire n_17001;
wire n_7908;
wire n_7974;
wire n_7551;
wire n_11980;
wire n_11255;
wire n_13592;
wire n_3858;
wire n_17224;
wire n_11720;
wire n_3502;
wire n_5461;
wire n_20269;
wire n_13874;
wire n_6482;
wire n_5147;
wire n_15506;
wire n_1355;
wire n_9810;
wire n_14469;
wire n_16201;
wire n_2562;
wire n_17690;
wire n_1522;
wire n_5755;
wire n_8043;
wire n_16377;
wire n_14492;
wire n_1548;
wire n_1155;
wire n_14134;
wire n_4944;
wire n_11990;
wire n_10103;
wire n_5245;
wire n_4343;
wire n_15457;
wire n_14345;
wire n_16847;
wire n_6841;
wire n_10153;
wire n_17622;
wire n_17952;
wire n_5054;
wire n_2962;
wire n_8171;
wire n_20437;
wire n_9006;
wire n_19641;
wire n_6774;
wire n_16964;
wire n_8600;
wire n_1925;
wire n_4407;
wire n_14816;
wire n_8710;
wire n_12806;
wire n_4045;
wire n_14302;
wire n_8549;
wire n_10172;
wire n_8054;
wire n_13904;
wire n_16614;
wire n_3258;
wire n_18694;
wire n_4524;
wire n_3143;
wire n_6020;
wire n_17045;
wire n_15784;
wire n_18613;
wire n_3149;
wire n_11969;
wire n_7914;
wire n_16388;
wire n_3365;
wire n_6521;
wire n_3379;
wire n_8857;
wire n_14243;
wire n_9040;
wire n_6162;
wire n_8010;
wire n_3939;
wire n_6432;
wire n_1375;
wire n_3972;
wire n_1650;
wire n_13574;
wire n_12762;
wire n_16740;
wire n_9830;
wire n_18870;
wire n_10761;
wire n_2761;
wire n_3776;
wire n_18781;
wire n_11579;
wire n_1019;
wire n_15303;
wire n_8291;
wire n_18017;
wire n_4170;
wire n_20143;
wire n_11535;
wire n_2845;
wire n_18400;
wire n_5173;
wire n_12975;
wire n_16291;
wire n_13850;
wire n_6740;
wire n_1113;
wire n_11510;
wire n_6315;
wire n_17866;
wire n_12736;
wire n_5283;
wire n_9111;
wire n_7156;
wire n_9163;
wire n_15461;
wire n_6910;
wire n_6262;
wire n_14800;
wire n_2827;
wire n_7703;
wire n_6319;
wire n_17352;
wire n_14888;
wire n_12350;
wire n_12542;
wire n_13860;
wire n_1879;
wire n_6536;
wire n_256;
wire n_6175;
wire n_7040;
wire n_8280;
wire n_12390;
wire n_367;
wire n_18898;
wire n_2569;
wire n_10235;
wire n_6978;
wire n_5351;
wire n_12805;
wire n_6093;
wire n_11649;
wire n_16306;
wire n_703;
wire n_18485;
wire n_9190;
wire n_6947;
wire n_14918;
wire n_5293;
wire n_8203;
wire n_6099;
wire n_1324;
wire n_1435;
wire n_20478;
wire n_3920;
wire n_4892;
wire n_6140;
wire n_15489;
wire n_19980;
wire n_12914;
wire n_17159;
wire n_17721;
wire n_9506;
wire n_18440;
wire n_6415;
wire n_4439;
wire n_18883;
wire n_20311;
wire n_16542;
wire n_15158;
wire n_10828;
wire n_18866;
wire n_12300;
wire n_15389;
wire n_7549;
wire n_17308;
wire n_17425;
wire n_11281;
wire n_13056;
wire n_16019;
wire n_17732;
wire n_12337;
wire n_18520;
wire n_13466;
wire n_15082;
wire n_8871;
wire n_11114;
wire n_19442;
wire n_8418;
wire n_7740;
wire n_20417;
wire n_3679;
wire n_5891;
wire n_13050;
wire n_10860;
wire n_18259;
wire n_17517;
wire n_4930;
wire n_16208;
wire n_19327;
wire n_15209;
wire n_12273;
wire n_8564;
wire n_11943;
wire n_6944;
wire n_9121;
wire n_12712;
wire n_360;
wire n_2149;
wire n_15078;
wire n_4557;
wire n_13012;
wire n_19895;
wire n_895;
wire n_8924;
wire n_20134;
wire n_20500;
wire n_12752;
wire n_6928;
wire n_4416;
wire n_10880;
wire n_15511;
wire n_4593;
wire n_4465;
wire n_3622;
wire n_19600;
wire n_18204;
wire n_20081;
wire n_4495;
wire n_14278;
wire n_5117;
wire n_12777;
wire n_14706;
wire n_8214;
wire n_5990;
wire n_20278;
wire n_20302;
wire n_7043;
wire n_11462;
wire n_11732;
wire n_5024;
wire n_4559;
wire n_18137;
wire n_12819;
wire n_10214;
wire n_8241;
wire n_838;
wire n_3336;
wire n_8442;
wire n_2952;
wire n_9572;
wire n_15282;
wire n_9229;
wire n_19505;
wire n_16812;
wire n_16038;
wire n_12237;
wire n_18350;
wire n_6134;
wire n_1656;
wire n_5803;
wire n_2112;
wire n_13372;
wire n_2430;
wire n_653;
wire n_11375;
wire n_11267;
wire n_9602;
wire n_9311;
wire n_4335;
wire n_19482;
wire n_2034;
wire n_576;
wire n_6593;
wire n_8630;
wire n_2683;
wire n_19432;
wire n_9884;
wire n_9876;
wire n_9260;
wire n_14534;
wire n_19832;
wire n_13630;
wire n_16535;
wire n_13700;
wire n_10406;
wire n_3204;
wire n_17859;
wire n_6746;
wire n_11985;
wire n_8447;
wire n_6443;
wire n_14290;
wire n_7980;
wire n_348;
wire n_8828;
wire n_18631;
wire n_17687;
wire n_19820;
wire n_390;
wire n_1148;
wire n_6749;
wire n_10965;
wire n_10798;
wire n_19657;
wire n_7732;
wire n_13325;
wire n_14850;
wire n_15135;
wire n_20338;
wire n_16196;
wire n_11911;
wire n_4265;
wire n_11442;
wire n_2950;
wire n_5634;
wire n_719;
wire n_18862;
wire n_14064;
wire n_14524;
wire n_1090;
wire n_8859;
wire n_16883;
wire n_11388;
wire n_11651;
wire n_1362;
wire n_17946;
wire n_10154;
wire n_18663;
wire n_7922;
wire n_17469;
wire n_15826;
wire n_5580;
wire n_1450;
wire n_19101;
wire n_10033;
wire n_1789;
wire n_17877;
wire n_8311;
wire n_12253;
wire n_15005;
wire n_11147;
wire n_12928;
wire n_9877;
wire n_8764;
wire n_19361;
wire n_16167;
wire n_2161;
wire n_19452;
wire n_12990;
wire n_20239;
wire n_14246;
wire n_5764;
wire n_6920;
wire n_19902;
wire n_11817;
wire n_8729;
wire n_10359;
wire n_3344;
wire n_2334;
wire n_20384;
wire n_14957;
wire n_5133;
wire n_1763;
wire n_6907;
wire n_13447;
wire n_7144;
wire n_16579;
wire n_11479;
wire n_11737;
wire n_8048;
wire n_635;
wire n_12028;
wire n_3786;
wire n_7072;
wire n_13095;
wire n_4254;
wire n_8253;
wire n_4303;
wire n_18592;
wire n_15032;
wire n_1158;
wire n_11600;
wire n_2248;
wire n_16607;
wire n_15085;
wire n_16390;
wire n_10722;
wire n_8088;
wire n_17855;
wire n_10666;
wire n_3147;
wire n_15440;
wire n_753;
wire n_3925;
wire n_3180;
wire n_8516;
wire n_8302;
wire n_17717;
wire n_20042;
wire n_15610;
wire n_359;
wire n_15329;
wire n_8167;
wire n_7859;
wire n_14315;
wire n_7872;
wire n_1479;
wire n_4768;
wire n_13858;
wire n_17913;
wire n_3717;
wire n_7480;
wire n_5410;
wire n_571;
wire n_2215;
wire n_16255;
wire n_8944;
wire n_1884;
wire n_10023;
wire n_10999;
wire n_665;
wire n_5156;
wire n_18716;
wire n_10410;
wire n_19732;
wire n_4447;
wire n_3445;
wire n_373;
wire n_16983;
wire n_8975;
wire n_1833;
wire n_17009;
wire n_19888;
wire n_11305;
wire n_17668;
wire n_9101;
wire n_15631;
wire n_14755;
wire n_8825;
wire n_12969;
wire n_1856;
wire n_12260;
wire n_12016;
wire n_8266;
wire n_5691;
wire n_8981;
wire n_4957;
wire n_17082;
wire n_165;
wire n_8771;
wire n_15750;
wire n_4039;
wire n_457;
wire n_3800;
wire n_4566;
wire n_12939;
wire n_20533;
wire n_20419;
wire n_15038;
wire n_17925;
wire n_10404;
wire n_8138;
wire n_6638;
wire n_12779;
wire n_17505;
wire n_17199;
wire n_2930;
wire n_15531;
wire n_13547;
wire n_12816;
wire n_9211;
wire n_8124;
wire n_9395;
wire n_7366;
wire n_5269;
wire n_17348;
wire n_1538;
wire n_8147;
wire n_5468;
wire n_4730;
wire n_8127;
wire n_9402;
wire n_14014;
wire n_10700;
wire n_17743;
wire n_10968;
wire n_3579;
wire n_14247;
wire n_3335;
wire n_9716;
wire n_4177;
wire n_3783;
wire n_700;
wire n_3178;
wire n_16155;
wire n_15418;
wire n_5256;
wire n_11970;
wire n_7918;
wire n_4168;
wire n_6651;
wire n_12308;
wire n_1923;
wire n_10783;
wire n_12163;
wire n_3952;
wire n_11523;
wire n_12944;
wire n_3911;
wire n_7472;
wire n_9737;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_14709;
wire n_10812;
wire n_12297;
wire n_13848;
wire n_6366;
wire n_19847;
wire n_2997;
wire n_10001;
wire n_13280;
wire n_12145;
wire n_11088;
wire n_5939;
wire n_5509;
wire n_8160;
wire n_20129;
wire n_3619;
wire n_11405;
wire n_19274;
wire n_1786;
wire n_13103;
wire n_18385;
wire n_15630;
wire n_4198;
wire n_1371;
wire n_10977;
wire n_2886;
wire n_11299;
wire n_10615;
wire n_1803;
wire n_11542;
wire n_4065;
wire n_229;
wire n_7647;
wire n_12426;
wire n_16222;
wire n_15442;
wire n_15068;
wire n_9054;
wire n_2470;
wire n_4446;
wire n_10532;
wire n_17776;
wire n_4417;
wire n_13995;
wire n_13073;
wire n_6728;
wire n_19907;
wire n_20139;
wire n_2286;
wire n_4743;
wire n_16029;
wire n_2018;
wire n_1903;
wire n_13556;
wire n_13367;
wire n_10771;
wire n_11441;
wire n_14203;
wire n_17269;
wire n_693;
wire n_1056;
wire n_19802;
wire n_12844;
wire n_5851;
wire n_7073;
wire n_9755;
wire n_5110;
wire n_10104;
wire n_772;
wire n_2806;
wire n_9117;
wire n_19426;
wire n_3028;
wire n_9381;
wire n_3076;
wire n_12049;
wire n_14498;
wire n_886;
wire n_343;
wire n_3624;
wire n_1820;
wire n_6549;
wire n_539;
wire n_19708;
wire n_20398;
wire n_6096;
wire n_7853;
wire n_12526;
wire n_2836;
wire n_8890;
wire n_16575;
wire n_7721;
wire n_7192;
wire n_19602;
wire n_20279;
wire n_11206;
wire n_11593;
wire n_15807;
wire n_3906;
wire n_11786;
wire n_12737;
wire n_4954;
wire n_17258;
wire n_15113;
wire n_9273;
wire n_2612;
wire n_8970;
wire n_16910;
wire n_2591;
wire n_1815;
wire n_10640;
wire n_2593;
wire n_10729;
wire n_14656;
wire n_20194;
wire n_16052;
wire n_20507;
wire n_14745;
wire n_20375;
wire n_19243;
wire n_4605;
wire n_7635;
wire n_19712;
wire n_11268;
wire n_17121;
wire n_14760;
wire n_20589;
wire n_3943;
wire n_11501;
wire n_7227;
wire n_13390;
wire n_8030;
wire n_6052;
wire n_8687;
wire n_13264;
wire n_5374;
wire n_12010;
wire n_1843;
wire n_9738;
wire n_12026;
wire n_4227;
wire n_521;
wire n_17481;
wire n_8633;
wire n_17645;
wire n_19999;
wire n_7689;
wire n_6511;
wire n_18470;
wire n_1309;
wire n_916;
wire n_4415;
wire n_7099;
wire n_1970;
wire n_14676;
wire n_6358;
wire n_2059;
wire n_2669;
wire n_18880;
wire n_11313;
wire n_10438;
wire n_6986;
wire n_8801;
wire n_3912;
wire n_3118;
wire n_1907;
wire n_2529;
wire n_16438;
wire n_860;
wire n_8219;
wire n_15373;
wire n_18580;
wire n_1302;
wire n_10575;
wire n_11028;
wire n_12171;
wire n_14193;
wire n_12935;
wire n_7827;
wire n_14906;
wire n_15211;
wire n_10760;
wire n_4792;
wire n_15334;
wire n_7731;
wire n_11527;
wire n_18404;
wire n_3514;
wire n_16486;
wire n_9535;
wire n_2654;
wire n_5302;
wire n_966;
wire n_12490;
wire n_3357;
wire n_692;
wire n_5781;
wire n_3895;
wire n_8486;
wire n_12829;
wire n_4118;
wire n_2176;
wire n_2459;
wire n_18662;
wire n_1111;
wire n_1251;
wire n_12739;
wire n_11610;
wire n_7132;
wire n_2711;
wire n_17021;
wire n_17710;
wire n_6663;
wire n_12609;
wire n_4441;
wire n_18248;
wire n_8155;
wire n_11360;
wire n_11868;
wire n_1664;
wire n_3022;
wire n_8098;
wire n_9191;
wire n_17791;
wire n_5654;
wire n_2345;
wire n_18202;
wire n_6376;
wire n_18141;
wire n_5113;
wire n_12888;
wire n_5479;
wire n_19407;
wire n_8485;
wire n_14852;
wire n_7001;
wire n_9650;
wire n_4822;
wire n_13070;
wire n_850;
wire n_5692;
wire n_8473;
wire n_13640;
wire n_14147;
wire n_14491;
wire n_15011;
wire n_17607;
wire n_3768;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_5441;
wire n_9664;
wire n_20367;
wire n_3785;
wire n_14928;
wire n_2602;
wire n_2980;
wire n_13778;
wire n_696;
wire n_9931;
wire n_16419;
wire n_16470;
wire n_1082;
wire n_1317;
wire n_16956;
wire n_3227;
wire n_4055;
wire n_14634;
wire n_2178;
wire n_10753;
wire n_13174;
wire n_7108;
wire n_14455;
wire n_1796;
wire n_17164;
wire n_11879;
wire n_2082;
wire n_7876;
wire n_17175;
wire n_9656;
wire n_3707;
wire n_8148;
wire n_8150;
wire n_3578;
wire n_909;
wire n_12596;
wire n_15398;
wire n_15593;
wire n_18175;
wire n_4925;
wire n_16424;
wire n_5415;
wire n_13945;
wire n_8986;
wire n_19367;
wire n_20137;
wire n_12697;
wire n_7260;
wire n_6409;
wire n_11939;
wire n_1634;
wire n_3252;
wire n_627;
wire n_14347;
wire n_7552;
wire n_19052;
wire n_17969;
wire n_12166;
wire n_2133;
wire n_1712;
wire n_1523;
wire n_10646;
wire n_15725;
wire n_1627;
wire n_11704;
wire n_20548;
wire n_17506;
wire n_18050;
wire n_8763;
wire n_5208;
wire n_8679;
wire n_7239;
wire n_15582;
wire n_16415;
wire n_9848;
wire n_14447;
wire n_11962;
wire n_5690;
wire n_9227;
wire n_7050;
wire n_17137;
wire n_2573;
wire n_2646;
wire n_6623;
wire n_13951;
wire n_13968;
wire n_10378;
wire n_16924;
wire n_1364;
wire n_13316;
wire n_10313;
wire n_13689;
wire n_8139;
wire n_17268;
wire n_18000;
wire n_19384;
wire n_3037;
wire n_19288;
wire n_3729;
wire n_19431;
wire n_10773;
wire n_18210;
wire n_2537;
wire n_8830;
wire n_4483;
wire n_5347;
wire n_14836;
wire n_12867;
wire n_4988;
wire n_15960;
wire n_7568;
wire n_15343;
wire n_6354;
wire n_6344;
wire n_12123;
wire n_9772;
wire n_18885;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_6021;
wire n_7949;
wire n_15370;
wire n_7724;
wire n_18001;
wire n_4284;
wire n_6305;
wire n_1947;
wire n_12547;
wire n_16148;
wire n_20557;
wire n_15577;
wire n_3426;
wire n_16550;
wire n_4971;
wire n_19066;
wire n_5857;
wire n_8646;
wire n_13415;
wire n_10259;
wire n_7107;
wire n_17111;
wire n_6457;
wire n_8597;
wire n_17951;
wire n_17379;
wire n_987;
wire n_7123;
wire n_5499;
wire n_720;
wire n_8117;
wire n_15169;
wire n_1707;
wire n_10213;
wire n_13888;
wire n_16592;
wire n_8208;
wire n_797;
wire n_2933;
wire n_19373;
wire n_1878;
wire n_20004;
wire n_8536;
wire n_17252;
wire n_9435;
wire n_7229;
wire n_8350;
wire n_16475;
wire n_5190;
wire n_13892;
wire n_16361;
wire n_14559;
wire n_16831;
wire n_4097;
wire n_1666;
wire n_19696;
wire n_5392;
wire n_17110;
wire n_14052;
wire n_14311;
wire n_13765;
wire n_10332;
wire n_7709;
wire n_15290;
wire n_11874;
wire n_13926;
wire n_10171;
wire n_15184;
wire n_1228;
wire n_5455;
wire n_18131;
wire n_5442;
wire n_6386;
wire n_12803;
wire n_5948;
wire n_19518;
wire n_5511;
wire n_2898;
wire n_6208;
wire n_6739;
wire n_15779;
wire n_8202;
wire n_15366;
wire n_3200;
wire n_12734;
wire n_3167;
wire n_7185;
wire n_6291;
wire n_11489;
wire n_10269;
wire n_19504;
wire n_12262;
wire n_14910;
wire n_14385;
wire n_14499;
wire n_8738;
wire n_9126;
wire n_15368;
wire n_19077;
wire n_11376;
wire n_9438;
wire n_18433;
wire n_7808;
wire n_6544;
wire n_9122;
wire n_14731;
wire n_20227;
wire n_20397;
wire n_683;
wire n_5140;
wire n_4992;
wire n_5197;
wire n_16337;
wire n_17691;
wire n_8721;
wire n_12820;
wire n_9912;
wire n_6356;
wire n_13558;
wire n_3577;
wire n_2432;
wire n_10148;
wire n_19491;
wire n_1363;
wire n_3641;
wire n_2218;
wire n_16890;
wire n_13890;
wire n_5481;
wire n_9264;
wire n_14483;
wire n_8326;
wire n_8670;
wire n_5308;
wire n_5184;
wire n_5794;
wire n_15179;
wire n_7638;
wire n_15724;
wire n_19303;
wire n_20412;
wire n_4053;
wire n_10234;
wire n_8836;
wire n_7019;
wire n_11325;
wire n_14838;
wire n_15207;
wire n_13521;
wire n_4167;
wire n_19788;
wire n_14926;
wire n_10731;
wire n_9878;
wire n_14591;
wire n_14363;
wire n_14576;
wire n_4431;
wire n_17797;
wire n_1125;
wire n_11498;
wire n_10513;
wire n_441;
wire n_7296;
wire n_4299;
wire n_7575;
wire n_3571;
wire n_7083;
wire n_1775;
wire n_7720;
wire n_11643;
wire n_1093;
wire n_6268;
wire n_5827;
wire n_5199;
wire n_6456;
wire n_11103;
wire n_16823;
wire n_16966;
wire n_14088;
wire n_5313;
wire n_17926;
wire n_13817;
wire n_3856;
wire n_9971;
wire n_19579;
wire n_3425;
wire n_10894;
wire n_14118;
wire n_18082;
wire n_9524;
wire n_20534;
wire n_6467;
wire n_9243;
wire n_9282;
wire n_1453;
wire n_6796;
wire n_19821;
wire n_18821;
wire n_12417;
wire n_4830;
wire n_13225;
wire n_20045;
wire n_17006;
wire n_1224;
wire n_10208;
wire n_20107;
wire n_3243;
wire n_1135;
wire n_2889;
wire n_10804;
wire n_6486;
wire n_3960;
wire n_17246;
wire n_17167;
wire n_20513;
wire n_18357;
wire n_8438;
wire n_13355;
wire n_18160;
wire n_4693;
wire n_18614;
wire n_20475;
wire n_10793;
wire n_2000;
wire n_14672;
wire n_4267;
wire n_15127;
wire n_6732;
wire n_2270;
wire n_12711;
wire n_20454;
wire n_12219;
wire n_906;
wire n_10440;
wire n_1733;
wire n_9695;
wire n_11306;
wire n_19169;
wire n_4609;
wire n_19813;
wire n_1687;
wire n_8757;
wire n_2328;
wire n_13035;
wire n_7020;
wire n_13021;
wire n_613;
wire n_12893;
wire n_8596;
wire n_3314;
wire n_3016;
wire n_11292;
wire n_20238;
wire n_554;
wire n_13502;
wire n_5223;
wire n_6298;
wire n_5474;
wire n_12289;
wire n_10813;
wire n_1889;
wire n_10757;
wire n_13046;
wire n_13935;
wire n_435;
wire n_16670;
wire n_762;
wire n_11431;
wire n_1778;
wire n_5287;
wire n_13646;
wire n_1079;
wire n_5083;
wire n_6007;
wire n_3338;
wire n_18186;
wire n_4217;
wire n_6197;
wire n_6658;
wire n_4906;
wire n_8834;
wire n_3636;
wire n_2327;
wire n_16429;
wire n_15262;
wire n_10822;
wire n_18773;
wire n_7104;
wire n_7467;
wire n_14609;
wire n_2597;
wire n_9534;
wire n_3194;
wire n_13380;
wire n_5771;
wire n_17369;
wire n_13053;
wire n_9792;
wire n_7513;
wire n_11836;
wire n_349;
wire n_6602;
wire n_10924;
wire n_17421;
wire n_11186;
wire n_9742;
wire n_6484;
wire n_19642;
wire n_3637;
wire n_12527;
wire n_4574;
wire n_19800;
wire n_1859;
wire n_9019;
wire n_13891;
wire n_1718;
wire n_8985;
wire n_7692;
wire n_19463;
wire n_12477;
wire n_4234;
wire n_14325;
wire n_15503;
wire n_10418;
wire n_1768;
wire n_19589;
wire n_3974;
wire n_10875;
wire n_1847;
wire n_3634;
wire n_11736;
wire n_7560;
wire n_16270;
wire n_14729;
wire n_11846;
wire n_1397;
wire n_12400;
wire n_901;
wire n_2755;
wire n_4660;
wire n_1623;
wire n_16861;
wire n_9145;
wire n_12092;
wire n_3112;
wire n_12295;
wire n_9754;
wire n_19549;
wire n_9315;
wire n_18483;
wire n_5428;
wire n_4151;
wire n_7451;
wire n_6734;
wire n_7476;
wire n_5570;
wire n_18096;
wire n_785;
wire n_7392;
wire n_7495;
wire n_5435;
wire n_9765;
wire n_3213;
wire n_3820;
wire n_5200;
wire n_6941;
wire n_1168;
wire n_5115;
wire n_1943;
wire n_5566;
wire n_7829;
wire n_3249;
wire n_8680;
wire n_2722;
wire n_20461;
wire n_4152;
wire n_16522;
wire n_20246;
wire n_10394;
wire n_11391;
wire n_15462;
wire n_20328;
wire n_5244;
wire n_12714;
wire n_16779;
wire n_5889;
wire n_19024;
wire n_5391;
wire n_1938;
wire n_9763;
wire n_11070;
wire n_13337;
wire n_15112;
wire n_18146;
wire n_3394;
wire n_9162;
wire n_19977;
wire n_1715;
wire n_14849;
wire n_1443;
wire n_1272;
wire n_16661;
wire n_5849;
wire n_11648;
wire n_4554;
wire n_19044;
wire n_10322;
wire n_7135;
wire n_8555;
wire n_10695;
wire n_8636;
wire n_7024;
wire n_15912;
wire n_16206;
wire n_19812;
wire n_8508;
wire n_19509;
wire n_18827;
wire n_16529;
wire n_1705;
wire n_3905;
wire n_8207;
wire n_11653;
wire n_4680;
wire n_3013;
wire n_20033;
wire n_11717;
wire n_15246;
wire n_14940;
wire n_6165;
wire n_19153;
wire n_17553;
wire n_15395;
wire n_12838;
wire n_2670;
wire n_19918;
wire n_18813;
wire n_13505;
wire n_5910;
wire n_12776;
wire n_1569;
wire n_19962;
wire n_7033;
wire n_13156;
wire n_15529;
wire n_10710;
wire n_5557;
wire n_411;
wire n_8850;
wire n_14647;
wire n_18384;
wire n_8002;
wire n_19610;
wire n_1795;
wire n_16722;
wire n_9090;
wire n_16412;
wire n_12008;
wire n_6119;
wire n_1545;
wire n_4145;
wire n_4821;
wire n_3121;
wire n_9261;
wire n_8301;
wire n_17453;
wire n_12223;
wire n_18706;
wire n_16758;
wire n_548;
wire n_10942;
wire n_19983;
wire n_11430;
wire n_13010;
wire n_19073;
wire n_345;
wire n_11239;
wire n_4943;
wire n_10953;
wire n_7842;
wire n_2629;
wire n_2172;
wire n_6202;
wire n_17831;
wire n_12898;
wire n_4682;
wire n_19523;
wire n_15540;
wire n_10343;
wire n_4942;
wire n_9258;
wire n_1086;
wire n_10286;
wire n_10371;
wire n_14990;
wire n_2561;
wire n_16691;
wire n_7236;
wire n_10257;
wire n_3305;
wire n_11219;
wire n_20232;
wire n_10047;
wire n_14541;
wire n_3267;
wire n_16186;
wire n_1914;
wire n_1318;
wire n_13766;
wire n_11226;
wire n_3005;
wire n_16989;
wire n_11413;
wire n_4840;
wire n_1029;
wire n_16617;
wire n_5320;
wire n_5353;
wire n_13710;
wire n_11232;
wire n_2417;
wire n_9105;
wire n_12080;
wire n_16261;
wire n_5093;
wire n_1556;
wire n_19512;
wire n_5979;
wire n_9668;
wire n_13335;
wire n_14022;
wire n_2083;
wire n_5517;
wire n_3207;
wire n_11276;
wire n_5605;
wire n_3401;
wire n_10744;
wire n_3242;
wire n_9870;
wire n_3613;
wire n_11334;
wire n_7678;
wire n_1045;
wire n_13075;
wire n_13736;
wire n_13129;
wire n_9178;
wire n_6063;
wire n_16118;
wire n_1325;
wire n_6504;
wire n_2923;
wire n_1727;
wire n_13586;
wire n_15813;
wire n_10597;
wire n_17382;
wire n_16281;
wire n_11827;
wire n_13049;
wire n_13961;
wire n_17413;
wire n_15745;
wire n_20400;
wire n_3814;
wire n_6003;
wire n_6684;
wire n_19084;
wire n_13063;
wire n_20057;
wire n_5451;
wire n_9323;
wire n_19728;
wire n_6961;
wire n_3543;
wire n_13252;
wire n_9922;
wire n_12024;
wire n_13084;
wire n_2903;
wire n_16622;
wire n_15374;
wire n_3808;
wire n_4365;
wire n_18123;
wire n_16440;
wire n_7929;
wire n_16821;
wire n_10572;
wire n_16431;
wire n_1007;
wire n_1929;
wire n_19272;
wire n_1592;
wire n_19455;
wire n_13985;
wire n_3758;
wire n_17594;
wire n_20411;
wire n_14124;
wire n_19119;
wire n_17658;
wire n_13552;
wire n_18086;
wire n_12681;
wire n_3343;
wire n_18419;
wire n_13022;
wire n_18583;
wire n_2752;
wire n_17047;
wire n_9513;
wire n_16447;
wire n_16124;
wire n_4885;
wire n_15446;
wire n_10555;
wire n_19179;
wire n_10314;
wire n_4550;
wire n_6988;
wire n_13656;
wire n_18967;
wire n_3658;
wire n_20585;
wire n_6834;
wire n_6817;
wire n_6927;
wire n_20017;
wire n_5209;
wire n_16841;
wire n_15470;
wire n_6215;
wire n_4212;
wire n_20316;
wire n_5699;
wire n_181;
wire n_5765;
wire n_15754;
wire n_17375;
wire n_7862;
wire n_16708;
wire n_17439;
wire n_10630;
wire n_17955;
wire n_8808;
wire n_10061;
wire n_300;
wire n_15599;
wire n_11865;
wire n_13024;
wire n_10694;
wire n_20499;
wire n_11041;
wire n_14490;
wire n_9708;
wire n_5064;
wire n_15479;
wire n_7119;
wire n_8889;
wire n_601;
wire n_13986;
wire n_9790;
wire n_11973;
wire n_5759;
wire n_13329;
wire n_7874;
wire n_8490;
wire n_10329;
wire n_9979;
wire n_8767;
wire n_13946;
wire n_9505;
wire n_2566;
wire n_15028;
wire n_2702;
wire n_7420;
wire n_7102;
wire n_13618;
wire n_19838;
wire n_4568;
wire n_10662;
wire n_5559;
wire n_18653;
wire n_17534;
wire n_14993;
wire n_14327;
wire n_8624;
wire n_11022;
wire n_10247;
wire n_5377;
wire n_1016;
wire n_8796;
wire n_4106;
wire n_1501;
wire n_17829;
wire n_10733;
wire n_10472;
wire n_12597;
wire n_13744;
wire n_12834;
wire n_10066;
wire n_17239;
wire n_14335;
wire n_6419;
wire n_3553;
wire n_18989;
wire n_2275;
wire n_15087;
wire n_2568;
wire n_2022;
wire n_3494;
wire n_6244;
wire n_6900;
wire n_9337;
wire n_15219;
wire n_908;
wire n_9432;
wire n_17295;
wire n_19563;
wire n_7705;
wire n_2106;
wire n_5350;
wire n_5470;
wire n_7932;
wire n_18331;
wire n_7058;
wire n_15009;
wire n_8262;
wire n_5700;
wire n_7981;
wire n_9874;
wire n_12588;
wire n_17203;
wire n_15648;
wire n_17548;
wire n_5874;
wire n_9231;
wire n_20230;
wire n_3328;
wire n_18612;
wire n_7973;
wire n_6815;
wire n_15634;
wire n_9569;
wire n_14823;
wire n_19938;
wire n_14691;
wire n_2530;
wire n_16908;
wire n_16508;
wire n_9719;
wire n_8358;
wire n_9552;
wire n_13822;
wire n_14948;
wire n_6317;
wire n_475;
wire n_492;
wire n_4012;
wire n_10756;
wire n_20333;
wire n_3645;
wire n_17099;
wire n_14387;
wire n_16572;
wire n_11797;
wire n_18889;
wire n_18933;
wire n_14106;
wire n_18788;
wire n_13616;
wire n_18667;
wire n_7820;
wire n_8881;
wire n_7844;
wire n_14301;
wire n_15468;
wire n_9633;
wire n_3422;
wire n_4845;
wire n_3086;
wire n_2033;
wire n_13627;
wire n_878;
wire n_19040;
wire n_5120;
wire n_13112;
wire n_10042;
wire n_10478;
wire n_16581;
wire n_981;
wire n_18597;
wire n_13163;
wire n_3702;
wire n_8754;
wire n_9847;
wire n_18098;
wire n_16968;
wire n_2233;
wire n_10367;
wire n_3233;
wire n_10867;
wire n_3310;
wire n_4061;
wire n_7460;
wire n_9519;
wire n_19735;
wire n_14814;
wire n_6367;
wire n_13564;
wire n_12671;
wire n_8714;
wire n_13260;
wire n_17302;
wire n_10085;
wire n_1051;
wire n_20023;
wire n_8182;
wire n_16165;
wire n_14090;
wire n_6056;
wire n_7200;
wire n_3206;
wire n_2363;
wire n_553;
wire n_15424;
wire n_4903;
wire n_17301;
wire n_15554;
wire n_15836;
wire n_15966;
wire n_16009;
wire n_15309;
wire n_14463;
wire n_2540;
wire n_973;
wire n_5743;
wire n_13503;
wire n_11152;
wire n_16318;
wire n_20182;
wire n_14166;
wire n_4522;
wire n_10122;
wire n_679;
wire n_9327;
wire n_16175;
wire n_5368;
wire n_4263;
wire n_14271;
wire n_7059;
wire n_915;
wire n_14425;
wire n_5971;
wire n_6327;
wire n_11964;
wire n_3155;
wire n_7826;
wire n_19078;
wire n_5933;
wire n_7076;
wire n_4780;
wire n_11403;
wire n_2697;
wire n_6866;
wire n_17108;
wire n_2512;
wire n_9387;
wire n_3039;
wire n_14596;
wire n_6514;
wire n_9794;
wire n_20571;
wire n_1322;
wire n_16387;
wire n_11142;
wire n_1958;
wire n_20147;
wire n_17434;
wire n_1197;
wire n_17509;
wire n_4984;
wire n_20261;
wire n_3420;
wire n_10862;
wire n_4283;
wire n_8911;
wire n_900;
wire n_8248;
wire n_11476;
wire n_2659;
wire n_13633;
wire n_14538;
wire n_2116;
wire n_19534;
wire n_1013;
wire n_17999;
wire n_11367;
wire n_15478;
wire n_2183;
wire n_16797;
wire n_12676;
wire n_20432;
wire n_18755;
wire n_3392;
wire n_13913;
wire n_19166;
wire n_8733;
wire n_6050;
wire n_7976;
wire n_13080;
wire n_13403;
wire n_17444;
wire n_1581;
wire n_1357;
wire n_14952;
wire n_1853;
wire n_10386;
wire n_12128;
wire n_14060;
wire n_14018;
wire n_15959;
wire n_5563;
wire n_1348;
wire n_11026;
wire n_13309;
wire n_15292;
wire n_11467;
wire n_12672;
wire n_12063;
wire n_8330;
wire n_1009;
wire n_15560;
wire n_1160;
wire n_15065;
wire n_5717;
wire n_1247;
wire n_6017;
wire n_9696;
wire n_20220;
wire n_15771;
wire n_15508;
wire n_20555;
wire n_471;
wire n_17990;
wire n_14148;
wire n_5720;
wire n_4702;
wire n_4895;
wire n_12924;
wire n_16331;
wire n_12732;
wire n_17171;
wire n_12649;
wire n_5898;
wire n_17458;
wire n_6858;
wire n_9464;
wire n_9252;
wire n_6649;
wire n_6283;
wire n_4026;
wire n_12843;
wire n_14279;
wire n_1140;
wire n_1670;
wire n_2344;
wire n_17856;
wire n_2365;
wire n_19573;
wire n_15687;
wire n_8540;
wire n_2447;
wire n_11248;
wire n_9915;
wire n_5940;
wire n_6089;
wire n_7588;
wire n_18480;
wire n_4969;
wire n_10017;
wire n_20540;
wire n_11141;
wire n_5105;
wire n_11093;
wire n_19556;
wire n_17716;
wire n_5263;
wire n_2510;
wire n_19873;
wire n_6713;
wire n_18750;
wire n_15968;
wire n_17893;
wire n_4602;
wire n_13181;
wire n_18303;
wire n_1163;
wire n_16487;
wire n_17592;
wire n_15047;
wire n_3122;
wire n_5567;
wire n_8343;
wire n_7593;
wire n_17156;
wire n_17908;
wire n_14085;
wire n_8068;
wire n_19599;
wire n_2173;
wire n_7764;
wire n_20357;
wire n_19634;
wire n_10196;
wire n_493;
wire n_14573;
wire n_17433;
wire n_19453;
wire n_20085;
wire n_2108;
wire n_8693;
wire n_6454;
wire n_12625;
wire n_12177;
wire n_7307;
wire n_14512;
wire n_1280;
wire n_6918;
wire n_16214;
wire n_13761;
wire n_19576;
wire n_3296;
wire n_19065;
wire n_16219;
wire n_17017;
wire n_14456;
wire n_13364;
wire n_11494;
wire n_14743;
wire n_10218;
wire n_18492;
wire n_3792;
wire n_4791;
wire n_19127;
wire n_14859;
wire n_8062;
wire n_11832;
wire n_6375;
wire n_12974;
wire n_13078;
wire n_1956;
wire n_7047;
wire n_6632;
wire n_4549;
wire n_17241;
wire n_15795;
wire n_10542;
wire n_16814;
wire n_4349;
wire n_10681;
wire n_15162;
wire n_9732;
wire n_16494;
wire n_13370;
wire n_11894;
wire n_10222;
wire n_10524;
wire n_6705;
wire n_17988;
wire n_8629;
wire n_818;
wire n_9517;
wire n_15237;
wire n_15862;
wire n_6591;
wire n_2207;
wire n_13643;
wire n_9780;
wire n_3482;
wire n_2198;
wire n_13607;
wire n_6289;
wire n_3272;
wire n_8524;
wire n_19355;
wire n_18907;
wire n_4393;
wire n_14114;
wire n_1068;
wire n_932;
wire n_14904;
wire n_3317;
wire n_3978;
wire n_5560;
wire n_6512;
wire n_4074;
wire n_4918;
wire n_13820;
wire n_4013;
wire n_6703;
wire n_12122;
wire n_13428;
wire n_354;
wire n_17958;
wire n_19667;
wire n_2941;
wire n_547;
wire n_17194;
wire n_19686;
wire n_6086;
wire n_20483;
wire n_16668;
wire n_4147;
wire n_4477;
wire n_18139;
wire n_3168;
wire n_12184;
wire n_10210;
wire n_1793;
wire n_5611;
wire n_12571;
wire n_6219;
wire n_11853;
wire n_19626;
wire n_16770;
wire n_4742;
wire n_9609;
wire n_10029;
wire n_1703;
wire n_6761;
wire n_8972;
wire n_19919;
wire n_11725;
wire n_13635;
wire n_10801;
wire n_9206;
wire n_3384;
wire n_18488;
wire n_15698;
wire n_1950;
wire n_6811;
wire n_16865;
wire n_18642;
wire n_11622;
wire n_4838;
wire n_12336;
wire n_18345;
wire n_19754;
wire n_12543;
wire n_16129;
wire n_347;
wire n_9705;
wire n_16585;
wire n_17490;
wire n_2965;
wire n_9624;
wire n_3861;
wire n_20306;
wire n_1977;
wire n_10389;
wire n_3891;
wire n_15688;
wire n_1655;
wire n_13677;
wire n_1886;
wire n_13757;
wire n_14036;
wire n_12463;
wire n_10990;
wire n_12263;
wire n_11640;
wire n_8982;
wire n_17899;
wire n_13910;
wire n_4673;
wire n_7086;
wire n_3415;
wire n_2947;
wire n_9532;
wire n_18195;
wire n_6601;
wire n_16247;
wire n_13196;
wire n_17482;
wire n_5088;
wire n_19261;
wire n_8034;
wire n_484;
wire n_15824;
wire n_5856;
wire n_9836;
wire n_2497;
wire n_11525;
wire n_11999;
wire n_10837;
wire n_3545;
wire n_18921;
wire n_20299;
wire n_10554;
wire n_3993;
wire n_8994;
wire n_17827;
wire n_8413;
wire n_4685;
wire n_19986;
wire n_10149;
wire n_19473;
wire n_19393;
wire n_2663;
wire n_5825;
wire n_20020;
wire n_2938;
wire n_3780;
wire n_15791;
wire n_12190;
wire n_15484;
wire n_15152;
wire n_19961;
wire n_11847;
wire n_11976;
wire n_20346;
wire n_12511;
wire n_2750;
wire n_11167;
wire n_2775;
wire n_8765;
wire n_3477;
wire n_2349;
wire n_2684;
wire n_8213;
wire n_1495;
wire n_14472;
wire n_10534;
wire n_11049;
wire n_14974;
wire n_8451;
wire n_19410;
wire n_1128;
wire n_12743;
wire n_16523;
wire n_8731;
wire n_8385;
wire n_4999;
wire n_15587;
wire n_4922;
wire n_7370;
wire n_15322;
wire n_13539;
wire n_9350;
wire n_18324;
wire n_19383;
wire n_17917;
wire n_7026;
wire n_7053;
wire n_14618;
wire n_9226;
wire n_1765;
wire n_2707;
wire n_18810;
wire n_10608;
wire n_16355;
wire n_7173;
wire n_7042;
wire n_17314;
wire n_718;
wire n_17915;
wire n_5331;
wire n_19225;
wire n_19011;
wire n_16774;
wire n_16436;
wire n_2089;
wire n_10638;
wire n_17923;
wire n_9112;
wire n_18582;
wire n_18970;
wire n_4216;
wire n_19284;
wire n_5797;
wire n_9235;
wire n_16570;
wire n_19124;
wire n_4240;
wire n_3491;
wire n_13852;
wire n_9333;
wire n_704;
wire n_4162;
wire n_17813;
wire n_14089;
wire n_15758;
wire n_1999;
wire n_2731;
wire n_622;
wire n_147;
wire n_3353;
wire n_11804;
wire n_14234;
wire n_3018;
wire n_14125;
wire n_5800;
wire n_6562;
wire n_12809;
wire n_18770;
wire n_4785;
wire n_2002;
wire n_2138;
wire n_2414;
wire n_1771;
wire n_11052;
wire n_3148;
wire n_17350;
wire n_18598;
wire n_6671;
wire n_13470;
wire n_6812;
wire n_12361;
wire n_4864;
wire n_19151;
wire n_9488;
wire n_5758;
wire n_10748;
wire n_13068;
wire n_19158;
wire n_3775;
wire n_18795;
wire n_1176;
wire n_20459;
wire n_7792;
wire n_15985;
wire n_8161;
wire n_18798;
wire n_5763;
wire n_10014;
wire n_15723;
wire n_16840;
wire n_6029;
wire n_18698;
wire n_10677;
wire n_18269;
wire n_5751;
wire n_15852;
wire n_18857;
wire n_19216;
wire n_12321;
wire n_5924;
wire n_11247;
wire n_290;
wire n_18581;
wire n_8384;
wire n_6445;
wire n_18079;
wire n_13106;
wire n_19863;
wire n_14294;
wire n_17609;
wire n_6701;
wire n_14862;
wire n_7380;
wire n_8736;
wire n_11514;
wire n_4497;
wire n_1568;
wire n_12470;
wire n_12994;
wire n_18604;
wire n_10215;
wire n_20005;
wire n_18768;
wire n_14059;
wire n_4871;
wire n_10834;
wire n_17632;
wire n_20257;
wire n_17611;
wire n_1665;
wire n_19341;
wire n_154;
wire n_12064;
wire n_2127;
wire n_12696;
wire n_18024;
wire n_15735;
wire n_11133;
wire n_5449;
wire n_20054;
wire n_17143;
wire n_18341;
wire n_10871;
wire n_16405;
wire n_5926;
wire n_2354;
wire n_5398;
wire n_4573;
wire n_14624;
wire n_16600;
wire n_15036;
wire n_17695;
wire n_18193;
wire n_19489;
wire n_11571;
wire n_14120;
wire n_13147;
wire n_8844;
wire n_7641;
wire n_6106;
wire n_3480;
wire n_1368;
wire n_14407;
wire n_14260;
wire n_16845;
wire n_18924;
wire n_17307;
wire n_7169;
wire n_10407;
wire n_19330;
wire n_14175;
wire n_11941;
wire n_4368;
wire n_15780;
wire n_18085;
wire n_1942;
wire n_3196;
wire n_15189;
wire n_8110;
wire n_5319;
wire n_9008;
wire n_12079;
wire n_15335;
wire n_399;
wire n_1440;
wire n_19147;
wire n_2063;
wire n_15227;
wire n_8805;
wire n_6014;
wire n_7209;
wire n_18908;
wire n_15026;
wire n_13895;
wire n_2475;
wire n_5181;
wire n_13222;
wire n_6979;
wire n_3144;
wire n_1268;
wire n_17284;
wire n_5583;
wire n_15987;
wire n_10462;
wire n_20440;
wire n_642;
wire n_3481;
wire n_11769;
wire n_8856;
wire n_19362;
wire n_303;
wire n_6142;
wire n_20582;
wire n_14901;
wire n_7769;
wire n_2374;
wire n_416;
wire n_17034;
wire n_10291;
wire n_4597;
wire n_18575;
wire n_18764;
wire n_3364;
wire n_17502;
wire n_14333;
wire n_7233;
wire n_8732;
wire n_13506;
wire n_7602;
wire n_18587;
wire n_9296;
wire n_7390;
wire n_10669;
wire n_19515;
wire n_8231;
wire n_20161;
wire n_13717;
wire n_5127;
wire n_2920;
wire n_7598;
wire n_12440;
wire n_19032;
wire n_8908;
wire n_1374;
wire n_2648;
wire n_16085;
wire n_1169;
wire n_6767;
wire n_12782;
wire n_3093;
wire n_10111;
wire n_19186;
wire n_19629;
wire n_15300;
wire n_6385;
wire n_11354;
wire n_20009;
wire n_17796;
wire n_7045;
wire n_3169;
wire n_8740;
wire n_11727;
wire n_6788;
wire n_12192;
wire n_2204;
wire n_177;
wire n_2087;
wire n_17342;
wire n_14465;
wire n_13412;
wire n_4422;
wire n_11749;
wire n_11300;
wire n_6143;
wire n_20569;
wire n_13457;
wire n_12551;
wire n_18066;
wire n_12497;
wire n_15043;
wire n_4632;
wire n_3084;
wire n_16602;
wire n_2343;
wire n_5967;
wire n_4963;
wire n_16864;
wire n_16761;
wire n_2942;
wire n_4966;
wire n_4714;
wire n_7679;
wire n_18133;
wire n_20529;
wire n_7936;
wire n_8966;
wire n_4847;
wire n_10287;
wire n_8538;
wire n_12101;
wire n_11145;
wire n_3586;
wire n_3653;
wire n_16684;
wire n_19594;
wire n_725;
wire n_10349;
wire n_4668;
wire n_5213;
wire n_16340;
wire n_7490;
wire n_7545;
wire n_1273;
wire n_7160;
wire n_9809;
wire n_10750;
wire n_617;
wire n_7295;
wire n_14338;
wire n_7348;
wire n_19071;
wire n_10673;
wire n_12460;
wire n_6681;
wire n_17554;
wire n_16071;
wire n_3991;
wire n_15394;
wire n_3516;
wire n_16875;
wire n_15941;
wire n_20439;
wire n_610;
wire n_9558;
wire n_11594;
wire n_8715;
wire n_12474;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_7162;
wire n_16655;
wire n_20272;
wire n_12346;
wire n_517;
wire n_18167;
wire n_4182;
wire n_667;
wire n_8371;
wire n_13916;
wire n_15195;
wire n_1279;
wire n_11458;
wire n_17056;
wire n_12244;
wire n_18753;
wire n_16188;
wire n_15644;
wire n_14255;
wire n_11670;
wire n_7681;
wire n_11504;
wire n_19972;
wire n_16850;
wire n_13981;
wire n_4637;
wire n_11516;
wire n_2412;
wire n_8392;
wire n_14659;
wire n_8095;
wire n_10830;
wire n_16868;
wire n_17644;
wire n_5118;
wire n_7503;
wire n_6854;
wire n_17254;
wire n_2757;
wire n_18733;
wire n_4977;
wire n_2716;
wire n_12953;
wire n_2452;
wire n_15224;
wire n_9215;
wire n_11406;
wire n_19835;
wire n_3043;
wire n_14963;
wire n_11047;
wire n_8050;
wire n_12817;
wire n_8399;
wire n_2543;
wire n_5090;
wire n_16916;
wire n_13866;
wire n_3177;
wire n_12435;
wire n_10946;
wire n_18106;
wire n_7065;
wire n_9216;
wire n_1262;
wire n_4835;
wire n_11961;
wire n_6122;
wire n_7911;
wire n_17486;
wire n_17504;
wire n_7330;
wire n_14605;
wire n_9202;
wire n_2373;
wire n_13543;
wire n_10351;
wire n_13772;
wire n_4734;
wire n_7493;
wire n_12940;
wire n_10460;
wire n_15487;
wire n_19221;
wire n_10334;
wire n_2244;
wire n_11614;
wire n_4290;
wire n_1684;
wire n_1352;
wire n_5407;
wire n_15242;
wire n_8422;
wire n_12224;
wire n_7088;
wire n_9394;
wire n_2704;
wire n_8878;
wire n_7440;
wire n_17681;
wire n_260;
wire n_17676;
wire n_14797;
wire n_9622;
wire n_14177;
wire n_14093;
wire n_3318;
wire n_14607;
wire n_10191;
wire n_4888;
wire n_17919;
wire n_776;
wire n_6000;
wire n_12679;
wire n_11168;
wire n_14921;
wire n_20406;
wire n_10911;
wire n_12756;
wire n_5294;
wire n_5004;
wire n_16097;
wire n_9845;
wire n_16147;
wire n_7374;
wire n_14389;
wire n_19514;
wire n_11937;
wire n_17277;
wire n_2229;
wire n_4527;
wire n_6046;
wire n_8251;
wire n_5323;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_14621;
wire n_3184;
wire n_18864;
wire n_20468;
wire n_3075;
wire n_17875;
wire n_11192;
wire n_4949;
wire n_6852;
wire n_8677;
wire n_9091;
wire n_17206;
wire n_13914;
wire n_14663;
wire n_16921;
wire n_17559;
wire n_2536;
wire n_9699;
wire n_13277;
wire n_12340;
wire n_18143;
wire n_16742;
wire n_18464;
wire n_13494;
wire n_5260;
wire n_9751;
wire n_20525;
wire n_5809;
wire n_10543;
wire n_7924;
wire n_17225;
wire n_20443;
wire n_560;
wire n_1321;
wire n_7659;
wire n_569;
wire n_3530;
wire n_20539;
wire n_16203;
wire n_8875;
wire n_20079;
wire n_9585;
wire n_7153;
wire n_11101;
wire n_1235;
wire n_12662;
wire n_1292;
wire n_15697;
wire n_17879;
wire n_18140;
wire n_9293;
wire n_12503;
wire n_18510;
wire n_15202;
wire n_18218;
wire n_12871;
wire n_13029;
wire n_10591;
wire n_11845;
wire n_18224;
wire n_16400;
wire n_2246;
wire n_4469;
wire n_20441;
wire n_431;
wire n_10809;
wire n_16934;
wire n_10899;
wire n_9639;
wire n_11898;
wire n_15250;
wire n_17193;
wire n_6711;
wire n_1941;
wire n_11997;
wire n_8946;
wire n_13090;
wire n_18984;
wire n_13541;
wire n_20092;
wire n_16958;
wire n_4924;
wire n_13908;
wire n_9646;
wire n_8017;
wire n_17396;
wire n_766;
wire n_1746;
wire n_7275;
wire n_8795;
wire n_7195;
wire n_11199;
wire n_17642;
wire n_11264;
wire n_19791;
wire n_2062;
wire n_4539;
wire n_6072;
wire n_7610;
wire n_12303;
wire n_9501;
wire n_11896;
wire n_16229;
wire n_10006;
wire n_11757;
wire n_2070;
wire n_18447;
wire n_12622;
wire n_6353;
wire n_4953;
wire n_12659;
wire n_2348;
wire n_6818;
wire n_391;
wire n_2066;
wire n_7539;
wire n_1476;
wire n_12629;
wire n_12868;
wire n_19263;
wire n_10275;
wire n_3458;
wire n_7775;
wire n_11392;
wire n_3190;
wire n_7930;
wire n_7661;
wire n_5383;
wire n_16498;
wire n_19673;
wire n_14165;
wire n_17309;
wire n_19413;
wire n_13787;
wire n_875;
wire n_1678;
wire n_13674;
wire n_18311;
wire n_13912;
wire n_10292;
wire n_7969;
wire n_6864;
wire n_11278;
wire n_14445;
wire n_3787;
wire n_7548;
wire n_16732;
wire n_4450;
wire n_6156;
wire n_12913;
wire n_7064;
wire n_19285;
wire n_16839;
wire n_16798;
wire n_12154;
wire n_8000;
wire n_14427;
wire n_5645;
wire n_3990;
wire n_18327;
wire n_6917;
wire n_6937;
wire n_1628;
wire n_20527;
wire n_9963;
wire n_988;
wire n_17211;
wire n_20337;
wire n_7324;
wire n_2507;
wire n_5878;
wire n_10152;
wire n_5671;
wire n_17568;
wire n_1536;
wire n_6301;
wire n_18061;
wire n_16815;
wire n_18022;
wire n_1132;
wire n_15570;
wire n_15562;
wire n_17207;
wire n_1327;
wire n_19000;
wire n_7729;
wire n_246;
wire n_19622;
wire n_1554;
wire n_4494;
wire n_6436;
wire n_16987;
wire n_18337;
wire n_2380;
wire n_20320;
wire n_6699;
wire n_12926;
wire n_14809;
wire n_4579;
wire n_14725;
wire n_16892;
wire n_4811;
wire n_19717;
wire n_6874;
wire n_6259;
wire n_9340;
wire n_16527;
wire n_17963;
wire n_6677;
wire n_12161;
wire n_3432;
wire n_11735;
wire n_20450;
wire n_4282;
wire n_1196;
wire n_8769;
wire n_6764;
wire n_10324;
wire n_11189;
wire n_8815;
wire n_12044;
wire n_748;
wire n_9303;
wire n_1785;
wire n_3057;
wire n_8261;
wire n_13104;
wire n_19730;
wire n_2287;
wire n_7139;
wire n_5727;
wire n_16819;
wire n_16612;
wire n_761;
wire n_5946;
wire n_20309;
wire n_3778;
wire n_9722;
wire n_12155;
wire n_15664;
wire n_4974;
wire n_12373;
wire n_5975;
wire n_19376;
wire n_14579;
wire n_17930;
wire n_4569;
wire n_8665;
wire n_15847;
wire n_5097;
wire n_7751;
wire n_2234;
wire n_18763;
wire n_20352;
wire n_14718;
wire n_4384;
wire n_19253;
wire n_2741;
wire n_3114;
wire n_18298;
wire n_888;
wire n_13116;
wire n_19781;
wire n_2203;
wire n_14589;
wire n_5246;
wire n_236;
wire n_12386;
wire n_14257;
wire n_16492;
wire n_16811;
wire n_3836;
wire n_8835;
wire n_18645;
wire n_20354;
wire n_10688;
wire n_16771;
wire n_1215;
wire n_12964;
wire n_20069;
wire n_16404;
wire n_15099;
wire n_20144;
wire n_779;
wire n_2205;
wire n_7579;
wire n_16874;
wire n_4025;
wire n_11687;
wire n_20157;
wire n_4121;
wire n_8870;
wire n_7155;
wire n_4313;
wire n_6475;
wire n_7699;
wire n_15951;
wire n_6103;
wire n_5546;
wire n_232;
wire n_6394;
wire n_8781;
wire n_18618;
wire n_14102;
wire n_20438;
wire n_17196;
wire n_4246;
wire n_12267;
wire n_15803;
wire n_8365;
wire n_3690;
wire n_2483;
wire n_4532;
wire n_13780;
wire n_16699;
wire n_19844;
wire n_7194;
wire n_4049;
wire n_6752;
wire n_6426;
wire n_984;
wire n_5626;
wire n_8025;
wire n_8502;
wire n_7612;
wire n_16999;
wire n_18843;
wire n_11120;
wire n_6350;
wire n_19702;
wire n_7736;
wire n_16040;
wire n_14259;
wire n_5921;
wire n_20030;
wire n_3596;
wire n_4537;
wire n_6159;
wire n_13360;
wire n_2429;
wire n_8479;
wire n_14214;
wire n_15558;
wire n_3521;
wire n_802;
wire n_17306;
wire n_6235;
wire n_17996;
wire n_2360;
wire n_12647;
wire n_7662;
wire n_15340;
wire n_16061;
wire n_7773;
wire n_5340;
wire n_3947;
wire n_16776;
wire n_13048;
wire n_13563;
wire n_17905;
wire n_7555;
wire n_1194;
wire n_4506;
wire n_19764;
wire n_2742;
wire n_3695;
wire n_12060;
wire n_3976;
wire n_18254;
wire n_10199;
wire n_8658;
wire n_11910;
wire n_15377;
wire n_15583;
wire n_13347;
wire n_5925;
wire n_2909;
wire n_8866;
wire n_8061;
wire n_5730;
wire n_16623;
wire n_17186;
wire n_13111;
wire n_15563;
wire n_10117;
wire n_12716;
wire n_467;
wire n_16341;
wire n_16679;
wire n_13456;
wire n_10198;
wire n_7157;
wire n_13237;
wire n_15448;
wire n_857;
wire n_7411;
wire n_19716;
wire n_16851;
wire n_2221;
wire n_588;
wire n_7871;
wire n_12051;
wire n_1010;
wire n_6477;
wire n_15298;
wire n_11533;
wire n_8652;
wire n_534;
wire n_7198;
wire n_1578;
wire n_9904;
wire n_17891;
wire n_19182;
wire n_1557;
wire n_3945;
wire n_6184;
wire n_730;
wire n_5817;
wire n_10973;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_4278;
wire n_5586;
wire n_11036;
wire n_3433;
wire n_17362;
wire n_4463;
wire n_10267;
wire n_10551;
wire n_18589;
wire n_17029;
wire n_3833;
wire n_2774;
wire n_17924;
wire n_18323;
wire n_13127;
wire n_18004;
wire n_4129;
wire n_11002;
wire n_19637;
wire n_5032;
wire n_14075;
wire n_9032;
wire n_6313;
wire n_18884;
wire n_16184;
wire n_3965;
wire n_7145;
wire n_12325;
wire n_9245;
wire n_5065;
wire n_9357;
wire n_3085;
wire n_19060;
wire n_5826;
wire n_15766;
wire n_18121;
wire n_2991;
wire n_16759;
wire n_14530;
wire n_17724;
wire n_19773;
wire n_7994;
wire n_14206;
wire n_17328;
wire n_4703;
wire n_7349;
wire n_9598;
wire n_14481;
wire n_17993;
wire n_15044;
wire n_12504;
wire n_12602;
wire n_12062;
wire n_15375;
wire n_16100;
wire n_12335;
wire n_12949;
wire n_13611;
wire n_801;
wire n_4452;
wire n_15268;
wire n_4649;
wire n_5315;
wire n_10487;
wire n_5362;
wire n_2157;
wire n_10960;
wire n_6141;
wire n_18540;
wire n_20409;
wire n_3849;
wire n_10931;
wire n_19831;
wire n_11574;
wire n_15049;
wire n_15181;
wire n_8168;
wire n_3257;
wire n_7190;
wire n_14870;
wire n_1387;
wire n_12322;
wire n_1151;
wire n_14196;
wire n_2317;
wire n_10236;
wire n_5524;
wire n_11776;
wire n_11205;
wire n_20169;
wire n_11650;
wire n_5818;
wire n_5963;
wire n_19197;
wire n_12179;
wire n_14439;
wire n_20229;
wire n_9896;
wire n_11856;
wire n_14825;
wire n_11536;
wire n_5950;
wire n_1192;
wire n_14914;
wire n_1844;
wire n_10283;
wire n_5057;
wire n_3030;
wire n_19865;
wire n_5838;
wire n_6324;
wire n_13437;
wire n_15623;
wire n_2838;
wire n_5325;
wire n_16696;
wire n_20516;
wire n_18865;
wire n_2926;
wire n_8411;
wire n_2019;
wire n_5102;
wire n_16733;
wire n_18799;
wire n_13221;
wire n_2074;
wire n_2919;
wire n_11163;
wire n_13657;
wire n_945;
wire n_14099;
wire n_15632;
wire n_16245;
wire n_11419;
wire n_12095;
wire n_9018;
wire n_13990;
wire n_16302;
wire n_13663;
wire n_6660;
wire n_13298;
wire n_9055;
wire n_4347;
wire n_14939;
wire n_11740;
wire n_17471;
wire n_8444;
wire n_20369;
wire n_17227;
wire n_5819;
wire n_2480;
wire n_7008;
wire n_12392;
wire n_11979;
wire n_7596;
wire n_20579;
wire n_6280;
wire n_18090;
wire n_18626;
wire n_2786;
wire n_10759;
wire n_9036;
wire n_9551;
wire n_13210;
wire n_19960;
wire n_18211;
wire n_8977;
wire n_20025;
wire n_15797;
wire n_9962;
wire n_2873;
wire n_11104;
wire n_3452;
wire n_3107;
wire n_11537;
wire n_13814;
wire n_18993;
wire n_12707;
wire n_14861;
wire n_7686;
wire n_1421;
wire n_15194;
wire n_1936;
wire n_5337;
wire n_18894;
wire n_15572;
wire n_12424;
wire n_1660;
wire n_3047;
wire n_11699;
wire n_8125;
wire n_14811;
wire n_17608;
wire n_10226;
wire n_6526;
wire n_1088;
wire n_17401;
wire n_7196;
wire n_3347;
wire n_907;
wire n_14864;
wire n_4110;
wire n_17936;
wire n_16643;
wire n_1658;
wire n_12107;
wire n_10161;
wire n_9842;
wire n_9614;
wire n_3999;
wire n_16024;
wire n_10699;
wire n_4751;
wire n_7846;
wire n_5151;
wire n_8598;
wire n_7256;
wire n_281;
wire n_16078;
wire n_7331;
wire n_13509;
wire n_17637;
wire n_5522;
wire n_5828;
wire n_7342;
wire n_14791;
wire n_14485;
wire n_10606;
wire n_11164;
wire n_4296;
wire n_12203;
wire n_7147;
wire n_5902;
wire n_512;
wire n_12359;
wire n_19175;
wire n_5063;
wire n_9037;
wire n_1328;
wire n_15983;
wire n_12548;
wire n_15874;
wire n_3900;
wire n_3732;
wire n_14461;
wire n_2832;
wire n_4226;
wire n_1762;
wire n_13958;
wire n_17619;
wire n_3980;
wire n_4366;
wire n_6863;
wire n_10012;
wire n_13754;
wire n_12985;
wire n_4445;
wire n_20087;
wire n_2692;
wire n_16191;
wire n_14171;
wire n_6768;
wire n_4456;
wire n_15212;
wire n_15977;
wire n_9128;
wire n_9872;
wire n_14380;
wire n_10310;
wire n_15896;
wire n_6151;
wire n_16843;
wire n_7110;
wire n_5476;
wire n_17273;
wire n_13920;
wire n_18119;
wire n_2922;
wire n_10097;
wire n_3882;
wire n_2068;
wire n_8915;
wire n_16509;
wire n_9866;
wire n_9858;
wire n_2072;
wire n_586;
wire n_423;
wire n_4375;
wire n_13977;
wire n_8727;
wire n_18494;
wire n_3935;
wire n_5130;
wire n_16538;
wire n_11662;
wire n_1726;
wire n_16992;
wire n_2878;
wire n_18065;
wire n_3012;
wire n_10266;
wire n_17949;
wire n_4877;
wire n_20099;
wire n_2641;
wire n_7734;
wire n_8955;
wire n_178;
wire n_20001;
wire n_17781;
wire n_12384;
wire n_15438;
wire n_11260;
wire n_3298;
wire n_11351;
wire n_4467;
wire n_195;
wire n_780;
wire n_15611;
wire n_14388;
wire n_12249;
wire n_2350;
wire n_14977;
wire n_10628;
wire n_13429;
wire n_4220;
wire n_11775;
wire n_5281;
wire n_7905;
wire n_10769;
wire n_10256;
wire n_1654;
wire n_13999;
wire n_14037;
wire n_11706;
wire n_11800;
wire n_18382;
wire n_1588;
wire n_11642;
wire n_20235;
wire n_4381;
wire n_11143;
wire n_17103;
wire n_11074;
wire n_6831;
wire n_16352;
wire n_18713;
wire n_18032;
wire n_11934;
wire n_4473;
wire n_6043;
wire n_687;
wire n_7677;
wire n_5457;
wire n_10396;
wire n_13919;
wire n_19357;
wire n_190;
wire n_13642;
wire n_8404;
wire n_8997;
wire n_6584;
wire n_11084;
wire n_1709;
wire n_10693;
wire n_2657;
wire n_15872;
wire n_13240;
wire n_20336;
wire n_949;
wire n_3500;
wire n_12578;
wire n_4589;
wire n_12194;
wire n_2972;
wire n_7519;
wire n_7400;
wire n_15649;
wire n_9724;
wire n_9281;
wire n_10101;
wire n_15863;
wire n_6581;
wire n_19690;
wire n_2279;
wire n_161;
wire n_7013;
wire n_14150;
wire n_12125;
wire n_7290;
wire n_18830;
wire n_595;
wire n_4921;
wire n_9687;
wire n_18052;
wire n_19108;
wire n_9426;
wire n_2712;
wire n_7889;
wire n_9102;
wire n_11526;
wire n_16115;
wire n_14128;
wire n_11851;
wire n_898;
wire n_18983;
wire n_17323;
wire n_6965;
wire n_9144;
wire n_18191;
wire n_7461;
wire n_15133;
wire n_16885;
wire n_4137;
wire n_9521;
wire n_15288;
wire n_16900;
wire n_13040;
wire n_963;
wire n_7278;
wire n_6509;
wire n_7454;
wire n_11253;
wire n_17102;
wire n_15527;
wire n_12861;
wire n_17443;
wire n_16146;
wire n_16654;
wire n_3400;
wire n_1521;
wire n_12918;
wire n_1366;
wire n_18332;
wire n_5501;
wire n_5342;
wire n_4345;
wire n_18145;
wire n_13353;
wire n_8648;
wire n_12388;
wire n_12102;
wire n_16991;
wire n_18051;
wire n_19051;
wire n_4664;
wire n_13716;
wire n_7069;
wire n_7904;
wire n_11691;
wire n_14408;
wire n_9410;
wire n_2643;
wire n_5748;
wire n_12865;
wire n_10712;
wire n_4713;
wire n_7168;
wire n_17604;
wire n_18765;
wire n_7970;
wire n_7091;
wire n_3166;
wire n_3435;
wire n_842;
wire n_10972;
wire n_6359;
wire n_1432;
wire n_20564;
wire n_10945;
wire n_8800;
wire n_10845;
wire n_8229;
wire n_18743;
wire n_14863;
wire n_5811;
wire n_6766;
wire n_1035;
wire n_7629;
wire n_9735;
wire n_18831;
wire n_5397;
wire n_20344;
wire n_20541;
wire n_14711;
wire n_9802;
wire n_1448;
wire n_14373;
wire n_8107;
wire n_12992;
wire n_11108;
wire n_11004;
wire n_2445;
wire n_6519;
wire n_15752;
wire n_11686;
wire n_6530;
wire n_4440;
wire n_10566;
wire n_17798;
wire n_19592;
wire n_16568;
wire n_17581;
wire n_18906;
wire n_12104;
wire n_17954;
wire n_6402;
wire n_12469;
wire n_19554;
wire n_15829;
wire n_19568;
wire n_7326;
wire n_17522;
wire n_7067;
wire n_14835;
wire n_15391;
wire n_16226;
wire n_14871;
wire n_8691;
wire n_14907;
wire n_3342;
wire n_6748;
wire n_11719;
wire n_19307;
wire n_16685;
wire n_19498;
wire n_3656;
wire n_16979;
wire n_1424;
wire n_18282;
wire n_15358;
wire n_14636;
wire n_1507;
wire n_2482;
wire n_8026;
wire n_9638;
wire n_16069;
wire n_7528;
wire n_20101;
wire n_8174;
wire n_13524;
wire n_912;
wire n_11175;
wire n_10040;
wire n_2661;
wire n_8861;
wire n_5359;
wire n_8644;
wire n_931;
wire n_1791;
wire n_12304;
wire n_15156;
wire n_1897;
wire n_2064;
wire n_7117;
wire n_13138;
wire n_18490;
wire n_6205;
wire n_20141;
wire n_7136;
wire n_6754;
wire n_12692;
wire n_1334;
wire n_7939;
wire n_13602;
wire n_17436;
wire n_16785;
wire n_9612;
wire n_10790;
wire n_14919;
wire n_16653;
wire n_6723;
wire n_9108;
wire n_16692;
wire n_6440;
wire n_7436;
wire n_14101;
wire n_9376;
wire n_8446;
wire n_17654;
wire n_3534;
wire n_20396;
wire n_12996;
wire n_15171;
wire n_19711;
wire n_13625;
wire n_12643;
wire n_3944;
wire n_6124;
wire n_7685;
wire n_7363;
wire n_8192;
wire n_19265;
wire n_1939;
wire n_8197;
wire n_2209;
wire n_6622;
wire n_11521;
wire n_20463;
wire n_12827;
wire n_12678;
wire n_15868;
wire n_1053;
wire n_17249;
wire n_9779;
wire n_7747;
wire n_8082;
wire n_8730;
wire n_15533;
wire n_266;
wire n_6528;
wire n_15165;
wire n_13475;
wire n_15079;
wire n_19822;
wire n_13859;
wire n_18640;
wire n_1745;
wire n_3479;
wire n_12713;
wire n_13144;
wire n_18129;
wire n_488;
wire n_19488;
wire n_10660;
wire n_7430;
wire n_18560;
wire n_9937;
wire n_5679;
wire n_7912;
wire n_5100;
wire n_16749;
wire n_5973;
wire n_8281;
wire n_20347;
wire n_4807;
wire n_1243;
wire n_301;
wire n_2928;
wire n_5166;
wire n_19437;
wire n_18876;
wire n_20174;
wire n_19430;
wire n_11428;
wire n_2822;
wire n_17626;
wire n_1281;
wire n_11677;
wire n_7281;
wire n_9717;
wire n_13577;
wire n_2572;
wire n_1520;
wire n_3126;
wire n_18523;
wire n_1419;
wire n_19176;
wire n_5688;
wire n_19970;
wire n_13769;
wire n_18044;
wire n_4676;
wire n_13672;
wire n_19036;
wire n_17600;
wire n_6763;
wire n_8956;
wire n_7858;
wire n_663;
wire n_4880;
wire n_20203;
wire n_6542;
wire n_15681;
wire n_2781;
wire n_4126;
wire n_17262;
wire n_1696;
wire n_6556;
wire n_20245;
wire n_12374;
wire n_4813;
wire n_5542;
wire n_1030;
wire n_8998;
wire n_10538;
wire n_1790;
wire n_4014;
wire n_13342;
wire n_18856;
wire n_9123;
wire n_17374;
wire n_6471;
wire n_5949;
wire n_15545;
wire n_4048;
wire n_14924;
wire n_4444;
wire n_11867;
wire n_12796;
wire n_3919;
wire n_16053;
wire n_19185;
wire n_15708;
wire n_19441;
wire n_11716;
wire n_8979;
wire n_7245;
wire n_18858;
wire n_6675;
wire n_6270;
wire n_18111;
wire n_6808;
wire n_2884;
wire n_16091;
wire n_20326;
wire n_11886;
wire n_7006;
wire n_16264;
wire n_14160;
wire n_6245;
wire n_14932;
wire n_17231;
wire n_3797;
wire n_10925;
wire n_20190;
wire n_4770;
wire n_11158;
wire n_9861;
wire n_15878;
wire n_2549;
wire n_4690;
wire n_14390;
wire n_18678;
wire n_8264;
wire n_7381;
wire n_16160;
wire n_12078;
wire n_15647;
wire n_9832;
wire n_19925;
wire n_20547;
wire n_6580;
wire n_18790;
wire n_9898;
wire n_5500;
wire n_6412;
wire n_18410;
wire n_19959;
wire n_183;
wire n_13293;
wire n_3967;
wire n_6437;
wire n_14381;
wire n_2526;
wire n_15709;
wire n_18590;
wire n_8408;
wire n_3277;
wire n_10661;
wire n_9495;
wire n_10028;
wire n_13878;
wire n_15000;
wire n_11771;
wire n_16870;
wire n_19082;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_13833;
wire n_16518;
wire n_1960;
wire n_2694;
wire n_1686;
wire n_9867;
wire n_6059;
wire n_14441;
wire n_9688;
wire n_5094;
wire n_10967;
wire n_7870;
wire n_3228;
wire n_18377;
wire n_3657;
wire n_20208;
wire n_1287;
wire n_6117;
wire n_11828;
wire n_12326;
wire n_1586;
wire n_14264;
wire n_19317;
wire n_14115;
wire n_16635;
wire n_3464;
wire n_380;
wire n_8963;
wire n_4380;
wire n_4996;
wire n_5247;
wire n_4398;
wire n_4193;
wire n_3570;
wire n_12309;
wire n_7399;
wire n_3828;
wire n_1539;
wire n_13953;
wire n_7482;
wire n_19830;
wire n_14847;
wire n_10312;
wire n_4090;
wire n_18308;
wire n_9223;
wire n_17465;
wire n_15930;
wire n_13226;
wire n_5931;
wire n_2371;
wire n_19416;
wire n_17943;
wire n_662;
wire n_16433;
wire n_3262;
wire n_11244;
wire n_4008;
wire n_18577;
wire n_14432;
wire n_1642;
wire n_10209;
wire n_13253;
wire n_4689;
wire n_8183;
wire n_19936;
wire n_16098;
wire n_4547;
wire n_11245;
wire n_13354;
wire n_6085;
wire n_12422;
wire n_15616;
wire n_17614;
wire n_3329;
wire n_14422;
wire n_9694;
wire n_3826;
wire n_16636;
wire n_9948;
wire n_14630;
wire n_17048;
wire n_3681;
wire n_18966;
wire n_19390;
wire n_19729;
wire n_10887;
wire n_16876;
wire n_5883;
wire n_6554;
wire n_12146;
wire n_5754;
wire n_6560;
wire n_14055;
wire n_1720;
wire n_12136;
wire n_17046;
wire n_16138;
wire n_12399;
wire n_942;
wire n_12342;
wire n_7414;
wire n_9744;
wire n_9548;
wire n_8973;
wire n_6448;
wire n_1964;
wire n_12378;
wire n_19155;
wire n_12533;
wire n_5434;
wire n_7431;
wire n_5934;
wire n_12178;
wire n_18871;
wire n_20192;
wire n_11346;
wire n_17210;
wire n_2626;
wire n_5880;
wire n_18206;
wire n_19851;
wire n_14810;
wire n_8249;
wire n_12257;
wire n_3528;
wire n_15770;
wire n_13394;
wire n_13391;
wire n_14680;
wire n_8234;
wire n_20442;
wire n_16835;
wire n_1066;
wire n_18438;
wire n_16863;
wire n_9280;
wire n_18285;
wire n_13263;
wire n_14877;
wire n_19815;
wire n_5145;
wire n_15203;
wire n_1229;
wire n_11491;
wire n_14048;
wire n_2427;
wire n_11772;
wire n_16063;
wire n_16237;
wire n_16112;
wire n_15891;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_12769;
wire n_4190;
wire n_5149;
wire n_12641;
wire n_10765;
wire n_3375;
wire n_15263;
wire n_11792;
wire n_20076;
wire n_18776;
wire n_2668;
wire n_8558;
wire n_10489;
wire n_12421;
wire n_2128;
wire n_7274;
wire n_10159;
wire n_14351;
wire n_7466;
wire n_1002;
wire n_13310;
wire n_2508;
wire n_11568;
wire n_2054;
wire n_7429;
wire n_11766;
wire n_11038;
wire n_13798;
wire n_16894;
wire n_18890;
wire n_17294;
wire n_16932;
wire n_15842;
wire n_14822;
wire n_2758;
wire n_8813;
wire n_10356;
wire n_17461;
wire n_18216;
wire n_10173;
wire n_20010;
wire n_4789;
wire n_19162;
wire n_12311;
wire n_14374;
wire n_2241;
wire n_6555;
wire n_9448;
wire n_14815;
wire n_10739;
wire n_8470;
wire n_1690;
wire n_5341;
wire n_16480;
wire n_4512;
wire n_20062;
wire n_1378;
wire n_17657;
wire n_14831;
wire n_11170;
wire n_17683;
wire n_11758;
wire n_1542;
wire n_9396;
wire n_19486;
wire n_14450;
wire n_7061;
wire n_12480;
wire n_14192;
wire n_1716;
wire n_278;
wire n_9053;
wire n_15504;
wire n_11893;
wire n_10573;
wire n_3303;
wire n_4324;
wire n_10850;
wire n_384;
wire n_9185;
wire n_19697;
wire n_13376;
wire n_2905;
wire n_8092;
wire n_13864;
wire n_3954;
wire n_15279;
wire n_11456;
wire n_10546;
wire n_5622;
wire n_3160;
wire n_6574;
wire n_20270;
wire n_6571;
wire n_17484;
wire n_143;
wire n_9151;
wire n_7824;
wire n_17202;
wire n_18080;
wire n_698;
wire n_20444;
wire n_13236;
wire n_3569;
wire n_14299;
wire n_7094;
wire n_2528;
wire n_16320;
wire n_4639;
wire n_7036;
wire n_13777;
wire n_19359;
wire n_20467;
wire n_1730;
wire n_814;
wire n_5779;
wire n_2020;
wire n_6260;
wire n_7413;
wire n_16803;
wire n_17229;
wire n_6286;
wire n_8267;
wire n_4023;
wire n_18929;
wire n_721;
wire n_7175;
wire n_6019;
wire n_4344;
wire n_9978;
wire n_11914;
wire n_9670;
wire n_3154;
wire n_19964;
wire n_9334;
wire n_15131;
wire n_20064;
wire n_3898;
wire n_12531;
wire n_4391;
wire n_11302;
wire n_946;
wire n_1303;
wire n_19931;
wire n_19006;
wire n_4095;
wire n_9413;
wire n_12727;
wire n_20043;
wire n_15509;
wire n_3551;
wire n_3064;
wire n_11707;
wire n_1689;
wire n_7697;
wire n_1944;
wire n_13835;
wire n_16260;
wire n_7547;
wire n_6013;
wire n_13815;
wire n_20515;
wire n_9557;
wire n_15957;
wire n_16319;
wire n_448;
wire n_3853;
wire n_17259;
wire n_20355;
wire n_14039;
wire n_6348;
wire n_6744;
wire n_18578;
wire n_8582;
wire n_6293;
wire n_5068;
wire n_234;
wire n_6049;
wire n_1460;
wire n_9762;
wire n_8957;
wire n_18646;
wire n_15793;
wire n_6558;
wire n_20323;
wire n_12227;
wire n_12258;
wire n_14117;
wire n_18209;
wire n_2437;
wire n_2444;
wire n_9271;
wire n_17747;
wire n_3035;
wire n_13688;
wire n_4166;
wire n_11396;
wire n_15196;
wire n_16176;
wire n_20207;
wire n_9483;
wire n_19649;
wire n_1058;
wire n_19435;
wire n_19769;
wire n_14754;
wire n_19768;
wire n_15020;
wire n_2934;
wire n_6091;
wire n_14252;
wire n_15830;
wire n_12583;
wire n_6551;
wire n_7691;
wire n_8747;
wire n_9539;
wire n_4817;
wire n_2014;
wire n_9385;
wire n_1584;
wire n_13462;
wire n_5381;
wire n_9785;
wire n_3468;
wire n_8922;
wire n_9027;
wire n_12750;
wire n_4383;
wire n_6995;
wire n_5696;
wire n_455;
wire n_4486;
wire n_19315;
wire n_9233;
wire n_20544;
wire n_3024;
wire n_16895;
wire n_10282;
wire n_17602;
wire n_4529;
wire n_500;
wire n_15142;
wire n_291;
wire n_10913;
wire n_18803;
wire n_18409;
wire n_17838;
wire n_15991;
wire n_5823;
wire n_13388;
wire n_2800;
wire n_13731;
wire n_10703;
wire n_9666;
wire n_14503;
wire n_12248;
wire n_8678;
wire n_10565;
wire n_10011;
wire n_17754;
wire n_14886;
wire n_7993;
wire n_20223;
wire n_7181;
wire n_9865;
wire n_3161;
wire n_2799;
wire n_14644;
wire n_11715;
wire n_7071;
wire n_15454;
wire n_15213;
wire n_10642;
wire n_756;
wire n_18859;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_19946;
wire n_18428;
wire n_12181;
wire n_18670;
wire n_14560;
wire n_17257;
wire n_19726;
wire n_3992;
wire n_14829;
wire n_11007;
wire n_15473;
wire n_249;
wire n_19864;
wire n_15584;
wire n_3125;
wire n_10316;
wire n_9795;
wire n_18386;
wire n_4684;
wire n_3116;
wire n_6429;
wire n_6407;
wire n_16515;
wire n_5027;
wire n_17914;
wire n_10479;
wire n_13660;
wire n_19280;
wire n_6801;
wire n_1921;
wire n_18099;
wire n_5630;
wire n_12738;
wire n_4057;
wire n_15062;
wire n_1170;
wire n_20402;
wire n_5379;
wire n_11599;
wire n_308;
wire n_3444;
wire n_6113;
wire n_10070;
wire n_16178;
wire n_1890;
wire n_20276;
wire n_18841;
wire n_2477;
wire n_17304;
wire n_18393;
wire n_14983;
wire n_2333;
wire n_8439;
wire n_18434;
wire n_9641;
wire n_1089;
wire n_12755;
wire n_18522;
wire n_12059;
wire n_18541;
wire n_18257;
wire n_15845;
wire n_5018;
wire n_6129;
wire n_6518;
wire n_20401;
wire n_9138;
wire n_18072;
wire n_18048;
wire n_7537;
wire n_10516;
wire n_8675;
wire n_1616;
wire n_15924;
wire n_17906;
wire n_12567;
wire n_9367;
wire n_15130;
wire n_4197;
wire n_4482;
wire n_2547;
wire n_2415;
wire n_11887;
wire n_17852;
wire n_17442;
wire n_10026;
wire n_9729;
wire n_5073;
wire n_827;
wire n_12471;
wire n_12451;
wire n_17243;
wire n_15740;
wire n_20048;
wire n_9411;
wire n_3660;
wire n_3766;
wire n_12507;
wire n_1027;
wire n_3266;
wire n_3574;
wire n_14564;
wire n_11277;
wire n_4907;
wire n_5077;
wire n_18416;
wire n_20133;
wire n_17606;
wire n_7410;
wire n_365;
wire n_8777;
wire n_2534;
wire n_4975;
wire n_13581;
wire n_2451;
wire n_12972;
wire n_13789;
wire n_4815;
wire n_14511;
wire n_13286;
wire n_9951;
wire n_396;
wire n_19023;
wire n_9424;
wire n_480;
wire n_4134;
wire n_10507;
wire n_11968;
wire n_19003;
wire n_1238;
wire n_4092;
wire n_10045;
wire n_20179;
wire n_11335;
wire n_18606;
wire n_13988;
wire n_4755;
wire n_4960;
wire n_1700;
wire n_15272;
wire n_4933;
wire n_17169;
wire n_13609;
wire n_4591;
wire n_5528;
wire n_16886;
wire n_5111;
wire n_13679;
wire n_11785;
wire n_873;
wire n_10417;
wire n_3946;
wire n_12841;
wire n_12855;
wire n_17370;
wire n_15834;
wire n_13276;
wire n_8938;
wire n_4474;
wire n_5665;
wire n_16058;
wire n_2509;
wire n_11801;
wire n_16994;
wire n_16519;
wire n_3757;
wire n_17810;
wire n_1704;
wire n_250;
wire n_4884;
wire n_14830;
wire n_7867;
wire n_14281;
wire n_14594;
wire n_18213;
wire n_6135;
wire n_17303;
wire n_20263;
wire n_3678;
wire n_6814;
wire n_10557;
wire n_8669;
wire n_7525;
wire n_19219;
wire n_7257;
wire n_9372;
wire n_4692;
wire n_6791;
wire n_616;
wire n_3165;
wire n_13704;
wire n_11915;
wire n_11016;
wire n_9326;
wire n_14976;
wire n_1902;
wire n_1735;
wire n_3890;
wire n_641;
wire n_3750;
wire n_7650;
wire n_17297;
wire n_19872;
wire n_13043;
wire n_4311;
wire n_4722;
wire n_17260;
wire n_12620;
wire n_12632;
wire n_20198;
wire n_20456;
wire n_6309;
wire n_19618;
wire n_11303;
wire n_405;
wire n_213;
wire n_6733;
wire n_19047;
wire n_20122;
wire n_1094;
wire n_5430;
wire n_5942;
wire n_9902;
wire n_4820;
wire n_19910;
wire n_9900;
wire n_17367;
wire n_18937;
wire n_15521;
wire n_18415;
wire n_7202;
wire n_12416;
wire n_8265;
wire n_4619;
wire n_5762;
wire n_11609;
wire n_1961;
wire n_18287;
wire n_16464;
wire n_5036;
wire n_4221;
wire n_19597;
wire n_3297;
wire n_12494;
wire n_10327;
wire n_13826;
wire n_7605;
wire n_11556;
wire n_15140;
wire n_11529;
wire n_10437;
wire n_10021;
wire n_16673;
wire n_9146;
wire n_15753;
wire n_2996;
wire n_8131;
wire n_8941;
wire n_5014;
wire n_17093;
wire n_17685;
wire n_16357;
wire n_12623;
wire n_11444;
wire n_659;
wire n_6269;
wire n_5233;
wire n_12213;
wire n_6654;
wire n_9358;
wire n_3164;
wire n_9565;
wire n_8257;
wire n_13072;
wire n_18120;
wire n_7726;
wire n_5436;
wire n_17026;
wire n_13839;
wire n_594;
wire n_6120;
wire n_6068;
wire n_4141;
wire n_13954;
wire n_8799;
wire n_2850;
wire n_572;
wire n_6641;
wire n_5789;
wire n_2104;
wire n_19215;
wire n_10124;
wire n_19595;
wire n_14689;
wire n_10245;
wire n_14132;
wire n_10905;
wire n_11235;
wire n_19020;
wire n_6399;
wire n_4499;
wire n_5195;
wire n_9563;
wire n_17077;
wire n_17702;
wire n_11166;
wire n_20310;
wire n_7031;
wire n_9285;
wire n_263;
wire n_18093;
wire n_16595;
wire n_7763;
wire n_1543;
wire n_8033;
wire n_1599;
wire n_15172;
wire n_4458;
wire n_19470;
wire n_19720;
wire n_5103;
wire n_8393;
wire n_16561;
wire n_10784;
wire n_1876;
wire n_4107;
wire n_8463;
wire n_8153;
wire n_10944;
wire n_10211;
wire n_18554;
wire n_18077;
wire n_12431;
wire n_11855;
wire n_6790;
wire n_3099;
wire n_17628;
wire n_13799;
wire n_16084;
wire n_13854;
wire n_18250;
wire n_19843;
wire n_15380;
wire n_2457;
wire n_6686;
wire n_15956;
wire n_4119;
wire n_18835;
wire n_20035;
wire n_11787;
wire n_5958;
wire n_16059;
wire n_8103;
wire n_2971;
wire n_20421;
wire n_715;
wire n_4526;
wire n_14752;
wire n_5792;
wire n_6183;
wire n_11544;
wire n_15447;
wire n_10730;
wire n_2028;
wire n_1069;
wire n_10564;
wire n_8682;
wire n_20307;
wire n_7655;
wire n_18276;
wire n_4485;
wire n_1504;
wire n_11509;
wire n_19191;
wire n_11960;
wire n_1801;
wire n_3917;
wire n_19905;
wire n_7878;
wire n_9514;
wire n_6210;
wire n_6500;
wire n_12465;
wire n_2206;
wire n_13532;
wire n_11029;
wire n_13118;
wire n_17390;
wire n_5739;
wire n_10951;
wire n_12152;
wire n_19415;
wire n_6785;
wire n_10454;
wire n_15401;
wire n_13339;
wire n_4940;
wire n_8039;
wire n_5757;
wire n_19323;
wire n_8916;
wire n_10087;
wire n_3510;
wire n_10146;
wire n_12959;
wire n_9946;
wire n_9885;
wire n_6849;
wire n_20482;
wire n_8162;
wire n_18263;
wire n_7457;
wire n_19982;
wire n_8744;
wire n_5488;
wire n_10701;
wire n_3827;
wire n_891;
wire n_2067;
wire n_7752;
wire n_15775;
wire n_4245;
wire n_17346;
wire n_8286;
wire n_9015;
wire n_20002;
wire n_6452;
wire n_16408;
wire n_20362;
wire n_1008;
wire n_6611;
wire n_4560;
wire n_18828;
wire n_4899;
wire n_18297;
wire n_5471;
wire n_11433;
wire n_10592;
wire n_5164;
wire n_18130;
wire n_7207;
wire n_8218;
wire n_17978;
wire n_1767;
wire n_8537;
wire n_10126;
wire n_14421;
wire n_15890;
wire n_4663;
wire n_2893;
wire n_13653;
wire n_5484;
wire n_12566;
wire n_6227;
wire n_13680;
wire n_3421;
wire n_16077;
wire n_9066;
wire n_10302;
wire n_12546;
wire n_13058;
wire n_18342;
wire n_12036;
wire n_17650;
wire n_8782;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_12911;
wire n_15715;
wire n_9857;
wire n_12781;
wire n_10057;
wire n_10882;
wire n_894;
wire n_9338;
wire n_353;
wire n_8144;
wire n_10435;
wire n_9542;
wire n_10921;
wire n_7171;
wire n_12061;
wire n_3922;
wire n_14585;
wire n_11085;
wire n_16541;
wire n_7068;
wire n_13649;
wire n_10609;
wire n_14804;
wire n_2554;
wire n_20015;
wire n_9783;
wire n_13806;
wire n_19542;
wire n_4934;
wire n_9404;
wire n_9916;
wire n_12645;
wire n_5526;
wire n_18351;
wire n_16198;
wire n_14466;
wire n_7777;
wire n_12138;
wire n_2765;
wire n_5403;
wire n_2590;
wire n_7652;
wire n_10220;
wire n_3150;
wire n_11347;
wire n_17635;
wire n_4479;
wire n_2608;
wire n_10550;
wire n_14673;
wire n_12365;
wire n_1959;
wire n_3133;
wire n_20334;
wire n_13738;
wire n_14972;
wire n_765;
wire n_1492;
wire n_16996;
wire n_9306;
wire n_14138;
wire n_1340;
wire n_10232;
wire n_10461;
wire n_14586;
wire n_7966;
wire n_8591;
wire n_8811;
wire n_19188;
wire n_1277;
wire n_14031;
wire n_5242;
wire n_10326;
wire n_8417;
wire n_2675;
wire n_5631;
wire n_19978;
wire n_6008;
wire n_3887;
wire n_12487;
wire n_7997;
wire n_6420;
wire n_20518;
wire n_4587;
wire n_1577;
wire n_12288;
wire n_17300;
wire n_1117;
wire n_12130;
wire n_13120;
wire n_19825;
wire n_3223;
wire n_16299;
wire n_12704;
wire n_12271;
wire n_7680;
wire n_15190;
wire n_16909;
wire n_12958;
wire n_8172;
wire n_19848;
wire n_19559;
wire n_9502;
wire n_6447;
wire n_5981;
wire n_3788;
wire n_4891;
wire n_19923;
wire n_14761;
wire n_6751;
wire n_2718;
wire n_15243;
wire n_20090;
wire n_1384;
wire n_11087;
wire n_11477;
wire n_3325;
wire n_2238;
wire n_8375;
wire n_8612;
wire n_4624;
wire n_8345;
wire n_13725;
wire n_3600;
wire n_6741;
wire n_11773;
wire n_12608;
wire n_8459;
wire n_5015;
wire n_1178;
wire n_2338;
wire n_19414;
wire n_17551;
wire n_19417;
wire n_9164;
wire n_7183;
wire n_13197;
wire n_10878;
wire n_18408;
wire n_7140;
wire n_20284;
wire n_14860;
wire n_10450;
wire n_623;
wire n_19609;
wire n_11472;
wire n_9114;
wire n_11978;
wire n_8515;
wire n_10529;
wire n_1502;
wire n_14685;
wire n_5773;
wire n_5482;
wire n_14892;
wire n_8812;
wire n_14505;
wire n_12254;
wire n_9392;
wire n_1250;
wire n_14531;
wire n_3615;
wire n_11538;
wire n_3087;
wire n_2121;
wire n_9698;
wire n_13435;
wire n_15408;
wire n_15173;
wire n_4015;
wire n_477;
wire n_9644;
wire n_11353;
wire n_18745;
wire n_2213;
wire n_2389;
wire n_9499;
wire n_2892;
wire n_6647;
wire n_4120;
wire n_6275;
wire n_14771;
wire n_1564;
wire n_5296;
wire n_3718;
wire n_7750;
wire n_11597;
wire n_537;
wire n_15902;
wire n_6277;
wire n_1919;
wire n_3705;
wire n_3211;
wire n_546;
wire n_10920;
wire n_14398;
wire n_3582;
wire n_11126;
wire n_4223;
wire n_5674;
wire n_18453;
wire n_5282;
wire n_9409;
wire n_18629;
wire n_1060;
wire n_20565;
wire n_1951;
wire n_17814;
wire n_12555;
wire n_11646;
wire n_1223;
wire n_5121;
wire n_9768;
wire n_6070;
wire n_1286;
wire n_12980;
wire n_9881;
wire n_5013;
wire n_6807;
wire n_7251;
wire n_4489;
wire n_7254;
wire n_18178;
wire n_12973;
wire n_3163;
wire n_17313;
wire n_13123;
wire n_14669;
wire n_5589;
wire n_12234;
wire n_10776;
wire n_7882;
wire n_16348;
wire n_16514;
wire n_17704;
wire n_10848;
wire n_20216;
wire n_2585;
wire n_5628;
wire n_4825;
wire n_2352;
wire n_7765;
wire n_11482;
wire n_1625;
wire n_5006;
wire n_7816;
wire n_2226;
wire n_2801;
wire n_10164;
wire n_15809;
wire n_1901;
wire n_3869;
wire n_15579;
wire n_18549;
wire n_18084;
wire n_15585;
wire n_3753;
wire n_12033;
wire n_1892;
wire n_1614;
wire n_3742;
wire n_14376;
wire n_20102;
wire n_3260;
wire n_20173;
wire n_9595;
wire n_18978;
wire n_15555;
wire n_13923;
wire n_13051;
wire n_11524;
wire n_17220;
wire n_9265;
wire n_8239;
wire n_16114;
wire n_13330;
wire n_2159;
wire n_2315;
wire n_11228;
wire n_5273;
wire n_7898;
wire n_18286;
wire n_9789;
wire n_5936;
wire n_7646;
wire n_20166;
wire n_17537;
wire n_3220;
wire n_14627;
wire n_13699;
wire n_6069;
wire n_171;
wire n_169;
wire n_19940;
wire n_7665;
wire n_9354;
wire n_14026;
wire n_10501;
wire n_2379;
wire n_17782;
wire n_19687;
wire n_9436;
wire n_18157;
wire n_8489;
wire n_4067;
wire n_4357;
wire n_10350;
wire n_12730;
wire n_6887;
wire n_18926;
wire n_16123;
wire n_13152;
wire n_17221;
wire n_4374;
wire n_6637;
wire n_9238;
wire n_358;
wire n_6633;
wire n_2420;
wire n_11031;
wire n_3722;
wire n_186;
wire n_4400;
wire n_17365;
wire n_9839;
wire n_18479;
wire n_15704;
wire n_7900;
wire n_6569;
wire n_10807;
wire n_12478;
wire n_2538;
wire n_724;
wire n_3250;
wire n_17265;
wire n_13545;
wire n_557;
wire n_13760;
wire n_1871;
wire n_13883;
wire n_10511;
wire n_7576;
wire n_19499;
wire n_11023;
wire n_3651;
wire n_7313;
wire n_2102;
wire n_10873;
wire n_14484;
wire n_7676;
wire n_18956;
wire n_9017;
wire n_4304;
wire n_15726;
wire n_14307;
wire n_2544;
wire n_8865;
wire n_15302;
wire n_10337;
wire n_7779;
wire n_8999;
wire n_1206;
wire n_11626;
wire n_12148;
wire n_16872;
wire n_6479;
wire n_10791;
wire n_10506;
wire n_16312;
wire n_16204;
wire n_8820;
wire n_16793;
wire n_16443;
wire n_6090;
wire n_20071;
wire n_18456;
wire n_5515;
wire n_3131;
wire n_18281;
wire n_12132;
wire n_1298;
wire n_10593;
wire n_5862;
wire n_16801;
wire n_2088;
wire n_12182;
wire n_12043;
wire n_10636;
wire n_16478;
wire n_18489;
wire n_5697;
wire n_2401;
wire n_18723;
wire n_8992;
wire n_8880;
wire n_8690;
wire n_2900;
wire n_6234;
wire n_3994;
wire n_1497;
wire n_7818;
wire n_11721;
wire n_13573;
wire n_19019;
wire n_6608;
wire n_9109;
wire n_5498;
wire n_2571;
wire n_3138;
wire n_7896;
wire n_12482;
wire n_18839;
wire n_15208;
wire n_6860;
wire n_12137;
wire n_12306;
wire n_11328;
wire n_2988;
wire n_1350;
wire n_11200;
wire n_14442;
wire n_15210;
wire n_4109;
wire n_16536;
wire n_19917;
wire n_13418;
wire n_5175;
wire n_7996;
wire n_986;
wire n_10533;
wire n_460;
wire n_5987;
wire n_16681;
wire n_10176;
wire n_19707;
wire n_7517;
wire n_8080;
wire n_450;
wire n_4150;
wire n_12345;
wire n_13551;
wire n_19135;
wire n_19178;
wire n_16060;
wire n_8772;
wire n_8786;
wire n_15597;
wire n_4643;
wire n_12694;
wire n_8083;
wire n_20060;
wire n_10155;
wire n_1332;
wire n_9805;
wire n_19799;
wire n_13593;
wire n_8157;
wire n_2346;
wire n_19660;
wire n_936;
wire n_3821;
wire n_13902;
wire n_19792;
wire n_3676;
wire n_4896;
wire n_3675;
wire n_9110;
wire n_18358;
wire n_5904;
wire n_599;
wire n_14468;
wire n_6062;
wire n_12550;
wire n_13861;
wire n_13350;
wire n_10051;
wire n_4209;
wire n_10414;
wire n_8344;
wire n_17597;
wire n_1341;
wire n_8120;
wire n_3003;
wire n_9075;
wire n_12961;
wire n_18882;
wire n_11496;
wire n_4128;
wire n_12225;
wire n_20118;
wire n_4271;
wire n_2258;
wire n_8621;
wire n_12884;
wire n_325;
wire n_5845;
wire n_20350;
wire n_19171;
wire n_6246;
wire n_8868;
wire n_8134;
wire n_4716;
wire n_12207;
wire n_9975;
wire n_1782;
wire n_5600;
wire n_12011;
wire n_707;
wire n_6053;
wire n_7252;
wire n_3246;
wire n_20031;
wire n_6843;
wire n_4715;
wire n_10626;
wire n_6901;
wire n_19014;
wire n_13273;
wire n_4694;
wire n_18855;
wire n_8101;
wire n_19751;
wire n_5448;
wire n_19954;
wire n_6489;
wire n_7402;
wire n_737;
wire n_3517;
wire n_3893;
wire n_19552;
wire n_11273;
wire n_138;
wire n_19089;
wire n_19993;
wire n_16954;
wire n_12472;
wire n_19526;
wire n_14035;
wire n_13218;
wire n_9081;
wire n_333;
wire n_4084;
wire n_9236;
wire n_6844;
wire n_11762;
wire n_459;
wire n_4850;
wire n_10156;
wire n_9607;
wire n_2840;
wire n_6779;
wire n_10774;
wire n_12332;
wire n_7216;
wire n_3855;
wire n_15990;
wire n_15364;
wire n_3091;
wire n_6543;
wire n_19585;
wire n_6178;
wire n_9621;
wire n_3398;
wire n_5685;
wire n_18075;
wire n_2793;
wire n_4235;
wire n_16117;
wire n_10398;
wire n_17947;
wire n_16459;
wire n_774;
wire n_17987;
wire n_18165;
wire n_15661;
wire n_20185;
wire n_17932;
wire n_7706;
wire n_1860;
wire n_5016;
wire n_20304;
wire n_479;
wire n_6458;
wire n_7642;
wire n_1777;
wire n_12506;
wire n_18356;
wire n_3308;
wire n_12718;
wire n_1600;
wire n_2253;
wire n_12638;
wire n_14116;
wire n_20391;
wire n_4799;
wire n_2261;
wire n_18710;
wire n_2516;
wire n_16453;
wire n_16645;
wire n_1177;
wire n_10470;
wire n_20156;
wire n_15034;
wire n_19808;
wire n_14240;
wire n_14504;
wire n_13449;
wire n_12747;
wire n_10625;
wire n_12561;
wire n_18420;
wire n_5514;
wire n_8388;
wire n_18469;
wire n_14730;
wire n_18732;
wire n_9589;
wire n_4543;
wire n_15110;
wire n_10445;
wire n_8988;
wire n_15025;
wire n_19329;
wire n_18161;
wire n_12900;
wire n_18761;
wire n_8569;
wire n_14598;
wire n_3255;
wire n_1401;
wire n_10679;
wire n_1516;
wire n_11323;
wire n_10799;
wire n_2029;
wire n_5890;
wire n_17228;
wire n_1394;
wire n_10585;
wire n_18519;
wire n_13696;
wire n_12948;
wire n_7931;
wire n_13322;
wire n_9092;
wire n_10034;
wire n_935;
wire n_9451;
wire n_11148;
wire n_18729;
wire n_13934;
wire n_6899;
wire n_19880;
wire n_7373;
wire n_7895;
wire n_676;
wire n_15331;
wire n_17109;
wire n_832;
wire n_13254;
wire n_3049;
wire n_15191;
wire n_17617;
wire n_8951;
wire n_5389;
wire n_5142;
wire n_18783;
wire n_15676;
wire n_17044;
wire n_9011;
wire n_7613;
wire n_3541;
wire n_6101;
wire n_14440;
wire n_7556;
wire n_5935;
wire n_10528;
wire n_372;
wire n_20168;
wire n_314;
wire n_13875;
wire n_17319;
wire n_17774;
wire n_338;
wire n_19255;
wire n_14076;
wire n_506;
wire n_11220;
wire n_17709;
wire n_9012;
wire n_2396;
wire n_18150;
wire n_2450;
wire n_14638;
wire n_2284;
wire n_19803;
wire n_7238;
wire n_2769;
wire n_14936;
wire n_16469;
wire n_8047;
wire n_11596;
wire n_6273;
wire n_5663;
wire n_525;
wire n_7572;
wire n_11955;
wire n_20535;
wire n_1677;
wire n_18818;
wire n_16156;
wire n_11654;
wire n_18361;
wire n_12982;
wire n_4160;
wire n_4231;
wire n_11619;
wire n_10649;
wire n_2779;
wire n_5203;
wire n_19638;
wire n_6311;
wire n_7590;
wire n_5162;
wire n_1464;
wire n_5285;
wire n_2721;
wire n_12275;
wire n_13742;
wire n_270;
wire n_15177;
wire n_12376;
wire n_563;
wire n_13114;
wire n_8583;
wire n_4521;
wire n_10447;
wire n_15063;
wire n_7176;
wire n_9353;
wire n_13054;
wire n_8948;
wire n_5715;
wire n_8295;
wire n_498;
wire n_5395;
wire n_10522;
wire n_13793;
wire n_11782;
wire n_16532;
wire n_20590;
wire n_1693;
wire n_16618;
wire n_10278;
wire n_15384;
wire n_13882;
wire n_9750;
wire n_9749;
wire n_14139;
wire n_2915;
wire n_15686;
wire n_9263;
wire n_11082;
wire n_1989;
wire n_15950;
wire n_2802;
wire n_19724;
wire n_6181;
wire n_7447;
wire n_17998;
wire n_19156;
wire n_18928;
wire n_12721;
wire n_18301;
wire n_5672;
wire n_16008;
wire n_11730;
wire n_3098;
wire n_6924;
wire n_9804;
wire n_1851;
wire n_9304;
wire n_5799;
wire n_8380;
wire n_12039;
wire n_3123;
wire n_3380;
wire n_5617;
wire n_10377;
wire n_9926;
wire n_570;
wire n_15161;
wire n_620;
wire n_2523;
wire n_10858;
wire n_5450;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_16303;
wire n_9843;
wire n_3130;
wire n_16559;
wire n_1710;
wire n_13320;
wire n_1301;
wire n_6683;
wire n_10683;
wire n_2282;
wire n_9921;
wire n_19606;
wire n_6229;
wire n_1609;
wire n_13488;
wire n_15907;
wire n_7286;
wire n_13668;
wire n_13016;
wire n_6177;
wire n_16961;
wire n_14708;
wire n_2867;
wire n_2726;
wire n_17293;
wire n_12048;
wire n_5982;
wire n_10930;
wire n_17972;
wire n_8749;
wire n_18264;
wire n_2662;
wire n_12057;
wire n_6696;
wire n_17590;
wire n_9527;
wire n_16450;
wire n_19651;
wire n_2795;
wire n_14875;
wire n_15860;
wire n_3472;
wire n_15056;
wire n_18352;
wire n_19460;
wire n_17288;
wire n_5376;
wire n_16197;
wire n_14003;
wire n_5106;
wire n_9511;
wire n_6730;
wire n_17822;
wire n_13670;
wire n_11254;
wire n_15023;
wire n_11617;
wire n_18184;
wire n_5561;
wire n_404;
wire n_158;
wire n_18436;
wire n_6170;
wire n_9459;
wire n_14185;
wire n_6094;
wire n_9098;
wire n_14953;
wire n_15604;
wire n_4826;
wire n_16000;
wire n_3903;
wire n_12360;
wire n_9268;
wire n_17116;
wire n_20497;
wire n_15431;
wire n_3854;
wire n_3235;
wire n_8673;
wire n_18702;
wire n_19174;
wire n_5378;
wire n_10456;
wire n_3673;
wire n_13186;
wire n_18824;
wire n_5916;
wire n_15655;
wire n_11907;
wire n_3094;
wire n_10627;
wire n_10475;
wire n_965;
wire n_1428;
wire n_20373;
wire n_15430;
wire n_1576;
wire n_2077;
wire n_20578;
wire n_8581;
wire n_15732;
wire n_12457;
wire n_16070;
wire n_16045;
wire n_4951;
wire n_17772;
wire n_540;
wire n_14170;
wire n_3070;
wire n_13496;
wire n_8058;
wire n_9308;
wire n_3504;
wire n_11838;
wire n_10508;
wire n_18008;
wire n_10811;
wire n_18696;
wire n_8333;
wire n_17152;
wire n_7619;
wire n_6985;
wire n_18551;
wire n_7170;
wire n_13853;
wire n_8823;
wire n_11457;
wire n_12751;
wire n_15284;
wire n_3054;
wire n_5399;
wire n_20374;
wire n_4620;
wire n_5421;
wire n_4127;
wire n_17901;
wire n_15443;
wire n_5206;
wire n_18228;
wire n_17833;
wire n_18471;
wire n_4517;
wire n_16852;
wire n_18817;
wire n_6916;
wire n_15524;
wire n_2260;
wire n_10725;
wire n_7845;
wire n_12688;
wire n_5550;
wire n_18354;
wire n_8290;
wire n_7536;
wire n_1743;
wire n_18152;
wire n_6230;
wire n_16108;
wire n_11107;
wire n_2956;
wire n_5573;
wire n_1553;
wire n_12757;
wire n_14379;
wire n_8840;
wire n_16284;
wire n_16001;
wire n_18873;
wire n_13189;
wire n_5881;
wire n_18915;
wire n_2382;
wire n_3754;
wire n_19492;
wire n_12328;
wire n_415;
wire n_9083;
wire n_17271;
wire n_383;
wire n_2974;
wire n_4213;
wire n_200;
wire n_6483;
wire n_10994;
wire n_14004;
wire n_17023;
wire n_5863;
wire n_2645;
wire n_16221;
wire n_3904;
wire n_8036;
wire n_11485;
wire n_1444;
wire n_7300;
wire n_6975;
wire n_14666;
wire n_1263;
wire n_13605;
wire n_17387;
wire n_11048;
wire n_4733;
wire n_14237;
wire n_6729;
wire n_4764;
wire n_1261;
wire n_3879;
wire n_11240;
wire n_13841;
wire n_3080;
wire n_11634;
wire n_12580;
wire n_10013;
wire n_17166;
wire n_2865;
wire n_16119;
wire n_6076;
wire n_8933;
wire n_19344;
wire n_15876;
wire n_18819;
wire n_15231;
wire n_11287;
wire n_943;
wire n_9774;
wire n_4879;
wire n_6390;
wire n_19846;
wire n_13409;
wire n_6665;
wire n_8797;
wire n_10723;
wire n_9720;
wire n_15727;
wire n_10169;
wire n_12690;
wire n_7563;
wire n_12475;
wire n_1345;
wire n_4556;
wire n_11765;
wire n_8434;
wire n_13405;
wire n_12302;
wire n_10477;
wire n_19510;
wire n_4117;
wire n_14414;
wire n_15565;
wire n_5995;
wire n_17823;
wire n_2378;
wire n_5905;
wire n_9149;
wire n_2655;
wire n_7035;
wire n_6193;
wire n_1467;
wire n_4250;
wire n_16858;
wire n_16980;
wire n_224;
wire n_3963;
wire n_9345;
wire n_11550;
wire n_17315;
wire n_7527;
wire n_13061;
wire n_9682;
wire n_2214;
wire n_17719;
wire n_6582;
wire n_18432;
wire n_12545;
wire n_20390;
wire n_18320;
wire n_1230;
wire n_3850;
wire n_18078;
wire n_9924;
wire n_14744;
wire n_15091;
wire n_5525;
wire n_17527;
wire n_163;
wire n_1644;
wire n_12753;
wire n_2277;
wire n_7090;
wire n_9254;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_11641;
wire n_7415;
wire n_11211;
wire n_13375;
wire n_13691;
wire n_824;
wire n_6745;
wire n_6972;
wire n_18526;
wire n_16913;
wire n_16663;
wire n_11857;
wire n_395;
wire n_6240;
wire n_13482;
wire n_18069;
wire n_5297;
wire n_15778;
wire n_7121;
wire n_9469;
wire n_15869;
wire n_2961;
wire n_15598;
wire n_15988;
wire n_16593;
wire n_6515;
wire n_483;
wire n_16604;
wire n_2546;
wire n_13873;
wire n_15805;
wire n_476;
wire n_1957;
wire n_17836;
wire n_4732;
wire n_18769;
wire n_11201;
wire n_10531;
wire n_14964;
wire n_8918;
wire n_12878;
wire n_19273;
wire n_8932;
wire n_17756;
wire n_4581;
wire n_16603;
wire n_9249;
wire n_2143;
wire n_8180;
wire n_20191;
wire n_15580;
wire n_9444;
wire n_10772;
wire n_2031;
wire n_7114;
wire n_4878;
wire n_15984;
wire n_6770;
wire n_20237;
wire n_20124;
wire n_17730;
wire n_15151;
wire n_16626;
wire n_5639;
wire n_487;
wire n_8943;
wire n_14767;
wire n_18463;
wire n_20343;
wire n_4503;
wire n_14773;
wire n_10127;
wire n_13654;
wire n_5361;
wire n_11814;
wire n_12255;
wire n_4199;
wire n_1912;
wire n_9723;
wire n_19446;
wire n_19669;
wire n_1982;
wire n_3872;
wire n_1312;
wire n_19834;
wire n_19577;
wire n_5330;
wire n_7199;
wire n_10039;
wire n_10854;
wire n_11358;
wire n_13366;
wire n_247;
wire n_5892;
wire n_7940;
wire n_16467;
wire n_6782;
wire n_18746;
wire n_2008;
wire n_2192;
wire n_328;
wire n_17669;
wire n_1386;
wire n_6503;
wire n_19423;
wire n_12017;
wire n_17357;
wire n_15381;
wire n_18477;
wire n_11958;
wire n_6621;
wire n_15624;
wire n_16103;
wire n_19041;
wire n_16460;
wire n_690;
wire n_8271;
wire n_4800;
wire n_1157;
wire n_20303;
wire n_12728;
wire n_1752;
wire n_16651;
wire n_4958;
wire n_6783;
wire n_19963;
wire n_12259;
wire n_8699;
wire n_16305;
wire n_19409;
wire n_2963;
wire n_19932;
wire n_15861;
wire n_3873;
wire n_8225;
wire n_9536;
wire n_14250;
wire n_16818;
wire n_16573;
wire n_18671;
wire n_16562;
wire n_6296;
wire n_7708;
wire n_11671;
wire n_10328;
wire n_5968;
wire n_2644;
wire n_3326;
wire n_6497;
wire n_15705;
wire n_2411;
wire n_16816;
wire n_7333;
wire n_15376;
wire n_8546;
wire n_10963;
wire n_16358;
wire n_18035;
wire n_7371;
wire n_17547;
wire n_8152;
wire n_15050;
wire n_10826;
wire n_7463;
wire n_8525;
wire n_17767;
wire n_18680;
wire n_283;
wire n_12160;
wire n_590;
wire n_9620;
wire n_1990;
wire n_3805;
wire n_5205;
wire n_17145;
wire n_11119;
wire n_7954;
wire n_1465;
wire n_2622;
wire n_7951;
wire n_8096;
wire n_13901;
wire n_7231;
wire n_5080;
wire n_3128;
wire n_15252;
wire n_18043;
wire n_20465;
wire n_16238;
wire n_5372;
wire n_14050;
wire n_15763;
wire n_17983;
wire n_2691;
wire n_15317;
wire n_7772;
wire n_2690;
wire n_14197;
wire n_18159;
wire n_19364;
wire n_8996;
wire n_12070;
wire n_9714;
wire n_3078;
wire n_14898;
wire n_15672;
wire n_20532;
wire n_3793;
wire n_15920;
wire n_11928;
wire n_5071;
wire n_14395;
wire n_5801;
wire n_13528;
wire n_6047;
wire n_8292;
wire n_8601;
wire n_9377;
wire n_11932;
wire n_6970;
wire n_19328;
wire n_1308;
wire n_13027;
wire n_20342;
wire n_12607;
wire n_7272;
wire n_15782;
wire n_19553;
wire n_12075;
wire n_4540;
wire n_13489;
wire n_2097;
wire n_18887;
wire n_3499;
wire n_19693;
wire n_19797;
wire n_13877;
wire n_1005;
wire n_6209;
wire n_11922;
wire n_14020;
wire n_1469;
wire n_12358;
wire n_7408;
wire n_2650;
wire n_10488;
wire n_8969;
wire n_14187;
wire n_11577;
wire n_17840;
wire n_16914;
wire n_18513;
wire n_153;
wire n_3348;
wire n_19165;
wire n_17907;
wire n_11475;
wire n_9048;
wire n_5228;
wire n_10274;
wire n_1723;
wire n_189;
wire n_6694;
wire n_15318;
wire n_9168;
wire n_14220;
wire n_13837;
wire n_2335;
wire n_18570;
wire n_529;
wire n_5507;
wire n_5569;
wire n_15559;
wire n_16871;
wire n_14221;
wire n_13964;
wire n_10832;
wire n_3173;
wire n_18829;
wire n_6856;
wire n_1049;
wire n_6466;
wire n_16039;
wire n_7864;
wire n_18295;
wire n_6727;
wire n_14360;
wire n_10584;
wire n_1717;
wire n_2449;
wire n_3880;
wire n_13601;
wire n_17457;
wire n_17115;
wire n_19281;
wire n_18155;
wire n_4545;
wire n_272;
wire n_6820;
wire n_2896;
wire n_2639;
wire n_17083;
wire n_458;
wire n_5490;
wire n_19007;
wire n_4771;
wire n_13392;
wire n_5836;
wire n_17563;
wire n_9169;
wire n_252;
wire n_5834;
wire n_3191;
wire n_10229;
wire n_5584;
wire n_7512;
wire n_3561;
wire n_19008;
wire n_18401;
wire n_6469;
wire n_6700;
wire n_20494;
wire n_3032;
wire n_6223;
wire n_11398;
wire n_8798;
wire n_9600;
wire n_2877;
wire n_8085;
wire n_11274;
wire n_1021;
wire n_8123;
wire n_811;
wire n_17997;
wire n_12512;
wire n_9927;
wire n_5497;
wire n_16973;
wire n_15657;
wire n_17571;
wire n_3598;
wire n_7127;
wire n_831;
wire n_15513;
wire n_8666;
wire n_2435;
wire n_12284;
wire n_18322;
wire n_1382;
wire n_7801;
wire n_9155;
wire n_1483;
wire n_10416;
wire n_15837;
wire n_1372;
wire n_14370;
wire n_1719;
wire n_7959;
wire n_13430;
wire n_1427;
wire n_2745;
wire n_14525;
wire n_7735;
wire n_8004;
wire n_6667;
wire n_10583;
wire n_10806;
wire n_2323;
wire n_162;
wire n_5234;
wire n_7546;
wire n_6272;
wire n_14274;
wire n_6588;
wire n_3265;
wire n_3755;
wire n_4042;
wire n_18125;
wire n_15403;
wire n_13081;
wire n_15602;
wire n_12252;
wire n_16743;
wire n_10439;
wire n_12627;
wire n_19378;
wire n_16730;
wire n_15637;
wire n_14272;
wire n_11237;
wire n_2410;
wire n_20012;
wire n_18868;
wire n_6222;
wire n_15012;
wire n_20451;
wire n_1783;
wire n_4176;
wire n_14551;
wire n_15720;
wire n_11181;
wire n_13651;
wire n_7521;
wire n_12968;
wire n_10663;
wire n_15517;
wire n_3894;
wire n_13974;
wire n_12277;
wire n_14917;
wire n_3127;
wire n_3623;
wire n_5312;
wire n_16075;
wire n_6625;
wire n_15680;
wire n_2502;
wire n_3646;
wire n_17441;
wire n_14855;
wire n_16757;
wire n_2783;
wire n_8487;
wire n_4034;
wire n_18601;
wire n_1470;
wire n_8141;
wire n_4887;
wire n_14058;
wire n_11020;
wire n_13141;
wire n_16461;
wire n_14065;
wire n_11920;
wire n_19756;
wire n_17299;
wire n_3862;
wire n_14366;
wire n_10481;
wire n_19250;
wire n_6876;
wire n_16022;
wire n_5049;
wire n_19001;
wire n_19627;
wire n_9573;
wire n_5846;
wire n_7636;
wire n_9799;
wire n_17235;
wire n_5592;
wire n_6954;
wire n_6938;
wire n_1855;
wire n_3051;
wire n_15143;
wire n_11198;
wire n_18932;
wire n_18346;
wire n_18238;
wire n_385;
wire n_1439;
wire n_2859;
wire n_1331;
wire n_19794;
wire n_5157;
wire n_3525;
wire n_2100;
wire n_11840;
wire n_13157;
wire n_1134;
wire n_10261;
wire n_4003;
wire n_5708;
wire n_3751;
wire n_4894;
wire n_14084;
wire n_4113;
wire n_5649;
wire n_9827;
wire n_13334;
wire n_10907;
wire n_4983;
wire n_14002;
wire n_19842;
wire n_19892;
wire n_419;
wire n_7214;
wire n_3907;
wire n_16205;
wire n_13399;
wire n_1254;
wire n_19984;
wire n_7075;
wire n_19503;
wire n_14697;
wire n_7124;
wire n_13967;
wire n_3291;
wire n_20506;
wire n_2304;
wire n_7799;
wire n_5698;
wire n_11092;
wire n_14310;
wire n_5084;
wire n_15792;
wire n_15281;
wire n_15675;
wire n_8917;
wire n_15515;
wire n_9647;
wire n_15106;
wire n_4710;
wire n_12067;
wire n_9214;
wire n_17030;
wire n_19537;
wire n_4101;
wire n_7776;
wire n_19621;
wire n_14309;
wire n_9864;
wire n_16256;
wire n_3236;
wire n_17416;
wire n_16741;
wire n_923;
wire n_11770;
wire n_19201;
wire n_13996;
wire n_19904;
wire n_19853;
wire n_17944;
wire n_17679;
wire n_9000;
wire n_18442;
wire n_18505;
wire n_10864;
wire n_18412;
wire n_14704;
wire n_8307;
wire n_9383;
wire n_17692;
wire n_4611;
wire n_15258;
wire n_2337;
wire n_12174;
wire n_16322;
wire n_15220;
wire n_6400;
wire n_19611;
wire n_16304;
wire n_18417;
wire n_7543;
wire n_13504;
wire n_16787;
wire n_13169;
wire n_7877;
wire n_9672;
wire n_15291;
wire n_8855;
wire n_18375;
wire n_8885;
wire n_5486;
wire n_15345;
wire n_137;
wire n_1596;
wire n_5092;
wire n_14721;
wire n_1734;
wire n_3172;
wire n_13265;
wire n_4832;
wire n_2902;
wire n_12153;
wire n_7284;
wire n_7264;
wire n_13666;
wire n_19192;
wire n_6537;
wire n_20408;
wire n_10702;
wire n_13730;
wire n_3536;
wire n_12405;
wire n_2894;
wire n_3710;
wire n_4195;
wire n_10319;
wire n_9654;
wire n_8802;
wire n_9859;
wire n_5240;
wire n_2225;
wire n_6092;
wire n_6241;
wire n_1692;
wire n_8667;
wire n_18996;
wire n_2006;
wire n_3402;
wire n_8121;
wire n_9645;
wire n_7754;
wire n_15549;
wire n_18777;
wire n_2789;
wire n_12792;
wire n_1828;
wire n_19661;
wire n_9796;
wire n_8320;
wire n_18219;
wire n_18231;
wire n_4862;
wire n_15889;
wire n_2376;
wire n_12438;
wire n_11830;
wire n_8766;
wire n_16665;
wire n_16173;
wire n_9165;
wire n_2700;
wire n_19555;
wire n_1041;
wire n_12539;
wire n_565;
wire n_5965;
wire n_9596;
wire n_13652;
wire n_13703;
wire n_18461;
wire n_14369;
wire n_1062;
wire n_7240;
wire n_15354;
wire n_10476;
wire n_9966;
wire n_16794;
wire n_1222;
wire n_2635;
wire n_11486;
wire n_15999;
wire n_15280;
wire n_12677;
wire n_4321;
wire n_7237;
wire n_17867;
wire n_16456;
wire n_6877;
wire n_12873;
wire n_16364;
wire n_6949;
wire n_20531;
wire n_19356;
wire n_17036;
wire n_19698;
wire n_806;
wire n_13401;
wire n_584;
wire n_12276;
wire n_9893;
wire n_14122;
wire n_17565;
wire n_8126;
wire n_15819;
wire n_10362;
wire n_9239;
wire n_3930;
wire n_4757;
wire n_15603;
wire n_12352;
wire n_17267;
wire n_2809;
wire n_18528;
wire n_787;
wire n_10099;
wire n_9961;
wire n_16833;
wire n_14895;
wire n_7163;
wire n_1528;
wire n_1146;
wire n_16582;
wire n_18028;
wire n_2021;
wire n_15270;
wire n_17964;
wire n_10181;
wire n_15670;
wire n_19974;
wire n_4604;
wire n_5724;
wire n_7201;
wire n_3157;
wire n_16825;
wire n_20274;
wire n_2422;
wire n_10949;
wire n_3457;
wire n_3762;
wire n_18197;
wire n_3411;
wire n_4519;
wire n_5355;
wire n_13969;
wire n_16548;
wire n_5186;
wire n_1498;
wire n_12693;
wire n_6792;
wire n_1210;
wire n_9316;
wire n_5438;
wire n_13259;
wire n_1269;
wire n_19164;
wire n_14954;
wire n_12648;
wire n_655;
wire n_4726;
wire n_6045;
wire n_1872;
wire n_9914;
wire n_8132;
wire n_19541;
wire n_20433;
wire n_10917;
wire n_16050;
wire n_3761;
wire n_18006;
wire n_7821;
wire n_12407;
wire n_11284;
wire n_20100;
wire n_14668;
wire n_14776;
wire n_10458;
wire n_2041;
wire n_11656;
wire n_13134;
wire n_10271;
wire n_15415;
wire n_20315;
wire n_16808;
wire n_18902;
wire n_1098;
wire n_5746;
wire n_6673;
wire n_20026;
wire n_18207;
wire n_11909;
wire n_12637;
wire n_7887;
wire n_398;
wire n_6060;
wire n_15414;
wire n_15783;
wire n_3726;
wire n_12009;
wire n_2369;
wire n_13612;
wire n_19388;
wire n_10648;
wire n_2587;
wire n_7550;
wire n_17498;
wire n_15077;
wire n_3199;
wire n_12414;
wire n_9760;
wire n_10690;
wire n_15733;
wire n_15864;
wire n_14207;
wire n_1953;
wire n_19080;
wire n_19736;
wire n_13863;
wire n_14305;
wire n_9863;
wire n_15330;
wire n_10500;
wire n_5432;
wire n_15261;
wire n_11929;
wire n_11075;
wire n_7851;
wire n_16605;
wire n_20372;
wire n_9791;
wire n_19228;
wire n_5453;
wire n_4900;
wire n_11177;
wire n_19761;
wire n_13667;
wire n_18056;
wire n_5842;
wire n_13126;
wire n_7798;
wire n_5253;
wire n_10857;
wire n_18491;
wire n_11310;
wire n_13275;
wire n_11165;
wire n_14411;
wire n_20503;
wire n_12823;
wire n_2953;
wire n_15412;
wire n_4295;
wire n_5943;
wire n_20331;
wire n_12193;
wire n_2500;
wire n_1729;
wire n_6088;
wire n_5777;
wire n_15257;
wire n_19701;
wire n_8528;
wire n_8204;
wire n_11733;
wire n_15646;
wire n_1389;
wire n_18214;
wire n_7100;
wire n_3583;
wire n_3860;
wire n_18347;
wire n_14738;
wire n_12242;
wire n_5610;
wire n_3015;
wire n_20108;
wire n_13796;
wire n_10502;
wire n_15522;
wire n_17577;
wire n_17874;
wire n_6722;
wire n_17892;
wire n_7622;
wire n_11123;
wire n_8512;
wire n_14464;
wire n_387;
wire n_744;
wire n_971;
wire n_8635;
wire n_3241;
wire n_2906;
wire n_4342;
wire n_10855;
wire n_7995;
wire n_6114;
wire n_1205;
wire n_15535;
wire n_16633;
wire n_7831;
wire n_10227;
wire n_10574;
wire n_19271;
wire n_2180;
wire n_16323;
wire n_2858;
wire n_18624;
wire n_6201;
wire n_12218;
wire n_5737;
wire n_3604;
wire n_12343;
wire n_4373;
wire n_8919;
wire n_17014;
wire n_12316;
wire n_14937;
wire n_14454;
wire n_4711;
wire n_11478;
wire n_16067;
wire n_3068;
wire n_15650;
wire n_12236;
wire n_12902;
wire n_16230;
wire n_7784;
wire n_9272;
wire n_5768;
wire n_13038;
wire n_2465;
wire n_12892;
wire n_17768;
wire n_3811;
wire n_11294;
wire n_910;
wire n_15667;
wire n_3486;
wire n_4086;
wire n_19861;
wire n_10289;
wire n_6565;
wire n_6942;
wire n_11819;
wire n_19389;
wire n_2032;
wire n_4812;
wire n_13420;
wire n_6862;
wire n_5858;
wire n_17200;
wire n_15053;
wire n_13005;
wire n_708;
wire n_14805;
wire n_20575;
wire n_6037;
wire n_2312;
wire n_11844;
wire n_1266;
wire n_15390;
wire n_6635;
wire n_185;
wire n_13184;
wire n_1276;
wire n_13535;
wire n_14982;
wire n_12247;
wire n_14770;
wire n_11100;
wire n_298;
wire n_1582;
wire n_5588;
wire n_3286;
wire n_19350;
wire n_7167;
wire n_6480;
wire n_15105;
wire n_5075;
wire n_3682;
wire n_18927;
wire n_3771;
wire n_18383;
wire n_12765;
wire n_7865;
wire n_15690;
wire n_9289;
wire n_11315;
wire n_6561;
wire n_12706;
wire n_19949;
wire n_11153;
wire n_17128;
wire n_859;
wire n_406;
wire n_6875;
wire n_10934;
wire n_1770;
wire n_10197;
wire n_18999;
wire n_3285;
wire n_19584;
wire n_11949;
wire n_8402;
wire n_9690;
wire n_2071;
wire n_11746;
wire n_9371;
wire n_19689;
wire n_19990;
wire n_16837;
wire n_20095;
wire n_7267;
wire n_4599;
wire n_12315;
wire n_18668;
wire n_5222;
wire n_7850;
wire n_14100;
wire n_12998;
wire n_7812;
wire n_13143;
wire n_9080;
wire n_14549;
wire n_8133;
wire n_6176;
wire n_14717;
wire n_3881;
wire n_16426;
wire n_14459;
wire n_4508;
wire n_11530;
wire n_13411;
wire n_7056;
wire n_8193;
wire n_12445;
wire n_12856;
wire n_19520;
wire n_7813;
wire n_7514;
wire n_18734;
wire n_7649;
wire n_12525;
wire n_16116;
wire n_1039;
wire n_6078;
wire n_2043;
wire n_1480;
wire n_15823;
wire n_5832;
wire n_13758;
wire n_1305;
wire n_7688;
wire n_4562;
wire n_16820;
wire n_3383;
wire n_12357;
wire n_8707;
wire n_9208;
wire n_11791;
wire n_19525;
wire n_7611;
wire n_19778;
wire n_17218;
wire n_15216;
wire n_11848;
wire n_3610;
wire n_11632;
wire n_15352;
wire n_7795;
wire n_12180;
wire n_2065;
wire n_15608;
wire n_10935;
wire n_20044;
wire n_2001;
wire n_7723;
wire n_11621;
wire n_19448;
wire n_225;
wire n_16171;
wire n_3555;
wire n_7450;
wire n_11667;
wire n_17311;
wire n_7362;
wire n_17455;
wire n_12208;
wire n_1131;
wire n_3110;
wire n_14565;
wire n_17248;
wire n_11298;
wire n_15796;
wire n_1888;
wire n_8993;
wire n_6204;
wire n_13314;
wire n_670;
wire n_11741;
wire n_3908;
wire n_15537;
wire n_3467;
wire n_12773;
wire n_9044;
wire n_12381;
wire n_19885;
wire n_19302;
wire n_18174;
wire n_14883;
wire n_17024;
wire n_6451;
wire n_9813;
wire n_1226;
wire n_3740;
wire n_18482;
wire n_3186;
wire n_640;
wire n_20217;
wire n_17322;
wire n_9244;
wire n_15304;
wire n_7049;
wire n_15271;
wire n_2632;
wire n_14865;
wire n_8278;
wire n_11644;
wire n_6345;
wire n_15893;
wire n_9094;
wire n_15432;
wire n_13108;
wire n_364;
wire n_5782;
wire n_5041;
wire n_13170;
wire n_1915;
wire n_4275;
wire n_14471;
wire n_11357;
wire n_19387;
wire n_4425;
wire n_9985;
wire n_4449;
wire n_12089;
wire n_20104;
wire n_7057;
wire n_17888;
wire n_11959;
wire n_19586;
wire n_1612;
wire n_4809;
wire n_12987;
wire n_8529;
wire n_625;
wire n_10254;
wire n_18625;
wire n_14715;
wire n_15970;
wire n_11208;
wire n_15978;
wire n_12452;
wire n_20495;
wire n_15961;
wire n_8574;
wire n_1038;
wire n_12292;
wire n_4241;
wire n_12818;
wire n_11420;
wire n_12500;
wire n_8044;
wire n_16330;
wire n_9439;
wire n_1380;
wire n_15239;
wire n_2557;
wire n_11630;
wire n_2405;
wire n_19759;
wire n_15444;
wire n_15289;
wire n_13172;
wire n_2336;
wire n_16234;
wire n_2521;
wire n_9120;
wire n_17335;
wire n_17610;
wire n_19522;
wire n_424;
wire n_12168;
wire n_16496;
wire n_8903;
wire n_141;
wire n_1985;
wire n_16057;
wire n_16401;
wire n_4531;
wire n_3282;
wire n_15781;
wire n_14448;
wire n_1532;
wire n_11017;
wire n_7247;
wire n_14622;
wire n_4666;
wire n_7893;
wire n_6213;
wire n_19924;
wire n_3031;
wire n_14739;
wire n_16649;
wire n_12613;
wire n_14365;
wire n_9325;
wire n_16448;
wire n_4555;
wire n_17173;
wire n_9384;
wire n_6216;
wire n_7340;
wire n_12695;
wire n_15467;
wire n_4308;
wire n_14219;
wire n_3463;
wire n_11576;
wire n_1954;
wire n_2729;
wire n_2582;
wire n_1798;
wire n_3998;
wire n_12006;
wire n_2495;
wire n_10128;
wire n_371;
wire n_18319;
wire n_12246;
wire n_18220;
wire n_9955;
wire n_19477;
wire n_3829;
wire n_9007;
wire n_10143;
wire n_1471;
wire n_18715;
wire n_3655;
wire n_17884;
wire n_3825;
wire n_2880;
wire n_13085;
wire n_19260;
wire n_7780;
wire n_20413;
wire n_8452;
wire n_11518;
wire n_5670;
wire n_8557;
wire n_10303;
wire n_16189;
wire n_15097;
wire n_18892;
wire n_11252;
wire n_8012;
wire n_1445;
wire n_1526;
wire n_17055;
wire n_1978;
wire n_6472;
wire n_18067;
wire n_574;
wire n_8114;
wire n_4202;
wire n_16227;
wire n_5879;
wire n_14563;
wire n_4403;
wire n_5238;
wire n_16329;
wire n_11256;
wire n_6166;
wire n_12370;
wire n_9136;
wire n_12860;
wire n_16278;
wire n_473;
wire n_17404;
wire n_559;
wire n_19635;
wire n_7063;
wire n_14768;
wire n_4139;
wire n_13885;
wire n_20364;
wire n_1986;
wire n_13631;
wire n_18103;
wire n_6081;
wire n_16746;
wire n_15929;
wire n_6724;
wire n_813;
wire n_11336;
wire n_12758;
wire n_17410;
wire n_19248;
wire n_11849;
wire n_3910;
wire n_9476;
wire n_9204;
wire n_12142;
wire n_9689;
wire n_16711;
wire n_10659;
wire n_7585;
wire n_4948;
wire n_5268;
wire n_6946;
wire n_3319;
wire n_12983;
wire n_3748;
wire n_6424;
wire n_11210;
wire n_7599;
wire n_16271;
wire n_15541;
wire n_13980;
wire n_16366;
wire n_982;
wire n_11191;
wire n_10547;
wire n_6778;
wire n_17359;
wire n_13205;
wire n_1697;
wire n_979;
wire n_5544;
wire n_5067;
wire n_15283;
wire n_12396;
wire n_15407;
wire n_7614;
wire n_19381;
wire n_1278;
wire n_7839;
wire n_9837;
wire n_634;
wire n_10896;
wire n_136;
wire n_17761;
wire n_4130;
wire n_10562;
wire n_16042;
wire n_5941;
wire n_2009;
wire n_14417;
wire n_3601;
wire n_6340;
wire n_10054;
wire n_10355;
wire n_1289;
wire n_16893;
wire n_3055;
wire n_6706;
wire n_3966;
wire n_13034;
wire n_1014;
wire n_16828;
wire n_10007;
wire n_882;
wire n_11751;
wire n_17550;
wire n_3746;
wire n_17185;
wire n_20286;
wire n_14637;
wire n_11495;
wire n_4478;
wire n_1662;
wire n_17015;
wire n_7372;
wire n_19617;
wire n_2818;
wire n_17980;
wire n_674;
wire n_3921;
wire n_17535;
wire n_16822;
wire n_10704;
wire n_11520;
wire n_1927;
wire n_19614;
wire n_12169;
wire n_16788;
wire n_15088;
wire n_17976;
wire n_702;
wire n_4965;
wire n_16383;
wire n_17538;
wire n_11012;
wire n_6111;
wire n_11502;
wire n_15348;
wire n_11631;
wire n_13588;
wire n_13570;
wire n_2193;
wire n_4523;
wire n_20176;
wire n_6011;
wire n_20038;
wire n_11842;
wire n_14710;
wire n_3153;
wire n_877;
wire n_13737;
wire n_16590;
wire n_728;
wire n_18188;
wire n_4607;
wire n_16640;
wire n_11389;
wire n_7226;
wire n_9013;
wire n_18373;
wire n_4041;
wire n_9634;
wire n_17846;
wire n_5876;
wire n_10916;
wire n_8584;
wire n_11557;
wire n_17113;
wire n_16748;
wire n_15363;
wire n_7810;
wire n_14955;
wire n_9364;
wire n_8228;
wire n_1825;
wire n_16015;
wire n_170;
wire n_15642;
wire n_1412;
wire n_10929;
wire n_18854;
wire n_19372;
wire n_13862;
wire n_8100;
wire n_13446;
wire n_13086;
wire n_8091;
wire n_5837;
wire n_148;
wire n_4675;
wire n_17155;
wire n_5491;
wire n_2987;
wire n_20236;
wire n_5496;
wire n_5802;
wire n_14965;
wire n_13887;
wire n_12787;
wire n_12799;
wire n_4002;
wire n_5178;
wire n_9317;
wire n_12657;
wire n_9769;
wire n_15205;
wire n_8158;
wire n_1295;
wire n_8469;
wire n_18718;
wire n_18481;
wire n_10102;
wire n_5983;
wire n_3146;
wire n_1438;
wire n_3953;
wire n_11825;
wire n_1100;
wire n_14354;
wire n_7684;
wire n_15532;
wire n_5604;
wire n_673;
wire n_16083;
wire n_10589;
wire n_11611;
wire n_6642;
wire n_6847;
wire n_10707;
wire n_865;
wire n_4191;
wire n_18221;
wire n_12408;
wire n_16287;
wire n_16169;
wire n_19314;
wire n_17556;
wire n_2341;
wire n_10110;
wire n_11230;
wire n_11688;
wire n_4350;
wire n_12715;
wire n_12434;
wire n_11709;
wire n_14328;
wire n_6095;
wire n_17049;
wire n_18938;
wire n_16540;
wire n_14429;
wire n_12979;
wire n_16901;
wire n_6559;
wire n_3924;
wire n_15799;
wire n_19733;
wire n_17195;
wire n_19050;
wire n_4621;
wire n_510;
wire n_1488;
wire n_2148;
wire n_5565;
wire n_14270;
wire n_15238;
wire n_2339;
wire n_10190;
wire n_19656;
wire n_5984;
wire n_6287;
wire n_13614;
wire n_8347;
wire n_17703;
wire n_19440;
wire n_1776;
wire n_1766;
wire n_14208;
wire n_9330;
wire n_20399;
wire n_4021;
wire n_3014;
wire n_15693;
wire n_12029;
wire n_4103;
wire n_9523;
wire n_14584;
wire n_4022;
wire n_19636;
wire n_10060;
wire n_18192;
wire n_9686;
wire n_4481;
wire n_20434;
wire n_17130;
wire n_19375;
wire n_1304;
wire n_10162;
wire n_4669;
wire n_15002;
wire n_9964;
wire n_17515;
wire n_13842;
wire n_7510;
wire n_6662;
wire n_11291;
wire n_13107;
wire n_5603;
wire n_9154;
wire n_14501;
wire n_3312;
wire n_7109;
wire n_2936;
wire n_3224;
wire n_8822;
wire n_14790;
wire n_1087;
wire n_17204;
wire n_12187;
wire n_657;
wire n_19662;
wire n_20121;
wire n_18772;
wire n_1505;
wire n_7253;
wire n_3129;
wire n_17201;
wire n_8476;
wire n_17745;
wire n_11927;
wire n_16674;
wire n_16326;
wire n_16571;
wire n_8359;
wire n_4484;
wire n_15808;
wire n_16497;
wire n_16752;
wire n_14574;
wire n_526;
wire n_14451;
wire n_2251;
wire n_9455;
wire n_8708;
wire n_14092;
wire n_2837;
wire n_4883;
wire n_14509;
wire n_11882;
wire n_17649;
wire n_11647;
wire n_15027;
wire n_15404;
wire n_10706;
wire n_3341;
wire n_19129;
wire n_8872;
wire n_20120;
wire n_19746;
wire n_3559;
wire n_8238;
wire n_15465;
wire n_20318;
wire n_11222;
wire n_9200;
wire n_16279;
wire n_5146;
wire n_3056;
wire n_745;
wire n_15858;
wire n_3447;
wire n_3971;
wire n_716;
wire n_1774;
wire n_18946;
wire n_2589;
wire n_4535;
wire n_14765;
wire n_7704;
wire n_18893;
wire n_16170;
wire n_14995;
wire n_6302;
wire n_2442;
wire n_17479;
wire n_7203;
wire n_11259;
wire n_7670;
wire n_18258;
wire n_16010;
wire n_14434;
wire n_9673;
wire n_20252;
wire n_2545;
wire n_8642;
wire n_11875;
wire n_18567;
wire n_12111;
wire n_8912;
wire n_19067;
wire n_1314;
wire n_864;
wire n_14275;
wire n_19309;
wire n_12903;
wire n_6343;
wire n_12593;
wire n_20051;
wire n_5270;
wire n_1534;
wire n_17849;
wire n_20588;
wire n_11602;
wire n_15689;
wire n_19850;
wire n_12413;
wire n_17474;
wire n_723;
wire n_13813;
wire n_16190;
wire n_18315;
wire n_8111;
wire n_10432;
wire n_19227;
wire n_16888;
wire n_8056;
wire n_18376;
wire n_3287;
wire n_9674;
wire n_2357;
wire n_6433;
wire n_18253;
wire n_15469;
wire n_17140;
wire n_18407;
wire n_1681;
wire n_520;
wire n_18816;
wire n_4020;
wire n_13636;
wire n_19332;
wire n_19456;
wire n_5220;
wire n_18920;
wire n_11341;
wire n_10787;
wire n_13256;
wire n_14567;
wire n_6870;
wire n_6221;
wire n_16308;
wire n_6279;
wire n_13905;
wire n_12290;
wire n_20558;
wire n_7881;
wire n_9369;
wire n_18896;
wire n_16986;
wire n_17872;
wire n_6071;
wire n_9583;
wire n_19422;
wire n_19858;
wire n_15119;
wire n_19117;
wire n_12150;
wire n_1617;
wire n_3370;
wire n_335;
wire n_15256;
wire n_18366;
wire n_8090;
wire n_8053;
wire n_10184;
wire n_15982;
wire n_274;
wire n_19643;
wire n_18647;
wire n_15452;
wire n_1267;
wire n_1806;
wire n_13615;
wire n_15625;
wire n_2023;
wire n_12633;
wire n_14779;
wire n_496;
wire n_15114;
wire n_4614;
wire n_3360;
wire n_10277;
wire n_17934;
wire n_3956;
wire n_8163;
wire n_16632;
wire n_16028;
wire n_19862;
wire n_10948;
wire n_10525;
wire n_14287;
wire n_9507;
wire n_11528;
wire n_15296;
wire n_15828;
wire n_18107;
wire n_19211;
wire n_3870;
wire n_16126;
wire n_18102;
wire n_19699;
wire n_18545;
wire n_16168;
wire n_15915;
wire n_793;
wire n_10049;
wire n_3749;
wire n_15551;
wire n_9457;
wire n_5780;
wire n_5037;
wire n_16738;
wire n_316;
wire n_6084;
wire n_11039;
wire n_14342;
wire n_2555;
wire n_13693;
wire n_18992;
wire n_12606;
wire n_10900;
wire n_2201;
wire n_14107;
wire n_14781;
wire n_13333;
wire n_13229;
wire n_994;
wire n_17336;
wire n_11380;
wire n_15737;
wire n_19567;
wire n_10792;
wire n_15573;
wire n_13296;
wire n_14611;
wire n_3448;
wire n_17863;
wire n_1036;
wire n_20165;
wire n_1661;
wire n_20196;
wire n_5360;
wire n_17088;
wire n_19100;
wire n_15051;
wire n_6548;
wire n_20383;
wire n_3926;
wire n_6993;
wire n_1095;
wire n_15916;
wire n_4405;
wire n_16468;
wire n_10241;
wire n_19598;
wire n_15639;
wire n_3670;
wire n_179;
wire n_4667;
wire n_8702;
wire n_17158;
wire n_8116;
wire n_1115;
wire n_8195;
wire n_7946;
wire n_14069;
wire n_18452;
wire n_19786;
wire n_1409;
wire n_9991;
wire n_11366;
wire n_11872;
wire n_19901;
wire n_10823;
wire n_19685;
wire n_14766;
wire n_11106;
wire n_1126;
wire n_14592;
wire n_15109;
wire n_11132;
wire n_17625;
wire n_18546;
wire n_18034;
wire n_3635;
wire n_18181;
wire n_17126;
wire n_10824;
wire n_4155;
wire n_19566;
wire n_16216;
wire n_19398;
wire n_14277;
wire n_19565;
wire n_13493;
wire n_16389;
wire n_9047;
wire n_12842;
wire n_18569;
wire n_12481;
wire n_18168;
wire n_11316;
wire n_9599;
wire n_11559;
wire n_9072;
wire n_19811;
wire n_4929;
wire n_9428;
wire n_10340;
wire n_17463;
wire n_15817;
wire n_15344;
wire n_2220;
wire n_2577;
wire n_13669;
wire n_17245;
wire n_3529;
wire n_17179;
wire n_11109;
wire n_13840;
wire n_16601;
wire n_20199;
wire n_11591;
wire n_19710;
wire n_14251;
wire n_11225;
wire n_6765;
wire n_4565;
wire n_4159;
wire n_8883;
wire n_10634;
wire n_4586;
wire n_11058;
wire n_15888;
wire n_1608;
wire n_7336;
wire n_11471;
wire n_7446;
wire n_3628;
wire n_14679;
wire n_10961;
wire n_7357;
wire n_1491;
wire n_20301;
wire n_17064;
wire n_8737;
wire n_13925;
wire n_18334;
wire n_10379;
wire n_16704;
wire n_2586;
wire n_18223;
wire n_13368;
wire n_14507;
wire n_9484;
wire n_10989;
wire n_17725;
wire n_10939;
wire n_19557;
wire n_1046;
wire n_2560;
wire n_1145;
wire n_11144;
wire n_14857;
wire n_6406;
wire n_14034;
wire n_10962;
wire n_11128;
wire n_15677;
wire n_10721;
wire n_8593;
wire n_12007;
wire n_11025;
wire n_5062;
wire n_15901;
wire n_321;
wire n_13481;
wire n_12018;
wire n_3588;
wire n_18040;
wire n_17393;
wire n_14457;
wire n_16931;
wire n_12872;
wire n_18189;
wire n_6492;
wire n_14517;
wire n_2288;
wire n_11460;
wire n_13713;
wire n_12372;
wire n_13608;
wire n_7046;
wire n_19059;
wire n_10956;
wire n_2642;
wire n_7468;
wire n_2383;
wire n_18785;
wire n_14934;
wire n_19663;
wire n_2351;
wire n_18844;
wire n_5069;
wire n_12453;
wire n_12572;
wire n_19968;
wire n_2986;
wire n_19752;
wire n_17870;
wire n_139;
wire n_15652;
wire n_3489;
wire n_19466;
wire n_16713;
wire n_14578;
wire n_15653;
wire n_5914;
wire n_12955;
wire n_9321;
wire n_16856;
wire n_18555;
wire n_1282;
wire n_15016;
wire n_2567;
wire n_18493;
wire n_275;
wire n_3377;
wire n_9161;
wire n_2869;
wire n_7836;
wire n_10737;
wire n_17910;
wire n_17750;
wire n_346;
wire n_15865;
wire n_13448;
wire n_16928;
wire n_5813;
wire n_13767;
wire n_790;
wire n_2611;
wire n_2901;
wire n_11055;
wire n_4358;
wire n_16616;
wire n_14832;
wire n_10982;
wire n_5616;
wire n_5805;
wire n_17599;
wire n_14571;
wire n_6631;
wire n_12369;
wire n_7577;
wire n_7308;
wire n_5169;
wire n_8927;
wire n_17985;
wire n_16396;
wire n_17531;
wire n_15155;
wire n_12686;
wire n_6228;
wire n_19336;
wire n_5416;
wire n_14881;
wire n_18588;
wire n_14527;
wire n_12822;
wire n_13307;
wire n_7279;
wire n_17460;
wire n_13312;
wire n_11761;
wire n_9984;
wire n_8474;
wire n_3524;
wire n_489;
wire n_2885;
wire n_10600;
wire n_6102;
wire n_636;
wire n_10833;
wire n_18329;
wire n_18649;
wire n_13023;
wire n_20382;
wire n_19343;
wire n_1607;
wire n_1454;
wire n_15315;
wire n_19210;
wire n_11185;
wire n_13440;
wire n_869;
wire n_1154;
wire n_13436;
wire n_19615;
wire n_19133;
wire n_16982;
wire n_846;
wire n_841;
wire n_508;
wire n_11081;
wire n_16687;
wire n_1562;
wire n_14858;
wire n_8787;
wire n_13911;
wire n_5051;
wire n_17544;
wire n_5587;
wire n_20241;
wire n_10941;
wire n_14617;
wire n_9816;
wire n_17132;
wire n_14263;
wire n_661;
wire n_8605;
wire n_10358;
wire n_3565;
wire n_17593;
wire n_9944;
wire n_6998;
wire n_16158;
wire n_4173;
wire n_20105;
wire n_12338;
wire n_7615;
wire n_5651;
wire n_9605;
wire n_1217;
wire n_7591;
wire n_11404;
wire n_16488;
wire n_20584;
wire n_15994;
wire n_15685;
wire n_9788;
wire n_16273;
wire n_10785;
wire n_18262;
wire n_13872;
wire n_17646;
wire n_12341;
wire n_18389;
wire n_5412;
wire n_14475;
wire n_10815;
wire n_1120;
wire n_555;
wire n_8784;
wire n_7382;
wire n_2048;
wire n_13955;
wire n_176;
wire n_17708;
wire n_14400;
wire n_4857;
wire n_16725;
wire n_16904;
wire n_16432;
wire n_12085;
wire n_2883;
wire n_18190;
wire n_13554;
wire n_18421;
wire n_863;
wire n_6780;
wire n_11582;
wire n_20083;
wire n_3268;
wire n_1147;
wire n_1754;
wire n_11705;
wire n_3701;
wire n_7673;
wire n_1812;
wire n_6830;
wire n_17391;
wire n_19782;
wire n_17682;
wire n_7282;
wire n_9968;
wire n_11474;
wire n_10657;
wire n_13595;
wire n_5997;
wire n_2492;
wire n_10687;
wire n_13283;
wire n_19543;
wire n_15615;
wire n_12110;
wire n_8363;
wire n_5119;
wire n_19445;
wire n_17802;
wire n_9669;
wire n_17775;
wire n_6510;
wire n_8282;
wire n_5938;
wire n_15972;
wire n_6237;
wire n_12216;
wire n_12040;
wire n_11752;
wire n_17446;
wire n_2117;
wire n_18573;
wire n_14975;
wire n_7581;
wire n_6360;
wire n_17960;
wire n_15217;
wire n_4858;
wire n_13308;
wire n_19049;
wire n_9952;
wire n_15323;
wire n_12183;
wire n_19857;
wire n_10668;
wire n_9256;
wire n_5750;
wire n_4823;
wire n_4309;
wire n_839;
wire n_14007;
wire n_7346;
wire n_1537;
wire n_13373;
wire n_4243;
wire n_7428;
wire n_12221;
wire n_5666;
wire n_9195;
wire n_16236;
wire n_17787;
wire n_7283;
wire n_4142;
wire n_6314;
wire n_10632;
wire n_18861;
wire n_9623;
wire n_3796;
wire n_6964;
wire n_3408;
wire n_19027;
wire n_19561;
wire n_1184;
wire n_18912;
wire n_19322;
wire n_16702;
wire n_1525;
wire n_2594;
wire n_11329;
wire n_6495;
wire n_5994;
wire n_17280;
wire n_13241;
wire n_4244;
wire n_2147;
wire n_9516;
wire n_16027;
wire n_2503;
wire n_8976;
wire n_17844;
wire n_18136;
wire n_10130;
wire n_11661;
wire n_9222;
wire n_8435;
wire n_8882;
wire n_16391;
wire n_4787;
wire n_15949;
wire n_10622;
wire n_5633;
wire n_19840;
wire n_5664;
wire n_6797;
wire n_15673;
wire n_14012;
wire n_8759;
wire n_16941;
wire n_7177;
wire n_357;
wire n_13066;
wire n_13665;
wire n_12993;
wire n_19604;
wire n_11314;
wire n_17784;
wire n_2681;
wire n_15678;
wire n_13083;
wire n_8235;
wire n_3764;
wire n_19093;
wire n_16164;
wire n_6152;
wire n_16444;
wire n_4075;
wire n_9820;
wire n_14071;
wire n_12749;
wire n_2303;
wire n_1619;
wire n_8448;
wire n_4538;
wire n_12066;
wire n_6513;
wire n_2367;
wire n_1034;
wire n_15908;
wire n_754;
wire n_11184;
wire n_11945;
wire n_11368;
wire n_6330;
wire n_17842;
wire n_19628;
wire n_8457;
wire n_19200;
wire n_18605;
wire n_18837;
wire n_9339;
wire n_14312;
wire n_9601;
wire n_15045;
wire n_11409;
wire n_18995;
wire n_2107;
wire n_2040;
wire n_20393;
wire n_18737;
wire n_12437;
wire n_5624;
wire n_10840;
wire n_6263;
wire n_10515;
wire n_15501;
wire n_6490;
wire n_15751;
wire n_11605;
wire n_1861;
wire n_10242;
wire n_10144;
wire n_9684;
wire n_15741;
wire n_16195;
wire n_14793;
wire n_18754;
wire n_13472;
wire n_2162;
wire n_15596;
wire n_207;
wire n_4763;
wire n_3587;
wire n_205;
wire n_18316;
wire n_6038;
wire n_15379;
wire n_16272;
wire n_14884;
wire n_3162;
wire n_8964;
wire n_16629;
wire n_1899;
wire n_9814;
wire n_4804;
wire n_5619;
wire n_5859;
wire n_14423;
wire n_16280;
wire n_16414;
wire n_4500;
wire n_13443;
wire n_4433;
wire n_5644;
wire n_2813;
wire n_14626;
wire n_20058;
wire n_2027;
wire n_2091;
wire n_8960;
wire n_19899;
wire n_5030;
wire n_15402;
wire n_20563;
wire n_4194;
wire n_18026;
wire n_8443;
wire n_7715;
wire n_2419;
wire n_8683;
wire n_18558;
wire n_5683;
wire n_6349;
wire n_10510;
wire n_3182;
wire n_5756;
wire n_15306;
wire n_15981;
wire n_19994;
wire n_16367;

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_48),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_4),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_20),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_44),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_71),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_53),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_79),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_129),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_61),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_96),
.Y(n_146)
);

BUFx10_ASAP7_75t_L g147 ( 
.A(n_109),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_45),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_126),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_123),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_83),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_2),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_19),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_104),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_86),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_82),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_131),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_77),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_89),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_84),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_21),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_59),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_52),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_112),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_65),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_73),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_127),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_97),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_74),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_36),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_43),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_33),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_125),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_122),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_16),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_13),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_3),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_5),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_114),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_72),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_37),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_101),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_130),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_29),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_41),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_28),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_8),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_15),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_91),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_76),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_124),
.Y(n_191)
);

BUFx10_ASAP7_75t_L g192 ( 
.A(n_133),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_87),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_100),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_94),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_10),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_107),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_22),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_80),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_47),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_0),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_116),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_39),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_68),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_105),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_78),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_35),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_103),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_17),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_12),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_57),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_56),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_7),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_49),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_46),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_24),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_54),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_34),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_92),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_1),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_23),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_0),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_99),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_132),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_18),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_51),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_119),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_6),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_42),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_60),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_75),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_81),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_64),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_38),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_88),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_9),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_90),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_118),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_32),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_58),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_26),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_108),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_110),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_27),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_98),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_106),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_121),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_128),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_69),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_30),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_111),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_95),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_134),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_14),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_40),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_115),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_55),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_50),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_93),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_113),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_11),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_66),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_63),
.Y(n_263)
);

BUFx5_ASAP7_75t_L g264 ( 
.A(n_70),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_62),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_102),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_135),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_67),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_85),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_144),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_148),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_151),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_136),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_137),
.Y(n_274)
);

BUFx5_ASAP7_75t_L g275 ( 
.A(n_159),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_141),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_140),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_201),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_152),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_163),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_145),
.B(n_1),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_153),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_154),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_165),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_155),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_156),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_161),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_172),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_162),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_166),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_167),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_176),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_177),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_143),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_264),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_182),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_157),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_168),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_169),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_185),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_187),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_170),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_188),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_173),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_174),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_194),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_204),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_175),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_178),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_220),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_147),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_206),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_270),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_310),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_277),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_271),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_272),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_L g318 ( 
.A(n_273),
.B(n_191),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_274),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_276),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_311),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_280),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_284),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_279),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_288),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_292),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_293),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_296),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_275),
.Y(n_329)
);

NOR2xp67_ASAP7_75t_L g330 ( 
.A(n_282),
.B(n_138),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_300),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_283),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_301),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_285),
.B(n_193),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_281),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_303),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_306),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_307),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_294),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_286),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_287),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_289),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_312),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_295),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_290),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_297),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_291),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_275),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_298),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_299),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_275),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_275),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_278),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_275),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_302),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_304),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_305),
.Y(n_357)
);

CKINVDCx14_ASAP7_75t_R g358 ( 
.A(n_278),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_308),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_309),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_313),
.Y(n_361)
);

AND2x6_ASAP7_75t_L g362 ( 
.A(n_356),
.B(n_164),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_316),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_322),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_323),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_325),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_326),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_330),
.B(n_158),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_317),
.B(n_246),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_344),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_327),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_331),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_334),
.B(n_259),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_335),
.A2(n_234),
.B1(n_243),
.B2(n_224),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_333),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_360),
.B(n_314),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_347),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_359),
.A2(n_171),
.B1(n_247),
.B2(n_222),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_328),
.B(n_142),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_336),
.Y(n_380)
);

OA21x2_ASAP7_75t_L g381 ( 
.A1(n_351),
.A2(n_195),
.B(n_213),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_337),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_338),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_321),
.Y(n_384)
);

AOI22x1_ASAP7_75t_SL g385 ( 
.A1(n_315),
.A2(n_248),
.B1(n_150),
.B2(n_149),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_318),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_348),
.B(n_160),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_319),
.B(n_146),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_348),
.B(n_189),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_343),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_352),
.B(n_179),
.Y(n_391)
);

INVx5_ASAP7_75t_L g392 ( 
.A(n_329),
.Y(n_392)
);

AOI22x1_ASAP7_75t_SL g393 ( 
.A1(n_339),
.A2(n_260),
.B1(n_268),
.B2(n_267),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_354),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_320),
.Y(n_395)
);

CKINVDCx8_ASAP7_75t_R g396 ( 
.A(n_324),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_332),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_340),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_341),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_342),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_358),
.B(n_147),
.Y(n_401)
);

OA21x2_ASAP7_75t_L g402 ( 
.A1(n_345),
.A2(n_230),
.B(n_235),
.Y(n_402)
);

OAI21x1_ASAP7_75t_L g403 ( 
.A1(n_349),
.A2(n_228),
.B(n_252),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_350),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_355),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_357),
.A2(n_223),
.B1(n_266),
.B2(n_265),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_353),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_346),
.B(n_269),
.Y(n_408)
);

AND2x6_ASAP7_75t_L g409 ( 
.A(n_356),
.B(n_196),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_344),
.Y(n_410)
);

INVx6_ASAP7_75t_L g411 ( 
.A(n_315),
.Y(n_411)
);

BUFx8_ASAP7_75t_SL g412 ( 
.A(n_315),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_321),
.B(n_221),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_344),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_330),
.B(n_219),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_313),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_319),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_344),
.Y(n_418)
);

NOR2x1_ASAP7_75t_L g419 ( 
.A(n_330),
.B(n_217),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_334),
.A2(n_214),
.B1(n_263),
.B2(n_262),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_321),
.B(n_255),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_313),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_334),
.A2(n_218),
.B1(n_261),
.B2(n_256),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_330),
.B(n_216),
.Y(n_424)
);

BUFx8_ASAP7_75t_L g425 ( 
.A(n_356),
.Y(n_425)
);

OAI21x1_ASAP7_75t_L g426 ( 
.A1(n_348),
.A2(n_233),
.B(n_251),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_315),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_344),
.Y(n_428)
);

AND2x6_ASAP7_75t_L g429 ( 
.A(n_356),
.B(n_225),
.Y(n_429)
);

OA21x2_ASAP7_75t_L g430 ( 
.A1(n_351),
.A2(n_212),
.B(n_236),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_313),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_313),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_321),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_344),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_315),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_313),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_330),
.B(n_205),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_334),
.A2(n_215),
.B1(n_254),
.B2(n_253),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_321),
.Y(n_439)
);

OA21x2_ASAP7_75t_L g440 ( 
.A1(n_351),
.A2(n_227),
.B(n_211),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_313),
.Y(n_441)
);

INVx5_ASAP7_75t_L g442 ( 
.A(n_358),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_344),
.Y(n_443)
);

INVx5_ASAP7_75t_L g444 ( 
.A(n_358),
.Y(n_444)
);

CKINVDCx6p67_ASAP7_75t_R g445 ( 
.A(n_359),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_315),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_330),
.B(n_200),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_313),
.Y(n_448)
);

AO22x1_ASAP7_75t_L g449 ( 
.A1(n_334),
.A2(n_240),
.B1(n_209),
.B2(n_257),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_313),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_321),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_313),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_344),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_313),
.Y(n_454)
);

NOR2x1_ASAP7_75t_L g455 ( 
.A(n_330),
.B(n_242),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_344),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_313),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_344),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_334),
.B(n_210),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_344),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_344),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_321),
.B(n_208),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_344),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_313),
.Y(n_464)
);

OA21x2_ASAP7_75t_L g465 ( 
.A1(n_351),
.A2(n_198),
.B(n_250),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_313),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_347),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_321),
.B(n_192),
.Y(n_468)
);

AND2x6_ASAP7_75t_L g469 ( 
.A(n_356),
.B(n_225),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_335),
.A2(n_203),
.B1(n_244),
.B2(n_241),
.Y(n_470)
);

INVx5_ASAP7_75t_L g471 ( 
.A(n_358),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_334),
.B(n_207),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_315),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_335),
.A2(n_199),
.B1(n_239),
.B2(n_238),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_321),
.B(n_192),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_313),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_330),
.B(n_184),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_359),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_313),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_313),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_334),
.B(n_197),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_314),
.A2(n_226),
.B1(n_245),
.B2(n_237),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_321),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_344),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_313),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_359),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_313),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_344),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_313),
.Y(n_489)
);

AND2x6_ASAP7_75t_L g490 ( 
.A(n_356),
.B(n_242),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_344),
.Y(n_491)
);

BUFx8_ASAP7_75t_L g492 ( 
.A(n_356),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_334),
.B(n_202),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_364),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_370),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_361),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_371),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_459),
.B(n_180),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_365),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_366),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_373),
.B(n_186),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_410),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_414),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_382),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_367),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g506 ( 
.A(n_446),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_472),
.B(n_229),
.Y(n_507)
);

CKINVDCx6p67_ASAP7_75t_R g508 ( 
.A(n_442),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_422),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_431),
.Y(n_510)
);

OA21x2_ASAP7_75t_L g511 ( 
.A1(n_426),
.A2(n_249),
.B(n_232),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_473),
.Y(n_512)
);

NAND2xp33_ASAP7_75t_SL g513 ( 
.A(n_388),
.B(n_190),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_493),
.B(n_231),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_372),
.B(n_183),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_390),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_433),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_418),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_394),
.B(n_264),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_387),
.B(n_264),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_389),
.B(n_264),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_432),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_428),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_436),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_434),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_448),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_384),
.B(n_264),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_441),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_443),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_453),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_467),
.B(n_181),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_454),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_480),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_487),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_376),
.B(n_181),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_380),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_439),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_451),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_468),
.B(n_475),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_450),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_401),
.B(n_181),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_383),
.B(n_363),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_456),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_458),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_460),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_461),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_463),
.Y(n_547)
);

NAND2xp33_ASAP7_75t_L g548 ( 
.A(n_362),
.B(n_225),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_484),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_488),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_391),
.B(n_139),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_452),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_491),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_375),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_411),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_416),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_457),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_464),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_412),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_413),
.B(n_139),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_466),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_476),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_479),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_483),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_485),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_489),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_392),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_377),
.B(n_139),
.Y(n_568)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_445),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_392),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_405),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_403),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_430),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_402),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_379),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_478),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_369),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_486),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_397),
.B(n_242),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_462),
.Y(n_580)
);

BUFx8_ASAP7_75t_L g581 ( 
.A(n_395),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_421),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_440),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_381),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_465),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_368),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_386),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_455),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_407),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_427),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_449),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_419),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_482),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_481),
.A2(n_257),
.B1(n_258),
.B2(n_117),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_420),
.B(n_257),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_398),
.B(n_258),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_470),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_474),
.Y(n_598)
);

AND2x2_ASAP7_75t_SL g599 ( 
.A(n_435),
.B(n_258),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_396),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_399),
.B(n_25),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_415),
.B(n_31),
.Y(n_602)
);

AND2x6_ASAP7_75t_L g603 ( 
.A(n_404),
.B(n_408),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_429),
.Y(n_604)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_374),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_429),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_469),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_469),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_490),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_444),
.B(n_471),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_490),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_400),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_362),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_424),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_423),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_438),
.Y(n_616)
);

CKINVDCx11_ASAP7_75t_R g617 ( 
.A(n_417),
.Y(n_617)
);

AND3x1_ASAP7_75t_L g618 ( 
.A(n_406),
.B(n_385),
.C(n_393),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_437),
.B(n_447),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_477),
.B(n_409),
.Y(n_620)
);

OA21x2_ASAP7_75t_L g621 ( 
.A1(n_409),
.A2(n_378),
.B(n_425),
.Y(n_621)
);

INVx6_ASAP7_75t_L g622 ( 
.A(n_492),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_364),
.Y(n_623)
);

BUFx2_ASAP7_75t_L g624 ( 
.A(n_446),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_370),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_361),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_370),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_370),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_433),
.Y(n_629)
);

OR2x2_ASAP7_75t_L g630 ( 
.A(n_369),
.B(n_335),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_361),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_373),
.B(n_384),
.Y(n_632)
);

OA21x2_ASAP7_75t_L g633 ( 
.A1(n_426),
.A2(n_394),
.B(n_391),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_361),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_370),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_361),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_412),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_373),
.B(n_376),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_372),
.B(n_380),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_433),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_433),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_361),
.Y(n_642)
);

OA21x2_ASAP7_75t_L g643 ( 
.A1(n_426),
.A2(n_394),
.B(n_391),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_364),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_459),
.B(n_472),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_364),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_361),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_370),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_361),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_364),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_370),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_370),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_459),
.B(n_472),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_361),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_373),
.B(n_384),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_361),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_370),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_373),
.B(n_376),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_370),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_361),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_370),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_364),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_361),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_361),
.Y(n_664)
);

NAND2x1_ASAP7_75t_L g665 ( 
.A(n_394),
.B(n_381),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_361),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_361),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_370),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_SL g669 ( 
.A1(n_374),
.A2(n_294),
.B1(n_297),
.B2(n_277),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_370),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_384),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_361),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_373),
.B(n_459),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_361),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_412),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g676 ( 
.A(n_446),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_361),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_370),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_373),
.B(n_376),
.Y(n_679)
);

BUFx6f_ASAP7_75t_SL g680 ( 
.A(n_478),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_361),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_361),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_361),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_433),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_373),
.B(n_384),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_372),
.B(n_380),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_459),
.B(n_472),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_364),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_364),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_370),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_370),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_373),
.B(n_376),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_370),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_364),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_361),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_361),
.Y(n_696)
);

BUFx2_ASAP7_75t_L g697 ( 
.A(n_446),
.Y(n_697)
);

NAND2xp33_ASAP7_75t_SL g698 ( 
.A(n_388),
.B(n_467),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_364),
.Y(n_699)
);

OAI21x1_ASAP7_75t_L g700 ( 
.A1(n_426),
.A2(n_394),
.B(n_391),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_373),
.A2(n_376),
.B1(n_472),
.B2(n_459),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_411),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_364),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_370),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_459),
.B(n_472),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_361),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_361),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_361),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_433),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_361),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_361),
.Y(n_711)
);

AND2x6_ASAP7_75t_L g712 ( 
.A(n_376),
.B(n_397),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_370),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_370),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_361),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_361),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_361),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_364),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_361),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_361),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_361),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_370),
.Y(n_722)
);

BUFx2_ASAP7_75t_L g723 ( 
.A(n_446),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_373),
.B(n_376),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_361),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_361),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_373),
.A2(n_376),
.B1(n_472),
.B2(n_459),
.Y(n_727)
);

NAND2xp33_ASAP7_75t_L g728 ( 
.A(n_362),
.B(n_409),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_433),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_384),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_364),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_370),
.Y(n_732)
);

BUFx2_ASAP7_75t_L g733 ( 
.A(n_446),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_364),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_361),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_364),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_373),
.B(n_376),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_370),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_SL g739 ( 
.A(n_396),
.B(n_442),
.Y(n_739)
);

INVx6_ASAP7_75t_L g740 ( 
.A(n_411),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_361),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_370),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_364),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_459),
.B(n_472),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_361),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_370),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_361),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_364),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_361),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_433),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_372),
.B(n_380),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_361),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_412),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_459),
.B(n_472),
.Y(n_754)
);

OA21x2_ASAP7_75t_L g755 ( 
.A1(n_426),
.A2(n_394),
.B(n_391),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_361),
.Y(n_756)
);

AND2x2_ASAP7_75t_SL g757 ( 
.A(n_373),
.B(n_401),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_361),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_370),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_459),
.B(n_472),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_370),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_361),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_373),
.B(n_384),
.Y(n_763)
);

INVxp67_ASAP7_75t_L g764 ( 
.A(n_468),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_364),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_361),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_446),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_361),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_459),
.B(n_472),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_361),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_364),
.Y(n_771)
);

AND3x1_ASAP7_75t_L g772 ( 
.A(n_373),
.B(n_334),
.C(n_376),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_373),
.A2(n_376),
.B1(n_472),
.B2(n_459),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_459),
.B(n_472),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_361),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_459),
.B(n_472),
.Y(n_776)
);

OAI21x1_ASAP7_75t_L g777 ( 
.A1(n_426),
.A2(n_394),
.B(n_391),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_361),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_433),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_370),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_364),
.Y(n_781)
);

BUFx2_ASAP7_75t_L g782 ( 
.A(n_446),
.Y(n_782)
);

BUFx2_ASAP7_75t_L g783 ( 
.A(n_446),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_459),
.B(n_472),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_433),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_373),
.B(n_376),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_SL g787 ( 
.A(n_396),
.B(n_442),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_373),
.B(n_459),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_459),
.B(n_472),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_370),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_364),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_361),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_370),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_370),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_370),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_364),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_459),
.B(n_472),
.Y(n_797)
);

AND2x6_ASAP7_75t_L g798 ( 
.A(n_376),
.B(n_397),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_373),
.B(n_384),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_372),
.B(n_380),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_373),
.B(n_384),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_364),
.Y(n_802)
);

BUFx2_ASAP7_75t_L g803 ( 
.A(n_446),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_361),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_361),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_370),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_373),
.B(n_459),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_364),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_370),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_364),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_671),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_673),
.B(n_788),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_496),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_807),
.B(n_701),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_617),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_499),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_494),
.Y(n_817)
);

INVx4_ASAP7_75t_L g818 ( 
.A(n_571),
.Y(n_818)
);

INVx4_ASAP7_75t_L g819 ( 
.A(n_571),
.Y(n_819)
);

INVx4_ASAP7_75t_L g820 ( 
.A(n_600),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_727),
.B(n_773),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_645),
.B(n_653),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_555),
.B(n_702),
.Y(n_823)
);

INVxp67_ASAP7_75t_SL g824 ( 
.A(n_494),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_500),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_687),
.B(n_705),
.Y(n_826)
);

INVx1_ASAP7_75t_SL g827 ( 
.A(n_730),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_505),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_744),
.B(n_754),
.Y(n_829)
);

AO22x2_ASAP7_75t_L g830 ( 
.A1(n_605),
.A2(n_597),
.B1(n_598),
.B2(n_638),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_497),
.B(n_526),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_509),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_510),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_522),
.Y(n_834)
);

OR2x2_ASAP7_75t_L g835 ( 
.A(n_630),
.B(n_632),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_497),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_760),
.B(n_769),
.Y(n_837)
);

AND2x6_ASAP7_75t_L g838 ( 
.A(n_539),
.B(n_585),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_655),
.B(n_685),
.Y(n_839)
);

NOR2x1p5_ASAP7_75t_L g840 ( 
.A(n_508),
.B(n_600),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_774),
.B(n_776),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_784),
.B(n_789),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_528),
.Y(n_843)
);

NAND2xp33_ASAP7_75t_L g844 ( 
.A(n_797),
.B(n_613),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_532),
.Y(n_845)
);

OR2x2_ASAP7_75t_L g846 ( 
.A(n_763),
.B(n_799),
.Y(n_846)
);

INVx5_ASAP7_75t_L g847 ( 
.A(n_610),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_533),
.Y(n_848)
);

BUFx10_ASAP7_75t_L g849 ( 
.A(n_680),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_534),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_626),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_631),
.Y(n_852)
);

INVx5_ASAP7_75t_L g853 ( 
.A(n_578),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_578),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_501),
.B(n_575),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_634),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_517),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_801),
.B(n_757),
.Y(n_858)
);

INVx4_ASAP7_75t_L g859 ( 
.A(n_526),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_636),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_577),
.B(n_658),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_642),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_740),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_679),
.B(n_692),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_772),
.A2(n_737),
.B1(n_786),
.B2(n_724),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_647),
.Y(n_866)
);

XOR2xp5_ASAP7_75t_L g867 ( 
.A(n_669),
.B(n_590),
.Y(n_867)
);

BUFx10_ASAP7_75t_L g868 ( 
.A(n_637),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_531),
.B(n_764),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_649),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_654),
.Y(n_871)
);

INVx4_ASAP7_75t_L g872 ( 
.A(n_540),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_615),
.B(n_616),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_656),
.Y(n_874)
);

INVx6_ASAP7_75t_L g875 ( 
.A(n_581),
.Y(n_875)
);

INVx8_ASAP7_75t_L g876 ( 
.A(n_540),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_593),
.B(n_537),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_660),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_663),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_664),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_614),
.B(n_498),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_666),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_538),
.B(n_564),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_667),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_586),
.B(n_601),
.Y(n_885)
);

BUFx2_ASAP7_75t_L g886 ( 
.A(n_506),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_629),
.B(n_640),
.Y(n_887)
);

NAND2xp33_ASAP7_75t_L g888 ( 
.A(n_613),
.B(n_712),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_672),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_595),
.A2(n_574),
.B1(n_677),
.B2(n_674),
.Y(n_890)
);

AND2x2_ASAP7_75t_SL g891 ( 
.A(n_599),
.B(n_512),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_641),
.B(n_684),
.Y(n_892)
);

OR2x2_ASAP7_75t_L g893 ( 
.A(n_709),
.B(n_729),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_681),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_682),
.Y(n_895)
);

BUFx3_ASAP7_75t_L g896 ( 
.A(n_563),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_563),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_568),
.B(n_750),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_683),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_695),
.Y(n_900)
);

INVx4_ASAP7_75t_L g901 ( 
.A(n_566),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_696),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_706),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_707),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_566),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_708),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_507),
.B(n_514),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_574),
.A2(n_719),
.B1(n_720),
.B2(n_717),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_710),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_711),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_715),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_716),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_721),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_779),
.B(n_785),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_644),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_725),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_726),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_735),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_542),
.B(n_554),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_644),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_662),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_587),
.B(n_576),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_741),
.Y(n_923)
);

INVx4_ASAP7_75t_L g924 ( 
.A(n_662),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_688),
.B(n_694),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_619),
.A2(n_589),
.B1(n_804),
.B2(n_792),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_745),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_747),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_688),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_694),
.Y(n_930)
);

AND3x1_ASAP7_75t_L g931 ( 
.A(n_527),
.B(n_787),
.C(n_739),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_L g932 ( 
.A1(n_749),
.A2(n_805),
.B1(n_752),
.B2(n_778),
.Y(n_932)
);

XNOR2xp5_ASAP7_75t_L g933 ( 
.A(n_624),
.B(n_676),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_712),
.B(n_798),
.Y(n_934)
);

NAND3xp33_ASAP7_75t_L g935 ( 
.A(n_756),
.B(n_762),
.C(n_758),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_703),
.B(n_731),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_766),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_703),
.Y(n_938)
);

BUFx3_ASAP7_75t_L g939 ( 
.A(n_731),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_734),
.B(n_736),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_768),
.Y(n_941)
);

INVx5_ASAP7_75t_L g942 ( 
.A(n_622),
.Y(n_942)
);

INVx5_ASAP7_75t_L g943 ( 
.A(n_609),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_770),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_734),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_775),
.Y(n_946)
);

BUFx2_ASAP7_75t_L g947 ( 
.A(n_697),
.Y(n_947)
);

OR2x6_ASAP7_75t_L g948 ( 
.A(n_723),
.B(n_733),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_736),
.B(n_743),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_712),
.B(n_798),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_536),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_743),
.B(n_748),
.Y(n_952)
);

CKINVDCx6p67_ASAP7_75t_R g953 ( 
.A(n_559),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_798),
.B(n_535),
.Y(n_954)
);

INVxp33_ASAP7_75t_L g955 ( 
.A(n_612),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_748),
.B(n_765),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_767),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_556),
.B(n_557),
.Y(n_958)
);

INVx5_ASAP7_75t_L g959 ( 
.A(n_609),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_765),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_541),
.B(n_620),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_L g962 ( 
.A1(n_572),
.A2(n_583),
.B1(n_591),
.B2(n_573),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_545),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_771),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_782),
.Y(n_965)
);

INVx5_ASAP7_75t_L g966 ( 
.A(n_611),
.Y(n_966)
);

INVx4_ASAP7_75t_L g967 ( 
.A(n_771),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_495),
.B(n_502),
.Y(n_968)
);

OAI21xp33_ASAP7_75t_SL g969 ( 
.A1(n_584),
.A2(n_592),
.B(n_521),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_547),
.Y(n_970)
);

OR2x2_ASAP7_75t_L g971 ( 
.A(n_783),
.B(n_803),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_503),
.B(n_518),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_550),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_781),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_781),
.B(n_802),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_802),
.B(n_808),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_808),
.B(n_504),
.Y(n_977)
);

NAND2xp33_ASAP7_75t_SL g978 ( 
.A(n_611),
.B(n_604),
.Y(n_978)
);

AND2x2_ASAP7_75t_SL g979 ( 
.A(n_618),
.B(n_621),
.Y(n_979)
);

INVx6_ASAP7_75t_L g980 ( 
.A(n_579),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_596),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_523),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_553),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_516),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_525),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_529),
.Y(n_986)
);

INVx2_ASAP7_75t_SL g987 ( 
.A(n_560),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_569),
.Y(n_988)
);

OR2x6_ASAP7_75t_L g989 ( 
.A(n_580),
.B(n_524),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_530),
.B(n_543),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_544),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_552),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_546),
.B(n_549),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_639),
.B(n_686),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_625),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_751),
.B(n_800),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_627),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_628),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_635),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_582),
.B(n_698),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_648),
.B(n_651),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_588),
.B(n_652),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_657),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_623),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_646),
.B(n_689),
.Y(n_1005)
);

NOR2x1p5_ASAP7_75t_L g1006 ( 
.A(n_675),
.B(n_753),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_659),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_650),
.B(n_810),
.Y(n_1008)
);

INVx5_ASAP7_75t_L g1009 ( 
.A(n_603),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_809),
.B(n_690),
.Y(n_1010)
);

NAND2xp33_ASAP7_75t_L g1011 ( 
.A(n_603),
.B(n_572),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_661),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_806),
.B(n_691),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_699),
.B(n_796),
.Y(n_1014)
);

AND2x2_ASAP7_75t_SL g1015 ( 
.A(n_728),
.B(n_548),
.Y(n_1015)
);

CKINVDCx6p67_ASAP7_75t_R g1016 ( 
.A(n_603),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_718),
.Y(n_1017)
);

AND3x2_ASAP7_75t_L g1018 ( 
.A(n_606),
.B(n_608),
.C(n_607),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_668),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_520),
.A2(n_594),
.B1(n_746),
.B2(n_742),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_670),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_678),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_693),
.B(n_704),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_713),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_714),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_722),
.B(n_795),
.Y(n_1026)
);

INVx4_ASAP7_75t_L g1027 ( 
.A(n_791),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_732),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_794),
.B(n_793),
.Y(n_1029)
);

INVx2_ASAP7_75t_SL g1030 ( 
.A(n_515),
.Y(n_1030)
);

OR2x2_ASAP7_75t_L g1031 ( 
.A(n_558),
.B(n_561),
.Y(n_1031)
);

CKINVDCx16_ASAP7_75t_R g1032 ( 
.A(n_513),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_738),
.B(n_790),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_759),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_761),
.B(n_780),
.Y(n_1035)
);

OR2x6_ASAP7_75t_L g1036 ( 
.A(n_562),
.B(n_565),
.Y(n_1036)
);

BUFx3_ASAP7_75t_L g1037 ( 
.A(n_567),
.Y(n_1037)
);

INVx1_ASAP7_75t_SL g1038 ( 
.A(n_570),
.Y(n_1038)
);

INVx5_ASAP7_75t_L g1039 ( 
.A(n_519),
.Y(n_1039)
);

INVxp33_ASAP7_75t_L g1040 ( 
.A(n_551),
.Y(n_1040)
);

NAND2xp33_ASAP7_75t_L g1041 ( 
.A(n_602),
.B(n_665),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_633),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_643),
.B(n_755),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_700),
.B(n_777),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_511),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_571),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_496),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_571),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_496),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_673),
.B(n_788),
.Y(n_1050)
);

CKINVDCx8_ASAP7_75t_R g1051 ( 
.A(n_600),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_496),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_496),
.Y(n_1053)
);

BUFx3_ASAP7_75t_L g1054 ( 
.A(n_571),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_496),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_671),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_496),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_496),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_632),
.B(n_655),
.Y(n_1059)
);

AND2x6_ASAP7_75t_L g1060 ( 
.A(n_539),
.B(n_585),
.Y(n_1060)
);

OR2x6_ASAP7_75t_L g1061 ( 
.A(n_571),
.B(n_600),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_496),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_494),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_496),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_496),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_673),
.A2(n_807),
.B1(n_788),
.B2(n_769),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_673),
.B(n_788),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_494),
.Y(n_1068)
);

INVx5_ASAP7_75t_L g1069 ( 
.A(n_600),
.Y(n_1069)
);

INVx4_ASAP7_75t_L g1070 ( 
.A(n_571),
.Y(n_1070)
);

INVx4_ASAP7_75t_L g1071 ( 
.A(n_571),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_673),
.B(n_788),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_496),
.Y(n_1073)
);

NAND2xp33_ASAP7_75t_L g1074 ( 
.A(n_645),
.B(n_653),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_496),
.Y(n_1075)
);

INVx3_ASAP7_75t_L g1076 ( 
.A(n_494),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_496),
.Y(n_1077)
);

INVx8_ASAP7_75t_L g1078 ( 
.A(n_680),
.Y(n_1078)
);

INVx4_ASAP7_75t_L g1079 ( 
.A(n_571),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_632),
.B(n_655),
.Y(n_1080)
);

AOI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_673),
.A2(n_788),
.B1(n_807),
.B2(n_653),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_496),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_496),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_496),
.Y(n_1084)
);

NAND2xp33_ASAP7_75t_R g1085 ( 
.A(n_673),
.B(n_807),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_673),
.B(n_807),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_673),
.B(n_788),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_496),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_673),
.A2(n_788),
.B1(n_807),
.B2(n_653),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_673),
.B(n_788),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_571),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_571),
.B(n_555),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_632),
.B(n_655),
.Y(n_1093)
);

INVx4_ASAP7_75t_L g1094 ( 
.A(n_571),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_496),
.Y(n_1095)
);

OAI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_701),
.A2(n_773),
.B1(n_727),
.B2(n_645),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_673),
.B(n_807),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_632),
.B(n_655),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_673),
.B(n_788),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_496),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_673),
.B(n_788),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_496),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_673),
.B(n_788),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_496),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_671),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_673),
.B(n_807),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_673),
.B(n_807),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_673),
.B(n_807),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_571),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_673),
.B(n_807),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_673),
.B(n_807),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_673),
.B(n_788),
.Y(n_1112)
);

OAI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_701),
.A2(n_773),
.B1(n_727),
.B2(n_645),
.Y(n_1113)
);

CKINVDCx20_ASAP7_75t_R g1114 ( 
.A(n_617),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_496),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_496),
.Y(n_1116)
);

CKINVDCx20_ASAP7_75t_R g1117 ( 
.A(n_617),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_496),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_496),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_496),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_496),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_571),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_632),
.B(n_655),
.Y(n_1123)
);

NAND3xp33_ASAP7_75t_L g1124 ( 
.A(n_673),
.B(n_807),
.C(n_788),
.Y(n_1124)
);

OR2x2_ASAP7_75t_L g1125 ( 
.A(n_630),
.B(n_671),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_496),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_496),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_617),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_494),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_673),
.B(n_807),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_673),
.B(n_788),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_496),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_496),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_496),
.Y(n_1134)
);

INVx4_ASAP7_75t_L g1135 ( 
.A(n_571),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_673),
.A2(n_807),
.B1(n_788),
.B2(n_769),
.Y(n_1136)
);

OR2x6_ASAP7_75t_L g1137 ( 
.A(n_571),
.B(n_600),
.Y(n_1137)
);

OAI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_701),
.A2(n_773),
.B1(n_727),
.B2(n_645),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_673),
.B(n_788),
.Y(n_1139)
);

INVx1_ASAP7_75t_SL g1140 ( 
.A(n_671),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_673),
.B(n_788),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_673),
.B(n_788),
.Y(n_1142)
);

NOR2x1p5_ASAP7_75t_L g1143 ( 
.A(n_508),
.B(n_571),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_673),
.B(n_807),
.Y(n_1144)
);

OAI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_701),
.A2(n_773),
.B1(n_727),
.B2(n_645),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_673),
.B(n_807),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_571),
.Y(n_1147)
);

INVx4_ASAP7_75t_L g1148 ( 
.A(n_571),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_496),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_571),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_632),
.B(n_655),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_496),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_673),
.B(n_788),
.Y(n_1153)
);

CKINVDCx20_ASAP7_75t_R g1154 ( 
.A(n_617),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_673),
.A2(n_807),
.B1(n_788),
.B2(n_769),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_496),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_673),
.B(n_807),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_496),
.Y(n_1158)
);

OR2x2_ASAP7_75t_L g1159 ( 
.A(n_630),
.B(n_671),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_673),
.B(n_807),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_496),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_494),
.Y(n_1162)
);

INVx1_ASAP7_75t_SL g1163 ( 
.A(n_671),
.Y(n_1163)
);

INVxp67_ASAP7_75t_SL g1164 ( 
.A(n_494),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_496),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_632),
.B(n_655),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_673),
.B(n_788),
.Y(n_1167)
);

AND2x6_ASAP7_75t_L g1168 ( 
.A(n_539),
.B(n_585),
.Y(n_1168)
);

OR2x6_ASAP7_75t_L g1169 ( 
.A(n_571),
.B(n_600),
.Y(n_1169)
);

INVxp33_ASAP7_75t_L g1170 ( 
.A(n_517),
.Y(n_1170)
);

OR2x6_ASAP7_75t_L g1171 ( 
.A(n_571),
.B(n_600),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_496),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_494),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_496),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_496),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_632),
.B(n_655),
.Y(n_1176)
);

CKINVDCx14_ASAP7_75t_R g1177 ( 
.A(n_669),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_571),
.Y(n_1178)
);

AND2x6_ASAP7_75t_L g1179 ( 
.A(n_539),
.B(n_585),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_673),
.B(n_807),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_496),
.Y(n_1181)
);

NAND3xp33_ASAP7_75t_L g1182 ( 
.A(n_673),
.B(n_807),
.C(n_788),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_496),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_496),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_496),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_496),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_496),
.Y(n_1187)
);

INVx2_ASAP7_75t_SL g1188 ( 
.A(n_494),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_496),
.Y(n_1189)
);

OR2x6_ASAP7_75t_L g1190 ( 
.A(n_571),
.B(n_600),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_673),
.B(n_807),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_496),
.Y(n_1192)
);

XNOR2xp5_ASAP7_75t_L g1193 ( 
.A(n_669),
.B(n_315),
.Y(n_1193)
);

INVx2_ASAP7_75t_SL g1194 ( 
.A(n_494),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_496),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_673),
.B(n_807),
.Y(n_1196)
);

NAND2xp33_ASAP7_75t_L g1197 ( 
.A(n_645),
.B(n_653),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_673),
.A2(n_788),
.B1(n_807),
.B2(n_653),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_496),
.Y(n_1199)
);

NAND2x1p5_ASAP7_75t_L g1200 ( 
.A(n_571),
.B(n_494),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_496),
.Y(n_1201)
);

INVx6_ASAP7_75t_L g1202 ( 
.A(n_571),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_496),
.Y(n_1203)
);

INVxp67_ASAP7_75t_SL g1204 ( 
.A(n_494),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_673),
.A2(n_807),
.B1(n_788),
.B2(n_769),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_496),
.Y(n_1206)
);

AO22x2_ASAP7_75t_L g1207 ( 
.A1(n_605),
.A2(n_598),
.B1(n_597),
.B2(n_638),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_673),
.B(n_807),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_673),
.A2(n_807),
.B1(n_788),
.B2(n_769),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_496),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_494),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_496),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_494),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_673),
.B(n_788),
.Y(n_1214)
);

OR2x6_ASAP7_75t_L g1215 ( 
.A(n_571),
.B(n_600),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_673),
.B(n_807),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_496),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_673),
.B(n_788),
.Y(n_1218)
);

OAI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_701),
.A2(n_773),
.B1(n_727),
.B2(n_645),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_494),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_496),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_496),
.Y(n_1222)
);

OR2x6_ASAP7_75t_L g1223 ( 
.A(n_571),
.B(n_600),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_496),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_496),
.Y(n_1225)
);

NOR2x1p5_ASAP7_75t_L g1226 ( 
.A(n_508),
.B(n_571),
.Y(n_1226)
);

BUFx4f_ASAP7_75t_L g1227 ( 
.A(n_508),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_671),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_571),
.Y(n_1229)
);

INVxp67_ASAP7_75t_SL g1230 ( 
.A(n_494),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_496),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_494),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_496),
.Y(n_1233)
);

AND3x1_ASAP7_75t_L g1234 ( 
.A(n_597),
.B(n_373),
.C(n_598),
.Y(n_1234)
);

INVxp67_ASAP7_75t_SL g1235 ( 
.A(n_494),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_496),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_496),
.Y(n_1237)
);

INVx3_ASAP7_75t_L g1238 ( 
.A(n_494),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_496),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_496),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_673),
.B(n_807),
.Y(n_1241)
);

INVx4_ASAP7_75t_L g1242 ( 
.A(n_571),
.Y(n_1242)
);

INVx3_ASAP7_75t_L g1243 ( 
.A(n_494),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_496),
.Y(n_1244)
);

NAND2xp33_ASAP7_75t_L g1245 ( 
.A(n_645),
.B(n_653),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_673),
.B(n_788),
.Y(n_1246)
);

NOR2x1p5_ASAP7_75t_L g1247 ( 
.A(n_508),
.B(n_571),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_494),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_496),
.Y(n_1249)
);

OAI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_701),
.A2(n_773),
.B1(n_727),
.B2(n_645),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_571),
.B(n_555),
.Y(n_1251)
);

BUFx4f_ASAP7_75t_L g1252 ( 
.A(n_508),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_673),
.B(n_788),
.Y(n_1253)
);

INVx3_ASAP7_75t_L g1254 ( 
.A(n_494),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_673),
.B(n_788),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_496),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_673),
.B(n_788),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_496),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_673),
.B(n_807),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_673),
.B(n_788),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_673),
.B(n_807),
.Y(n_1261)
);

INVx6_ASAP7_75t_L g1262 ( 
.A(n_571),
.Y(n_1262)
);

OR2x6_ASAP7_75t_L g1263 ( 
.A(n_571),
.B(n_600),
.Y(n_1263)
);

INVx2_ASAP7_75t_SL g1264 ( 
.A(n_494),
.Y(n_1264)
);

NAND3xp33_ASAP7_75t_L g1265 ( 
.A(n_673),
.B(n_807),
.C(n_788),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_673),
.B(n_807),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_571),
.Y(n_1267)
);

BUFx8_ASAP7_75t_SL g1268 ( 
.A(n_637),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_571),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_571),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_571),
.Y(n_1271)
);

BUFx5_ASAP7_75t_L g1272 ( 
.A(n_838),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_813),
.Y(n_1273)
);

AND2x4_ASAP7_75t_L g1274 ( 
.A(n_853),
.B(n_1092),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_839),
.B(n_1059),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_829),
.B(n_841),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_816),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1087),
.B(n_1090),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1101),
.B(n_1141),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1142),
.B(n_1167),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1246),
.B(n_1086),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1097),
.B(n_1106),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_825),
.Y(n_1284)
);

OR2x2_ASAP7_75t_L g1285 ( 
.A(n_1107),
.B(n_1108),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_834),
.Y(n_1286)
);

BUFx3_ASAP7_75t_L g1287 ( 
.A(n_853),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1110),
.B(n_1111),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_848),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_SL g1290 ( 
.A(n_1251),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1130),
.B(n_1144),
.Y(n_1291)
);

NOR2xp67_ASAP7_75t_L g1292 ( 
.A(n_1069),
.B(n_820),
.Y(n_1292)
);

NAND2xp33_ASAP7_75t_L g1293 ( 
.A(n_1066),
.B(n_1136),
.Y(n_1293)
);

INVx8_ASAP7_75t_L g1294 ( 
.A(n_876),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_828),
.Y(n_1295)
);

NOR3xp33_ASAP7_75t_L g1296 ( 
.A(n_1124),
.B(n_1265),
.C(n_1182),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1080),
.B(n_1093),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_832),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1098),
.B(n_1123),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1146),
.B(n_1157),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_833),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_852),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1160),
.B(n_1180),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1191),
.B(n_1196),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1208),
.B(n_1216),
.Y(n_1305)
);

INVxp33_ASAP7_75t_L g1306 ( 
.A(n_1125),
.Y(n_1306)
);

AOI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1085),
.A2(n_1081),
.B1(n_1198),
.B2(n_1089),
.Y(n_1307)
);

INVxp67_ASAP7_75t_SL g1308 ( 
.A(n_1241),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1259),
.B(n_1261),
.Y(n_1309)
);

NOR3xp33_ASAP7_75t_L g1310 ( 
.A(n_1266),
.B(n_1113),
.C(n_1096),
.Y(n_1310)
);

NOR3xp33_ASAP7_75t_L g1311 ( 
.A(n_1138),
.B(n_1219),
.C(n_1145),
.Y(n_1311)
);

AND2x2_ASAP7_75t_SL g1312 ( 
.A(n_891),
.B(n_1155),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_812),
.B(n_1050),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1250),
.B(n_1205),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_843),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_860),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_845),
.Y(n_1317)
);

NOR3xp33_ASAP7_75t_L g1318 ( 
.A(n_821),
.B(n_814),
.C(n_1099),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_862),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_871),
.Y(n_1320)
);

INVxp67_ASAP7_75t_SL g1321 ( 
.A(n_826),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1209),
.A2(n_1112),
.B1(n_1131),
.B2(n_1103),
.Y(n_1322)
);

BUFx12f_ASAP7_75t_L g1323 ( 
.A(n_849),
.Y(n_1323)
);

NOR3xp33_ASAP7_75t_L g1324 ( 
.A(n_1139),
.B(n_1214),
.C(n_1153),
.Y(n_1324)
);

AND2x4_ASAP7_75t_L g1325 ( 
.A(n_863),
.B(n_823),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_874),
.Y(n_1326)
);

NOR3xp33_ASAP7_75t_L g1327 ( 
.A(n_1218),
.B(n_1255),
.C(n_1253),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_842),
.B(n_1257),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1260),
.B(n_822),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_855),
.B(n_837),
.Y(n_1330)
);

INVxp33_ASAP7_75t_L g1331 ( 
.A(n_1159),
.Y(n_1331)
);

NOR3xp33_ASAP7_75t_L g1332 ( 
.A(n_835),
.B(n_885),
.C(n_922),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_846),
.B(n_1151),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_878),
.Y(n_1334)
);

NOR2x1_ASAP7_75t_L g1335 ( 
.A(n_1006),
.B(n_818),
.Y(n_1335)
);

INVx2_ASAP7_75t_SL g1336 ( 
.A(n_1202),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_879),
.Y(n_1337)
);

NOR3xp33_ASAP7_75t_L g1338 ( 
.A(n_1166),
.B(n_1176),
.C(n_858),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1074),
.B(n_1197),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1245),
.B(n_881),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_864),
.B(n_861),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_865),
.B(n_1170),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_850),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_851),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_931),
.B(n_1234),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_856),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_898),
.B(n_869),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_827),
.B(n_1140),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_1163),
.B(n_857),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_880),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_893),
.B(n_883),
.Y(n_1351)
);

INVxp33_ASAP7_75t_L g1352 ( 
.A(n_887),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_907),
.B(n_961),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_892),
.B(n_914),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_926),
.B(n_873),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_866),
.Y(n_1356)
);

NOR3xp33_ASAP7_75t_L g1357 ( 
.A(n_811),
.B(n_1105),
.C(n_1056),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1228),
.B(n_877),
.Y(n_1358)
);

NOR3xp33_ASAP7_75t_L g1359 ( 
.A(n_1032),
.B(n_947),
.C(n_886),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_955),
.B(n_934),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_882),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_870),
.B(n_884),
.Y(n_1362)
);

CKINVDCx20_ASAP7_75t_R g1363 ( 
.A(n_1268),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_950),
.B(n_971),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_889),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_894),
.B(n_895),
.Y(n_1366)
);

INVx2_ASAP7_75t_SL g1367 ( 
.A(n_1262),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_L g1368 ( 
.A(n_957),
.B(n_965),
.Y(n_1368)
);

BUFx5_ASAP7_75t_L g1369 ( 
.A(n_838),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_844),
.B(n_988),
.Y(n_1370)
);

INVxp67_ASAP7_75t_L g1371 ( 
.A(n_1091),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_830),
.A2(n_1207),
.B1(n_899),
.B2(n_909),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_900),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1009),
.B(n_890),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_903),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_902),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_904),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_906),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_819),
.B(n_1070),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_SL g1380 ( 
.A(n_1009),
.B(n_911),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_1091),
.Y(n_1381)
);

BUFx3_ASAP7_75t_L g1382 ( 
.A(n_1109),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_910),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1061),
.Y(n_1384)
);

BUFx6f_ASAP7_75t_SL g1385 ( 
.A(n_1061),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1071),
.B(n_1079),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_912),
.B(n_916),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_L g1388 ( 
.A(n_1094),
.B(n_1135),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_923),
.B(n_927),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_928),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_937),
.B(n_1047),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_913),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1049),
.B(n_1052),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1053),
.B(n_1055),
.Y(n_1394)
);

NOR3xp33_ASAP7_75t_L g1395 ( 
.A(n_1177),
.B(n_1000),
.C(n_996),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1057),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1062),
.B(n_1064),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_917),
.B(n_918),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1065),
.B(n_1073),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1075),
.B(n_1077),
.Y(n_1400)
);

INVxp67_ASAP7_75t_L g1401 ( 
.A(n_1109),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1084),
.B(n_1095),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_SL g1403 ( 
.A1(n_979),
.A2(n_1030),
.B1(n_854),
.B2(n_944),
.Y(n_1403)
);

NOR2xp67_ASAP7_75t_L g1404 ( 
.A(n_1069),
.B(n_942),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_941),
.Y(n_1405)
);

NAND2xp33_ASAP7_75t_L g1406 ( 
.A(n_838),
.B(n_1060),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1100),
.B(n_1102),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_SL g1408 ( 
.A(n_946),
.B(n_1058),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1148),
.B(n_1242),
.Y(n_1409)
);

INVx2_ASAP7_75t_SL g1410 ( 
.A(n_1122),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1115),
.Y(n_1411)
);

NOR2xp67_ASAP7_75t_L g1412 ( 
.A(n_942),
.B(n_847),
.Y(n_1412)
);

BUFx6f_ASAP7_75t_SL g1413 ( 
.A(n_1137),
.Y(n_1413)
);

NOR3xp33_ASAP7_75t_L g1414 ( 
.A(n_994),
.B(n_935),
.C(n_888),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1116),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1118),
.B(n_1119),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1082),
.Y(n_1417)
);

NAND2xp33_ASAP7_75t_L g1418 ( 
.A(n_1060),
.B(n_1168),
.Y(n_1418)
);

INVx2_ASAP7_75t_SL g1419 ( 
.A(n_1122),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1147),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1083),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1088),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1126),
.B(n_1133),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1149),
.B(n_1152),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1158),
.Y(n_1425)
);

NAND2xp33_ASAP7_75t_L g1426 ( 
.A(n_1060),
.B(n_1168),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1038),
.B(n_1040),
.Y(n_1427)
);

INVx2_ASAP7_75t_SL g1428 ( 
.A(n_1147),
.Y(n_1428)
);

NAND2xp33_ASAP7_75t_L g1429 ( 
.A(n_1168),
.B(n_1179),
.Y(n_1429)
);

INVxp33_ASAP7_75t_L g1430 ( 
.A(n_933),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1161),
.B(n_1172),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1181),
.Y(n_1432)
);

NAND2xp33_ASAP7_75t_L g1433 ( 
.A(n_1179),
.B(n_908),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1271),
.B(n_1178),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1104),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1178),
.B(n_1271),
.Y(n_1436)
);

NOR3xp33_ASAP7_75t_L g1437 ( 
.A(n_1027),
.B(n_919),
.C(n_987),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1186),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1189),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1195),
.B(n_1203),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_SL g1441 ( 
.A(n_1120),
.B(n_1121),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1127),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1212),
.B(n_1217),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1222),
.Y(n_1444)
);

INVx1_ASAP7_75t_SL g1445 ( 
.A(n_1046),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1236),
.B(n_1237),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1132),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1267),
.B(n_1134),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_SL g1449 ( 
.A(n_1156),
.B(n_1165),
.Y(n_1449)
);

A2O1A1Ixp33_ASAP7_75t_L g1450 ( 
.A1(n_1174),
.A2(n_1210),
.B(n_1175),
.C(n_1183),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1240),
.B(n_1244),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1137),
.B(n_1169),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_SL g1453 ( 
.A(n_1184),
.B(n_1185),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1267),
.B(n_1187),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1192),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1256),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1199),
.B(n_1201),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_SL g1458 ( 
.A(n_1206),
.B(n_1221),
.Y(n_1458)
);

INVxp67_ASAP7_75t_L g1459 ( 
.A(n_1169),
.Y(n_1459)
);

BUFx12f_ASAP7_75t_SL g1460 ( 
.A(n_1171),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1224),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1225),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_SL g1463 ( 
.A(n_1231),
.B(n_1233),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1239),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1249),
.B(n_1258),
.Y(n_1465)
);

A2O1A1Ixp33_ASAP7_75t_L g1466 ( 
.A1(n_969),
.A2(n_993),
.B(n_958),
.C(n_954),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_L g1467 ( 
.A(n_854),
.B(n_1048),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_951),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_982),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1054),
.B(n_1150),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_963),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1171),
.B(n_1190),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_876),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_932),
.B(n_970),
.Y(n_1474)
);

NAND2xp33_ASAP7_75t_L g1475 ( 
.A(n_1179),
.B(n_962),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_SL g1476 ( 
.A(n_847),
.B(n_921),
.Y(n_1476)
);

NOR2xp67_ASAP7_75t_L g1477 ( 
.A(n_859),
.B(n_872),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_973),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_983),
.B(n_995),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_SL g1480 ( 
.A(n_921),
.B(n_929),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_998),
.B(n_999),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_929),
.B(n_831),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1022),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1229),
.B(n_1269),
.Y(n_1484)
);

BUFx6f_ASAP7_75t_L g1485 ( 
.A(n_1190),
.Y(n_1485)
);

NAND3xp33_ASAP7_75t_L g1486 ( 
.A(n_1193),
.B(n_1031),
.C(n_985),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1024),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_SL g1488 ( 
.A(n_1025),
.B(n_1028),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1270),
.B(n_867),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_901),
.B(n_924),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_968),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_SL g1492 ( 
.A(n_1215),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_972),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_990),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_967),
.B(n_824),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1164),
.B(n_1204),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_1051),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1215),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_986),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_SL g1500 ( 
.A(n_815),
.B(n_1128),
.Y(n_1500)
);

BUFx6f_ASAP7_75t_L g1501 ( 
.A(n_1223),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_L g1502 ( 
.A(n_1230),
.B(n_1235),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1001),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_991),
.B(n_997),
.Y(n_1504)
);

INVxp33_ASAP7_75t_L g1505 ( 
.A(n_1200),
.Y(n_1505)
);

AND2x6_ASAP7_75t_L g1506 ( 
.A(n_1003),
.B(n_1007),
.Y(n_1506)
);

XNOR2xp5_ASAP7_75t_L g1507 ( 
.A(n_840),
.B(n_948),
.Y(n_1507)
);

INVx1_ASAP7_75t_SL g1508 ( 
.A(n_1223),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1012),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1019),
.B(n_1021),
.Y(n_1510)
);

NOR2x1p5_ASAP7_75t_L g1511 ( 
.A(n_953),
.B(n_1016),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1034),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1002),
.B(n_836),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_897),
.B(n_905),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1023),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_930),
.B(n_938),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1263),
.B(n_1005),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1026),
.Y(n_1518)
);

A2O1A1Ixp33_ASAP7_75t_L g1519 ( 
.A1(n_1033),
.A2(n_1035),
.B(n_1015),
.C(n_1020),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1010),
.Y(n_1520)
);

NOR3xp33_ASAP7_75t_L g1521 ( 
.A(n_981),
.B(n_992),
.C(n_1004),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1039),
.B(n_1013),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1029),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1037),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1008),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1039),
.B(n_1042),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1017),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_960),
.B(n_1254),
.Y(n_1528)
);

NAND2xp33_ASAP7_75t_L g1529 ( 
.A(n_943),
.B(n_966),
.Y(n_1529)
);

CKINVDCx20_ASAP7_75t_R g1530 ( 
.A(n_1114),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_SL g1531 ( 
.A(n_943),
.B(n_959),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1014),
.Y(n_1532)
);

INVx2_ASAP7_75t_SL g1533 ( 
.A(n_1263),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_964),
.B(n_1248),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1063),
.B(n_1243),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1018),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1068),
.B(n_1213),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_R g1538 ( 
.A(n_1117),
.B(n_1154),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_L g1539 ( 
.A(n_1076),
.B(n_1211),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_925),
.Y(n_1540)
);

OR2x6_ASAP7_75t_L g1541 ( 
.A(n_1078),
.B(n_1247),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1036),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_936),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_SL g1544 ( 
.A(n_959),
.B(n_966),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_940),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1036),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1162),
.B(n_1238),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1011),
.A2(n_1045),
.B1(n_980),
.B2(n_978),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_949),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_L g1550 ( 
.A(n_1173),
.B(n_1232),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1220),
.B(n_817),
.Y(n_1551)
);

INVx2_ASAP7_75t_SL g1552 ( 
.A(n_896),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_SL g1553 ( 
.A(n_977),
.B(n_1264),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_915),
.Y(n_1554)
);

BUFx3_ASAP7_75t_L g1555 ( 
.A(n_939),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_952),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_945),
.B(n_989),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_920),
.B(n_1188),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_974),
.B(n_1129),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1194),
.B(n_984),
.Y(n_1560)
);

NAND2xp33_ASAP7_75t_L g1561 ( 
.A(n_1078),
.B(n_1226),
.Y(n_1561)
);

BUFx6f_ASAP7_75t_L g1562 ( 
.A(n_1227),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_989),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_956),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_SL g1565 ( 
.A(n_975),
.B(n_976),
.Y(n_1565)
);

BUFx6f_ASAP7_75t_L g1566 ( 
.A(n_1252),
.Y(n_1566)
);

BUFx3_ASAP7_75t_L g1567 ( 
.A(n_948),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_868),
.B(n_1043),
.Y(n_1568)
);

NOR3xp33_ASAP7_75t_L g1569 ( 
.A(n_1041),
.B(n_1044),
.C(n_1143),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_875),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_813),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_839),
.B(n_1059),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_813),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_816),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_813),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_813),
.Y(n_1577)
);

BUFx5_ASAP7_75t_L g1578 ( 
.A(n_838),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_L g1579 ( 
.A(n_1091),
.Y(n_1579)
);

NAND3xp33_ASAP7_75t_L g1580 ( 
.A(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_829),
.B(n_841),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_829),
.B(n_841),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_813),
.Y(n_1583)
);

BUFx6f_ASAP7_75t_SL g1584 ( 
.A(n_1092),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_829),
.B(n_841),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_829),
.B(n_841),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_L g1587 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_829),
.B(n_841),
.Y(n_1589)
);

INVxp67_ASAP7_75t_L g1590 ( 
.A(n_811),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_853),
.B(n_1092),
.Y(n_1591)
);

INVxp67_ASAP7_75t_SL g1592 ( 
.A(n_1067),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_813),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_813),
.Y(n_1594)
);

BUFx5_ASAP7_75t_L g1595 ( 
.A(n_838),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_829),
.B(n_841),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_829),
.B(n_841),
.Y(n_1597)
);

NAND3xp33_ASAP7_75t_L g1598 ( 
.A(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_SL g1601 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_SL g1602 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1602)
);

BUFx6f_ASAP7_75t_L g1603 ( 
.A(n_1091),
.Y(n_1603)
);

CKINVDCx20_ASAP7_75t_R g1604 ( 
.A(n_1268),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_SL g1605 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_1091),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_816),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_813),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_816),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_813),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_813),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_816),
.Y(n_1614)
);

BUFx5_ASAP7_75t_L g1615 ( 
.A(n_838),
.Y(n_1615)
);

NOR3xp33_ASAP7_75t_L g1616 ( 
.A(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_SL g1617 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1617)
);

INVx1_ASAP7_75t_SL g1618 ( 
.A(n_811),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_839),
.B(n_1059),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_813),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_816),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_SL g1624 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_816),
.Y(n_1625)
);

INVxp67_ASAP7_75t_L g1626 ( 
.A(n_811),
.Y(n_1626)
);

NOR3xp33_ASAP7_75t_L g1627 ( 
.A(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_1627)
);

BUFx6f_ASAP7_75t_L g1628 ( 
.A(n_1091),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1067),
.A2(n_1072),
.B1(n_1090),
.B2(n_1087),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_839),
.B(n_1059),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_816),
.Y(n_1631)
);

OAI221xp5_ASAP7_75t_L g1632 ( 
.A1(n_1067),
.A2(n_1087),
.B1(n_1101),
.B2(n_1090),
.C(n_1072),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_829),
.B(n_841),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_853),
.B(n_1092),
.Y(n_1634)
);

INVx2_ASAP7_75t_SL g1635 ( 
.A(n_853),
.Y(n_1635)
);

OAI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1081),
.A2(n_1089),
.B1(n_1198),
.B2(n_1136),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_816),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_SL g1638 ( 
.A(n_820),
.B(n_396),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_L g1639 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_813),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_SL g1641 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1641)
);

BUFx3_ASAP7_75t_L g1642 ( 
.A(n_853),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_813),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_829),
.B(n_841),
.Y(n_1644)
);

BUFx6f_ASAP7_75t_L g1645 ( 
.A(n_1091),
.Y(n_1645)
);

INVxp67_ASAP7_75t_SL g1646 ( 
.A(n_1067),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_813),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_816),
.Y(n_1648)
);

NOR3xp33_ASAP7_75t_L g1649 ( 
.A(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_SL g1650 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1651)
);

NOR3xp33_ASAP7_75t_L g1652 ( 
.A(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_SL g1653 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1653)
);

INVx3_ASAP7_75t_L g1654 ( 
.A(n_854),
.Y(n_1654)
);

INVxp33_ASAP7_75t_L g1655 ( 
.A(n_1125),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_816),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_813),
.Y(n_1657)
);

INVx2_ASAP7_75t_SL g1658 ( 
.A(n_853),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_829),
.B(n_841),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_829),
.B(n_841),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_813),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1268),
.Y(n_1662)
);

AO221x1_ASAP7_75t_L g1663 ( 
.A1(n_1096),
.A2(n_1113),
.B1(n_1219),
.B2(n_1145),
.C(n_1138),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_813),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_816),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1666)
);

NAND2xp33_ASAP7_75t_L g1667 ( 
.A(n_1066),
.B(n_1136),
.Y(n_1667)
);

BUFx3_ASAP7_75t_L g1668 ( 
.A(n_853),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_829),
.B(n_841),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_813),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_816),
.Y(n_1671)
);

INVxp67_ASAP7_75t_SL g1672 ( 
.A(n_1067),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_813),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_SL g1674 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1674)
);

INVx2_ASAP7_75t_SL g1675 ( 
.A(n_853),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_SL g1676 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_816),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_816),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_813),
.Y(n_1679)
);

INVx3_ASAP7_75t_L g1680 ( 
.A(n_854),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_813),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_SL g1682 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_816),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_813),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_829),
.B(n_841),
.Y(n_1685)
);

NAND3xp33_ASAP7_75t_L g1686 ( 
.A(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_829),
.B(n_841),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_813),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_829),
.B(n_841),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_813),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_829),
.B(n_841),
.Y(n_1691)
);

NOR2x1p5_ASAP7_75t_L g1692 ( 
.A(n_820),
.B(n_508),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_829),
.B(n_841),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_813),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_SL g1695 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_816),
.Y(n_1696)
);

INVxp67_ASAP7_75t_SL g1697 ( 
.A(n_1067),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_829),
.B(n_841),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_816),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_829),
.B(n_841),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_SL g1701 ( 
.A1(n_1067),
.A2(n_1087),
.B1(n_1090),
.B2(n_1072),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1702)
);

INVx3_ASAP7_75t_L g1703 ( 
.A(n_854),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_829),
.B(n_841),
.Y(n_1704)
);

BUFx6f_ASAP7_75t_L g1705 ( 
.A(n_1091),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_SL g1706 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_829),
.B(n_841),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_816),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_L g1712 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_SL g1713 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_816),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_829),
.B(n_841),
.Y(n_1715)
);

INVx2_ASAP7_75t_SL g1716 ( 
.A(n_853),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_829),
.B(n_841),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_816),
.Y(n_1718)
);

A2O1A1Ixp33_ASAP7_75t_L g1719 ( 
.A1(n_1067),
.A2(n_1087),
.B(n_1090),
.C(n_1072),
.Y(n_1719)
);

NOR2xp67_ASAP7_75t_L g1720 ( 
.A(n_1069),
.B(n_853),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_816),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_813),
.Y(n_1722)
);

INVx2_ASAP7_75t_SL g1723 ( 
.A(n_853),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_829),
.B(n_841),
.Y(n_1724)
);

INVx2_ASAP7_75t_SL g1725 ( 
.A(n_853),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_816),
.Y(n_1726)
);

INVxp67_ASAP7_75t_L g1727 ( 
.A(n_811),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_829),
.B(n_841),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_829),
.B(n_841),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_813),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_816),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_829),
.B(n_841),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_829),
.B(n_841),
.Y(n_1734)
);

BUFx6f_ASAP7_75t_L g1735 ( 
.A(n_1091),
.Y(n_1735)
);

INVx8_ASAP7_75t_L g1736 ( 
.A(n_876),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1737)
);

INVxp33_ASAP7_75t_L g1738 ( 
.A(n_1125),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_813),
.Y(n_1740)
);

NAND3xp33_ASAP7_75t_SL g1741 ( 
.A(n_1081),
.B(n_1198),
.C(n_1089),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_813),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_829),
.B(n_841),
.Y(n_1743)
);

BUFx6f_ASAP7_75t_L g1744 ( 
.A(n_1091),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_L g1745 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1745)
);

AND2x2_ASAP7_75t_SL g1746 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_816),
.Y(n_1747)
);

INVx2_ASAP7_75t_SL g1748 ( 
.A(n_853),
.Y(n_1748)
);

INVxp67_ASAP7_75t_L g1749 ( 
.A(n_811),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_829),
.B(n_841),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1751)
);

OA21x2_ASAP7_75t_L g1752 ( 
.A1(n_1043),
.A2(n_585),
.B(n_1042),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_1268),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_813),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_829),
.B(n_841),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_SL g1756 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_813),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_L g1758 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1758)
);

XNOR2xp5_ASAP7_75t_L g1759 ( 
.A(n_1193),
.B(n_315),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_813),
.Y(n_1760)
);

NOR3xp33_ASAP7_75t_L g1761 ( 
.A(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_1761)
);

AOI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1067),
.A2(n_1087),
.B1(n_1090),
.B2(n_1072),
.Y(n_1762)
);

BUFx3_ASAP7_75t_L g1763 ( 
.A(n_853),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_813),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_839),
.B(n_1059),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_813),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_L g1767 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_813),
.Y(n_1768)
);

BUFx5_ASAP7_75t_L g1769 ( 
.A(n_838),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_829),
.B(n_841),
.Y(n_1770)
);

INVxp67_ASAP7_75t_SL g1771 ( 
.A(n_1067),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_813),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_816),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_829),
.B(n_841),
.Y(n_1774)
);

BUFx3_ASAP7_75t_L g1775 ( 
.A(n_853),
.Y(n_1775)
);

NOR3xp33_ASAP7_75t_L g1776 ( 
.A(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_829),
.B(n_841),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_SL g1778 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1778)
);

A2O1A1Ixp33_ASAP7_75t_L g1779 ( 
.A1(n_1067),
.A2(n_1087),
.B(n_1090),
.C(n_1072),
.Y(n_1779)
);

HB1xp67_ASAP7_75t_L g1780 ( 
.A(n_811),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_829),
.B(n_841),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_829),
.B(n_841),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_829),
.B(n_841),
.Y(n_1783)
);

BUFx6f_ASAP7_75t_L g1784 ( 
.A(n_1091),
.Y(n_1784)
);

BUFx6f_ASAP7_75t_L g1785 ( 
.A(n_1091),
.Y(n_1785)
);

NOR2xp67_ASAP7_75t_L g1786 ( 
.A(n_1069),
.B(n_853),
.Y(n_1786)
);

NAND3xp33_ASAP7_75t_L g1787 ( 
.A(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_829),
.B(n_841),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1789)
);

OAI21xp33_ASAP7_75t_L g1790 ( 
.A1(n_1067),
.A2(n_1087),
.B(n_1072),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_816),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_829),
.B(n_841),
.Y(n_1792)
);

BUFx6f_ASAP7_75t_L g1793 ( 
.A(n_1091),
.Y(n_1793)
);

NOR2xp67_ASAP7_75t_L g1794 ( 
.A(n_1069),
.B(n_853),
.Y(n_1794)
);

INVx2_ASAP7_75t_SL g1795 ( 
.A(n_853),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_816),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_816),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_829),
.B(n_841),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_829),
.B(n_841),
.Y(n_1800)
);

BUFx6f_ASAP7_75t_L g1801 ( 
.A(n_1091),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_829),
.B(n_841),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_813),
.Y(n_1803)
);

OAI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_829),
.A2(n_788),
.B(n_673),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_816),
.Y(n_1805)
);

XNOR2xp5_ASAP7_75t_L g1806 ( 
.A(n_1193),
.B(n_315),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_829),
.B(n_841),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_816),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_SL g1809 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_813),
.Y(n_1810)
);

BUFx6f_ASAP7_75t_L g1811 ( 
.A(n_1091),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_816),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_829),
.B(n_841),
.Y(n_1813)
);

NOR3xp33_ASAP7_75t_L g1814 ( 
.A(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_1814)
);

AND2x6_ASAP7_75t_SL g1815 ( 
.A(n_1061),
.B(n_1137),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_829),
.B(n_841),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_816),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_813),
.Y(n_1818)
);

INVx1_ASAP7_75t_SL g1819 ( 
.A(n_811),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_813),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_813),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_829),
.B(n_841),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_SL g1823 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_829),
.B(n_841),
.Y(n_1824)
);

AND2x4_ASAP7_75t_L g1825 ( 
.A(n_853),
.B(n_1092),
.Y(n_1825)
);

INVxp33_ASAP7_75t_L g1826 ( 
.A(n_1125),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_816),
.Y(n_1827)
);

INVxp67_ASAP7_75t_L g1828 ( 
.A(n_811),
.Y(n_1828)
);

INVx2_ASAP7_75t_SL g1829 ( 
.A(n_853),
.Y(n_1829)
);

NOR2x1p5_ASAP7_75t_L g1830 ( 
.A(n_820),
.B(n_508),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_816),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_SL g1832 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_829),
.B(n_841),
.Y(n_1833)
);

NOR2xp33_ASAP7_75t_L g1834 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1834)
);

AO221x1_ASAP7_75t_L g1835 ( 
.A1(n_1096),
.A2(n_1113),
.B1(n_1219),
.B2(n_1145),
.C(n_1138),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_SL g1836 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1836)
);

AND2x6_ASAP7_75t_L g1837 ( 
.A(n_934),
.B(n_950),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_813),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_829),
.B(n_841),
.Y(n_1839)
);

NAND3xp33_ASAP7_75t_L g1840 ( 
.A(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_816),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_SL g1842 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_829),
.B(n_841),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_SL g1844 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_SL g1845 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1845)
);

XNOR2xp5_ASAP7_75t_L g1846 ( 
.A(n_1193),
.B(n_315),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_813),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_829),
.B(n_841),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_829),
.B(n_841),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_816),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_816),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_SL g1852 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1852)
);

NOR3xp33_ASAP7_75t_L g1853 ( 
.A(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_829),
.B(n_841),
.Y(n_1855)
);

INVx4_ASAP7_75t_L g1856 ( 
.A(n_853),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_L g1858 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1858)
);

INVx2_ASAP7_75t_SL g1859 ( 
.A(n_853),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_829),
.B(n_841),
.Y(n_1860)
);

NOR3xp33_ASAP7_75t_L g1861 ( 
.A(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_1861)
);

NAND3xp33_ASAP7_75t_L g1862 ( 
.A(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_829),
.B(n_841),
.Y(n_1863)
);

NOR2xp67_ASAP7_75t_L g1864 ( 
.A(n_1069),
.B(n_853),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_813),
.Y(n_1865)
);

A2O1A1Ixp33_ASAP7_75t_L g1866 ( 
.A1(n_1067),
.A2(n_1087),
.B(n_1090),
.C(n_1072),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_829),
.B(n_841),
.Y(n_1867)
);

BUFx6f_ASAP7_75t_L g1868 ( 
.A(n_1091),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_SL g1869 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1869)
);

INVxp67_ASAP7_75t_SL g1870 ( 
.A(n_1067),
.Y(n_1870)
);

NOR2xp33_ASAP7_75t_L g1871 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1871)
);

BUFx6f_ASAP7_75t_L g1872 ( 
.A(n_1091),
.Y(n_1872)
);

INVx2_ASAP7_75t_SL g1873 ( 
.A(n_853),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_829),
.B(n_841),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_813),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_813),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_813),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_SL g1878 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1878)
);

INVx1_ASAP7_75t_SL g1879 ( 
.A(n_811),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_829),
.B(n_841),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_L g1881 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1881)
);

INVxp67_ASAP7_75t_L g1882 ( 
.A(n_811),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_829),
.B(n_841),
.Y(n_1884)
);

INVxp67_ASAP7_75t_L g1885 ( 
.A(n_811),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_813),
.Y(n_1886)
);

INVx2_ASAP7_75t_SL g1887 ( 
.A(n_853),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_829),
.B(n_841),
.Y(n_1888)
);

BUFx6f_ASAP7_75t_L g1889 ( 
.A(n_1091),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_SL g1890 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_816),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1892)
);

BUFx6f_ASAP7_75t_L g1893 ( 
.A(n_1091),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_829),
.B(n_841),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_829),
.B(n_841),
.Y(n_1895)
);

NAND2xp33_ASAP7_75t_SL g1896 ( 
.A(n_1086),
.B(n_1097),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_813),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_816),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_829),
.B(n_841),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_829),
.B(n_841),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_829),
.B(n_841),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_L g1902 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1902)
);

AOI21x1_ASAP7_75t_L g1903 ( 
.A1(n_954),
.A2(n_1045),
.B(n_585),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_813),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_SL g1905 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_829),
.B(n_841),
.Y(n_1906)
);

INVx4_ASAP7_75t_SL g1907 ( 
.A(n_1202),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_816),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_839),
.B(n_1059),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_816),
.Y(n_1910)
);

NOR2xp33_ASAP7_75t_L g1911 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1911)
);

NOR2xp67_ASAP7_75t_L g1912 ( 
.A(n_1069),
.B(n_853),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_816),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_829),
.B(n_841),
.Y(n_1914)
);

INVxp33_ASAP7_75t_L g1915 ( 
.A(n_1125),
.Y(n_1915)
);

NAND3xp33_ASAP7_75t_L g1916 ( 
.A(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_829),
.B(n_841),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_816),
.Y(n_1918)
);

BUFx6f_ASAP7_75t_L g1919 ( 
.A(n_1091),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_SL g1920 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1920)
);

NOR2xp67_ASAP7_75t_L g1921 ( 
.A(n_1069),
.B(n_853),
.Y(n_1921)
);

NOR2xp33_ASAP7_75t_L g1922 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_816),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_SL g1924 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_SL g1925 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_SL g1926 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1926)
);

AOI221xp5_ASAP7_75t_L g1927 ( 
.A1(n_1067),
.A2(n_1072),
.B1(n_1101),
.B2(n_1090),
.C(n_1087),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_L g1928 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1928)
);

NOR2xp33_ASAP7_75t_L g1929 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1929)
);

INVx3_ASAP7_75t_L g1930 ( 
.A(n_854),
.Y(n_1930)
);

NOR2xp33_ASAP7_75t_SL g1931 ( 
.A(n_820),
.B(n_396),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_829),
.B(n_841),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_813),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_813),
.Y(n_1934)
);

NOR2xp33_ASAP7_75t_L g1935 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_L g1936 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_813),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_829),
.B(n_841),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_829),
.B(n_841),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_816),
.Y(n_1940)
);

NOR2xp33_ASAP7_75t_SL g1941 ( 
.A(n_820),
.B(n_396),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_SL g1942 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_829),
.B(n_841),
.Y(n_1944)
);

NAND3xp33_ASAP7_75t_L g1945 ( 
.A(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1946)
);

AO221x1_ASAP7_75t_L g1947 ( 
.A1(n_1096),
.A2(n_1113),
.B1(n_1219),
.B2(n_1145),
.C(n_1138),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_829),
.B(n_841),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_SL g1949 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_SL g1950 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1950)
);

INVxp67_ASAP7_75t_L g1951 ( 
.A(n_811),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_813),
.Y(n_1952)
);

NOR2xp67_ASAP7_75t_L g1953 ( 
.A(n_1069),
.B(n_853),
.Y(n_1953)
);

NAND2xp33_ASAP7_75t_L g1954 ( 
.A(n_1066),
.B(n_1136),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_SL g1955 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_829),
.B(n_841),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_816),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_813),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_816),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_SL g1960 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_SL g1961 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1961)
);

NOR2xp33_ASAP7_75t_L g1962 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_813),
.Y(n_1963)
);

INVxp67_ASAP7_75t_L g1964 ( 
.A(n_811),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_816),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_829),
.B(n_841),
.Y(n_1966)
);

BUFx2_ASAP7_75t_L g1967 ( 
.A(n_811),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_829),
.B(n_841),
.Y(n_1968)
);

AOI221xp5_ASAP7_75t_L g1969 ( 
.A1(n_1067),
.A2(n_1072),
.B1(n_1101),
.B2(n_1090),
.C(n_1087),
.Y(n_1969)
);

NOR3xp33_ASAP7_75t_L g1970 ( 
.A(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_1970)
);

INVxp33_ASAP7_75t_L g1971 ( 
.A(n_1125),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_829),
.B(n_841),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_L g1973 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1973)
);

NOR2xp33_ASAP7_75t_L g1974 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1974)
);

INVx2_ASAP7_75t_SL g1975 ( 
.A(n_853),
.Y(n_1975)
);

INVxp67_ASAP7_75t_L g1976 ( 
.A(n_811),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_SL g1977 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1977)
);

NOR2xp67_ASAP7_75t_L g1978 ( 
.A(n_1069),
.B(n_853),
.Y(n_1978)
);

XOR2xp5_ASAP7_75t_L g1979 ( 
.A(n_933),
.B(n_446),
.Y(n_1979)
);

NOR2xp67_ASAP7_75t_L g1980 ( 
.A(n_1069),
.B(n_853),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_SL g1981 ( 
.A(n_1081),
.B(n_1089),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_813),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_816),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_829),
.B(n_841),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_829),
.B(n_841),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_816),
.Y(n_1986)
);

NAND3xp33_ASAP7_75t_SL g1987 ( 
.A(n_1804),
.B(n_1969),
.C(n_1927),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_SL g1988 ( 
.A(n_1636),
.B(n_1310),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1277),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1275),
.B(n_1297),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1276),
.B(n_1581),
.Y(n_1991)
);

BUFx2_ASAP7_75t_L g1992 ( 
.A(n_1967),
.Y(n_1992)
);

AOI22xp5_ASAP7_75t_L g1993 ( 
.A1(n_1280),
.A2(n_1587),
.B1(n_1599),
.B2(n_1588),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1284),
.Y(n_1994)
);

AND2x6_ASAP7_75t_SL g1995 ( 
.A(n_1489),
.B(n_1541),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1295),
.Y(n_1996)
);

NOR2xp33_ASAP7_75t_SL g1997 ( 
.A(n_1662),
.B(n_1753),
.Y(n_1997)
);

INVx2_ASAP7_75t_SL g1998 ( 
.A(n_1294),
.Y(n_1998)
);

AND2x4_ASAP7_75t_L g1999 ( 
.A(n_1335),
.B(n_1395),
.Y(n_1999)
);

NOR2xp33_ASAP7_75t_SL g2000 ( 
.A(n_1638),
.B(n_1931),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1582),
.B(n_1585),
.Y(n_2001)
);

AOI22xp33_ASAP7_75t_L g2002 ( 
.A1(n_1311),
.A2(n_1741),
.B1(n_1627),
.B2(n_1649),
.Y(n_2002)
);

O2A1O1Ixp33_ASAP7_75t_L g2003 ( 
.A1(n_1719),
.A2(n_1779),
.B(n_1866),
.C(n_1632),
.Y(n_2003)
);

OAI221xp5_ASAP7_75t_L g2004 ( 
.A1(n_1629),
.A2(n_1701),
.B1(n_1762),
.B2(n_1619),
.C(n_1620),
.Y(n_2004)
);

AOI21xp5_ASAP7_75t_L g2005 ( 
.A1(n_1321),
.A2(n_1353),
.B(n_1340),
.Y(n_2005)
);

NAND3xp33_ASAP7_75t_SL g2006 ( 
.A(n_1616),
.B(n_1761),
.C(n_1652),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1298),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1586),
.B(n_1589),
.Y(n_2008)
);

INVx5_ASAP7_75t_L g2009 ( 
.A(n_1506),
.Y(n_2009)
);

AOI22xp33_ASAP7_75t_L g2010 ( 
.A1(n_1776),
.A2(n_1853),
.B1(n_1861),
.B2(n_1814),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1596),
.B(n_1597),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1633),
.B(n_1644),
.Y(n_2012)
);

AOI22xp5_ASAP7_75t_L g2013 ( 
.A1(n_1609),
.A2(n_1611),
.B1(n_1651),
.B2(n_1639),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1659),
.B(n_1660),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1669),
.B(n_1685),
.Y(n_2015)
);

AOI22xp33_ASAP7_75t_L g2016 ( 
.A1(n_1970),
.A2(n_1293),
.B1(n_1954),
.B2(n_1667),
.Y(n_2016)
);

AOI22xp5_ASAP7_75t_L g2017 ( 
.A1(n_1666),
.A2(n_1702),
.B1(n_1711),
.B2(n_1707),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1687),
.B(n_1689),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1301),
.Y(n_2019)
);

CKINVDCx5p33_ASAP7_75t_R g2020 ( 
.A(n_1538),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_SL g2021 ( 
.A(n_1318),
.B(n_1307),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1691),
.B(n_1693),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1299),
.B(n_1572),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_SL g2024 ( 
.A(n_1314),
.B(n_1574),
.Y(n_2024)
);

NOR2xp33_ASAP7_75t_L g2025 ( 
.A(n_1712),
.B(n_1737),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1698),
.B(n_1700),
.Y(n_2026)
);

NAND2x1_ASAP7_75t_L g2027 ( 
.A(n_1506),
.B(n_1837),
.Y(n_2027)
);

INVx3_ASAP7_75t_L g2028 ( 
.A(n_1506),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1315),
.Y(n_2029)
);

NOR2xp33_ASAP7_75t_L g2030 ( 
.A(n_1739),
.B(n_1745),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1317),
.Y(n_2031)
);

AOI22xp5_ASAP7_75t_L g2032 ( 
.A1(n_1751),
.A2(n_1758),
.B1(n_1789),
.B2(n_1767),
.Y(n_2032)
);

NOR2xp67_ASAP7_75t_L g2033 ( 
.A(n_1349),
.B(n_1486),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1343),
.Y(n_2034)
);

NOR2xp67_ASAP7_75t_L g2035 ( 
.A(n_1348),
.B(n_1856),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1704),
.B(n_1709),
.Y(n_2036)
);

AND2x4_ASAP7_75t_L g2037 ( 
.A(n_1517),
.B(n_1563),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1344),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1715),
.B(n_1717),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1346),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1724),
.B(n_1728),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1729),
.B(n_1733),
.Y(n_2042)
);

AOI22xp5_ASAP7_75t_L g2043 ( 
.A1(n_1797),
.A2(n_1834),
.B1(n_1857),
.B2(n_1854),
.Y(n_2043)
);

NOR2xp33_ASAP7_75t_L g2044 ( 
.A(n_1858),
.B(n_1871),
.Y(n_2044)
);

NOR2xp33_ASAP7_75t_L g2045 ( 
.A(n_1881),
.B(n_1883),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1734),
.B(n_1743),
.Y(n_2046)
);

NOR2xp33_ASAP7_75t_L g2047 ( 
.A(n_1902),
.B(n_1911),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1356),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1621),
.B(n_1630),
.Y(n_2049)
);

AOI22xp33_ASAP7_75t_L g2050 ( 
.A1(n_1600),
.A2(n_1602),
.B1(n_1605),
.B2(n_1601),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1750),
.B(n_1755),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1770),
.B(n_1774),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1777),
.B(n_1781),
.Y(n_2053)
);

BUFx6f_ASAP7_75t_L g2054 ( 
.A(n_1381),
.Y(n_2054)
);

AOI22xp33_ASAP7_75t_L g2055 ( 
.A1(n_1617),
.A2(n_1641),
.B1(n_1650),
.B2(n_1624),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1365),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1373),
.Y(n_2057)
);

INVxp67_ASAP7_75t_L g2058 ( 
.A(n_1780),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1375),
.Y(n_2059)
);

NOR2xp33_ASAP7_75t_L g2060 ( 
.A(n_1922),
.B(n_1928),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1782),
.B(n_1783),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_1765),
.B(n_1909),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1788),
.B(n_1792),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1377),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_SL g2065 ( 
.A(n_1746),
.B(n_1358),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_1592),
.B(n_1646),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1799),
.B(n_1800),
.Y(n_2067)
);

INVxp67_ASAP7_75t_L g2068 ( 
.A(n_1351),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_SL g2069 ( 
.A(n_1354),
.B(n_1352),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1802),
.B(n_1807),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_SL g2071 ( 
.A(n_1332),
.B(n_1333),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1378),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1813),
.B(n_1816),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_SL g2074 ( 
.A(n_1580),
.B(n_1598),
.Y(n_2074)
);

NAND2xp33_ASAP7_75t_L g2075 ( 
.A(n_1822),
.B(n_1824),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1833),
.B(n_1839),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1843),
.B(n_1848),
.Y(n_2077)
);

AOI22xp5_ASAP7_75t_L g2078 ( 
.A1(n_1929),
.A2(n_1935),
.B1(n_1943),
.B2(n_1936),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_SL g2079 ( 
.A(n_1686),
.B(n_1787),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1849),
.B(n_1855),
.Y(n_2080)
);

INVx3_ASAP7_75t_L g2081 ( 
.A(n_1272),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_1672),
.B(n_1697),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_1771),
.B(n_1870),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_1962),
.B(n_1973),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1860),
.B(n_1863),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1867),
.B(n_1874),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1383),
.Y(n_2087)
);

AOI22xp5_ASAP7_75t_L g2088 ( 
.A1(n_1974),
.A2(n_1282),
.B1(n_1790),
.B2(n_1840),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1880),
.B(n_1884),
.Y(n_2089)
);

NAND2x1_ASAP7_75t_L g2090 ( 
.A(n_1837),
.B(n_1461),
.Y(n_2090)
);

NOR2xp33_ASAP7_75t_L g2091 ( 
.A(n_1278),
.B(n_1279),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1390),
.Y(n_2092)
);

NAND2xp33_ASAP7_75t_L g2093 ( 
.A(n_1888),
.B(n_1894),
.Y(n_2093)
);

INVx2_ASAP7_75t_SL g2094 ( 
.A(n_1294),
.Y(n_2094)
);

NOR2xp33_ASAP7_75t_L g2095 ( 
.A(n_1281),
.B(n_1862),
.Y(n_2095)
);

NOR2xp33_ASAP7_75t_L g2096 ( 
.A(n_1916),
.B(n_1945),
.Y(n_2096)
);

INVx2_ASAP7_75t_SL g2097 ( 
.A(n_1736),
.Y(n_2097)
);

INVx5_ASAP7_75t_L g2098 ( 
.A(n_1837),
.Y(n_2098)
);

NAND2xp33_ASAP7_75t_L g2099 ( 
.A(n_1895),
.B(n_1899),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1396),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_SL g2101 ( 
.A(n_1653),
.B(n_1674),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1900),
.B(n_1901),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1411),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_1906),
.B(n_1914),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1917),
.B(n_1932),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1938),
.B(n_1939),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_1347),
.B(n_1308),
.Y(n_2107)
);

CKINVDCx5p33_ASAP7_75t_R g2108 ( 
.A(n_1363),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_1415),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_1944),
.B(n_1948),
.Y(n_2110)
);

AND3x1_ASAP7_75t_L g2111 ( 
.A(n_1359),
.B(n_1357),
.C(n_1368),
.Y(n_2111)
);

AOI22xp5_ASAP7_75t_L g2112 ( 
.A1(n_1338),
.A2(n_1966),
.B1(n_1968),
.B2(n_1956),
.Y(n_2112)
);

BUFx3_ASAP7_75t_L g2113 ( 
.A(n_1736),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1425),
.Y(n_2114)
);

INVx2_ASAP7_75t_SL g2115 ( 
.A(n_1287),
.Y(n_2115)
);

NOR3xp33_ASAP7_75t_L g2116 ( 
.A(n_1676),
.B(n_1695),
.C(n_1682),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_1972),
.B(n_1984),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1432),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_1985),
.B(n_1283),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_SL g2120 ( 
.A(n_1312),
.B(n_1291),
.Y(n_2120)
);

AOI22xp33_ASAP7_75t_L g2121 ( 
.A1(n_1706),
.A2(n_1713),
.B1(n_1730),
.B2(n_1708),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_1285),
.B(n_1288),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1300),
.B(n_1303),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1304),
.B(n_1305),
.Y(n_2124)
);

BUFx6f_ASAP7_75t_SL g2125 ( 
.A(n_1452),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1309),
.B(n_1328),
.Y(n_2126)
);

AOI22xp33_ASAP7_75t_L g2127 ( 
.A1(n_1756),
.A2(n_1809),
.B1(n_1823),
.B2(n_1778),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1330),
.B(n_1341),
.Y(n_2128)
);

NAND2x1p5_ASAP7_75t_L g2129 ( 
.A(n_1374),
.B(n_1380),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1438),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1439),
.Y(n_2131)
);

NAND2xp33_ASAP7_75t_L g2132 ( 
.A(n_1324),
.B(n_1327),
.Y(n_2132)
);

INVx2_ASAP7_75t_SL g2133 ( 
.A(n_1642),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1444),
.Y(n_2134)
);

NOR2xp33_ASAP7_75t_L g2135 ( 
.A(n_1832),
.B(n_1836),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1456),
.Y(n_2136)
);

INVx2_ASAP7_75t_SL g2137 ( 
.A(n_1668),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_1842),
.B(n_1844),
.Y(n_2138)
);

AOI22xp33_ASAP7_75t_SL g2139 ( 
.A1(n_1663),
.A2(n_1835),
.B1(n_1947),
.B2(n_1342),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_1845),
.B(n_1852),
.Y(n_2140)
);

AND2x4_ASAP7_75t_L g2141 ( 
.A(n_1274),
.B(n_1591),
.Y(n_2141)
);

INVx2_ASAP7_75t_SL g2142 ( 
.A(n_1763),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_1364),
.B(n_1322),
.Y(n_2143)
);

OR2x2_ASAP7_75t_L g2144 ( 
.A(n_1618),
.B(n_1819),
.Y(n_2144)
);

OAI22xp5_ASAP7_75t_L g2145 ( 
.A1(n_1869),
.A2(n_1890),
.B1(n_1892),
.B2(n_1878),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_1905),
.B(n_1920),
.Y(n_2146)
);

BUFx2_ASAP7_75t_L g2147 ( 
.A(n_1460),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1924),
.B(n_1925),
.Y(n_2148)
);

AND2x4_ASAP7_75t_L g2149 ( 
.A(n_1634),
.B(n_1825),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1575),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1926),
.B(n_1942),
.Y(n_2151)
);

INVxp67_ASAP7_75t_SL g2152 ( 
.A(n_1590),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1946),
.B(n_1949),
.Y(n_2153)
);

INVx8_ASAP7_75t_L g2154 ( 
.A(n_1290),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_SL g2155 ( 
.A(n_1950),
.B(n_1955),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1960),
.B(n_1961),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_1607),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1610),
.Y(n_2158)
);

INVx4_ASAP7_75t_L g2159 ( 
.A(n_1907),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_1977),
.B(n_1981),
.Y(n_2160)
);

AOI22xp5_ASAP7_75t_L g2161 ( 
.A1(n_1296),
.A2(n_1896),
.B1(n_1360),
.B2(n_1313),
.Y(n_2161)
);

INVx2_ASAP7_75t_SL g2162 ( 
.A(n_1775),
.Y(n_2162)
);

BUFx3_ASAP7_75t_L g2163 ( 
.A(n_1325),
.Y(n_2163)
);

NOR2xp33_ASAP7_75t_L g2164 ( 
.A(n_1306),
.B(n_1331),
.Y(n_2164)
);

INVx2_ASAP7_75t_SL g2165 ( 
.A(n_1381),
.Y(n_2165)
);

AOI22xp33_ASAP7_75t_L g2166 ( 
.A1(n_1355),
.A2(n_1345),
.B1(n_1414),
.B2(n_1329),
.Y(n_2166)
);

AOI21xp5_ASAP7_75t_L g2167 ( 
.A1(n_1466),
.A2(n_1339),
.B(n_1519),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_SL g2168 ( 
.A(n_1403),
.B(n_1474),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_SL g2169 ( 
.A(n_1526),
.B(n_1372),
.Y(n_2169)
);

NOR2xp33_ASAP7_75t_L g2170 ( 
.A(n_1655),
.B(n_1738),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1614),
.Y(n_2171)
);

NOR2xp33_ASAP7_75t_R g2172 ( 
.A(n_1497),
.B(n_1941),
.Y(n_2172)
);

AND2x6_ASAP7_75t_SL g2173 ( 
.A(n_1541),
.B(n_1470),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1623),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_1625),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_1491),
.B(n_1493),
.Y(n_2176)
);

BUFx8_ASAP7_75t_L g2177 ( 
.A(n_1385),
.Y(n_2177)
);

NOR2xp33_ASAP7_75t_L g2178 ( 
.A(n_1826),
.B(n_1915),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_1971),
.B(n_1879),
.Y(n_2179)
);

BUFx6f_ASAP7_75t_SL g2180 ( 
.A(n_1562),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_1631),
.Y(n_2181)
);

BUFx3_ASAP7_75t_L g2182 ( 
.A(n_1382),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_1494),
.B(n_1503),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_1518),
.B(n_1515),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_SL g2185 ( 
.A(n_1272),
.B(n_1369),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_1465),
.B(n_1362),
.Y(n_2186)
);

OAI22xp5_ASAP7_75t_L g2187 ( 
.A1(n_1366),
.A2(n_1389),
.B1(n_1391),
.B2(n_1387),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_SL g2188 ( 
.A(n_1272),
.B(n_1369),
.Y(n_2188)
);

AOI22xp5_ASAP7_75t_L g2189 ( 
.A1(n_1370),
.A2(n_1427),
.B1(n_1806),
.B2(n_1759),
.Y(n_2189)
);

NAND2x1p5_ASAP7_75t_L g2190 ( 
.A(n_1637),
.B(n_1648),
.Y(n_2190)
);

NAND3xp33_ASAP7_75t_L g2191 ( 
.A(n_1568),
.B(n_1569),
.C(n_1626),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_SL g2192 ( 
.A(n_1272),
.B(n_1369),
.Y(n_2192)
);

AOI22xp33_ASAP7_75t_L g2193 ( 
.A1(n_1468),
.A2(n_1471),
.B1(n_1478),
.B2(n_1656),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_SL g2194 ( 
.A(n_1369),
.B(n_1578),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_SL g2195 ( 
.A(n_1578),
.B(n_1595),
.Y(n_2195)
);

AND2x4_ASAP7_75t_L g2196 ( 
.A(n_1542),
.B(n_1546),
.Y(n_2196)
);

BUFx3_ASAP7_75t_L g2197 ( 
.A(n_1420),
.Y(n_2197)
);

INVx8_ASAP7_75t_L g2198 ( 
.A(n_1584),
.Y(n_2198)
);

AOI22xp33_ASAP7_75t_L g2199 ( 
.A1(n_1665),
.A2(n_1677),
.B1(n_1678),
.B2(n_1671),
.Y(n_2199)
);

OAI22xp5_ASAP7_75t_L g2200 ( 
.A1(n_1393),
.A2(n_1397),
.B1(n_1399),
.B2(n_1394),
.Y(n_2200)
);

INVxp67_ASAP7_75t_L g2201 ( 
.A(n_1484),
.Y(n_2201)
);

NOR2xp33_ASAP7_75t_L g2202 ( 
.A(n_1430),
.B(n_1727),
.Y(n_2202)
);

OAI22xp33_ASAP7_75t_L g2203 ( 
.A1(n_1400),
.A2(n_1407),
.B1(n_1416),
.B2(n_1402),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_1423),
.B(n_1424),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_1431),
.B(n_1440),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_1443),
.B(n_1446),
.Y(n_2206)
);

INVxp67_ASAP7_75t_L g2207 ( 
.A(n_1467),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_1451),
.B(n_1683),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_1696),
.B(n_1699),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_SL g2210 ( 
.A(n_1578),
.B(n_1595),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_1710),
.Y(n_2211)
);

NOR2xp33_ASAP7_75t_L g2212 ( 
.A(n_1749),
.B(n_1828),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_1714),
.B(n_1718),
.Y(n_2213)
);

AOI22xp33_ASAP7_75t_L g2214 ( 
.A1(n_1721),
.A2(n_1732),
.B1(n_1747),
.B2(n_1726),
.Y(n_2214)
);

INVx1_ASAP7_75t_SL g2215 ( 
.A(n_1445),
.Y(n_2215)
);

NOR2xp33_ASAP7_75t_L g2216 ( 
.A(n_1882),
.B(n_1885),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_1525),
.B(n_1532),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_1773),
.Y(n_2218)
);

NOR2xp33_ASAP7_75t_SL g2219 ( 
.A(n_1604),
.B(n_1404),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_1791),
.B(n_1796),
.Y(n_2220)
);

AOI21xp5_ASAP7_75t_L g2221 ( 
.A1(n_1433),
.A2(n_1475),
.B(n_1418),
.Y(n_2221)
);

O2A1O1Ixp5_ASAP7_75t_L g2222 ( 
.A1(n_1903),
.A2(n_1565),
.B(n_1522),
.C(n_1408),
.Y(n_2222)
);

AND2x6_ASAP7_75t_SL g2223 ( 
.A(n_1472),
.B(n_1557),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_1798),
.B(n_1805),
.Y(n_2224)
);

NOR3xp33_ASAP7_75t_L g2225 ( 
.A(n_1437),
.B(n_1495),
.C(n_1951),
.Y(n_2225)
);

BUFx6f_ASAP7_75t_L g2226 ( 
.A(n_1579),
.Y(n_2226)
);

AOI21xp5_ASAP7_75t_L g2227 ( 
.A1(n_1406),
.A2(n_1429),
.B(n_1426),
.Y(n_2227)
);

A2O1A1Ixp33_ASAP7_75t_L g2228 ( 
.A1(n_1450),
.A2(n_1523),
.B(n_1520),
.C(n_1513),
.Y(n_2228)
);

BUFx2_ASAP7_75t_L g2229 ( 
.A(n_1964),
.Y(n_2229)
);

A2O1A1Ixp33_ASAP7_75t_SL g2230 ( 
.A1(n_1448),
.A2(n_1454),
.B(n_1548),
.C(n_1502),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_1808),
.B(n_1812),
.Y(n_2231)
);

OA22x2_ASAP7_75t_L g2232 ( 
.A1(n_1540),
.A2(n_1545),
.B1(n_1549),
.B2(n_1543),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1817),
.Y(n_2233)
);

INVx4_ASAP7_75t_L g2234 ( 
.A(n_1907),
.Y(n_2234)
);

NOR2xp33_ASAP7_75t_L g2235 ( 
.A(n_1976),
.B(n_1979),
.Y(n_2235)
);

A2O1A1Ixp33_ASAP7_75t_SL g2236 ( 
.A1(n_1496),
.A2(n_1509),
.B(n_1512),
.C(n_1499),
.Y(n_2236)
);

AOI22xp5_ASAP7_75t_L g2237 ( 
.A1(n_1846),
.A2(n_1521),
.B1(n_1500),
.B2(n_1386),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_SL g2238 ( 
.A(n_1524),
.B(n_1485),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_SL g2239 ( 
.A(n_1485),
.B(n_1501),
.Y(n_2239)
);

AND2x4_ASAP7_75t_L g2240 ( 
.A(n_1477),
.B(n_1527),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_1827),
.B(n_1831),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_SL g2242 ( 
.A(n_1501),
.B(n_1292),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_1841),
.B(n_1850),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_1851),
.Y(n_2244)
);

AND2x4_ASAP7_75t_L g2245 ( 
.A(n_1273),
.B(n_1286),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_SL g2246 ( 
.A(n_1720),
.B(n_1786),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_1891),
.B(n_1898),
.Y(n_2247)
);

BUFx6f_ASAP7_75t_L g2248 ( 
.A(n_1579),
.Y(n_2248)
);

AOI22xp5_ASAP7_75t_L g2249 ( 
.A1(n_1379),
.A2(n_1409),
.B1(n_1490),
.B2(n_1388),
.Y(n_2249)
);

NAND2xp33_ASAP7_75t_SL g2250 ( 
.A(n_1413),
.B(n_1492),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_1289),
.B(n_1302),
.Y(n_2251)
);

INVx3_ASAP7_75t_L g2252 ( 
.A(n_1578),
.Y(n_2252)
);

INVx2_ASAP7_75t_SL g2253 ( 
.A(n_1603),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_1908),
.Y(n_2254)
);

INVx2_ASAP7_75t_L g2255 ( 
.A(n_1910),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1913),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_1918),
.B(n_1923),
.Y(n_2257)
);

NOR2xp33_ASAP7_75t_L g2258 ( 
.A(n_1556),
.B(n_1564),
.Y(n_2258)
);

AOI22xp33_ASAP7_75t_L g2259 ( 
.A1(n_1940),
.A2(n_1959),
.B1(n_1965),
.B2(n_1957),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_1983),
.B(n_1986),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_1457),
.B(n_1316),
.Y(n_2261)
);

NOR2xp33_ASAP7_75t_L g2262 ( 
.A(n_1398),
.B(n_1441),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_1319),
.B(n_1320),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_SL g2264 ( 
.A(n_1595),
.B(n_1615),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1326),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_SL g2266 ( 
.A(n_1595),
.B(n_1615),
.Y(n_2266)
);

AOI21xp5_ASAP7_75t_L g2267 ( 
.A1(n_1449),
.A2(n_1458),
.B(n_1453),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1479),
.Y(n_2268)
);

NOR2xp33_ASAP7_75t_L g2269 ( 
.A(n_1463),
.B(n_1334),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1504),
.Y(n_2270)
);

BUFx3_ASAP7_75t_L g2271 ( 
.A(n_1603),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_1337),
.B(n_1350),
.Y(n_2272)
);

AND2x4_ASAP7_75t_L g2273 ( 
.A(n_1361),
.B(n_1376),
.Y(n_2273)
);

NOR2xp33_ASAP7_75t_L g2274 ( 
.A(n_1392),
.B(n_1405),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_SL g2275 ( 
.A(n_1615),
.B(n_1769),
.Y(n_2275)
);

NOR2xp33_ASAP7_75t_L g2276 ( 
.A(n_1417),
.B(n_1421),
.Y(n_2276)
);

AOI22xp33_ASAP7_75t_SL g2277 ( 
.A1(n_1567),
.A2(n_1529),
.B1(n_1561),
.B2(n_1384),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_1422),
.B(n_1435),
.Y(n_2278)
);

AOI22xp5_ASAP7_75t_L g2279 ( 
.A1(n_1514),
.A2(n_1550),
.B1(n_1539),
.B2(n_1516),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_SL g2280 ( 
.A(n_1615),
.B(n_1769),
.Y(n_2280)
);

AND2x6_ASAP7_75t_SL g2281 ( 
.A(n_1434),
.B(n_1436),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_SL g2282 ( 
.A(n_1769),
.B(n_1510),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_1442),
.B(n_1447),
.Y(n_2283)
);

OAI22xp5_ASAP7_75t_L g2284 ( 
.A1(n_1455),
.A2(n_1982),
.B1(n_1571),
.B2(n_1573),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1462),
.Y(n_2285)
);

BUFx3_ASAP7_75t_L g2286 ( 
.A(n_1606),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_1464),
.B(n_1576),
.Y(n_2287)
);

AOI22xp33_ASAP7_75t_SL g2288 ( 
.A1(n_1508),
.A2(n_1498),
.B1(n_1533),
.B2(n_1536),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_1577),
.B(n_1583),
.Y(n_2289)
);

AOI22xp33_ASAP7_75t_L g2290 ( 
.A1(n_1593),
.A2(n_1694),
.B1(n_1963),
.B2(n_1958),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_1594),
.B(n_1608),
.Y(n_2291)
);

AOI22xp5_ASAP7_75t_L g2292 ( 
.A1(n_1528),
.A2(n_1535),
.B1(n_1459),
.B2(n_1818),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_1612),
.B(n_1613),
.Y(n_2293)
);

OAI22xp33_ASAP7_75t_L g2294 ( 
.A1(n_1622),
.A2(n_1821),
.B1(n_1740),
.B2(n_1722),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_1640),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_1643),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_1647),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_1657),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_1661),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_1664),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_1670),
.B(n_1673),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_1679),
.B(n_1681),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_SL g2303 ( 
.A(n_1769),
.B(n_1684),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_1688),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_1690),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_1731),
.Y(n_2306)
);

BUFx3_ASAP7_75t_L g2307 ( 
.A(n_1606),
.Y(n_2307)
);

CKINVDCx5p33_ASAP7_75t_R g2308 ( 
.A(n_1530),
.Y(n_2308)
);

AOI22xp5_ASAP7_75t_L g2309 ( 
.A1(n_1742),
.A2(n_1847),
.B1(n_1838),
.B2(n_1820),
.Y(n_2309)
);

BUFx6f_ASAP7_75t_L g2310 ( 
.A(n_1628),
.Y(n_2310)
);

O2A1O1Ixp5_ASAP7_75t_L g2311 ( 
.A1(n_1488),
.A2(n_1865),
.B(n_1897),
.C(n_1875),
.Y(n_2311)
);

AND2x6_ASAP7_75t_SL g2312 ( 
.A(n_1559),
.B(n_1558),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_SL g2313 ( 
.A(n_1754),
.B(n_1757),
.Y(n_2313)
);

OAI22xp5_ASAP7_75t_L g2314 ( 
.A1(n_1760),
.A2(n_1904),
.B1(n_1764),
.B2(n_1766),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_1768),
.B(n_1772),
.Y(n_2315)
);

AOI22xp33_ASAP7_75t_L g2316 ( 
.A1(n_1803),
.A2(n_1877),
.B1(n_1952),
.B2(n_1937),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_1810),
.Y(n_2317)
);

NOR2xp33_ASAP7_75t_L g2318 ( 
.A(n_1876),
.B(n_1886),
.Y(n_2318)
);

NOR2xp33_ASAP7_75t_L g2319 ( 
.A(n_1933),
.B(n_1934),
.Y(n_2319)
);

AO22x1_ASAP7_75t_L g2320 ( 
.A1(n_1505),
.A2(n_1675),
.B1(n_1748),
.B2(n_1725),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_1469),
.B(n_1483),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_1487),
.B(n_1481),
.Y(n_2322)
);

INVx2_ASAP7_75t_SL g2323 ( 
.A(n_1628),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_SL g2324 ( 
.A(n_1412),
.B(n_1794),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_1534),
.Y(n_2325)
);

AOI22xp5_ASAP7_75t_L g2326 ( 
.A1(n_1507),
.A2(n_1553),
.B1(n_1978),
.B2(n_1980),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_1537),
.Y(n_2327)
);

CKINVDCx5p33_ASAP7_75t_R g2328 ( 
.A(n_1570),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_1547),
.Y(n_2329)
);

NOR2xp33_ASAP7_75t_L g2330 ( 
.A(n_1371),
.B(n_1401),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_1752),
.B(n_1703),
.Y(n_2331)
);

AOI22xp5_ASAP7_75t_L g2332 ( 
.A1(n_1864),
.A2(n_1953),
.B1(n_1921),
.B2(n_1912),
.Y(n_2332)
);

OR2x6_ASAP7_75t_L g2333 ( 
.A(n_1511),
.B(n_1476),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_1551),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_1752),
.B(n_1680),
.Y(n_2335)
);

NOR2xp33_ASAP7_75t_L g2336 ( 
.A(n_1482),
.B(n_1480),
.Y(n_2336)
);

AOI22xp33_ASAP7_75t_L g2337 ( 
.A1(n_1560),
.A2(n_1930),
.B1(n_1654),
.B2(n_1692),
.Y(n_2337)
);

CKINVDCx5p33_ASAP7_75t_R g2338 ( 
.A(n_1323),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_1552),
.B(n_1428),
.Y(n_2339)
);

AND2x2_ASAP7_75t_L g2340 ( 
.A(n_1554),
.B(n_1555),
.Y(n_2340)
);

NAND2x1p5_ASAP7_75t_L g2341 ( 
.A(n_1531),
.B(n_1544),
.Y(n_2341)
);

NOR2xp33_ASAP7_75t_L g2342 ( 
.A(n_1645),
.B(n_1793),
.Y(n_2342)
);

NOR2x1p5_ASAP7_75t_L g2343 ( 
.A(n_1562),
.B(n_1566),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_1410),
.B(n_1419),
.Y(n_2344)
);

NAND3xp33_ASAP7_75t_L g2345 ( 
.A(n_1566),
.B(n_1975),
.C(n_1795),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_SL g2346 ( 
.A(n_1645),
.B(n_1801),
.Y(n_2346)
);

AND2x4_ASAP7_75t_L g2347 ( 
.A(n_1473),
.B(n_1336),
.Y(n_2347)
);

INVx4_ASAP7_75t_L g2348 ( 
.A(n_1705),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_1705),
.B(n_1811),
.Y(n_2349)
);

AOI22xp5_ASAP7_75t_L g2350 ( 
.A1(n_1830),
.A2(n_1723),
.B1(n_1635),
.B2(n_1658),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_1735),
.Y(n_2351)
);

AND2x4_ASAP7_75t_L g2352 ( 
.A(n_1367),
.B(n_1716),
.Y(n_2352)
);

NAND3xp33_ASAP7_75t_SL g2353 ( 
.A(n_1815),
.B(n_1859),
.C(n_1887),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_1735),
.B(n_1744),
.Y(n_2354)
);

NOR2xp33_ASAP7_75t_L g2355 ( 
.A(n_1744),
.B(n_1784),
.Y(n_2355)
);

AOI22xp33_ASAP7_75t_L g2356 ( 
.A1(n_1784),
.A2(n_1785),
.B1(n_1793),
.B2(n_1801),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_1785),
.B(n_1811),
.Y(n_2357)
);

AOI22xp33_ASAP7_75t_L g2358 ( 
.A1(n_1868),
.A2(n_1872),
.B1(n_1889),
.B2(n_1893),
.Y(n_2358)
);

A2O1A1Ixp33_ASAP7_75t_L g2359 ( 
.A1(n_1829),
.A2(n_1873),
.B(n_1872),
.C(n_1868),
.Y(n_2359)
);

A2O1A1Ixp33_ASAP7_75t_L g2360 ( 
.A1(n_1889),
.A2(n_1893),
.B(n_1919),
.C(n_1067),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_1919),
.B(n_1067),
.Y(n_2361)
);

NOR2xp33_ASAP7_75t_L g2362 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_SL g2363 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_1277),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2366)
);

AOI22xp33_ASAP7_75t_L g2367 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2367)
);

INVxp67_ASAP7_75t_L g2368 ( 
.A(n_1349),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2370)
);

BUFx6f_ASAP7_75t_L g2371 ( 
.A(n_1381),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_SL g2372 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2372)
);

NOR2xp33_ASAP7_75t_L g2373 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2373)
);

OAI21xp5_ASAP7_75t_L g2374 ( 
.A1(n_1804),
.A2(n_788),
.B(n_673),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_1277),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_1277),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_SL g2378 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_SL g2380 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2382)
);

A2O1A1Ixp33_ASAP7_75t_L g2383 ( 
.A1(n_1804),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_1277),
.Y(n_2385)
);

A2O1A1Ixp33_ASAP7_75t_L g2386 ( 
.A1(n_1804),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_2386)
);

NOR2xp33_ASAP7_75t_L g2387 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_1277),
.Y(n_2388)
);

NOR2xp33_ASAP7_75t_L g2389 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2389)
);

AOI22xp5_ASAP7_75t_L g2390 ( 
.A1(n_1280),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2390)
);

OR2x2_ASAP7_75t_L g2391 ( 
.A(n_1285),
.B(n_846),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2392)
);

O2A1O1Ixp5_ASAP7_75t_L g2393 ( 
.A1(n_1804),
.A2(n_788),
.B(n_807),
.C(n_673),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2395)
);

AND2x2_ASAP7_75t_L g2396 ( 
.A(n_1275),
.B(n_839),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_SL g2397 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2397)
);

NOR2xp33_ASAP7_75t_L g2398 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_SL g2400 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_1277),
.Y(n_2401)
);

NOR2xp33_ASAP7_75t_L g2402 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2402)
);

INVx2_ASAP7_75t_SL g2403 ( 
.A(n_1294),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_SL g2404 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2405)
);

INVx2_ASAP7_75t_L g2406 ( 
.A(n_1277),
.Y(n_2406)
);

O2A1O1Ixp33_ASAP7_75t_L g2407 ( 
.A1(n_1804),
.A2(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_2407)
);

INVx2_ASAP7_75t_SL g2408 ( 
.A(n_1294),
.Y(n_2408)
);

BUFx8_ASAP7_75t_L g2409 ( 
.A(n_1385),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2410)
);

BUFx2_ASAP7_75t_L g2411 ( 
.A(n_1967),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_1277),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_1277),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2415)
);

NOR3xp33_ASAP7_75t_L g2416 ( 
.A(n_1804),
.B(n_1072),
.C(n_1067),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2417)
);

AND2x6_ASAP7_75t_SL g2418 ( 
.A(n_1489),
.B(n_1541),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_SL g2419 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2419)
);

NOR2xp33_ASAP7_75t_L g2420 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2420)
);

AOI22xp33_ASAP7_75t_L g2421 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2421)
);

BUFx6f_ASAP7_75t_L g2422 ( 
.A(n_1381),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2423)
);

O2A1O1Ixp5_ASAP7_75t_L g2424 ( 
.A1(n_1804),
.A2(n_788),
.B(n_807),
.C(n_673),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_1277),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_SL g2427 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_SL g2428 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2428)
);

NOR2xp33_ASAP7_75t_L g2429 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2429)
);

NOR3xp33_ASAP7_75t_L g2430 ( 
.A(n_1804),
.B(n_1072),
.C(n_1067),
.Y(n_2430)
);

NOR2xp33_ASAP7_75t_L g2431 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_1277),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2435)
);

AND2x2_ASAP7_75t_L g2436 ( 
.A(n_1275),
.B(n_839),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_1277),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_SL g2439 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_1277),
.Y(n_2440)
);

INVx4_ASAP7_75t_L g2441 ( 
.A(n_1294),
.Y(n_2441)
);

BUFx3_ASAP7_75t_L g2442 ( 
.A(n_1294),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_1277),
.Y(n_2444)
);

CKINVDCx5p33_ASAP7_75t_R g2445 ( 
.A(n_1538),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_1277),
.Y(n_2447)
);

CKINVDCx5p33_ASAP7_75t_R g2448 ( 
.A(n_1538),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_1277),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_1277),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_SL g2451 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2451)
);

NOR2xp67_ASAP7_75t_L g2452 ( 
.A(n_1349),
.B(n_853),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2454)
);

NOR2xp33_ASAP7_75t_L g2455 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_1277),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2458)
);

AND2x2_ASAP7_75t_L g2459 ( 
.A(n_1275),
.B(n_839),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_1277),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_1277),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_L g2463 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2464)
);

AND2x6_ASAP7_75t_SL g2465 ( 
.A(n_1489),
.B(n_1541),
.Y(n_2465)
);

AOI22xp33_ASAP7_75t_L g2466 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2466)
);

AOI22xp33_ASAP7_75t_L g2467 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2467)
);

NOR2xp33_ASAP7_75t_L g2468 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_L g2470 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2470)
);

NOR2xp33_ASAP7_75t_L g2471 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_1277),
.Y(n_2472)
);

INVx2_ASAP7_75t_L g2473 ( 
.A(n_1277),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_L g2474 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_L g2475 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_1277),
.Y(n_2476)
);

NOR2xp33_ASAP7_75t_L g2477 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2478)
);

NOR2xp33_ASAP7_75t_L g2479 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2479)
);

CKINVDCx16_ASAP7_75t_R g2480 ( 
.A(n_1538),
.Y(n_2480)
);

INVxp67_ASAP7_75t_L g2481 ( 
.A(n_1349),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2482)
);

NOR2xp33_ASAP7_75t_L g2483 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2483)
);

AOI22xp5_ASAP7_75t_L g2484 ( 
.A1(n_1280),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2484)
);

INVx2_ASAP7_75t_SL g2485 ( 
.A(n_1294),
.Y(n_2485)
);

AOI22xp33_ASAP7_75t_L g2486 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2486)
);

O2A1O1Ixp33_ASAP7_75t_L g2487 ( 
.A1(n_1804),
.A2(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_1277),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2489)
);

NAND2xp33_ASAP7_75t_L g2490 ( 
.A(n_1804),
.B(n_1066),
.Y(n_2490)
);

AND2x2_ASAP7_75t_L g2491 ( 
.A(n_1275),
.B(n_839),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_1277),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_1277),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2496)
);

AND2x6_ASAP7_75t_SL g2497 ( 
.A(n_1489),
.B(n_1541),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_1277),
.Y(n_2498)
);

AND2x2_ASAP7_75t_L g2499 ( 
.A(n_1275),
.B(n_839),
.Y(n_2499)
);

INVx2_ASAP7_75t_SL g2500 ( 
.A(n_1294),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2501)
);

INVx2_ASAP7_75t_SL g2502 ( 
.A(n_1294),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_L g2503 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2503)
);

AND2x2_ASAP7_75t_L g2504 ( 
.A(n_1275),
.B(n_839),
.Y(n_2504)
);

AOI22xp33_ASAP7_75t_L g2505 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2505)
);

OR2x6_ASAP7_75t_L g2506 ( 
.A(n_1294),
.B(n_1736),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_SL g2510 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_1277),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2512)
);

BUFx6f_ASAP7_75t_L g2513 ( 
.A(n_1381),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_SL g2514 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2514)
);

INVx2_ASAP7_75t_L g2515 ( 
.A(n_1277),
.Y(n_2515)
);

AO22x1_ASAP7_75t_L g2516 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2516)
);

INVx2_ASAP7_75t_L g2517 ( 
.A(n_1277),
.Y(n_2517)
);

CKINVDCx5p33_ASAP7_75t_R g2518 ( 
.A(n_1538),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_1277),
.Y(n_2519)
);

AND2x2_ASAP7_75t_L g2520 ( 
.A(n_1275),
.B(n_839),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_1277),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_1277),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2525)
);

NAND3xp33_ASAP7_75t_L g2526 ( 
.A(n_1804),
.B(n_1072),
.C(n_1067),
.Y(n_2526)
);

AND2x2_ASAP7_75t_L g2527 ( 
.A(n_1275),
.B(n_839),
.Y(n_2527)
);

AND2x6_ASAP7_75t_SL g2528 ( 
.A(n_1489),
.B(n_1541),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_1277),
.Y(n_2529)
);

AND2x6_ASAP7_75t_SL g2530 ( 
.A(n_1489),
.B(n_1541),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2531)
);

AND2x2_ASAP7_75t_L g2532 ( 
.A(n_1275),
.B(n_839),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_1277),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_SL g2535 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2537)
);

A2O1A1Ixp33_ASAP7_75t_L g2538 ( 
.A1(n_1804),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_2538)
);

OAI22xp33_ASAP7_75t_L g2539 ( 
.A1(n_1804),
.A2(n_1089),
.B1(n_1198),
.B2(n_1081),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_1277),
.Y(n_2540)
);

AOI22xp5_ASAP7_75t_L g2541 ( 
.A1(n_1280),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2541)
);

NOR2xp33_ASAP7_75t_L g2542 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_SL g2543 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2543)
);

OR2x6_ASAP7_75t_L g2544 ( 
.A(n_1294),
.B(n_1736),
.Y(n_2544)
);

A2O1A1Ixp33_ASAP7_75t_L g2545 ( 
.A1(n_1804),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_SL g2546 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_1277),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_SL g2548 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2548)
);

AND2x2_ASAP7_75t_SL g2549 ( 
.A(n_1311),
.B(n_1067),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_SL g2550 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2551)
);

AND2x2_ASAP7_75t_L g2552 ( 
.A(n_1275),
.B(n_839),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_SL g2554 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2554)
);

AND2x6_ASAP7_75t_SL g2555 ( 
.A(n_1489),
.B(n_1541),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2556)
);

OR2x6_ASAP7_75t_L g2557 ( 
.A(n_1294),
.B(n_1736),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_1277),
.Y(n_2558)
);

AND2x6_ASAP7_75t_SL g2559 ( 
.A(n_1489),
.B(n_1541),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_1277),
.Y(n_2560)
);

AOI22xp33_ASAP7_75t_L g2561 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2561)
);

BUFx6f_ASAP7_75t_L g2562 ( 
.A(n_1381),
.Y(n_2562)
);

CKINVDCx5p33_ASAP7_75t_R g2563 ( 
.A(n_1538),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_1275),
.B(n_839),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2565)
);

AND2x6_ASAP7_75t_L g2566 ( 
.A(n_1339),
.B(n_934),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2567)
);

AOI21xp5_ASAP7_75t_L g2568 ( 
.A1(n_1804),
.A2(n_907),
.B(n_653),
.Y(n_2568)
);

OAI21xp5_ASAP7_75t_L g2569 ( 
.A1(n_1804),
.A2(n_788),
.B(n_673),
.Y(n_2569)
);

AOI22xp33_ASAP7_75t_L g2570 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2570)
);

AOI22xp5_ASAP7_75t_L g2571 ( 
.A1(n_1280),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_1277),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_1277),
.Y(n_2573)
);

INVx2_ASAP7_75t_SL g2574 ( 
.A(n_1294),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_L g2575 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2575)
);

NOR3xp33_ASAP7_75t_L g2576 ( 
.A(n_1804),
.B(n_1072),
.C(n_1067),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_SL g2577 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_SL g2578 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_L g2579 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2579)
);

AOI22xp33_ASAP7_75t_L g2580 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_1277),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2582)
);

NAND2x1_ASAP7_75t_L g2583 ( 
.A(n_1506),
.B(n_1837),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2584)
);

NOR2xp67_ASAP7_75t_L g2585 ( 
.A(n_1349),
.B(n_853),
.Y(n_2585)
);

AOI21xp5_ASAP7_75t_L g2586 ( 
.A1(n_1804),
.A2(n_907),
.B(n_653),
.Y(n_2586)
);

INVx2_ASAP7_75t_L g2587 ( 
.A(n_1277),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_SL g2588 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2588)
);

AOI22xp5_ASAP7_75t_L g2589 ( 
.A1(n_1280),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_SL g2590 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_SL g2591 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2591)
);

INVx2_ASAP7_75t_L g2592 ( 
.A(n_1277),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_1277),
.Y(n_2593)
);

NAND2xp33_ASAP7_75t_L g2594 ( 
.A(n_1804),
.B(n_1066),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_1277),
.Y(n_2595)
);

AOI22xp33_ASAP7_75t_L g2596 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2596)
);

NOR2xp33_ASAP7_75t_L g2597 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_SL g2598 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_1277),
.Y(n_2599)
);

O2A1O1Ixp33_ASAP7_75t_L g2600 ( 
.A1(n_1804),
.A2(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2601)
);

AND2x6_ASAP7_75t_SL g2602 ( 
.A(n_1489),
.B(n_1541),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2603)
);

NOR3xp33_ASAP7_75t_L g2604 ( 
.A(n_1804),
.B(n_1072),
.C(n_1067),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_L g2605 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_SL g2606 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2607)
);

NOR2xp33_ASAP7_75t_L g2608 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_1277),
.Y(n_2609)
);

NOR2xp33_ASAP7_75t_L g2610 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_L g2611 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2611)
);

AOI22xp5_ASAP7_75t_L g2612 ( 
.A1(n_1280),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2612)
);

AOI21xp5_ASAP7_75t_L g2613 ( 
.A1(n_1804),
.A2(n_907),
.B(n_653),
.Y(n_2613)
);

BUFx5_ASAP7_75t_L g2614 ( 
.A(n_1837),
.Y(n_2614)
);

OR2x2_ASAP7_75t_L g2615 ( 
.A(n_1285),
.B(n_846),
.Y(n_2615)
);

AOI22xp33_ASAP7_75t_L g2616 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_1277),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_1277),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_L g2622 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_SL g2623 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2624)
);

INVxp67_ASAP7_75t_L g2625 ( 
.A(n_1349),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_L g2626 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2626)
);

NOR2xp33_ASAP7_75t_L g2627 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2627)
);

AOI22xp33_ASAP7_75t_L g2628 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2628)
);

AOI22xp5_ASAP7_75t_L g2629 ( 
.A1(n_1280),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2629)
);

NOR2xp33_ASAP7_75t_L g2630 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2630)
);

NAND2x1p5_ASAP7_75t_L g2631 ( 
.A(n_1374),
.B(n_1009),
.Y(n_2631)
);

AND2x6_ASAP7_75t_SL g2632 ( 
.A(n_1489),
.B(n_1541),
.Y(n_2632)
);

AND2x2_ASAP7_75t_L g2633 ( 
.A(n_1275),
.B(n_839),
.Y(n_2633)
);

NOR2xp33_ASAP7_75t_L g2634 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2634)
);

CKINVDCx5p33_ASAP7_75t_R g2635 ( 
.A(n_1538),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_1277),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_L g2638 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_1277),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2641)
);

OR2x2_ASAP7_75t_L g2642 ( 
.A(n_1285),
.B(n_846),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_L g2643 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_1277),
.Y(n_2645)
);

AOI22xp5_ASAP7_75t_L g2646 ( 
.A1(n_1280),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_1277),
.Y(n_2648)
);

INVx2_ASAP7_75t_L g2649 ( 
.A(n_1277),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_1277),
.Y(n_2650)
);

NOR2xp33_ASAP7_75t_L g2651 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2651)
);

NOR2xp33_ASAP7_75t_L g2652 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2654)
);

AOI22xp33_ASAP7_75t_L g2655 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2655)
);

AND2x6_ASAP7_75t_SL g2656 ( 
.A(n_1489),
.B(n_1541),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_1277),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_SL g2659 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2659)
);

NAND2x1p5_ASAP7_75t_L g2660 ( 
.A(n_1374),
.B(n_1009),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_L g2661 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2661)
);

NOR3xp33_ASAP7_75t_L g2662 ( 
.A(n_1804),
.B(n_1072),
.C(n_1067),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_L g2665 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2665)
);

AND2x2_ASAP7_75t_L g2666 ( 
.A(n_1275),
.B(n_839),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2667)
);

BUFx6f_ASAP7_75t_L g2668 ( 
.A(n_1381),
.Y(n_2668)
);

BUFx3_ASAP7_75t_L g2669 ( 
.A(n_1294),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_1277),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_L g2671 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_1277),
.Y(n_2672)
);

BUFx3_ASAP7_75t_L g2673 ( 
.A(n_1294),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_L g2674 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_SL g2675 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_SL g2676 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2676)
);

AOI22xp33_ASAP7_75t_L g2677 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2678)
);

BUFx6f_ASAP7_75t_L g2679 ( 
.A(n_1381),
.Y(n_2679)
);

OR2x2_ASAP7_75t_L g2680 ( 
.A(n_1285),
.B(n_846),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_1277),
.Y(n_2681)
);

INVx2_ASAP7_75t_SL g2682 ( 
.A(n_1294),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_SL g2683 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_1277),
.Y(n_2685)
);

AOI22xp33_ASAP7_75t_L g2686 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2686)
);

INVx2_ASAP7_75t_L g2687 ( 
.A(n_1277),
.Y(n_2687)
);

NOR2xp67_ASAP7_75t_L g2688 ( 
.A(n_1349),
.B(n_853),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_1277),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_1277),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_1277),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_SL g2693 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2693)
);

NOR2xp33_ASAP7_75t_L g2694 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2694)
);

BUFx2_ASAP7_75t_L g2695 ( 
.A(n_1967),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_1277),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2697)
);

NOR2xp33_ASAP7_75t_L g2698 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2698)
);

AOI22xp33_ASAP7_75t_L g2699 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_1277),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_1277),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_1277),
.Y(n_2702)
);

AOI22xp33_ASAP7_75t_SL g2703 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_1277),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2705)
);

BUFx2_ASAP7_75t_L g2706 ( 
.A(n_1967),
.Y(n_2706)
);

AOI22xp33_ASAP7_75t_L g2707 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2707)
);

BUFx6f_ASAP7_75t_L g2708 ( 
.A(n_1381),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_1277),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2710)
);

AOI22xp33_ASAP7_75t_L g2711 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2711)
);

AOI21xp5_ASAP7_75t_L g2712 ( 
.A1(n_1804),
.A2(n_907),
.B(n_653),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_1277),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_SL g2714 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2714)
);

A2O1A1Ixp33_ASAP7_75t_L g2715 ( 
.A1(n_1804),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_2715)
);

AND2x2_ASAP7_75t_L g2716 ( 
.A(n_1275),
.B(n_839),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2717)
);

AOI22xp33_ASAP7_75t_L g2718 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2718)
);

INVx8_ASAP7_75t_L g2719 ( 
.A(n_1294),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_1277),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_1277),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_L g2723 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2723)
);

AND2x2_ASAP7_75t_L g2724 ( 
.A(n_1275),
.B(n_839),
.Y(n_2724)
);

BUFx4f_ASAP7_75t_L g2725 ( 
.A(n_1562),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_1277),
.Y(n_2726)
);

NOR2xp33_ASAP7_75t_L g2727 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2727)
);

AOI22xp33_ASAP7_75t_L g2728 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2728)
);

INVx2_ASAP7_75t_L g2729 ( 
.A(n_1277),
.Y(n_2729)
);

O2A1O1Ixp33_ASAP7_75t_L g2730 ( 
.A1(n_1804),
.A2(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_L g2731 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2731)
);

AND2x2_ASAP7_75t_L g2732 ( 
.A(n_1275),
.B(n_839),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_1277),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2735)
);

AND2x2_ASAP7_75t_L g2736 ( 
.A(n_1275),
.B(n_839),
.Y(n_2736)
);

OAI21xp5_ASAP7_75t_L g2737 ( 
.A1(n_1804),
.A2(n_788),
.B(n_673),
.Y(n_2737)
);

NOR2x1p5_ASAP7_75t_L g2738 ( 
.A(n_1497),
.B(n_820),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_1277),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_1277),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_1277),
.Y(n_2741)
);

NOR2xp33_ASAP7_75t_L g2742 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2742)
);

INVx5_ASAP7_75t_L g2743 ( 
.A(n_1506),
.Y(n_2743)
);

AND2x2_ASAP7_75t_L g2744 ( 
.A(n_1275),
.B(n_839),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2745)
);

NOR2xp33_ASAP7_75t_L g2746 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_1277),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_SL g2748 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2748)
);

OAI22xp5_ASAP7_75t_L g2749 ( 
.A1(n_1804),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2751)
);

AND2x2_ASAP7_75t_L g2752 ( 
.A(n_1275),
.B(n_839),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2753)
);

NOR2xp33_ASAP7_75t_L g2754 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_1277),
.Y(n_2755)
);

OR2x2_ASAP7_75t_SL g2756 ( 
.A(n_1580),
.B(n_1124),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_1277),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_SL g2759 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2759)
);

HB1xp67_ASAP7_75t_L g2760 ( 
.A(n_1780),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2762)
);

AOI22xp33_ASAP7_75t_L g2763 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2763)
);

NOR2xp33_ASAP7_75t_L g2764 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_1277),
.Y(n_2765)
);

NOR3xp33_ASAP7_75t_L g2766 ( 
.A(n_1804),
.B(n_1072),
.C(n_1067),
.Y(n_2766)
);

NAND2x1_ASAP7_75t_L g2767 ( 
.A(n_1506),
.B(n_1837),
.Y(n_2767)
);

AND2x2_ASAP7_75t_L g2768 ( 
.A(n_1275),
.B(n_839),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_1277),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_1277),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_SL g2772 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2772)
);

NOR2xp33_ASAP7_75t_L g2773 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2773)
);

INVx2_ASAP7_75t_L g2774 ( 
.A(n_1277),
.Y(n_2774)
);

O2A1O1Ixp33_ASAP7_75t_L g2775 ( 
.A1(n_1804),
.A2(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_2775)
);

AOI22xp5_ASAP7_75t_L g2776 ( 
.A1(n_1280),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_SL g2777 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2777)
);

NOR2xp33_ASAP7_75t_L g2778 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_1277),
.Y(n_2779)
);

AND2x2_ASAP7_75t_SL g2780 ( 
.A(n_1311),
.B(n_1067),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_1277),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_1277),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_1277),
.Y(n_2783)
);

OAI22xp5_ASAP7_75t_L g2784 ( 
.A1(n_1804),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_L g2785 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2785)
);

INVx2_ASAP7_75t_L g2786 ( 
.A(n_1277),
.Y(n_2786)
);

NOR2xp33_ASAP7_75t_L g2787 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2787)
);

INVx2_ASAP7_75t_L g2788 ( 
.A(n_1277),
.Y(n_2788)
);

OAI22xp5_ASAP7_75t_L g2789 ( 
.A1(n_1804),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_L g2791 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_1277),
.Y(n_2792)
);

NOR2xp33_ASAP7_75t_L g2793 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2794)
);

AND2x2_ASAP7_75t_SL g2795 ( 
.A(n_1311),
.B(n_1067),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_1277),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_SL g2797 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2797)
);

BUFx6f_ASAP7_75t_L g2798 ( 
.A(n_1381),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2799)
);

INVx8_ASAP7_75t_L g2800 ( 
.A(n_1294),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_SL g2801 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2801)
);

A2O1A1Ixp33_ASAP7_75t_L g2802 ( 
.A1(n_1804),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_2802)
);

INVx2_ASAP7_75t_L g2803 ( 
.A(n_1277),
.Y(n_2803)
);

NOR2xp33_ASAP7_75t_L g2804 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_L g2805 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2805)
);

AOI22xp33_ASAP7_75t_L g2806 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_1277),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_1277),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_1277),
.Y(n_2809)
);

AND2x2_ASAP7_75t_L g2810 ( 
.A(n_1275),
.B(n_839),
.Y(n_2810)
);

OR2x2_ASAP7_75t_L g2811 ( 
.A(n_1285),
.B(n_846),
.Y(n_2811)
);

BUFx12f_ASAP7_75t_L g2812 ( 
.A(n_1497),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2813)
);

AOI22xp33_ASAP7_75t_L g2814 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_1277),
.Y(n_2815)
);

AOI22xp33_ASAP7_75t_L g2816 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2816)
);

INVx3_ASAP7_75t_L g2817 ( 
.A(n_1506),
.Y(n_2817)
);

O2A1O1Ixp33_ASAP7_75t_L g2818 ( 
.A1(n_1804),
.A2(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_1277),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_1277),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2822)
);

NOR2xp33_ASAP7_75t_L g2823 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2823)
);

NOR2xp67_ASAP7_75t_L g2824 ( 
.A(n_1349),
.B(n_853),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2825)
);

BUFx6f_ASAP7_75t_L g2826 ( 
.A(n_1381),
.Y(n_2826)
);

INVx2_ASAP7_75t_L g2827 ( 
.A(n_1277),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_SL g2828 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2828)
);

O2A1O1Ixp5_ASAP7_75t_L g2829 ( 
.A1(n_1804),
.A2(n_788),
.B(n_807),
.C(n_673),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2831)
);

CKINVDCx5p33_ASAP7_75t_R g2832 ( 
.A(n_1538),
.Y(n_2832)
);

AOI22xp5_ASAP7_75t_L g2833 ( 
.A1(n_1280),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2833)
);

INVx3_ASAP7_75t_L g2834 ( 
.A(n_1506),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2835)
);

INVxp67_ASAP7_75t_L g2836 ( 
.A(n_1349),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_L g2837 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2837)
);

BUFx6f_ASAP7_75t_L g2838 ( 
.A(n_1381),
.Y(n_2838)
);

O2A1O1Ixp5_ASAP7_75t_L g2839 ( 
.A1(n_1804),
.A2(n_788),
.B(n_807),
.C(n_673),
.Y(n_2839)
);

OAI21xp5_ASAP7_75t_L g2840 ( 
.A1(n_1804),
.A2(n_788),
.B(n_673),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_1277),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_1277),
.Y(n_2843)
);

NOR2xp33_ASAP7_75t_L g2844 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2844)
);

NAND2xp33_ASAP7_75t_L g2845 ( 
.A(n_1804),
.B(n_1066),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_1277),
.Y(n_2847)
);

AOI22xp33_ASAP7_75t_L g2848 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2848)
);

AOI22xp33_ASAP7_75t_SL g2849 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_SL g2851 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2851)
);

NAND2xp33_ASAP7_75t_L g2852 ( 
.A(n_1804),
.B(n_1066),
.Y(n_2852)
);

AOI22xp5_ASAP7_75t_L g2853 ( 
.A1(n_1280),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_SL g2856 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2856)
);

INVx2_ASAP7_75t_L g2857 ( 
.A(n_1277),
.Y(n_2857)
);

AOI22xp5_ASAP7_75t_L g2858 ( 
.A1(n_1280),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2858)
);

INVx2_ASAP7_75t_SL g2859 ( 
.A(n_1294),
.Y(n_2859)
);

NAND2xp33_ASAP7_75t_SL g2860 ( 
.A(n_1276),
.B(n_1581),
.Y(n_2860)
);

INVx2_ASAP7_75t_SL g2861 ( 
.A(n_1294),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_1277),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_1277),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_1277),
.Y(n_2864)
);

A2O1A1Ixp33_ASAP7_75t_L g2865 ( 
.A1(n_1804),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_2865)
);

OR2x2_ASAP7_75t_L g2866 ( 
.A(n_1285),
.B(n_846),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_SL g2867 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_1277),
.Y(n_2868)
);

NOR2xp33_ASAP7_75t_L g2869 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2869)
);

NOR2xp33_ASAP7_75t_L g2870 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_1277),
.Y(n_2871)
);

AOI22xp33_ASAP7_75t_L g2872 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2873)
);

INVx5_ASAP7_75t_L g2874 ( 
.A(n_1506),
.Y(n_2874)
);

O2A1O1Ixp33_ASAP7_75t_L g2875 ( 
.A1(n_1804),
.A2(n_1067),
.B(n_1087),
.C(n_1072),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_1277),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2877)
);

NOR2x2_ASAP7_75t_L g2878 ( 
.A(n_1524),
.B(n_948),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_1277),
.Y(n_2879)
);

NOR2xp33_ASAP7_75t_L g2880 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2880)
);

AOI22xp33_ASAP7_75t_L g2881 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_SL g2883 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2883)
);

NOR2x1p5_ASAP7_75t_L g2884 ( 
.A(n_1497),
.B(n_820),
.Y(n_2884)
);

BUFx3_ASAP7_75t_L g2885 ( 
.A(n_1294),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2886)
);

AOI22xp33_ASAP7_75t_L g2887 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2887)
);

NOR2xp33_ASAP7_75t_L g2888 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_1277),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_SL g2890 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2890)
);

AOI21xp5_ASAP7_75t_L g2891 ( 
.A1(n_1804),
.A2(n_907),
.B(n_653),
.Y(n_2891)
);

A2O1A1Ixp33_ASAP7_75t_L g2892 ( 
.A1(n_1804),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_2892)
);

INVx2_ASAP7_75t_SL g2893 ( 
.A(n_1294),
.Y(n_2893)
);

OAI22xp5_ASAP7_75t_L g2894 ( 
.A1(n_1804),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_2894)
);

O2A1O1Ixp5_ASAP7_75t_L g2895 ( 
.A1(n_1804),
.A2(n_788),
.B(n_807),
.C(n_673),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2896)
);

INVx2_ASAP7_75t_SL g2897 ( 
.A(n_1294),
.Y(n_2897)
);

AND2x4_ASAP7_75t_L g2898 ( 
.A(n_1335),
.B(n_1395),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2899)
);

AOI22xp33_ASAP7_75t_SL g2900 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_L g2901 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2901)
);

O2A1O1Ixp5_ASAP7_75t_L g2902 ( 
.A1(n_1804),
.A2(n_788),
.B(n_807),
.C(n_673),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_L g2903 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_SL g2904 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_1277),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_1277),
.Y(n_2906)
);

AND2x6_ASAP7_75t_SL g2907 ( 
.A(n_1489),
.B(n_1541),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_L g2908 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2908)
);

INVx2_ASAP7_75t_L g2909 ( 
.A(n_1277),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_SL g2910 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2910)
);

NAND2xp33_ASAP7_75t_L g2911 ( 
.A(n_1804),
.B(n_1066),
.Y(n_2911)
);

AND2x4_ASAP7_75t_L g2912 ( 
.A(n_1335),
.B(n_1395),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_1277),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2914)
);

OAI22xp5_ASAP7_75t_L g2915 ( 
.A1(n_1804),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_2915)
);

NOR3xp33_ASAP7_75t_L g2916 ( 
.A(n_1804),
.B(n_1072),
.C(n_1067),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_SL g2917 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2918)
);

NOR2xp33_ASAP7_75t_L g2919 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_SL g2920 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2920)
);

INVx2_ASAP7_75t_SL g2921 ( 
.A(n_1294),
.Y(n_2921)
);

NAND3xp33_ASAP7_75t_L g2922 ( 
.A(n_1804),
.B(n_1072),
.C(n_1067),
.Y(n_2922)
);

AOI22xp33_ASAP7_75t_L g2923 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2923)
);

INVx2_ASAP7_75t_SL g2924 ( 
.A(n_1294),
.Y(n_2924)
);

NAND2xp5_ASAP7_75t_L g2925 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2925)
);

AOI21xp5_ASAP7_75t_L g2926 ( 
.A1(n_1804),
.A2(n_907),
.B(n_653),
.Y(n_2926)
);

AND2x2_ASAP7_75t_SL g2927 ( 
.A(n_1311),
.B(n_1067),
.Y(n_2927)
);

AND2x6_ASAP7_75t_SL g2928 ( 
.A(n_1489),
.B(n_1541),
.Y(n_2928)
);

INVx2_ASAP7_75t_SL g2929 ( 
.A(n_1294),
.Y(n_2929)
);

AOI22xp33_ASAP7_75t_L g2930 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2930)
);

NOR2xp33_ASAP7_75t_L g2931 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2931)
);

NAND2xp5_ASAP7_75t_L g2932 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2932)
);

NOR2xp33_ASAP7_75t_L g2933 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2934)
);

NOR2xp33_ASAP7_75t_L g2935 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2935)
);

INVxp67_ASAP7_75t_L g2936 ( 
.A(n_1349),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_SL g2937 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2937)
);

NAND2x1p5_ASAP7_75t_L g2938 ( 
.A(n_1374),
.B(n_1009),
.Y(n_2938)
);

OR2x2_ASAP7_75t_L g2939 ( 
.A(n_1285),
.B(n_846),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_1277),
.Y(n_2940)
);

NOR2xp33_ASAP7_75t_L g2941 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_SL g2943 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_SL g2944 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2944)
);

AOI22xp33_ASAP7_75t_L g2945 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2945)
);

OAI21xp5_ASAP7_75t_L g2946 ( 
.A1(n_1804),
.A2(n_788),
.B(n_673),
.Y(n_2946)
);

BUFx12f_ASAP7_75t_L g2947 ( 
.A(n_1497),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2948)
);

NOR2xp33_ASAP7_75t_L g2949 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2949)
);

INVx2_ASAP7_75t_SL g2950 ( 
.A(n_1294),
.Y(n_2950)
);

NOR2xp33_ASAP7_75t_L g2951 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_SL g2952 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2952)
);

INVx2_ASAP7_75t_L g2953 ( 
.A(n_1277),
.Y(n_2953)
);

NOR2xp33_ASAP7_75t_L g2954 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2954)
);

AND2x2_ASAP7_75t_L g2955 ( 
.A(n_1275),
.B(n_839),
.Y(n_2955)
);

INVx2_ASAP7_75t_L g2956 ( 
.A(n_1277),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_1277),
.Y(n_2957)
);

AO22x1_ASAP7_75t_L g2958 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_SL g2959 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_1277),
.Y(n_2960)
);

AOI22xp33_ASAP7_75t_L g2961 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_L g2962 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_1277),
.Y(n_2963)
);

AOI21xp5_ASAP7_75t_L g2964 ( 
.A1(n_1804),
.A2(n_907),
.B(n_653),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2966)
);

CKINVDCx5p33_ASAP7_75t_R g2967 ( 
.A(n_1538),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_SL g2968 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_1277),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_L g2971 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2971)
);

AOI22xp33_ASAP7_75t_L g2972 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2972)
);

OAI21xp33_ASAP7_75t_L g2973 ( 
.A1(n_1804),
.A2(n_1072),
.B(n_1067),
.Y(n_2973)
);

OAI22xp5_ASAP7_75t_L g2974 ( 
.A1(n_1804),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_L g2975 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2975)
);

NAND2xp33_ASAP7_75t_L g2976 ( 
.A(n_1804),
.B(n_1066),
.Y(n_2976)
);

AND2x6_ASAP7_75t_L g2977 ( 
.A(n_1339),
.B(n_934),
.Y(n_2977)
);

AOI22xp33_ASAP7_75t_L g2978 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_L g2979 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2979)
);

AND2x6_ASAP7_75t_SL g2980 ( 
.A(n_1489),
.B(n_1541),
.Y(n_2980)
);

AOI22xp33_ASAP7_75t_L g2981 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_1277),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_1277),
.Y(n_2983)
);

NOR2xp33_ASAP7_75t_L g2984 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2984)
);

NOR2xp33_ASAP7_75t_L g2985 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_SL g2986 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_1277),
.Y(n_2987)
);

INVxp67_ASAP7_75t_L g2988 ( 
.A(n_1349),
.Y(n_2988)
);

NOR2xp33_ASAP7_75t_L g2989 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2989)
);

INVx2_ASAP7_75t_L g2990 ( 
.A(n_1277),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_SL g2991 ( 
.A(n_1804),
.B(n_1067),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_1276),
.B(n_1067),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_1277),
.Y(n_2994)
);

AND2x4_ASAP7_75t_L g2995 ( 
.A(n_1335),
.B(n_1395),
.Y(n_2995)
);

INVx2_ASAP7_75t_SL g2996 ( 
.A(n_1294),
.Y(n_2996)
);

NOR2xp33_ASAP7_75t_L g2997 ( 
.A(n_1632),
.B(n_1067),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_1277),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_SL g2999 ( 
.A(n_1804),
.B(n_1096),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3000)
);

NAND2xp5_ASAP7_75t_SL g3001 ( 
.A(n_1804),
.B(n_1096),
.Y(n_3001)
);

INVx3_ASAP7_75t_L g3002 ( 
.A(n_1506),
.Y(n_3002)
);

INVxp67_ASAP7_75t_SL g3003 ( 
.A(n_1276),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_1277),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_L g3006 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3007)
);

NAND2xp5_ASAP7_75t_SL g3008 ( 
.A(n_1804),
.B(n_1096),
.Y(n_3008)
);

BUFx8_ASAP7_75t_L g3009 ( 
.A(n_1385),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3010)
);

NOR2x2_ASAP7_75t_L g3011 ( 
.A(n_1524),
.B(n_948),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_1277),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_L g3013 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3013)
);

OAI22xp5_ASAP7_75t_L g3014 ( 
.A1(n_1804),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_3014)
);

INVx2_ASAP7_75t_SL g3015 ( 
.A(n_1294),
.Y(n_3015)
);

NOR3x1_ASAP7_75t_L g3016 ( 
.A(n_1632),
.B(n_1182),
.C(n_1124),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_1277),
.Y(n_3017)
);

AND2x4_ASAP7_75t_L g3018 ( 
.A(n_1335),
.B(n_1395),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3019)
);

AND2x4_ASAP7_75t_L g3020 ( 
.A(n_1335),
.B(n_1395),
.Y(n_3020)
);

INVx5_ASAP7_75t_L g3021 ( 
.A(n_1506),
.Y(n_3021)
);

NOR2xp33_ASAP7_75t_L g3022 ( 
.A(n_1632),
.B(n_1067),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3023)
);

NAND3xp33_ASAP7_75t_L g3024 ( 
.A(n_1804),
.B(n_1072),
.C(n_1067),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_1277),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_L g3026 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_1277),
.Y(n_3027)
);

AOI22xp33_ASAP7_75t_L g3028 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_3028)
);

AOI21xp5_ASAP7_75t_L g3029 ( 
.A1(n_1804),
.A2(n_907),
.B(n_653),
.Y(n_3029)
);

OR2x2_ASAP7_75t_L g3030 ( 
.A(n_1285),
.B(n_846),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_SL g3031 ( 
.A(n_1804),
.B(n_1096),
.Y(n_3031)
);

BUFx3_ASAP7_75t_L g3032 ( 
.A(n_1294),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3033)
);

INVx2_ASAP7_75t_L g3034 ( 
.A(n_1277),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3035)
);

BUFx8_ASAP7_75t_L g3036 ( 
.A(n_1385),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_SL g3038 ( 
.A(n_1804),
.B(n_1067),
.Y(n_3038)
);

NOR2xp33_ASAP7_75t_L g3039 ( 
.A(n_1632),
.B(n_1067),
.Y(n_3039)
);

OAI221xp5_ASAP7_75t_L g3040 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1090),
.B2(n_1087),
.C(n_1067),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_SL g3041 ( 
.A(n_1804),
.B(n_1067),
.Y(n_3041)
);

NAND3xp33_ASAP7_75t_SL g3042 ( 
.A(n_1804),
.B(n_1072),
.C(n_1067),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3043)
);

BUFx2_ASAP7_75t_SL g3044 ( 
.A(n_1404),
.Y(n_3044)
);

A2O1A1Ixp33_ASAP7_75t_L g3045 ( 
.A1(n_1804),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_3045)
);

AOI22xp5_ASAP7_75t_L g3046 ( 
.A1(n_1280),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_3046)
);

AOI22xp33_ASAP7_75t_L g3047 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_3047)
);

NAND3xp33_ASAP7_75t_L g3048 ( 
.A(n_1804),
.B(n_1072),
.C(n_1067),
.Y(n_3048)
);

XOR2x2_ASAP7_75t_L g3049 ( 
.A(n_1759),
.B(n_1193),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_1277),
.Y(n_3050)
);

AOI22xp5_ASAP7_75t_L g3051 ( 
.A1(n_1280),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_3051)
);

INVx2_ASAP7_75t_SL g3052 ( 
.A(n_1294),
.Y(n_3052)
);

OAI22xp5_ASAP7_75t_SL g3053 ( 
.A1(n_1701),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_3053)
);

INVx3_ASAP7_75t_L g3054 ( 
.A(n_1506),
.Y(n_3054)
);

BUFx2_ASAP7_75t_SL g3055 ( 
.A(n_1404),
.Y(n_3055)
);

NOR2xp33_ASAP7_75t_L g3056 ( 
.A(n_1632),
.B(n_1067),
.Y(n_3056)
);

INVx2_ASAP7_75t_L g3057 ( 
.A(n_1277),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_SL g3058 ( 
.A(n_1804),
.B(n_1096),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_L g3059 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3059)
);

NOR2xp33_ASAP7_75t_L g3060 ( 
.A(n_1632),
.B(n_1067),
.Y(n_3060)
);

NAND2xp5_ASAP7_75t_L g3061 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_SL g3062 ( 
.A(n_1804),
.B(n_1096),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_1277),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_1277),
.Y(n_3064)
);

NAND2xp33_ASAP7_75t_L g3065 ( 
.A(n_1804),
.B(n_1066),
.Y(n_3065)
);

AOI22xp33_ASAP7_75t_L g3066 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_3066)
);

OAI22xp33_ASAP7_75t_L g3067 ( 
.A1(n_1804),
.A2(n_1089),
.B1(n_1198),
.B2(n_1081),
.Y(n_3067)
);

AND2x4_ASAP7_75t_SL g3068 ( 
.A(n_1274),
.B(n_854),
.Y(n_3068)
);

HB1xp67_ASAP7_75t_L g3069 ( 
.A(n_1780),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_L g3070 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3072)
);

INVxp67_ASAP7_75t_L g3073 ( 
.A(n_1349),
.Y(n_3073)
);

NOR2xp33_ASAP7_75t_L g3074 ( 
.A(n_1632),
.B(n_1067),
.Y(n_3074)
);

AOI21xp5_ASAP7_75t_L g3075 ( 
.A1(n_1804),
.A2(n_907),
.B(n_653),
.Y(n_3075)
);

INVxp67_ASAP7_75t_SL g3076 ( 
.A(n_1276),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_SL g3077 ( 
.A(n_1804),
.B(n_1096),
.Y(n_3077)
);

NOR2xp33_ASAP7_75t_L g3078 ( 
.A(n_1632),
.B(n_1067),
.Y(n_3078)
);

BUFx2_ASAP7_75t_L g3079 ( 
.A(n_1967),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_SL g3081 ( 
.A(n_1804),
.B(n_1096),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_SL g3082 ( 
.A(n_1804),
.B(n_1096),
.Y(n_3082)
);

NOR2x2_ASAP7_75t_L g3083 ( 
.A(n_1524),
.B(n_948),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_L g3084 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_L g3085 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_SL g3086 ( 
.A(n_1804),
.B(n_1096),
.Y(n_3086)
);

INVx2_ASAP7_75t_SL g3087 ( 
.A(n_1294),
.Y(n_3087)
);

NOR2xp33_ASAP7_75t_L g3088 ( 
.A(n_1632),
.B(n_1067),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_SL g3089 ( 
.A(n_1804),
.B(n_1096),
.Y(n_3089)
);

A2O1A1Ixp33_ASAP7_75t_L g3090 ( 
.A1(n_1804),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_L g3091 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3091)
);

OAI22xp5_ASAP7_75t_L g3092 ( 
.A1(n_1804),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_3092)
);

OAI221xp5_ASAP7_75t_L g3093 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1090),
.B2(n_1087),
.C(n_1067),
.Y(n_3093)
);

AOI22x1_ASAP7_75t_SL g3094 ( 
.A1(n_1363),
.A2(n_1604),
.B1(n_1753),
.B2(n_1662),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3096)
);

NOR2xp33_ASAP7_75t_SL g3097 ( 
.A(n_1662),
.B(n_396),
.Y(n_3097)
);

AOI22xp33_ASAP7_75t_L g3098 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_1277),
.Y(n_3099)
);

HB1xp67_ASAP7_75t_L g3100 ( 
.A(n_1780),
.Y(n_3100)
);

AOI22xp33_ASAP7_75t_L g3101 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_1277),
.Y(n_3102)
);

INVx2_ASAP7_75t_L g3103 ( 
.A(n_1277),
.Y(n_3103)
);

NOR2xp33_ASAP7_75t_L g3104 ( 
.A(n_1632),
.B(n_1067),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_L g3105 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3105)
);

OR2x2_ASAP7_75t_L g3106 ( 
.A(n_1285),
.B(n_846),
.Y(n_3106)
);

NAND2xp33_ASAP7_75t_L g3107 ( 
.A(n_1804),
.B(n_1066),
.Y(n_3107)
);

AOI22xp5_ASAP7_75t_L g3108 ( 
.A1(n_1280),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_1277),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_1277),
.Y(n_3110)
);

INVx2_ASAP7_75t_L g3111 ( 
.A(n_1277),
.Y(n_3111)
);

AND2x6_ASAP7_75t_L g3112 ( 
.A(n_1339),
.B(n_934),
.Y(n_3112)
);

INVx5_ASAP7_75t_L g3113 ( 
.A(n_1506),
.Y(n_3113)
);

BUFx6f_ASAP7_75t_L g3114 ( 
.A(n_1381),
.Y(n_3114)
);

AOI22xp5_ASAP7_75t_L g3115 ( 
.A1(n_1280),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_3115)
);

INVx2_ASAP7_75t_L g3116 ( 
.A(n_1277),
.Y(n_3116)
);

NOR2xp33_ASAP7_75t_L g3117 ( 
.A(n_1632),
.B(n_1067),
.Y(n_3117)
);

AO22x1_ASAP7_75t_L g3118 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_L g3119 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3119)
);

INVx2_ASAP7_75t_L g3120 ( 
.A(n_1277),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_SL g3121 ( 
.A(n_1804),
.B(n_1067),
.Y(n_3121)
);

AND2x6_ASAP7_75t_SL g3122 ( 
.A(n_1489),
.B(n_1541),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_L g3123 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3124)
);

HB1xp67_ASAP7_75t_L g3125 ( 
.A(n_1780),
.Y(n_3125)
);

NOR2xp67_ASAP7_75t_L g3126 ( 
.A(n_1349),
.B(n_853),
.Y(n_3126)
);

A2O1A1Ixp33_ASAP7_75t_L g3127 ( 
.A1(n_1804),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_3127)
);

NOR2xp33_ASAP7_75t_L g3128 ( 
.A(n_1632),
.B(n_1067),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_1277),
.Y(n_3129)
);

AND2x6_ASAP7_75t_SL g3130 ( 
.A(n_1489),
.B(n_1541),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_1277),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_SL g3132 ( 
.A(n_1804),
.B(n_1096),
.Y(n_3132)
);

AND2x4_ASAP7_75t_L g3133 ( 
.A(n_1335),
.B(n_1395),
.Y(n_3133)
);

INVx2_ASAP7_75t_L g3134 ( 
.A(n_1277),
.Y(n_3134)
);

AOI22xp33_ASAP7_75t_L g3135 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_L g3137 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3137)
);

AND2x2_ASAP7_75t_L g3138 ( 
.A(n_1275),
.B(n_839),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3140)
);

BUFx3_ASAP7_75t_L g3141 ( 
.A(n_1294),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_SL g3144 ( 
.A(n_1804),
.B(n_1096),
.Y(n_3144)
);

NOR2x2_ASAP7_75t_L g3145 ( 
.A(n_1524),
.B(n_948),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_L g3146 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3146)
);

INVx8_ASAP7_75t_L g3147 ( 
.A(n_1294),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_L g3148 ( 
.A(n_1276),
.B(n_1067),
.Y(n_3148)
);

INVx2_ASAP7_75t_L g3149 ( 
.A(n_1277),
.Y(n_3149)
);

INVx2_ASAP7_75t_L g3150 ( 
.A(n_1277),
.Y(n_3150)
);

AOI22xp33_ASAP7_75t_L g3151 ( 
.A1(n_1804),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_3151)
);

BUFx2_ASAP7_75t_L g3152 ( 
.A(n_1967),
.Y(n_3152)
);

OAI22xp5_ASAP7_75t_L g3153 ( 
.A1(n_1804),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_SL g3154 ( 
.A(n_1804),
.B(n_1096),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_SL g3155 ( 
.A(n_1804),
.B(n_1067),
.Y(n_3155)
);

NAND2xp5_ASAP7_75t_L g3156 ( 
.A(n_2135),
.B(n_2050),
.Y(n_3156)
);

AND2x2_ASAP7_75t_L g3157 ( 
.A(n_2549),
.B(n_2780),
.Y(n_3157)
);

AOI21xp5_ASAP7_75t_L g3158 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3158)
);

CKINVDCx6p67_ASAP7_75t_R g3159 ( 
.A(n_2180),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_SL g3160 ( 
.A(n_2374),
.B(n_2569),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2232),
.Y(n_3161)
);

OAI21xp5_ASAP7_75t_L g3162 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_3162)
);

NOR2xp33_ASAP7_75t_L g3163 ( 
.A(n_2025),
.B(n_2030),
.Y(n_3163)
);

AOI22xp5_ASAP7_75t_L g3164 ( 
.A1(n_3053),
.A2(n_1987),
.B1(n_2784),
.B2(n_2749),
.Y(n_3164)
);

OAI21xp5_ASAP7_75t_L g3165 ( 
.A1(n_2839),
.A2(n_2902),
.B(n_2895),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_2091),
.B(n_2365),
.Y(n_3166)
);

AOI21xp5_ASAP7_75t_L g3167 ( 
.A1(n_2712),
.A2(n_2926),
.B(n_2891),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2232),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_2091),
.B(n_2366),
.Y(n_3169)
);

INVx2_ASAP7_75t_L g3170 ( 
.A(n_1988),
.Y(n_3170)
);

AOI21xp5_ASAP7_75t_L g3171 ( 
.A1(n_2964),
.A2(n_3075),
.B(n_3029),
.Y(n_3171)
);

INVx2_ASAP7_75t_SL g3172 ( 
.A(n_2054),
.Y(n_3172)
);

A2O1A1Ixp33_ASAP7_75t_L g3173 ( 
.A1(n_2737),
.A2(n_2946),
.B(n_2840),
.C(n_2487),
.Y(n_3173)
);

INVxp67_ASAP7_75t_L g3174 ( 
.A(n_2760),
.Y(n_3174)
);

AOI21xp5_ASAP7_75t_L g3175 ( 
.A1(n_2005),
.A2(n_1988),
.B(n_3154),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_L g3176 ( 
.A(n_2135),
.B(n_2050),
.Y(n_3176)
);

AOI21xp5_ASAP7_75t_L g3177 ( 
.A1(n_2550),
.A2(n_2714),
.B(n_2577),
.Y(n_3177)
);

NOR2xp33_ASAP7_75t_L g3178 ( 
.A(n_2025),
.B(n_2030),
.Y(n_3178)
);

BUFx2_ASAP7_75t_L g3179 ( 
.A(n_2760),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_L g3180 ( 
.A(n_2055),
.B(n_2121),
.Y(n_3180)
);

CKINVDCx6p67_ASAP7_75t_R g3181 ( 
.A(n_2180),
.Y(n_3181)
);

AOI22xp5_ASAP7_75t_L g3182 ( 
.A1(n_2789),
.A2(n_2915),
.B1(n_2974),
.B2(n_2894),
.Y(n_3182)
);

AOI21xp5_ASAP7_75t_L g3183 ( 
.A1(n_2588),
.A2(n_2748),
.B(n_2676),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_L g3184 ( 
.A(n_2055),
.B(n_2121),
.Y(n_3184)
);

O2A1O1Ixp5_ASAP7_75t_L g3185 ( 
.A1(n_2516),
.A2(n_3118),
.B(n_2958),
.C(n_3014),
.Y(n_3185)
);

AOI22xp5_ASAP7_75t_L g3186 ( 
.A1(n_3092),
.A2(n_3153),
.B1(n_2045),
.B2(n_2047),
.Y(n_3186)
);

INVxp67_ASAP7_75t_L g3187 ( 
.A(n_3069),
.Y(n_3187)
);

AOI21xp5_ASAP7_75t_L g3188 ( 
.A1(n_2548),
.A2(n_2777),
.B(n_2623),
.Y(n_3188)
);

AOI21xp5_ASAP7_75t_L g3189 ( 
.A1(n_2363),
.A2(n_2828),
.B(n_2550),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_SL g3190 ( 
.A(n_2112),
.B(n_2033),
.Y(n_3190)
);

NOR2xp33_ASAP7_75t_L g3191 ( 
.A(n_2044),
.B(n_2045),
.Y(n_3191)
);

NAND2xp5_ASAP7_75t_L g3192 ( 
.A(n_2127),
.B(n_2138),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_1989),
.Y(n_3193)
);

INVx11_ASAP7_75t_L g3194 ( 
.A(n_2177),
.Y(n_3194)
);

BUFx4f_ASAP7_75t_L g3195 ( 
.A(n_2566),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_L g3196 ( 
.A(n_2127),
.B(n_2140),
.Y(n_3196)
);

NOR3xp33_ASAP7_75t_L g3197 ( 
.A(n_3040),
.B(n_3093),
.C(n_2600),
.Y(n_3197)
);

OAI21xp5_ASAP7_75t_L g3198 ( 
.A1(n_2145),
.A2(n_2535),
.B(n_2363),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_1996),
.Y(n_3199)
);

A2O1A1Ixp33_ASAP7_75t_L g3200 ( 
.A1(n_2407),
.A2(n_2775),
.B(n_2818),
.C(n_2730),
.Y(n_3200)
);

NAND2xp33_ASAP7_75t_L g3201 ( 
.A(n_2416),
.B(n_2430),
.Y(n_3201)
);

AND2x4_ASAP7_75t_L g3202 ( 
.A(n_2098),
.B(n_2221),
.Y(n_3202)
);

AOI21x1_ASAP7_75t_L g3203 ( 
.A1(n_2167),
.A2(n_2024),
.B(n_2101),
.Y(n_3203)
);

INVx2_ASAP7_75t_L g3204 ( 
.A(n_2024),
.Y(n_3204)
);

OAI21xp5_ASAP7_75t_L g3205 ( 
.A1(n_2535),
.A2(n_2546),
.B(n_2543),
.Y(n_3205)
);

AOI21x1_ASAP7_75t_L g3206 ( 
.A1(n_2101),
.A2(n_2155),
.B(n_2021),
.Y(n_3206)
);

AOI21xp5_ASAP7_75t_L g3207 ( 
.A1(n_2543),
.A2(n_2676),
.B(n_2588),
.Y(n_3207)
);

AND2x4_ASAP7_75t_L g3208 ( 
.A(n_2098),
.B(n_2116),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_SL g3209 ( 
.A(n_2088),
.B(n_2703),
.Y(n_3209)
);

NOR3xp33_ASAP7_75t_L g3210 ( 
.A(n_2875),
.B(n_2004),
.C(n_3042),
.Y(n_3210)
);

AOI21xp5_ASAP7_75t_L g3211 ( 
.A1(n_2999),
.A2(n_3144),
.B(n_3077),
.Y(n_3211)
);

OAI21xp5_ASAP7_75t_L g3212 ( 
.A1(n_2546),
.A2(n_2554),
.B(n_2548),
.Y(n_3212)
);

BUFx8_ASAP7_75t_L g3213 ( 
.A(n_2125),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_2019),
.Y(n_3214)
);

O2A1O1Ixp5_ASAP7_75t_L g3215 ( 
.A1(n_3154),
.A2(n_2554),
.B(n_2578),
.C(n_2577),
.Y(n_3215)
);

AOI21xp5_ASAP7_75t_L g3216 ( 
.A1(n_2797),
.A2(n_3082),
.B(n_2883),
.Y(n_3216)
);

AO21x1_ASAP7_75t_L g3217 ( 
.A1(n_2578),
.A2(n_2591),
.B(n_2590),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_2146),
.B(n_2148),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_L g3219 ( 
.A(n_2151),
.B(n_2153),
.Y(n_3219)
);

NAND2xp33_ASAP7_75t_SL g3220 ( 
.A(n_2172),
.B(n_2159),
.Y(n_3220)
);

OAI21xp5_ASAP7_75t_L g3221 ( 
.A1(n_2590),
.A2(n_2598),
.B(n_2591),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_SL g3222 ( 
.A(n_2849),
.B(n_2900),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_2156),
.B(n_2160),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_L g3224 ( 
.A(n_2539),
.B(n_3067),
.Y(n_3224)
);

AOI21xp5_ASAP7_75t_L g3225 ( 
.A1(n_2598),
.A2(n_3144),
.B(n_2714),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_L g3226 ( 
.A(n_2539),
.B(n_3067),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_2031),
.Y(n_3227)
);

NAND2xp5_ASAP7_75t_SL g3228 ( 
.A(n_1993),
.B(n_2017),
.Y(n_3228)
);

AOI21xp5_ASAP7_75t_L g3229 ( 
.A1(n_2659),
.A2(n_2797),
.B(n_2693),
.Y(n_3229)
);

INVx4_ASAP7_75t_L g3230 ( 
.A(n_2009),
.Y(n_3230)
);

AOI21x1_ASAP7_75t_L g3231 ( 
.A1(n_2155),
.A2(n_2021),
.B(n_2606),
.Y(n_3231)
);

NOR3xp33_ASAP7_75t_L g3232 ( 
.A(n_2006),
.B(n_2922),
.C(n_2526),
.Y(n_3232)
);

O2A1O1Ixp33_ASAP7_75t_L g3233 ( 
.A1(n_2383),
.A2(n_2538),
.B(n_2545),
.C(n_2386),
.Y(n_3233)
);

INVx2_ASAP7_75t_L g3234 ( 
.A(n_2038),
.Y(n_3234)
);

NAND2xp5_ASAP7_75t_L g3235 ( 
.A(n_2369),
.B(n_2370),
.Y(n_3235)
);

INVx2_ASAP7_75t_L g3236 ( 
.A(n_2059),
.Y(n_3236)
);

A2O1A1Ixp33_ASAP7_75t_L g3237 ( 
.A1(n_2362),
.A2(n_2387),
.B(n_2389),
.C(n_2373),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_2072),
.Y(n_3238)
);

AOI21x1_ASAP7_75t_L g3239 ( 
.A1(n_2606),
.A2(n_2659),
.B(n_2623),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_2087),
.Y(n_3240)
);

AOI21xp5_ASAP7_75t_L g3241 ( 
.A1(n_2693),
.A2(n_3001),
.B(n_2683),
.Y(n_3241)
);

BUFx6f_ASAP7_75t_L g3242 ( 
.A(n_2098),
.Y(n_3242)
);

OAI21xp33_ASAP7_75t_L g3243 ( 
.A1(n_2390),
.A2(n_2541),
.B(n_2484),
.Y(n_3243)
);

AOI21xp5_ASAP7_75t_L g3244 ( 
.A1(n_2748),
.A2(n_2856),
.B(n_2828),
.Y(n_3244)
);

NOR2xp33_ASAP7_75t_L g3245 ( 
.A(n_2044),
.B(n_2047),
.Y(n_3245)
);

AO21x1_ASAP7_75t_L g3246 ( 
.A1(n_2675),
.A2(n_2759),
.B(n_2683),
.Y(n_3246)
);

AOI21xp5_ASAP7_75t_L g3247 ( 
.A1(n_3062),
.A2(n_3089),
.B(n_3081),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_L g3248 ( 
.A(n_2376),
.B(n_2379),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_L g3249 ( 
.A(n_2381),
.B(n_2382),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_2384),
.B(n_2392),
.Y(n_3250)
);

INVx1_ASAP7_75t_SL g3251 ( 
.A(n_2144),
.Y(n_3251)
);

O2A1O1Ixp33_ASAP7_75t_SL g3252 ( 
.A1(n_2715),
.A2(n_2865),
.B(n_2892),
.C(n_2802),
.Y(n_3252)
);

AOI21xp5_ASAP7_75t_L g3253 ( 
.A1(n_2801),
.A2(n_3008),
.B(n_2883),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_2092),
.Y(n_3254)
);

A2O1A1Ixp33_ASAP7_75t_L g3255 ( 
.A1(n_2362),
.A2(n_2387),
.B(n_2389),
.C(n_2373),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_2118),
.Y(n_3256)
);

NOR2xp33_ASAP7_75t_L g3257 ( 
.A(n_2060),
.B(n_2571),
.Y(n_3257)
);

AND2x2_ASAP7_75t_L g3258 ( 
.A(n_2780),
.B(n_2795),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_2150),
.Y(n_3259)
);

AOI21xp5_ASAP7_75t_L g3260 ( 
.A1(n_2867),
.A2(n_3089),
.B(n_3081),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_L g3261 ( 
.A(n_2394),
.B(n_2395),
.Y(n_3261)
);

INVx3_ASAP7_75t_L g3262 ( 
.A(n_2098),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_SL g3263 ( 
.A(n_2013),
.B(n_2032),
.Y(n_3263)
);

O2A1O1Ixp33_ASAP7_75t_L g3264 ( 
.A1(n_3045),
.A2(n_3127),
.B(n_3090),
.C(n_2402),
.Y(n_3264)
);

NAND2xp5_ASAP7_75t_L g3265 ( 
.A(n_2399),
.B(n_2405),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_L g3266 ( 
.A(n_2410),
.B(n_2413),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_2415),
.B(n_2417),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_2423),
.B(n_2426),
.Y(n_3268)
);

AOI21xp5_ASAP7_75t_L g3269 ( 
.A1(n_2772),
.A2(n_3062),
.B(n_3001),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_2432),
.B(n_2433),
.Y(n_3270)
);

OAI21xp33_ASAP7_75t_L g3271 ( 
.A1(n_2589),
.A2(n_2629),
.B(n_2612),
.Y(n_3271)
);

AOI21xp5_ASAP7_75t_L g3272 ( 
.A1(n_3031),
.A2(n_2772),
.B(n_2759),
.Y(n_3272)
);

NAND2xp5_ASAP7_75t_L g3273 ( 
.A(n_2435),
.B(n_2437),
.Y(n_3273)
);

O2A1O1Ixp33_ASAP7_75t_L g3274 ( 
.A1(n_2398),
.A2(n_2420),
.B(n_2429),
.C(n_2402),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_2171),
.Y(n_3275)
);

AND2x2_ASAP7_75t_L g3276 ( 
.A(n_2795),
.B(n_2927),
.Y(n_3276)
);

AND2x2_ASAP7_75t_L g3277 ( 
.A(n_2927),
.B(n_2016),
.Y(n_3277)
);

AOI21xp5_ASAP7_75t_L g3278 ( 
.A1(n_2999),
.A2(n_3082),
.B(n_2801),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_SL g3279 ( 
.A(n_2078),
.B(n_2043),
.Y(n_3279)
);

AOI21xp5_ASAP7_75t_L g3280 ( 
.A1(n_3086),
.A2(n_2851),
.B(n_2777),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_2443),
.B(n_2446),
.Y(n_3281)
);

BUFx6f_ASAP7_75t_L g3282 ( 
.A(n_2027),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_L g3283 ( 
.A(n_2453),
.B(n_2454),
.Y(n_3283)
);

AND2x2_ASAP7_75t_L g3284 ( 
.A(n_2002),
.B(n_2143),
.Y(n_3284)
);

INVx2_ASAP7_75t_SL g3285 ( 
.A(n_2054),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_SL g3286 ( 
.A(n_2576),
.B(n_2604),
.Y(n_3286)
);

INVxp67_ASAP7_75t_L g3287 ( 
.A(n_3069),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_2456),
.B(n_2458),
.Y(n_3288)
);

AOI21xp5_ASAP7_75t_L g3289 ( 
.A1(n_2851),
.A2(n_3008),
.B(n_2867),
.Y(n_3289)
);

OAI22xp5_ASAP7_75t_L g3290 ( 
.A1(n_2646),
.A2(n_2833),
.B1(n_2853),
.B2(n_2776),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_2174),
.Y(n_3291)
);

NAND2xp5_ASAP7_75t_L g3292 ( 
.A(n_2462),
.B(n_2463),
.Y(n_3292)
);

BUFx12f_ASAP7_75t_L g3293 ( 
.A(n_2328),
.Y(n_3293)
);

A2O1A1Ixp33_ASAP7_75t_L g3294 ( 
.A1(n_2398),
.A2(n_2429),
.B(n_2431),
.C(n_2420),
.Y(n_3294)
);

NOR2xp67_ASAP7_75t_L g3295 ( 
.A(n_2009),
.B(n_2743),
.Y(n_3295)
);

O2A1O1Ixp33_ASAP7_75t_L g3296 ( 
.A1(n_2431),
.A2(n_2468),
.B(n_2471),
.C(n_2455),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_2464),
.B(n_2469),
.Y(n_3297)
);

AOI22x1_ASAP7_75t_L g3298 ( 
.A1(n_3003),
.A2(n_3076),
.B1(n_2227),
.B2(n_2267),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_2470),
.B(n_2474),
.Y(n_3299)
);

NOR2xp33_ASAP7_75t_L g3300 ( 
.A(n_2060),
.B(n_2858),
.Y(n_3300)
);

NOR3xp33_ASAP7_75t_L g3301 ( 
.A(n_3024),
.B(n_3048),
.C(n_2973),
.Y(n_3301)
);

AOI21xp5_ASAP7_75t_L g3302 ( 
.A1(n_2856),
.A2(n_3077),
.B(n_2904),
.Y(n_3302)
);

OAI21xp5_ASAP7_75t_L g3303 ( 
.A1(n_2890),
.A2(n_3031),
.B(n_2904),
.Y(n_3303)
);

BUFx3_ASAP7_75t_L g3304 ( 
.A(n_2719),
.Y(n_3304)
);

OAI21xp5_ASAP7_75t_L g3305 ( 
.A1(n_2890),
.A2(n_3086),
.B(n_3058),
.Y(n_3305)
);

AOI21xp5_ASAP7_75t_L g3306 ( 
.A1(n_3058),
.A2(n_3132),
.B(n_2203),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_2475),
.B(n_2478),
.Y(n_3307)
);

AND2x2_ASAP7_75t_L g3308 ( 
.A(n_2002),
.B(n_2139),
.Y(n_3308)
);

AOI22xp5_ASAP7_75t_L g3309 ( 
.A1(n_2662),
.A2(n_2916),
.B1(n_2766),
.B2(n_2468),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_2482),
.B(n_2489),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_2492),
.B(n_2495),
.Y(n_3311)
);

OAI21xp5_ASAP7_75t_L g3312 ( 
.A1(n_3132),
.A2(n_2003),
.B(n_2455),
.Y(n_3312)
);

NOR2xp33_ASAP7_75t_L g3313 ( 
.A(n_3046),
.B(n_3051),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_2496),
.B(n_2501),
.Y(n_3314)
);

OAI22xp5_ASAP7_75t_L g3315 ( 
.A1(n_3108),
.A2(n_3115),
.B1(n_2421),
.B2(n_2466),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_2503),
.B(n_2507),
.Y(n_3316)
);

AOI21xp5_ASAP7_75t_L g3317 ( 
.A1(n_2203),
.A2(n_2093),
.B(n_2075),
.Y(n_3317)
);

NOR2xp33_ASAP7_75t_L g3318 ( 
.A(n_2471),
.B(n_2477),
.Y(n_3318)
);

INVx2_ASAP7_75t_L g3319 ( 
.A(n_2233),
.Y(n_3319)
);

NAND2xp5_ASAP7_75t_L g3320 ( 
.A(n_2508),
.B(n_2509),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_2244),
.Y(n_3321)
);

OAI21xp33_ASAP7_75t_L g3322 ( 
.A1(n_2477),
.A2(n_2483),
.B(n_2479),
.Y(n_3322)
);

OAI21xp5_ASAP7_75t_L g3323 ( 
.A1(n_2479),
.A2(n_2542),
.B(n_2483),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_2256),
.Y(n_3324)
);

OAI22xp5_ASAP7_75t_L g3325 ( 
.A1(n_2367),
.A2(n_2466),
.B1(n_2467),
.B2(n_2421),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_L g3326 ( 
.A(n_2512),
.B(n_2523),
.Y(n_3326)
);

A2O1A1Ixp33_ASAP7_75t_L g3327 ( 
.A1(n_2542),
.A2(n_2608),
.B(n_2610),
.C(n_2597),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_2364),
.Y(n_3328)
);

OA21x2_ASAP7_75t_L g3329 ( 
.A1(n_2168),
.A2(n_2222),
.B(n_2166),
.Y(n_3329)
);

INVx11_ASAP7_75t_L g3330 ( 
.A(n_2177),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_2375),
.Y(n_3331)
);

AOI21xp5_ASAP7_75t_L g3332 ( 
.A1(n_2099),
.A2(n_2860),
.B(n_2128),
.Y(n_3332)
);

NOR2xp33_ASAP7_75t_L g3333 ( 
.A(n_2597),
.B(n_2608),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_SL g3334 ( 
.A(n_2095),
.B(n_2123),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_L g3335 ( 
.A(n_2524),
.B(n_2525),
.Y(n_3335)
);

AOI21xp5_ASAP7_75t_L g3336 ( 
.A1(n_2490),
.A2(n_2845),
.B(n_2594),
.Y(n_3336)
);

BUFx12f_ASAP7_75t_L g3337 ( 
.A(n_2409),
.Y(n_3337)
);

AOI21xp5_ASAP7_75t_L g3338 ( 
.A1(n_2852),
.A2(n_2976),
.B(n_2911),
.Y(n_3338)
);

AOI21xp5_ASAP7_75t_L g3339 ( 
.A1(n_3065),
.A2(n_3107),
.B(n_3155),
.Y(n_3339)
);

OAI21xp33_ASAP7_75t_L g3340 ( 
.A1(n_2610),
.A2(n_2630),
.B(n_2627),
.Y(n_3340)
);

BUFx8_ASAP7_75t_SL g3341 ( 
.A(n_2308),
.Y(n_3341)
);

INVx1_ASAP7_75t_SL g3342 ( 
.A(n_3100),
.Y(n_3342)
);

INVx1_ASAP7_75t_SL g3343 ( 
.A(n_3100),
.Y(n_3343)
);

AOI22xp5_ASAP7_75t_L g3344 ( 
.A1(n_2627),
.A2(n_2634),
.B1(n_2651),
.B2(n_2630),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_L g3345 ( 
.A(n_2531),
.B(n_2533),
.Y(n_3345)
);

OAI21xp5_ASAP7_75t_L g3346 ( 
.A1(n_2634),
.A2(n_2652),
.B(n_2651),
.Y(n_3346)
);

NOR2x1_ASAP7_75t_L g3347 ( 
.A(n_2132),
.B(n_2191),
.Y(n_3347)
);

INVx1_ASAP7_75t_L g3348 ( 
.A(n_2385),
.Y(n_3348)
);

O2A1O1Ixp5_ASAP7_75t_L g3349 ( 
.A1(n_2652),
.A2(n_2694),
.B(n_2727),
.C(n_2698),
.Y(n_3349)
);

AO21x1_ASAP7_75t_L g3350 ( 
.A1(n_2168),
.A2(n_2698),
.B(n_2694),
.Y(n_3350)
);

INVx2_ASAP7_75t_L g3351 ( 
.A(n_2388),
.Y(n_3351)
);

AOI21xp5_ASAP7_75t_L g3352 ( 
.A1(n_2372),
.A2(n_2380),
.B(n_2378),
.Y(n_3352)
);

AOI21x1_ASAP7_75t_L g3353 ( 
.A1(n_2282),
.A2(n_2303),
.B(n_2079),
.Y(n_3353)
);

NOR2xp33_ASAP7_75t_L g3354 ( 
.A(n_2727),
.B(n_2742),
.Y(n_3354)
);

AND2x2_ASAP7_75t_L g3355 ( 
.A(n_2120),
.B(n_2166),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_2536),
.B(n_2537),
.Y(n_3356)
);

AOI21xp5_ASAP7_75t_L g3357 ( 
.A1(n_2397),
.A2(n_2404),
.B(n_2400),
.Y(n_3357)
);

NOR2xp33_ASAP7_75t_L g3358 ( 
.A(n_2742),
.B(n_2746),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_2551),
.B(n_2553),
.Y(n_3359)
);

OAI22xp5_ASAP7_75t_L g3360 ( 
.A1(n_3151),
.A2(n_2467),
.B1(n_2486),
.B2(n_2367),
.Y(n_3360)
);

AOI22xp33_ASAP7_75t_L g3361 ( 
.A1(n_2746),
.A2(n_2764),
.B1(n_2773),
.B2(n_2754),
.Y(n_3361)
);

OAI21xp5_ASAP7_75t_L g3362 ( 
.A1(n_2754),
.A2(n_2773),
.B(n_2764),
.Y(n_3362)
);

A2O1A1Ixp33_ASAP7_75t_L g3363 ( 
.A1(n_2778),
.A2(n_2793),
.B(n_2804),
.C(n_2787),
.Y(n_3363)
);

AND2x4_ASAP7_75t_SL g3364 ( 
.A(n_2028),
.B(n_2817),
.Y(n_3364)
);

NOR2x1_ASAP7_75t_L g3365 ( 
.A(n_2071),
.B(n_2074),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_L g3366 ( 
.A(n_2556),
.B(n_2565),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_2401),
.Y(n_3367)
);

O2A1O1Ixp33_ASAP7_75t_L g3368 ( 
.A1(n_2778),
.A2(n_2793),
.B(n_2804),
.C(n_2787),
.Y(n_3368)
);

OAI22xp5_ASAP7_75t_L g3369 ( 
.A1(n_3151),
.A2(n_2505),
.B1(n_2561),
.B2(n_2486),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_L g3370 ( 
.A(n_2567),
.B(n_2575),
.Y(n_3370)
);

A2O1A1Ixp33_ASAP7_75t_L g3371 ( 
.A1(n_2823),
.A2(n_2869),
.B(n_2870),
.C(n_2844),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_SL g3372 ( 
.A(n_2095),
.B(n_2124),
.Y(n_3372)
);

NOR3xp33_ASAP7_75t_L g3373 ( 
.A(n_2823),
.B(n_2869),
.C(n_2844),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_2579),
.B(n_2582),
.Y(n_3374)
);

AND2x2_ASAP7_75t_L g3375 ( 
.A(n_2870),
.B(n_2880),
.Y(n_3375)
);

NOR2xp67_ASAP7_75t_L g3376 ( 
.A(n_2009),
.B(n_2743),
.Y(n_3376)
);

AOI22xp33_ASAP7_75t_L g3377 ( 
.A1(n_2880),
.A2(n_2919),
.B1(n_2931),
.B2(n_2888),
.Y(n_3377)
);

BUFx6f_ASAP7_75t_L g3378 ( 
.A(n_2583),
.Y(n_3378)
);

OAI21xp5_ASAP7_75t_L g3379 ( 
.A1(n_2888),
.A2(n_2931),
.B(n_2919),
.Y(n_3379)
);

NOR2xp33_ASAP7_75t_L g3380 ( 
.A(n_2933),
.B(n_2935),
.Y(n_3380)
);

AOI21xp5_ASAP7_75t_L g3381 ( 
.A1(n_2419),
.A2(n_2428),
.B(n_2427),
.Y(n_3381)
);

AOI21xp5_ASAP7_75t_L g3382 ( 
.A1(n_2439),
.A2(n_2510),
.B(n_2451),
.Y(n_3382)
);

OAI22xp5_ASAP7_75t_L g3383 ( 
.A1(n_2505),
.A2(n_2570),
.B1(n_2580),
.B2(n_2561),
.Y(n_3383)
);

AOI22xp5_ASAP7_75t_L g3384 ( 
.A1(n_2933),
.A2(n_2941),
.B1(n_2949),
.B2(n_2935),
.Y(n_3384)
);

NAND2xp33_ASAP7_75t_L g3385 ( 
.A(n_2570),
.B(n_2580),
.Y(n_3385)
);

BUFx8_ASAP7_75t_L g3386 ( 
.A(n_2125),
.Y(n_3386)
);

INVx2_ASAP7_75t_L g3387 ( 
.A(n_2414),
.Y(n_3387)
);

AO21x1_ASAP7_75t_L g3388 ( 
.A1(n_2941),
.A2(n_2951),
.B(n_2949),
.Y(n_3388)
);

A2O1A1Ixp33_ASAP7_75t_L g3389 ( 
.A1(n_2951),
.A2(n_2984),
.B(n_2985),
.C(n_2954),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_2584),
.B(n_2601),
.Y(n_3390)
);

AOI21xp33_ASAP7_75t_L g3391 ( 
.A1(n_2954),
.A2(n_2985),
.B(n_2984),
.Y(n_3391)
);

A2O1A1Ixp33_ASAP7_75t_L g3392 ( 
.A1(n_2989),
.A2(n_3022),
.B(n_3039),
.C(n_2997),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_SL g3393 ( 
.A(n_2161),
.B(n_2119),
.Y(n_3393)
);

AOI21xp5_ASAP7_75t_L g3394 ( 
.A1(n_2514),
.A2(n_2917),
.B(n_2910),
.Y(n_3394)
);

OAI21xp5_ASAP7_75t_L g3395 ( 
.A1(n_2989),
.A2(n_3022),
.B(n_2997),
.Y(n_3395)
);

AOI21xp5_ASAP7_75t_L g3396 ( 
.A1(n_2920),
.A2(n_2943),
.B(n_2937),
.Y(n_3396)
);

AOI21xp5_ASAP7_75t_L g3397 ( 
.A1(n_2944),
.A2(n_2959),
.B(n_2952),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_2425),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_2603),
.B(n_2605),
.Y(n_3399)
);

OAI21xp33_ASAP7_75t_L g3400 ( 
.A1(n_3039),
.A2(n_3060),
.B(n_3056),
.Y(n_3400)
);

AOI21xp5_ASAP7_75t_L g3401 ( 
.A1(n_2968),
.A2(n_2991),
.B(n_2986),
.Y(n_3401)
);

CKINVDCx8_ASAP7_75t_R g3402 ( 
.A(n_2173),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_2607),
.B(n_2611),
.Y(n_3403)
);

AOI21xp5_ASAP7_75t_L g3404 ( 
.A1(n_3038),
.A2(n_3121),
.B(n_3041),
.Y(n_3404)
);

AND2x2_ASAP7_75t_SL g3405 ( 
.A(n_2596),
.B(n_2616),
.Y(n_3405)
);

AOI21xp5_ASAP7_75t_L g3406 ( 
.A1(n_2204),
.A2(n_2206),
.B(n_2205),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_2617),
.B(n_2620),
.Y(n_3407)
);

BUFx6f_ASAP7_75t_L g3408 ( 
.A(n_2767),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_2621),
.B(n_2622),
.Y(n_3409)
);

AOI21xp5_ASAP7_75t_L g3410 ( 
.A1(n_2187),
.A2(n_2200),
.B(n_2186),
.Y(n_3410)
);

NOR2xp67_ASAP7_75t_L g3411 ( 
.A(n_2009),
.B(n_2743),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_2434),
.Y(n_3412)
);

NOR2xp33_ASAP7_75t_L g3413 ( 
.A(n_3056),
.B(n_3060),
.Y(n_3413)
);

AOI21xp5_ASAP7_75t_L g3414 ( 
.A1(n_2126),
.A2(n_2282),
.B(n_2001),
.Y(n_3414)
);

NOR2x1p5_ASAP7_75t_L g3415 ( 
.A(n_2353),
.B(n_2090),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_L g3416 ( 
.A(n_2624),
.B(n_2626),
.Y(n_3416)
);

AOI21xp5_ASAP7_75t_L g3417 ( 
.A1(n_1991),
.A2(n_2011),
.B(n_2008),
.Y(n_3417)
);

AOI22xp5_ASAP7_75t_L g3418 ( 
.A1(n_3074),
.A2(n_3088),
.B1(n_3104),
.B2(n_3078),
.Y(n_3418)
);

NOR2x1_ASAP7_75t_L g3419 ( 
.A(n_2331),
.B(n_2335),
.Y(n_3419)
);

O2A1O1Ixp33_ASAP7_75t_L g3420 ( 
.A1(n_3074),
.A2(n_3088),
.B(n_3104),
.C(n_3078),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_2444),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_L g3422 ( 
.A(n_2636),
.B(n_2638),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_L g3423 ( 
.A(n_2640),
.B(n_2641),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_L g3424 ( 
.A(n_2643),
.B(n_2644),
.Y(n_3424)
);

AND2x2_ASAP7_75t_SL g3425 ( 
.A(n_2596),
.B(n_2616),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_2450),
.Y(n_3426)
);

AOI21xp33_ASAP7_75t_L g3427 ( 
.A1(n_3117),
.A2(n_3128),
.B(n_2655),
.Y(n_3427)
);

NOR2xp33_ASAP7_75t_L g3428 ( 
.A(n_3117),
.B(n_3128),
.Y(n_3428)
);

INVx5_ASAP7_75t_L g3429 ( 
.A(n_2743),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_2457),
.Y(n_3430)
);

BUFx4f_ASAP7_75t_L g3431 ( 
.A(n_2566),
.Y(n_3431)
);

OAI321xp33_ASAP7_75t_L g3432 ( 
.A1(n_2628),
.A2(n_2677),
.A3(n_2686),
.B1(n_2707),
.B2(n_2699),
.C(n_2655),
.Y(n_3432)
);

AOI22xp5_ASAP7_75t_L g3433 ( 
.A1(n_2628),
.A2(n_2686),
.B1(n_2699),
.B2(n_2677),
.Y(n_3433)
);

CKINVDCx5p33_ASAP7_75t_R g3434 ( 
.A(n_2172),
.Y(n_3434)
);

AND2x2_ASAP7_75t_L g3435 ( 
.A(n_2010),
.B(n_3016),
.Y(n_3435)
);

A2O1A1Ixp33_ASAP7_75t_L g3436 ( 
.A1(n_2707),
.A2(n_2711),
.B(n_2728),
.C(n_2718),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_2647),
.B(n_2653),
.Y(n_3437)
);

AOI21x1_ASAP7_75t_L g3438 ( 
.A1(n_2303),
.A2(n_2188),
.B(n_2185),
.Y(n_3438)
);

OAI21xp5_ASAP7_75t_L g3439 ( 
.A1(n_2711),
.A2(n_2728),
.B(n_2718),
.Y(n_3439)
);

AOI21xp5_ASAP7_75t_L g3440 ( 
.A1(n_2012),
.A2(n_2015),
.B(n_2014),
.Y(n_3440)
);

BUFx4f_ASAP7_75t_L g3441 ( 
.A(n_2566),
.Y(n_3441)
);

AOI21xp5_ASAP7_75t_L g3442 ( 
.A1(n_2018),
.A2(n_2026),
.B(n_2022),
.Y(n_3442)
);

OAI22xp5_ASAP7_75t_L g3443 ( 
.A1(n_2763),
.A2(n_2814),
.B1(n_2816),
.B2(n_2806),
.Y(n_3443)
);

OAI22xp5_ASAP7_75t_L g3444 ( 
.A1(n_2763),
.A2(n_2814),
.B1(n_2816),
.B2(n_2806),
.Y(n_3444)
);

OAI21xp5_ASAP7_75t_L g3445 ( 
.A1(n_2848),
.A2(n_2881),
.B(n_2872),
.Y(n_3445)
);

OAI22xp5_ASAP7_75t_L g3446 ( 
.A1(n_2848),
.A2(n_2881),
.B1(n_2887),
.B2(n_2872),
.Y(n_3446)
);

INVx1_ASAP7_75t_SL g3447 ( 
.A(n_3125),
.Y(n_3447)
);

AOI21xp5_ASAP7_75t_L g3448 ( 
.A1(n_2036),
.A2(n_2041),
.B(n_2039),
.Y(n_3448)
);

HB1xp67_ASAP7_75t_L g3449 ( 
.A(n_3125),
.Y(n_3449)
);

AOI21x1_ASAP7_75t_L g3450 ( 
.A1(n_2185),
.A2(n_2192),
.B(n_2188),
.Y(n_3450)
);

AOI21xp5_ASAP7_75t_L g3451 ( 
.A1(n_2042),
.A2(n_2051),
.B(n_2046),
.Y(n_3451)
);

AOI21xp5_ASAP7_75t_L g3452 ( 
.A1(n_2052),
.A2(n_2061),
.B(n_2053),
.Y(n_3452)
);

AOI21xp5_ASAP7_75t_L g3453 ( 
.A1(n_2063),
.A2(n_2070),
.B(n_2067),
.Y(n_3453)
);

OAI22xp5_ASAP7_75t_L g3454 ( 
.A1(n_2887),
.A2(n_2930),
.B1(n_2945),
.B2(n_2923),
.Y(n_3454)
);

BUFx4f_ASAP7_75t_L g3455 ( 
.A(n_2566),
.Y(n_3455)
);

NOR3xp33_ASAP7_75t_L g3456 ( 
.A(n_3142),
.B(n_3146),
.C(n_3143),
.Y(n_3456)
);

INVx1_ASAP7_75t_SL g3457 ( 
.A(n_1992),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_2476),
.Y(n_3458)
);

A2O1A1Ixp33_ASAP7_75t_L g3459 ( 
.A1(n_2923),
.A2(n_2945),
.B(n_2961),
.C(n_2930),
.Y(n_3459)
);

NAND2xp5_ASAP7_75t_L g3460 ( 
.A(n_2961),
.B(n_2972),
.Y(n_3460)
);

BUFx6f_ASAP7_75t_L g3461 ( 
.A(n_2874),
.Y(n_3461)
);

AOI21xp5_ASAP7_75t_L g3462 ( 
.A1(n_2073),
.A2(n_2077),
.B(n_2076),
.Y(n_3462)
);

INVx2_ASAP7_75t_L g3463 ( 
.A(n_2494),
.Y(n_3463)
);

OAI22xp5_ASAP7_75t_L g3464 ( 
.A1(n_2972),
.A2(n_2981),
.B1(n_3028),
.B2(n_2978),
.Y(n_3464)
);

AOI21xp5_ASAP7_75t_L g3465 ( 
.A1(n_2080),
.A2(n_2086),
.B(n_2085),
.Y(n_3465)
);

NAND2xp33_ASAP7_75t_L g3466 ( 
.A(n_2978),
.B(n_2981),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_L g3467 ( 
.A(n_3028),
.B(n_3047),
.Y(n_3467)
);

OAI21xp33_ASAP7_75t_L g3468 ( 
.A1(n_3047),
.A2(n_3098),
.B(n_3066),
.Y(n_3468)
);

OR2x2_ASAP7_75t_L g3469 ( 
.A(n_2391),
.B(n_2615),
.Y(n_3469)
);

AOI21xp5_ASAP7_75t_L g3470 ( 
.A1(n_2089),
.A2(n_2104),
.B(n_2102),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_SL g3471 ( 
.A(n_3066),
.B(n_3098),
.Y(n_3471)
);

AOI21xp5_ASAP7_75t_L g3472 ( 
.A1(n_2105),
.A2(n_2110),
.B(n_2106),
.Y(n_3472)
);

AOI21x1_ASAP7_75t_L g3473 ( 
.A1(n_2192),
.A2(n_2195),
.B(n_2194),
.Y(n_3473)
);

A2O1A1Ixp33_ASAP7_75t_L g3474 ( 
.A1(n_3101),
.A2(n_3135),
.B(n_2096),
.C(n_2010),
.Y(n_3474)
);

OAI21xp5_ASAP7_75t_L g3475 ( 
.A1(n_3101),
.A2(n_3135),
.B(n_2096),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_2498),
.Y(n_3476)
);

NOR2x1_ASAP7_75t_L g3477 ( 
.A(n_2194),
.B(n_2195),
.Y(n_3477)
);

INVx2_ASAP7_75t_L g3478 ( 
.A(n_2519),
.Y(n_3478)
);

OAI21xp5_ASAP7_75t_L g3479 ( 
.A1(n_2228),
.A2(n_2117),
.B(n_2658),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_L g3480 ( 
.A(n_2654),
.B(n_2661),
.Y(n_3480)
);

BUFx6f_ASAP7_75t_L g3481 ( 
.A(n_2874),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_2663),
.B(n_2664),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_2534),
.Y(n_3483)
);

A2O1A1Ixp33_ASAP7_75t_L g3484 ( 
.A1(n_2665),
.A2(n_2671),
.B(n_2674),
.C(n_2667),
.Y(n_3484)
);

INVx3_ASAP7_75t_L g3485 ( 
.A(n_2614),
.Y(n_3485)
);

AOI21xp5_ASAP7_75t_L g3486 ( 
.A1(n_2236),
.A2(n_2183),
.B(n_2176),
.Y(n_3486)
);

NOR2xp67_ASAP7_75t_L g3487 ( 
.A(n_2874),
.B(n_3021),
.Y(n_3487)
);

INVx3_ASAP7_75t_L g3488 ( 
.A(n_2614),
.Y(n_3488)
);

NOR2xp33_ASAP7_75t_L g3489 ( 
.A(n_2084),
.B(n_2678),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_L g3490 ( 
.A(n_2684),
.B(n_2690),
.Y(n_3490)
);

AOI21xp5_ASAP7_75t_L g3491 ( 
.A1(n_2236),
.A2(n_2264),
.B(n_2210),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_SL g3492 ( 
.A(n_2249),
.B(n_2000),
.Y(n_3492)
);

NOR2x1_ASAP7_75t_L g3493 ( 
.A(n_2210),
.B(n_2264),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_L g3494 ( 
.A(n_2697),
.B(n_2705),
.Y(n_3494)
);

OAI321xp33_ASAP7_75t_L g3495 ( 
.A1(n_3140),
.A2(n_3148),
.A3(n_2710),
.B1(n_2722),
.B2(n_2731),
.C(n_2723),
.Y(n_3495)
);

AOI21xp5_ASAP7_75t_L g3496 ( 
.A1(n_2266),
.A2(n_2280),
.B(n_2275),
.Y(n_3496)
);

AOI22xp5_ASAP7_75t_L g3497 ( 
.A1(n_2717),
.A2(n_2735),
.B1(n_2745),
.B2(n_2734),
.Y(n_3497)
);

NAND2x1p5_ASAP7_75t_L g3498 ( 
.A(n_2874),
.B(n_3021),
.Y(n_3498)
);

INVx1_ASAP7_75t_L g3499 ( 
.A(n_2540),
.Y(n_3499)
);

AOI22xp33_ASAP7_75t_L g3500 ( 
.A1(n_2069),
.A2(n_2169),
.B1(n_2751),
.B2(n_2750),
.Y(n_3500)
);

AOI21xp5_ASAP7_75t_L g3501 ( 
.A1(n_2266),
.A2(n_2280),
.B(n_2275),
.Y(n_3501)
);

OR2x2_ASAP7_75t_L g3502 ( 
.A(n_2642),
.B(n_2680),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_2753),
.B(n_2757),
.Y(n_3503)
);

AOI21xp5_ASAP7_75t_L g3504 ( 
.A1(n_3021),
.A2(n_3113),
.B(n_2230),
.Y(n_3504)
);

NOR3xp33_ASAP7_75t_L g3505 ( 
.A(n_2761),
.B(n_2769),
.C(n_2762),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_SL g3506 ( 
.A(n_2107),
.B(n_2065),
.Y(n_3506)
);

AOI21xp5_ASAP7_75t_L g3507 ( 
.A1(n_3021),
.A2(n_3113),
.B(n_2230),
.Y(n_3507)
);

NOR2xp33_ASAP7_75t_L g3508 ( 
.A(n_2785),
.B(n_2790),
.Y(n_3508)
);

OAI22xp5_ASAP7_75t_L g3509 ( 
.A1(n_2791),
.A2(n_2794),
.B1(n_2805),
.B2(n_2799),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_2572),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_2813),
.B(n_2819),
.Y(n_3511)
);

AOI21x1_ASAP7_75t_L g3512 ( 
.A1(n_2169),
.A2(n_2313),
.B(n_2284),
.Y(n_3512)
);

NOR2xp33_ASAP7_75t_SL g3513 ( 
.A(n_3113),
.B(n_2480),
.Y(n_3513)
);

INVx2_ASAP7_75t_L g3514 ( 
.A(n_2573),
.Y(n_3514)
);

AOI21xp5_ASAP7_75t_L g3515 ( 
.A1(n_3113),
.A2(n_2208),
.B(n_2822),
.Y(n_3515)
);

O2A1O1Ixp33_ASAP7_75t_L g3516 ( 
.A1(n_2825),
.A2(n_2830),
.B(n_2835),
.C(n_2831),
.Y(n_3516)
);

AND2x4_ASAP7_75t_L g3517 ( 
.A(n_2028),
.B(n_2817),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_L g3518 ( 
.A(n_2837),
.B(n_2841),
.Y(n_3518)
);

NOR2xp33_ASAP7_75t_L g3519 ( 
.A(n_2846),
.B(n_2850),
.Y(n_3519)
);

NOR2xp67_ASAP7_75t_L g3520 ( 
.A(n_2270),
.B(n_2309),
.Y(n_3520)
);

AND2x2_ASAP7_75t_SL g3521 ( 
.A(n_2854),
.B(n_2855),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_SL g3522 ( 
.A(n_2279),
.B(n_2068),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_L g3523 ( 
.A(n_2873),
.B(n_2877),
.Y(n_3523)
);

NAND3xp33_ASAP7_75t_L g3524 ( 
.A(n_2882),
.B(n_2896),
.C(n_2886),
.Y(n_3524)
);

AND2x2_ASAP7_75t_L g3525 ( 
.A(n_2122),
.B(n_1990),
.Y(n_3525)
);

INVxp67_ASAP7_75t_L g3526 ( 
.A(n_2212),
.Y(n_3526)
);

INVx1_ASAP7_75t_L g3527 ( 
.A(n_2581),
.Y(n_3527)
);

AOI21xp5_ASAP7_75t_L g3528 ( 
.A1(n_2899),
.A2(n_2903),
.B(n_2901),
.Y(n_3528)
);

AOI21x1_ASAP7_75t_L g3529 ( 
.A1(n_2313),
.A2(n_2314),
.B(n_2322),
.Y(n_3529)
);

AOI22xp5_ASAP7_75t_L g3530 ( 
.A1(n_2908),
.A2(n_2918),
.B1(n_2925),
.B2(n_2914),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_SL g3531 ( 
.A(n_2932),
.B(n_2934),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_L g3532 ( 
.A(n_2942),
.B(n_2948),
.Y(n_3532)
);

AOI21xp5_ASAP7_75t_L g3533 ( 
.A1(n_2962),
.A2(n_2966),
.B(n_2965),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_L g3534 ( 
.A(n_2970),
.B(n_2971),
.Y(n_3534)
);

AND2x4_ASAP7_75t_L g3535 ( 
.A(n_2834),
.B(n_3002),
.Y(n_3535)
);

BUFx3_ASAP7_75t_L g3536 ( 
.A(n_2719),
.Y(n_3536)
);

AND2x4_ASAP7_75t_L g3537 ( 
.A(n_2834),
.B(n_3002),
.Y(n_3537)
);

OAI22xp5_ASAP7_75t_L g3538 ( 
.A1(n_2975),
.A2(n_2979),
.B1(n_2993),
.B2(n_2992),
.Y(n_3538)
);

INVx2_ASAP7_75t_L g3539 ( 
.A(n_2593),
.Y(n_3539)
);

NAND2xp5_ASAP7_75t_L g3540 ( 
.A(n_3000),
.B(n_3005),
.Y(n_3540)
);

BUFx6f_ASAP7_75t_L g3541 ( 
.A(n_2566),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3006),
.B(n_3007),
.Y(n_3542)
);

AND2x2_ASAP7_75t_L g3543 ( 
.A(n_2023),
.B(n_2049),
.Y(n_3543)
);

OAI21xp33_ASAP7_75t_L g3544 ( 
.A1(n_3010),
.A2(n_3019),
.B(n_3013),
.Y(n_3544)
);

AOI21xp5_ASAP7_75t_L g3545 ( 
.A1(n_3023),
.A2(n_3033),
.B(n_3026),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_2599),
.Y(n_3546)
);

AOI21xp5_ASAP7_75t_L g3547 ( 
.A1(n_3035),
.A2(n_3043),
.B(n_3037),
.Y(n_3547)
);

AND2x2_ASAP7_75t_L g3548 ( 
.A(n_2062),
.B(n_2268),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_SL g3549 ( 
.A(n_3059),
.B(n_3061),
.Y(n_3549)
);

NOR2xp33_ASAP7_75t_L g3550 ( 
.A(n_3070),
.B(n_3071),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_SL g3551 ( 
.A(n_3072),
.B(n_3080),
.Y(n_3551)
);

AOI21xp5_ASAP7_75t_L g3552 ( 
.A1(n_3084),
.A2(n_3091),
.B(n_3085),
.Y(n_3552)
);

AOI21xp5_ASAP7_75t_L g3553 ( 
.A1(n_3095),
.A2(n_3105),
.B(n_3096),
.Y(n_3553)
);

AOI21xp5_ASAP7_75t_L g3554 ( 
.A1(n_3119),
.A2(n_3124),
.B(n_3123),
.Y(n_3554)
);

O2A1O1Ixp33_ASAP7_75t_L g3555 ( 
.A1(n_3136),
.A2(n_3139),
.B(n_3137),
.C(n_2360),
.Y(n_3555)
);

NOR2xp33_ASAP7_75t_SL g3556 ( 
.A(n_3097),
.B(n_2219),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_L g3557 ( 
.A(n_2184),
.B(n_2977),
.Y(n_3557)
);

OAI22xp5_ASAP7_75t_L g3558 ( 
.A1(n_2756),
.A2(n_2866),
.B1(n_2939),
.B2(n_2811),
.Y(n_3558)
);

BUFx6f_ASAP7_75t_L g3559 ( 
.A(n_2977),
.Y(n_3559)
);

INVx2_ASAP7_75t_L g3560 ( 
.A(n_2609),
.Y(n_3560)
);

BUFx6f_ASAP7_75t_L g3561 ( 
.A(n_2977),
.Y(n_3561)
);

NOR2x1_ASAP7_75t_L g3562 ( 
.A(n_2294),
.B(n_3054),
.Y(n_3562)
);

AOI21x1_ASAP7_75t_L g3563 ( 
.A1(n_2261),
.A2(n_2639),
.B(n_2619),
.Y(n_3563)
);

AOI21x1_ASAP7_75t_L g3564 ( 
.A1(n_2645),
.A2(n_2657),
.B(n_2648),
.Y(n_3564)
);

AOI21xp5_ASAP7_75t_L g3565 ( 
.A1(n_2294),
.A2(n_2262),
.B(n_2258),
.Y(n_3565)
);

AND2x2_ASAP7_75t_L g3566 ( 
.A(n_2396),
.B(n_2436),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_2977),
.B(n_3112),
.Y(n_3567)
);

BUFx6f_ASAP7_75t_L g3568 ( 
.A(n_2977),
.Y(n_3568)
);

OR2x2_ASAP7_75t_L g3569 ( 
.A(n_3030),
.B(n_3106),
.Y(n_3569)
);

NOR2xp33_ASAP7_75t_SL g3570 ( 
.A(n_2441),
.B(n_2020),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_SL g3571 ( 
.A(n_2066),
.B(n_2082),
.Y(n_3571)
);

NOR2xp33_ASAP7_75t_L g3572 ( 
.A(n_2368),
.B(n_2481),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3112),
.B(n_2083),
.Y(n_3573)
);

AOI21xp5_ASAP7_75t_L g3574 ( 
.A1(n_2262),
.A2(n_2258),
.B(n_2213),
.Y(n_3574)
);

AOI22xp33_ASAP7_75t_L g3575 ( 
.A1(n_2164),
.A2(n_2178),
.B1(n_2170),
.B2(n_3112),
.Y(n_3575)
);

AOI22xp5_ASAP7_75t_L g3576 ( 
.A1(n_2459),
.A2(n_2491),
.B1(n_2504),
.B2(n_2499),
.Y(n_3576)
);

NOR2xp33_ASAP7_75t_L g3577 ( 
.A(n_2625),
.B(n_2836),
.Y(n_3577)
);

AOI22xp5_ASAP7_75t_L g3578 ( 
.A1(n_2520),
.A2(n_2527),
.B1(n_2552),
.B2(n_2532),
.Y(n_3578)
);

AOI21xp5_ASAP7_75t_L g3579 ( 
.A1(n_2209),
.A2(n_2224),
.B(n_2220),
.Y(n_3579)
);

AOI21x1_ASAP7_75t_L g3580 ( 
.A1(n_2672),
.A2(n_2689),
.B(n_2685),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_3112),
.B(n_2691),
.Y(n_3581)
);

NOR2x1p5_ASAP7_75t_L g3582 ( 
.A(n_3054),
.B(n_1999),
.Y(n_3582)
);

AND2x4_ASAP7_75t_L g3583 ( 
.A(n_3112),
.B(n_2037),
.Y(n_3583)
);

INVxp67_ASAP7_75t_L g3584 ( 
.A(n_2212),
.Y(n_3584)
);

AOI21xp5_ASAP7_75t_L g3585 ( 
.A1(n_2231),
.A2(n_2243),
.B(n_2241),
.Y(n_3585)
);

A2O1A1Ixp33_ASAP7_75t_L g3586 ( 
.A1(n_2269),
.A2(n_2336),
.B(n_2276),
.C(n_2318),
.Y(n_3586)
);

AOI22xp5_ASAP7_75t_L g3587 ( 
.A1(n_2564),
.A2(n_2633),
.B1(n_2716),
.B2(n_2666),
.Y(n_3587)
);

AOI21xp5_ASAP7_75t_L g3588 ( 
.A1(n_2247),
.A2(n_2260),
.B(n_2257),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_SL g3589 ( 
.A(n_2189),
.B(n_2225),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_SL g3590 ( 
.A(n_2936),
.B(n_2988),
.Y(n_3590)
);

AOI21xp5_ASAP7_75t_L g3591 ( 
.A1(n_2269),
.A2(n_2311),
.B(n_2190),
.Y(n_3591)
);

AOI21xp5_ASAP7_75t_L g3592 ( 
.A1(n_2190),
.A2(n_2199),
.B(n_2193),
.Y(n_3592)
);

AND2x4_ASAP7_75t_L g3593 ( 
.A(n_2037),
.B(n_2196),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_2692),
.Y(n_3594)
);

AND2x4_ASAP7_75t_L g3595 ( 
.A(n_2196),
.B(n_2245),
.Y(n_3595)
);

O2A1O1Ixp33_ASAP7_75t_L g3596 ( 
.A1(n_3073),
.A2(n_2129),
.B(n_2361),
.C(n_2336),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_L g3597 ( 
.A(n_2696),
.B(n_2700),
.Y(n_3597)
);

AND2x4_ASAP7_75t_L g3598 ( 
.A(n_2245),
.B(n_2273),
.Y(n_3598)
);

INVx2_ASAP7_75t_L g3599 ( 
.A(n_2704),
.Y(n_3599)
);

OAI22xp5_ASAP7_75t_L g3600 ( 
.A1(n_2193),
.A2(n_2199),
.B1(n_2259),
.B2(n_2214),
.Y(n_3600)
);

OAI21xp5_ASAP7_75t_L g3601 ( 
.A1(n_2290),
.A2(n_2316),
.B(n_2276),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_L g3602 ( 
.A(n_2720),
.B(n_2726),
.Y(n_3602)
);

AOI21xp5_ASAP7_75t_L g3603 ( 
.A1(n_2214),
.A2(n_2259),
.B(n_2631),
.Y(n_3603)
);

O2A1O1Ixp33_ASAP7_75t_L g3604 ( 
.A1(n_2129),
.A2(n_2631),
.B(n_2938),
.C(n_2660),
.Y(n_3604)
);

AOI21xp5_ASAP7_75t_L g3605 ( 
.A1(n_2660),
.A2(n_2938),
.B(n_2318),
.Y(n_3605)
);

NOR2x2_ASAP7_75t_L g3606 ( 
.A(n_2333),
.B(n_2351),
.Y(n_3606)
);

OAI21xp5_ASAP7_75t_L g3607 ( 
.A1(n_2290),
.A2(n_2316),
.B(n_2274),
.Y(n_3607)
);

AOI21xp5_ASAP7_75t_L g3608 ( 
.A1(n_2274),
.A2(n_2319),
.B(n_2007),
.Y(n_3608)
);

O2A1O1Ixp5_ASAP7_75t_L g3609 ( 
.A1(n_1999),
.A2(n_2912),
.B(n_2995),
.C(n_2898),
.Y(n_3609)
);

OAI21xp33_ASAP7_75t_L g3610 ( 
.A1(n_2724),
.A2(n_2736),
.B(n_2732),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_2733),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_L g3612 ( 
.A(n_2740),
.B(n_2747),
.Y(n_3612)
);

AOI21xp5_ASAP7_75t_L g3613 ( 
.A1(n_2319),
.A2(n_2029),
.B(n_1994),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_L g3614 ( 
.A(n_2755),
.B(n_2758),
.Y(n_3614)
);

OAI22xp5_ASAP7_75t_L g3615 ( 
.A1(n_2771),
.A2(n_2781),
.B1(n_2782),
.B2(n_2779),
.Y(n_3615)
);

INVx11_ASAP7_75t_L g3616 ( 
.A(n_2409),
.Y(n_3616)
);

AOI21xp5_ASAP7_75t_L g3617 ( 
.A1(n_2034),
.A2(n_2048),
.B(n_2040),
.Y(n_3617)
);

NAND3xp33_ASAP7_75t_L g3618 ( 
.A(n_2164),
.B(n_2178),
.C(n_2170),
.Y(n_3618)
);

AND2x2_ASAP7_75t_L g3619 ( 
.A(n_2744),
.B(n_2752),
.Y(n_3619)
);

INVx2_ASAP7_75t_L g3620 ( 
.A(n_2796),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_2807),
.B(n_2808),
.Y(n_3621)
);

AOI21xp5_ASAP7_75t_L g3622 ( 
.A1(n_2056),
.A2(n_2064),
.B(n_2057),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_2809),
.Y(n_3623)
);

BUFx6f_ASAP7_75t_L g3624 ( 
.A(n_2898),
.Y(n_3624)
);

OAI321xp33_ASAP7_75t_L g3625 ( 
.A1(n_2341),
.A2(n_2955),
.A3(n_2810),
.B1(n_3138),
.B2(n_2768),
.C(n_2292),
.Y(n_3625)
);

AOI21xp5_ASAP7_75t_L g3626 ( 
.A1(n_2100),
.A2(n_2109),
.B(n_2103),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_2815),
.B(n_2820),
.Y(n_3627)
);

NOR2xp67_ASAP7_75t_L g3628 ( 
.A(n_2285),
.B(n_2296),
.Y(n_3628)
);

OAI21xp5_ASAP7_75t_L g3629 ( 
.A1(n_2298),
.A2(n_2300),
.B(n_2299),
.Y(n_3629)
);

AOI21xp5_ASAP7_75t_L g3630 ( 
.A1(n_2114),
.A2(n_2131),
.B(n_2130),
.Y(n_3630)
);

NAND2xp5_ASAP7_75t_L g3631 ( 
.A(n_2842),
.B(n_2847),
.Y(n_3631)
);

CKINVDCx6p67_ASAP7_75t_R g3632 ( 
.A(n_2159),
.Y(n_3632)
);

BUFx2_ASAP7_75t_L g3633 ( 
.A(n_3152),
.Y(n_3633)
);

AOI22xp33_ASAP7_75t_L g3634 ( 
.A1(n_2912),
.A2(n_3018),
.B1(n_3020),
.B2(n_2995),
.Y(n_3634)
);

NAND2xp5_ASAP7_75t_L g3635 ( 
.A(n_2862),
.B(n_2863),
.Y(n_3635)
);

O2A1O1Ixp5_ASAP7_75t_L g3636 ( 
.A1(n_3018),
.A2(n_3133),
.B(n_3020),
.C(n_2239),
.Y(n_3636)
);

AOI21xp33_ASAP7_75t_L g3637 ( 
.A1(n_2868),
.A2(n_2876),
.B(n_2871),
.Y(n_3637)
);

AOI21xp5_ASAP7_75t_L g3638 ( 
.A1(n_2134),
.A2(n_2157),
.B(n_2136),
.Y(n_3638)
);

OAI21xp5_ASAP7_75t_L g3639 ( 
.A1(n_2306),
.A2(n_2278),
.B(n_2272),
.Y(n_3639)
);

AOI21xp5_ASAP7_75t_L g3640 ( 
.A1(n_2158),
.A2(n_2181),
.B(n_2175),
.Y(n_3640)
);

HB1xp67_ASAP7_75t_L g3641 ( 
.A(n_2179),
.Y(n_3641)
);

OAI21xp5_ASAP7_75t_L g3642 ( 
.A1(n_2283),
.A2(n_2289),
.B(n_2287),
.Y(n_3642)
);

OAI21xp5_ASAP7_75t_L g3643 ( 
.A1(n_2291),
.A2(n_2301),
.B(n_2293),
.Y(n_3643)
);

AOI21xp5_ASAP7_75t_L g3644 ( 
.A1(n_2211),
.A2(n_2254),
.B(n_2218),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_L g3645 ( 
.A(n_2889),
.B(n_2905),
.Y(n_3645)
);

NAND2xp5_ASAP7_75t_L g3646 ( 
.A(n_2940),
.B(n_2957),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_L g3647 ( 
.A(n_2960),
.B(n_2969),
.Y(n_3647)
);

NAND2xp5_ASAP7_75t_L g3648 ( 
.A(n_2983),
.B(n_2987),
.Y(n_3648)
);

OAI22xp5_ASAP7_75t_L g3649 ( 
.A1(n_2998),
.A2(n_3012),
.B1(n_3017),
.B2(n_3004),
.Y(n_3649)
);

AOI21xp5_ASAP7_75t_L g3650 ( 
.A1(n_2255),
.A2(n_2406),
.B(n_2377),
.Y(n_3650)
);

NAND2xp5_ASAP7_75t_SL g3651 ( 
.A(n_2237),
.B(n_3133),
.Y(n_3651)
);

AND2x2_ASAP7_75t_L g3652 ( 
.A(n_2412),
.B(n_2438),
.Y(n_3652)
);

O2A1O1Ixp5_ASAP7_75t_L g3653 ( 
.A1(n_2320),
.A2(n_2238),
.B(n_2346),
.C(n_2324),
.Y(n_3653)
);

NOR2xp33_ASAP7_75t_SL g3654 ( 
.A(n_2441),
.B(n_2445),
.Y(n_3654)
);

NOR2xp33_ASAP7_75t_L g3655 ( 
.A(n_2202),
.B(n_2201),
.Y(n_3655)
);

OAI21xp33_ASAP7_75t_L g3656 ( 
.A1(n_3049),
.A2(n_2288),
.B(n_2217),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_3025),
.B(n_3027),
.Y(n_3657)
);

AOI21xp5_ASAP7_75t_L g3658 ( 
.A1(n_2440),
.A2(n_2449),
.B(n_2447),
.Y(n_3658)
);

A2O1A1Ixp33_ASAP7_75t_L g3659 ( 
.A1(n_2325),
.A2(n_2329),
.B(n_2327),
.C(n_2334),
.Y(n_3659)
);

OAI21xp5_ASAP7_75t_L g3660 ( 
.A1(n_2302),
.A2(n_2315),
.B(n_2321),
.Y(n_3660)
);

INVx2_ASAP7_75t_L g3661 ( 
.A(n_3050),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_SL g3662 ( 
.A(n_2111),
.B(n_2035),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_3063),
.B(n_3064),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_SL g3664 ( 
.A(n_2452),
.B(n_2585),
.Y(n_3664)
);

AOI21xp5_ASAP7_75t_L g3665 ( 
.A1(n_2460),
.A2(n_2472),
.B(n_2461),
.Y(n_3665)
);

INVx2_ASAP7_75t_L g3666 ( 
.A(n_3099),
.Y(n_3666)
);

OAI21xp5_ASAP7_75t_L g3667 ( 
.A1(n_3102),
.A2(n_3129),
.B(n_3109),
.Y(n_3667)
);

INVx4_ASAP7_75t_L g3668 ( 
.A(n_2614),
.Y(n_3668)
);

AOI221xp5_ASAP7_75t_SL g3669 ( 
.A1(n_2058),
.A2(n_3131),
.B1(n_2207),
.B2(n_2359),
.C(n_2650),
.Y(n_3669)
);

INVx2_ASAP7_75t_L g3670 ( 
.A(n_2473),
.Y(n_3670)
);

INVx3_ASAP7_75t_L g3671 ( 
.A(n_2614),
.Y(n_3671)
);

NAND3xp33_ASAP7_75t_L g3672 ( 
.A(n_2216),
.B(n_2152),
.C(n_2277),
.Y(n_3672)
);

NAND2xp5_ASAP7_75t_L g3673 ( 
.A(n_2488),
.B(n_2493),
.Y(n_3673)
);

A2O1A1Ixp33_ASAP7_75t_L g3674 ( 
.A1(n_2511),
.A2(n_3150),
.B(n_2515),
.C(n_2521),
.Y(n_3674)
);

NAND2xp33_ASAP7_75t_L g3675 ( 
.A(n_2719),
.B(n_2800),
.Y(n_3675)
);

OAI22xp5_ASAP7_75t_L g3676 ( 
.A1(n_2517),
.A2(n_2529),
.B1(n_2547),
.B2(n_2522),
.Y(n_3676)
);

AOI21xp5_ASAP7_75t_L g3677 ( 
.A1(n_2558),
.A2(n_2587),
.B(n_2560),
.Y(n_3677)
);

A2O1A1Ixp33_ASAP7_75t_L g3678 ( 
.A1(n_2592),
.A2(n_3149),
.B(n_2595),
.C(n_2618),
.Y(n_3678)
);

AOI21xp5_ASAP7_75t_L g3679 ( 
.A1(n_2637),
.A2(n_2670),
.B(n_2649),
.Y(n_3679)
);

AOI22xp5_ASAP7_75t_L g3680 ( 
.A1(n_2202),
.A2(n_2235),
.B1(n_2216),
.B2(n_2273),
.Y(n_3680)
);

AND2x2_ASAP7_75t_L g3681 ( 
.A(n_2681),
.B(n_2687),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_SL g3682 ( 
.A(n_2688),
.B(n_2824),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_L g3683 ( 
.A(n_2701),
.B(n_2702),
.Y(n_3683)
);

OAI21xp5_ASAP7_75t_L g3684 ( 
.A1(n_2709),
.A2(n_2721),
.B(n_2713),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_SL g3685 ( 
.A(n_3126),
.B(n_2326),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_SL g3686 ( 
.A(n_2235),
.B(n_2411),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_L g3687 ( 
.A(n_2729),
.B(n_2739),
.Y(n_3687)
);

INVx2_ASAP7_75t_L g3688 ( 
.A(n_2741),
.Y(n_3688)
);

O2A1O1Ixp5_ASAP7_75t_L g3689 ( 
.A1(n_2346),
.A2(n_2324),
.B(n_3134),
.C(n_3120),
.Y(n_3689)
);

AOI22xp5_ASAP7_75t_L g3690 ( 
.A1(n_2250),
.A2(n_2229),
.B1(n_2251),
.B2(n_2263),
.Y(n_3690)
);

A2O1A1Ixp33_ASAP7_75t_L g3691 ( 
.A1(n_2765),
.A2(n_2953),
.B(n_2770),
.C(n_2783),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_L g3692 ( 
.A(n_2774),
.B(n_2786),
.Y(n_3692)
);

AOI22xp5_ASAP7_75t_L g3693 ( 
.A1(n_2788),
.A2(n_2843),
.B1(n_2909),
.B2(n_3116),
.Y(n_3693)
);

AOI21x1_ASAP7_75t_L g3694 ( 
.A1(n_2792),
.A2(n_2821),
.B(n_2803),
.Y(n_3694)
);

AOI21xp5_ASAP7_75t_L g3695 ( 
.A1(n_2827),
.A2(n_2864),
.B(n_2857),
.Y(n_3695)
);

INVx4_ASAP7_75t_L g3696 ( 
.A(n_3147),
.Y(n_3696)
);

NAND2xp5_ASAP7_75t_L g3697 ( 
.A(n_2879),
.B(n_2906),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_L g3698 ( 
.A(n_2913),
.B(n_2956),
.Y(n_3698)
);

BUFx3_ASAP7_75t_L g3699 ( 
.A(n_2800),
.Y(n_3699)
);

AOI21xp5_ASAP7_75t_L g3700 ( 
.A1(n_2963),
.A2(n_2990),
.B(n_2982),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_L g3701 ( 
.A(n_2994),
.B(n_3034),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_L g3702 ( 
.A(n_3057),
.B(n_3103),
.Y(n_3702)
);

AND2x4_ASAP7_75t_L g3703 ( 
.A(n_3110),
.B(n_3111),
.Y(n_3703)
);

AOI21xp5_ASAP7_75t_L g3704 ( 
.A1(n_2265),
.A2(n_2297),
.B(n_2295),
.Y(n_3704)
);

AOI21x1_ASAP7_75t_L g3705 ( 
.A1(n_2304),
.A2(n_2317),
.B(n_2305),
.Y(n_3705)
);

O2A1O1Ixp33_ASAP7_75t_L g3706 ( 
.A1(n_2246),
.A2(n_2341),
.B(n_2242),
.C(n_2333),
.Y(n_3706)
);

AOI22xp33_ASAP7_75t_L g3707 ( 
.A1(n_2695),
.A2(n_3079),
.B1(n_2706),
.B2(n_2147),
.Y(n_3707)
);

AOI21xp33_ASAP7_75t_L g3708 ( 
.A1(n_2215),
.A2(n_2333),
.B(n_2330),
.Y(n_3708)
);

A2O1A1Ixp33_ASAP7_75t_L g3709 ( 
.A1(n_2240),
.A2(n_2337),
.B(n_2330),
.C(n_2350),
.Y(n_3709)
);

OAI22xp5_ASAP7_75t_L g3710 ( 
.A1(n_2356),
.A2(n_2358),
.B1(n_2337),
.B2(n_2332),
.Y(n_3710)
);

OAI22xp5_ASAP7_75t_L g3711 ( 
.A1(n_2356),
.A2(n_2358),
.B1(n_2506),
.B2(n_2544),
.Y(n_3711)
);

AOI21xp5_ASAP7_75t_L g3712 ( 
.A1(n_2240),
.A2(n_2544),
.B(n_2506),
.Y(n_3712)
);

AOI21xp5_ASAP7_75t_L g3713 ( 
.A1(n_2506),
.A2(n_2544),
.B(n_2557),
.Y(n_3713)
);

NAND2xp5_ASAP7_75t_SL g3714 ( 
.A(n_2448),
.B(n_2518),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_2223),
.B(n_2312),
.Y(n_3715)
);

INVx2_ASAP7_75t_L g3716 ( 
.A(n_2054),
.Y(n_3716)
);

AOI21xp5_ASAP7_75t_L g3717 ( 
.A1(n_2557),
.A2(n_3147),
.B(n_2800),
.Y(n_3717)
);

OAI22xp5_ASAP7_75t_L g3718 ( 
.A1(n_2557),
.A2(n_2345),
.B1(n_2422),
.B2(n_2838),
.Y(n_3718)
);

AOI21xp5_ASAP7_75t_L g3719 ( 
.A1(n_3147),
.A2(n_2339),
.B(n_2344),
.Y(n_3719)
);

AOI21x1_ASAP7_75t_L g3720 ( 
.A1(n_2349),
.A2(n_2357),
.B(n_2354),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_2281),
.B(n_2054),
.Y(n_3721)
);

AOI21xp5_ASAP7_75t_L g3722 ( 
.A1(n_3068),
.A2(n_2347),
.B(n_2725),
.Y(n_3722)
);

AOI21xp5_ASAP7_75t_L g3723 ( 
.A1(n_2347),
.A2(n_2725),
.B(n_2198),
.Y(n_3723)
);

AND2x2_ASAP7_75t_L g3724 ( 
.A(n_2226),
.B(n_2248),
.Y(n_3724)
);

INVx2_ASAP7_75t_L g3725 ( 
.A(n_2226),
.Y(n_3725)
);

NAND2xp5_ASAP7_75t_L g3726 ( 
.A(n_2226),
.B(n_2248),
.Y(n_3726)
);

AO21x1_ASAP7_75t_L g3727 ( 
.A1(n_2342),
.A2(n_2355),
.B(n_2348),
.Y(n_3727)
);

NOR2xp33_ASAP7_75t_L g3728 ( 
.A(n_2563),
.B(n_2635),
.Y(n_3728)
);

AOI22xp5_ASAP7_75t_L g3729 ( 
.A1(n_2832),
.A2(n_2967),
.B1(n_2738),
.B2(n_2884),
.Y(n_3729)
);

O2A1O1Ixp33_ASAP7_75t_L g3730 ( 
.A1(n_2115),
.A2(n_2162),
.B(n_2142),
.C(n_2137),
.Y(n_3730)
);

AOI21xp5_ASAP7_75t_L g3731 ( 
.A1(n_2154),
.A2(n_2198),
.B(n_2893),
.Y(n_3731)
);

INVx3_ASAP7_75t_L g3732 ( 
.A(n_2226),
.Y(n_3732)
);

A2O1A1Ixp33_ASAP7_75t_L g3733 ( 
.A1(n_2342),
.A2(n_2355),
.B(n_2861),
.C(n_1998),
.Y(n_3733)
);

INVx2_ASAP7_75t_L g3734 ( 
.A(n_2248),
.Y(n_3734)
);

INVx2_ASAP7_75t_L g3735 ( 
.A(n_2248),
.Y(n_3735)
);

BUFx2_ASAP7_75t_L g3736 ( 
.A(n_2878),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_2310),
.B(n_2371),
.Y(n_3737)
);

OAI21xp5_ASAP7_75t_L g3738 ( 
.A1(n_2094),
.A2(n_2574),
.B(n_2682),
.Y(n_3738)
);

NAND2xp5_ASAP7_75t_L g3739 ( 
.A(n_2310),
.B(n_2371),
.Y(n_3739)
);

AND2x4_ASAP7_75t_L g3740 ( 
.A(n_2113),
.B(n_2442),
.Y(n_3740)
);

AOI21xp5_ASAP7_75t_L g3741 ( 
.A1(n_2154),
.A2(n_2198),
.B(n_3015),
.Y(n_3741)
);

AOI22xp5_ASAP7_75t_L g3742 ( 
.A1(n_3009),
.A2(n_3036),
.B1(n_1997),
.B2(n_2154),
.Y(n_3742)
);

INVxp33_ASAP7_75t_L g3743 ( 
.A(n_2141),
.Y(n_3743)
);

AND2x2_ASAP7_75t_SL g3744 ( 
.A(n_2234),
.B(n_3011),
.Y(n_3744)
);

AOI21xp5_ASAP7_75t_L g3745 ( 
.A1(n_2097),
.A2(n_2996),
.B(n_2502),
.Y(n_3745)
);

NAND2xp5_ASAP7_75t_L g3746 ( 
.A(n_2310),
.B(n_2371),
.Y(n_3746)
);

OR2x2_ASAP7_75t_L g3747 ( 
.A(n_2163),
.B(n_2141),
.Y(n_3747)
);

O2A1O1Ixp33_ASAP7_75t_L g3748 ( 
.A1(n_2133),
.A2(n_3052),
.B(n_2897),
.C(n_2485),
.Y(n_3748)
);

NAND2xp5_ASAP7_75t_L g3749 ( 
.A(n_2310),
.B(n_2371),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_2422),
.Y(n_3750)
);

AOI21xp5_ASAP7_75t_L g3751 ( 
.A1(n_2403),
.A2(n_2500),
.B(n_2408),
.Y(n_3751)
);

OAI21xp5_ASAP7_75t_L g3752 ( 
.A1(n_2859),
.A2(n_3087),
.B(n_2921),
.Y(n_3752)
);

INVxp67_ASAP7_75t_SL g3753 ( 
.A(n_2422),
.Y(n_3753)
);

NAND2xp5_ASAP7_75t_L g3754 ( 
.A(n_2422),
.B(n_2668),
.Y(n_3754)
);

NAND2xp5_ASAP7_75t_L g3755 ( 
.A(n_2513),
.B(n_2668),
.Y(n_3755)
);

BUFx2_ASAP7_75t_L g3756 ( 
.A(n_3083),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_2513),
.Y(n_3757)
);

NOR3xp33_ASAP7_75t_L g3758 ( 
.A(n_2340),
.B(n_2234),
.C(n_2348),
.Y(n_3758)
);

BUFx8_ASAP7_75t_SL g3759 ( 
.A(n_2812),
.Y(n_3759)
);

NOR2xp67_ASAP7_75t_L g3760 ( 
.A(n_2924),
.B(n_2929),
.Y(n_3760)
);

AOI222xp33_ASAP7_75t_L g3761 ( 
.A1(n_3009),
.A2(n_3036),
.B1(n_2947),
.B2(n_2149),
.C1(n_2352),
.C2(n_2669),
.Y(n_3761)
);

AND2x4_ASAP7_75t_L g3762 ( 
.A(n_2673),
.B(n_2885),
.Y(n_3762)
);

BUFx6f_ASAP7_75t_L g3763 ( 
.A(n_2513),
.Y(n_3763)
);

NOR2xp33_ASAP7_75t_L g3764 ( 
.A(n_2149),
.B(n_2197),
.Y(n_3764)
);

AOI21xp5_ASAP7_75t_L g3765 ( 
.A1(n_2950),
.A2(n_2562),
.B(n_2668),
.Y(n_3765)
);

AOI21xp5_ASAP7_75t_L g3766 ( 
.A1(n_2513),
.A2(n_3114),
.B(n_2668),
.Y(n_3766)
);

OAI21xp5_ASAP7_75t_L g3767 ( 
.A1(n_2352),
.A2(n_2165),
.B(n_2323),
.Y(n_3767)
);

INVx2_ASAP7_75t_L g3768 ( 
.A(n_2562),
.Y(n_3768)
);

NOR2xp33_ASAP7_75t_L g3769 ( 
.A(n_2182),
.B(n_1995),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_SL g3770 ( 
.A(n_2562),
.B(n_2679),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_2562),
.Y(n_3771)
);

NAND2xp5_ASAP7_75t_L g3772 ( 
.A(n_2679),
.B(n_3114),
.Y(n_3772)
);

NAND2xp5_ASAP7_75t_L g3773 ( 
.A(n_2679),
.B(n_3114),
.Y(n_3773)
);

AOI22x1_ASAP7_75t_L g3774 ( 
.A1(n_3044),
.A2(n_3055),
.B1(n_3114),
.B2(n_2826),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_SL g3775 ( 
.A(n_2679),
.B(n_2708),
.Y(n_3775)
);

NOR2xp33_ASAP7_75t_R g3776 ( 
.A(n_2108),
.B(n_2338),
.Y(n_3776)
);

AOI21xp5_ASAP7_75t_L g3777 ( 
.A1(n_2708),
.A2(n_2838),
.B(n_2826),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_L g3778 ( 
.A(n_2708),
.B(n_2838),
.Y(n_3778)
);

NAND2xp5_ASAP7_75t_L g3779 ( 
.A(n_2708),
.B(n_2838),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_2798),
.B(n_2826),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_L g3781 ( 
.A(n_2798),
.B(n_2826),
.Y(n_3781)
);

NAND2xp33_ASAP7_75t_SL g3782 ( 
.A(n_2343),
.B(n_2798),
.Y(n_3782)
);

NAND2xp5_ASAP7_75t_L g3783 ( 
.A(n_2798),
.B(n_2253),
.Y(n_3783)
);

AOI21xp5_ASAP7_75t_L g3784 ( 
.A1(n_3145),
.A2(n_3141),
.B(n_3032),
.Y(n_3784)
);

NOR2xp33_ASAP7_75t_L g3785 ( 
.A(n_2418),
.B(n_2602),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_SL g3786 ( 
.A(n_2271),
.B(n_2286),
.Y(n_3786)
);

A2O1A1Ixp33_ASAP7_75t_L g3787 ( 
.A1(n_2307),
.A2(n_2465),
.B(n_2497),
.C(n_2528),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_L g3788 ( 
.A(n_2530),
.B(n_2555),
.Y(n_3788)
);

NAND2xp5_ASAP7_75t_L g3789 ( 
.A(n_2559),
.B(n_2632),
.Y(n_3789)
);

A2O1A1Ixp33_ASAP7_75t_L g3790 ( 
.A1(n_2656),
.A2(n_2907),
.B(n_2928),
.C(n_2980),
.Y(n_3790)
);

NOR2xp33_ASAP7_75t_L g3791 ( 
.A(n_3122),
.B(n_3130),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_3094),
.B(n_2135),
.Y(n_3792)
);

AOI21xp5_ASAP7_75t_L g3793 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3793)
);

OAI21xp5_ASAP7_75t_L g3794 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_3794)
);

NAND2xp5_ASAP7_75t_L g3795 ( 
.A(n_2135),
.B(n_2050),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_L g3796 ( 
.A(n_2135),
.B(n_2050),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_L g3797 ( 
.A(n_2135),
.B(n_2050),
.Y(n_3797)
);

NAND2xp5_ASAP7_75t_L g3798 ( 
.A(n_2135),
.B(n_2050),
.Y(n_3798)
);

AOI21xp5_ASAP7_75t_L g3799 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3799)
);

NAND2xp5_ASAP7_75t_L g3800 ( 
.A(n_2135),
.B(n_2050),
.Y(n_3800)
);

NOR2xp33_ASAP7_75t_L g3801 ( 
.A(n_2025),
.B(n_1067),
.Y(n_3801)
);

NOR2xp67_ASAP7_75t_L g3802 ( 
.A(n_2009),
.B(n_2743),
.Y(n_3802)
);

O2A1O1Ixp5_ASAP7_75t_L g3803 ( 
.A1(n_2393),
.A2(n_788),
.B(n_807),
.C(n_673),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_2232),
.Y(n_3804)
);

NOR2xp33_ASAP7_75t_L g3805 ( 
.A(n_2025),
.B(n_1067),
.Y(n_3805)
);

NAND2xp5_ASAP7_75t_L g3806 ( 
.A(n_2135),
.B(n_2050),
.Y(n_3806)
);

OAI22xp5_ASAP7_75t_L g3807 ( 
.A1(n_3040),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_3807)
);

AND2x2_ASAP7_75t_SL g3808 ( 
.A(n_2549),
.B(n_1311),
.Y(n_3808)
);

NAND2xp5_ASAP7_75t_L g3809 ( 
.A(n_2135),
.B(n_2050),
.Y(n_3809)
);

NAND2x1_ASAP7_75t_L g3810 ( 
.A(n_2081),
.B(n_2252),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_SL g3811 ( 
.A(n_2374),
.B(n_1096),
.Y(n_3811)
);

OAI21xp5_ASAP7_75t_L g3812 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_3812)
);

AND2x2_ASAP7_75t_SL g3813 ( 
.A(n_2549),
.B(n_1311),
.Y(n_3813)
);

AOI22xp5_ASAP7_75t_L g3814 ( 
.A1(n_3053),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_3814)
);

AOI21xp5_ASAP7_75t_L g3815 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3815)
);

AOI21xp5_ASAP7_75t_L g3816 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3816)
);

AOI21x1_ASAP7_75t_L g3817 ( 
.A1(n_1988),
.A2(n_2167),
.B(n_1903),
.Y(n_3817)
);

AOI21xp5_ASAP7_75t_L g3818 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3818)
);

NOR2xp33_ASAP7_75t_L g3819 ( 
.A(n_2025),
.B(n_1067),
.Y(n_3819)
);

A2O1A1Ixp33_ASAP7_75t_L g3820 ( 
.A1(n_2737),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_3820)
);

INVx4_ASAP7_75t_L g3821 ( 
.A(n_2009),
.Y(n_3821)
);

NAND2xp5_ASAP7_75t_L g3822 ( 
.A(n_2135),
.B(n_2050),
.Y(n_3822)
);

BUFx6f_ASAP7_75t_L g3823 ( 
.A(n_2098),
.Y(n_3823)
);

OAI21xp33_ASAP7_75t_L g3824 ( 
.A1(n_2374),
.A2(n_1072),
.B(n_1067),
.Y(n_3824)
);

AOI21xp5_ASAP7_75t_L g3825 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3825)
);

AOI21xp5_ASAP7_75t_L g3826 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3826)
);

INVx1_ASAP7_75t_L g3827 ( 
.A(n_2232),
.Y(n_3827)
);

NAND2xp5_ASAP7_75t_L g3828 ( 
.A(n_2135),
.B(n_2050),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_SL g3829 ( 
.A(n_2374),
.B(n_1096),
.Y(n_3829)
);

BUFx8_ASAP7_75t_L g3830 ( 
.A(n_2180),
.Y(n_3830)
);

INVxp67_ASAP7_75t_L g3831 ( 
.A(n_2760),
.Y(n_3831)
);

INVx1_ASAP7_75t_SL g3832 ( 
.A(n_2144),
.Y(n_3832)
);

BUFx4f_ASAP7_75t_L g3833 ( 
.A(n_2566),
.Y(n_3833)
);

AND2x2_ASAP7_75t_L g3834 ( 
.A(n_2549),
.B(n_2780),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_2232),
.Y(n_3835)
);

O2A1O1Ixp33_ASAP7_75t_L g3836 ( 
.A1(n_3040),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_SL g3837 ( 
.A(n_2374),
.B(n_1096),
.Y(n_3837)
);

NOR2xp33_ASAP7_75t_L g3838 ( 
.A(n_2025),
.B(n_1067),
.Y(n_3838)
);

OAI22xp5_ASAP7_75t_L g3839 ( 
.A1(n_3040),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_3839)
);

NAND2xp5_ASAP7_75t_L g3840 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3841)
);

NOR2x1_ASAP7_75t_R g3842 ( 
.A(n_2328),
.B(n_617),
.Y(n_3842)
);

AOI21xp5_ASAP7_75t_L g3843 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3843)
);

AOI21xp5_ASAP7_75t_L g3844 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3844)
);

AOI21xp5_ASAP7_75t_L g3845 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3845)
);

A2O1A1Ixp33_ASAP7_75t_L g3846 ( 
.A1(n_2737),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_3846)
);

O2A1O1Ixp33_ASAP7_75t_L g3847 ( 
.A1(n_3040),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_3847)
);

INVx1_ASAP7_75t_L g3848 ( 
.A(n_2232),
.Y(n_3848)
);

O2A1O1Ixp33_ASAP7_75t_SL g3849 ( 
.A1(n_2383),
.A2(n_1719),
.B(n_1866),
.C(n_1779),
.Y(n_3849)
);

AND2x4_ASAP7_75t_L g3850 ( 
.A(n_2098),
.B(n_2221),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_SL g3851 ( 
.A(n_2374),
.B(n_1096),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_L g3852 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3852)
);

AOI21x1_ASAP7_75t_L g3853 ( 
.A1(n_1988),
.A2(n_2167),
.B(n_1903),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_2232),
.Y(n_3854)
);

OAI21xp5_ASAP7_75t_L g3855 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_3855)
);

INVx11_ASAP7_75t_L g3856 ( 
.A(n_2177),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_L g3857 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_L g3858 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3858)
);

AND2x2_ASAP7_75t_L g3859 ( 
.A(n_2549),
.B(n_2780),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_2232),
.Y(n_3860)
);

AOI21xp5_ASAP7_75t_L g3861 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3861)
);

INVxp67_ASAP7_75t_L g3862 ( 
.A(n_2760),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_L g3863 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3863)
);

AOI21xp5_ASAP7_75t_L g3864 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3864)
);

BUFx6f_ASAP7_75t_L g3865 ( 
.A(n_2098),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_2232),
.Y(n_3866)
);

AOI21xp5_ASAP7_75t_L g3867 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3867)
);

NAND2xp5_ASAP7_75t_SL g3868 ( 
.A(n_2374),
.B(n_1096),
.Y(n_3868)
);

INVx1_ASAP7_75t_L g3869 ( 
.A(n_2232),
.Y(n_3869)
);

AOI21xp5_ASAP7_75t_L g3870 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3870)
);

AO21x1_ASAP7_75t_L g3871 ( 
.A1(n_1988),
.A2(n_2145),
.B(n_2363),
.Y(n_3871)
);

NAND2xp5_ASAP7_75t_L g3872 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3872)
);

AOI21xp5_ASAP7_75t_L g3873 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3873)
);

NAND2xp5_ASAP7_75t_L g3874 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3874)
);

OR2x6_ASAP7_75t_L g3875 ( 
.A(n_2167),
.B(n_2221),
.Y(n_3875)
);

A2O1A1Ixp33_ASAP7_75t_L g3876 ( 
.A1(n_2737),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_L g3877 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3877)
);

NAND2xp5_ASAP7_75t_L g3878 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_2232),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_L g3880 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3880)
);

AOI21xp5_ASAP7_75t_L g3881 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3881)
);

A2O1A1Ixp33_ASAP7_75t_L g3882 ( 
.A1(n_2737),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3883)
);

NAND2xp5_ASAP7_75t_SL g3884 ( 
.A(n_2374),
.B(n_1096),
.Y(n_3884)
);

INVx2_ASAP7_75t_SL g3885 ( 
.A(n_2054),
.Y(n_3885)
);

NAND2xp5_ASAP7_75t_L g3886 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3886)
);

O2A1O1Ixp33_ASAP7_75t_L g3887 ( 
.A1(n_3040),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_L g3888 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3888)
);

HB1xp67_ASAP7_75t_L g3889 ( 
.A(n_2144),
.Y(n_3889)
);

OAI22xp5_ASAP7_75t_L g3890 ( 
.A1(n_3040),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_3890)
);

NOR2xp33_ASAP7_75t_L g3891 ( 
.A(n_2025),
.B(n_1067),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_L g3892 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3892)
);

NAND2x1p5_ASAP7_75t_L g3893 ( 
.A(n_2098),
.B(n_2027),
.Y(n_3893)
);

OAI21xp5_ASAP7_75t_L g3894 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_3894)
);

NAND2xp5_ASAP7_75t_L g3895 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3895)
);

OAI21xp5_ASAP7_75t_L g3896 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_3896)
);

NAND2xp5_ASAP7_75t_L g3897 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3897)
);

AO21x1_ASAP7_75t_L g3898 ( 
.A1(n_1988),
.A2(n_2145),
.B(n_2363),
.Y(n_3898)
);

CKINVDCx5p33_ASAP7_75t_R g3899 ( 
.A(n_2328),
.Y(n_3899)
);

AOI21xp5_ASAP7_75t_L g3900 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3900)
);

INVx1_ASAP7_75t_SL g3901 ( 
.A(n_2144),
.Y(n_3901)
);

OAI21xp5_ASAP7_75t_L g3902 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_3902)
);

AOI21xp5_ASAP7_75t_L g3903 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3903)
);

NOR2xp33_ASAP7_75t_L g3904 ( 
.A(n_2025),
.B(n_1067),
.Y(n_3904)
);

A2O1A1Ixp33_ASAP7_75t_L g3905 ( 
.A1(n_2737),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_3905)
);

A2O1A1Ixp33_ASAP7_75t_L g3906 ( 
.A1(n_2737),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_3906)
);

AOI21xp5_ASAP7_75t_L g3907 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3907)
);

AOI21xp5_ASAP7_75t_L g3908 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3908)
);

AOI21xp5_ASAP7_75t_L g3909 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3909)
);

AO21x1_ASAP7_75t_L g3910 ( 
.A1(n_1988),
.A2(n_2145),
.B(n_2363),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_L g3911 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3911)
);

AND2x4_ASAP7_75t_L g3912 ( 
.A(n_2098),
.B(n_2221),
.Y(n_3912)
);

NAND2xp5_ASAP7_75t_L g3913 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3913)
);

INVx4_ASAP7_75t_L g3914 ( 
.A(n_2009),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_2232),
.Y(n_3915)
);

NAND2xp5_ASAP7_75t_L g3916 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3916)
);

AOI21xp5_ASAP7_75t_L g3917 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3917)
);

OR2x6_ASAP7_75t_L g3918 ( 
.A(n_2167),
.B(n_2221),
.Y(n_3918)
);

OAI21xp5_ASAP7_75t_L g3919 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_3919)
);

NOR2xp33_ASAP7_75t_L g3920 ( 
.A(n_2025),
.B(n_1067),
.Y(n_3920)
);

OAI22xp5_ASAP7_75t_L g3921 ( 
.A1(n_3040),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_3921)
);

AOI21xp5_ASAP7_75t_L g3922 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3922)
);

BUFx12f_ASAP7_75t_L g3923 ( 
.A(n_2328),
.Y(n_3923)
);

OAI21xp5_ASAP7_75t_L g3924 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_3924)
);

AND2x2_ASAP7_75t_SL g3925 ( 
.A(n_2549),
.B(n_1311),
.Y(n_3925)
);

AND2x2_ASAP7_75t_L g3926 ( 
.A(n_2549),
.B(n_2780),
.Y(n_3926)
);

NAND2xp5_ASAP7_75t_L g3927 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_SL g3928 ( 
.A(n_2374),
.B(n_1096),
.Y(n_3928)
);

BUFx6f_ASAP7_75t_L g3929 ( 
.A(n_2098),
.Y(n_3929)
);

AOI21xp5_ASAP7_75t_L g3930 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3930)
);

NAND2xp5_ASAP7_75t_SL g3931 ( 
.A(n_2374),
.B(n_1096),
.Y(n_3931)
);

OAI21xp33_ASAP7_75t_L g3932 ( 
.A1(n_2374),
.A2(n_1072),
.B(n_1067),
.Y(n_3932)
);

AOI21xp5_ASAP7_75t_L g3933 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3934)
);

BUFx6f_ASAP7_75t_L g3935 ( 
.A(n_2098),
.Y(n_3935)
);

AOI22xp5_ASAP7_75t_L g3936 ( 
.A1(n_3053),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_2232),
.Y(n_3937)
);

AOI21xp5_ASAP7_75t_L g3938 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3938)
);

BUFx4f_ASAP7_75t_L g3939 ( 
.A(n_2566),
.Y(n_3939)
);

NAND2xp5_ASAP7_75t_L g3940 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3940)
);

AOI21x1_ASAP7_75t_L g3941 ( 
.A1(n_1988),
.A2(n_2167),
.B(n_1903),
.Y(n_3941)
);

AOI21xp5_ASAP7_75t_L g3942 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3942)
);

NAND2xp5_ASAP7_75t_L g3943 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3943)
);

AOI21xp5_ASAP7_75t_L g3944 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3944)
);

NOR2xp33_ASAP7_75t_L g3945 ( 
.A(n_2025),
.B(n_1067),
.Y(n_3945)
);

NOR2xp33_ASAP7_75t_L g3946 ( 
.A(n_2025),
.B(n_1067),
.Y(n_3946)
);

AOI21x1_ASAP7_75t_L g3947 ( 
.A1(n_1988),
.A2(n_2167),
.B(n_1903),
.Y(n_3947)
);

AOI21xp5_ASAP7_75t_L g3948 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3948)
);

O2A1O1Ixp33_ASAP7_75t_L g3949 ( 
.A1(n_3040),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_3949)
);

BUFx6f_ASAP7_75t_L g3950 ( 
.A(n_2098),
.Y(n_3950)
);

AND2x4_ASAP7_75t_L g3951 ( 
.A(n_2098),
.B(n_2221),
.Y(n_3951)
);

NOR2xp33_ASAP7_75t_L g3952 ( 
.A(n_2025),
.B(n_1067),
.Y(n_3952)
);

AND2x2_ASAP7_75t_L g3953 ( 
.A(n_2549),
.B(n_2780),
.Y(n_3953)
);

NOR2xp33_ASAP7_75t_SL g3954 ( 
.A(n_3040),
.B(n_1067),
.Y(n_3954)
);

NAND2xp5_ASAP7_75t_L g3955 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3955)
);

OAI21xp5_ASAP7_75t_L g3956 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_3956)
);

NAND2xp5_ASAP7_75t_L g3957 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3957)
);

NAND2xp5_ASAP7_75t_SL g3958 ( 
.A(n_2374),
.B(n_1096),
.Y(n_3958)
);

AND2x2_ASAP7_75t_L g3959 ( 
.A(n_2549),
.B(n_2780),
.Y(n_3959)
);

O2A1O1Ixp33_ASAP7_75t_L g3960 ( 
.A1(n_3040),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_3960)
);

AOI21xp5_ASAP7_75t_L g3961 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_L g3962 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3962)
);

NAND2xp5_ASAP7_75t_L g3963 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3963)
);

AOI21xp5_ASAP7_75t_L g3964 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_2232),
.Y(n_3965)
);

A2O1A1Ixp33_ASAP7_75t_L g3966 ( 
.A1(n_2737),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_3966)
);

NAND2xp5_ASAP7_75t_L g3967 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_2232),
.Y(n_3968)
);

INVx4_ASAP7_75t_L g3969 ( 
.A(n_2009),
.Y(n_3969)
);

OAI21xp5_ASAP7_75t_L g3970 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_3970)
);

AOI21xp5_ASAP7_75t_L g3971 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3971)
);

NAND2xp5_ASAP7_75t_L g3972 ( 
.A(n_2091),
.B(n_1067),
.Y(n_3972)
);

INVx1_ASAP7_75t_L g3973 ( 
.A(n_2232),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_L g3974 ( 
.A(n_2135),
.B(n_2050),
.Y(n_3974)
);

NOR3xp33_ASAP7_75t_L g3975 ( 
.A(n_2829),
.B(n_788),
.C(n_673),
.Y(n_3975)
);

INVx2_ASAP7_75t_SL g3976 ( 
.A(n_2054),
.Y(n_3976)
);

CKINVDCx10_ASAP7_75t_R g3977 ( 
.A(n_2180),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_L g3978 ( 
.A(n_2135),
.B(n_2050),
.Y(n_3978)
);

OAI21xp5_ASAP7_75t_L g3979 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_3979)
);

OAI21xp5_ASAP7_75t_L g3980 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_3980)
);

NAND2xp5_ASAP7_75t_SL g3981 ( 
.A(n_2374),
.B(n_1096),
.Y(n_3981)
);

NAND2xp5_ASAP7_75t_L g3982 ( 
.A(n_2135),
.B(n_2050),
.Y(n_3982)
);

AOI22xp33_ASAP7_75t_L g3983 ( 
.A1(n_1987),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_3983)
);

AOI22xp5_ASAP7_75t_L g3984 ( 
.A1(n_3053),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_3984)
);

NOR3xp33_ASAP7_75t_L g3985 ( 
.A(n_2829),
.B(n_788),
.C(n_673),
.Y(n_3985)
);

INVx2_ASAP7_75t_SL g3986 ( 
.A(n_2054),
.Y(n_3986)
);

AOI22xp5_ASAP7_75t_L g3987 ( 
.A1(n_3053),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_3987)
);

INVx4_ASAP7_75t_L g3988 ( 
.A(n_2009),
.Y(n_3988)
);

AOI21xp5_ASAP7_75t_L g3989 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3989)
);

AOI21xp5_ASAP7_75t_L g3990 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3990)
);

NAND2xp5_ASAP7_75t_L g3991 ( 
.A(n_2135),
.B(n_2050),
.Y(n_3991)
);

NOR2xp33_ASAP7_75t_L g3992 ( 
.A(n_2025),
.B(n_1067),
.Y(n_3992)
);

AOI21xp5_ASAP7_75t_L g3993 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3993)
);

AOI21xp5_ASAP7_75t_L g3994 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3994)
);

NOR2xp33_ASAP7_75t_L g3995 ( 
.A(n_2025),
.B(n_1067),
.Y(n_3995)
);

NOR2x1_ASAP7_75t_R g3996 ( 
.A(n_2328),
.B(n_617),
.Y(n_3996)
);

NAND2xp5_ASAP7_75t_SL g3997 ( 
.A(n_2374),
.B(n_1096),
.Y(n_3997)
);

AOI21xp5_ASAP7_75t_L g3998 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3998)
);

AOI21xp5_ASAP7_75t_L g3999 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_2232),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_L g4001 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4001)
);

AOI21xp5_ASAP7_75t_L g4002 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_2232),
.Y(n_4003)
);

BUFx3_ASAP7_75t_L g4004 ( 
.A(n_2719),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_SL g4005 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4005)
);

INVx1_ASAP7_75t_L g4006 ( 
.A(n_2232),
.Y(n_4006)
);

NAND2xp5_ASAP7_75t_SL g4007 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4007)
);

AOI21xp5_ASAP7_75t_L g4008 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4008)
);

AO21x1_ASAP7_75t_L g4009 ( 
.A1(n_1988),
.A2(n_2145),
.B(n_2363),
.Y(n_4009)
);

AOI21xp5_ASAP7_75t_L g4010 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4010)
);

NAND2xp5_ASAP7_75t_L g4011 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4011)
);

OAI21xp33_ASAP7_75t_L g4012 ( 
.A1(n_2374),
.A2(n_1072),
.B(n_1067),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_L g4013 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4013)
);

OAI21xp5_ASAP7_75t_L g4014 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4014)
);

AOI21xp5_ASAP7_75t_L g4015 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4015)
);

AOI21xp5_ASAP7_75t_L g4016 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4016)
);

NAND2xp5_ASAP7_75t_SL g4017 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4017)
);

AOI22xp33_ASAP7_75t_L g4018 ( 
.A1(n_1987),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_4018)
);

AOI21x1_ASAP7_75t_L g4019 ( 
.A1(n_1988),
.A2(n_2167),
.B(n_1903),
.Y(n_4019)
);

AND2x2_ASAP7_75t_L g4020 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4020)
);

INVx2_ASAP7_75t_SL g4021 ( 
.A(n_2054),
.Y(n_4021)
);

INVx1_ASAP7_75t_L g4022 ( 
.A(n_2232),
.Y(n_4022)
);

NAND2xp5_ASAP7_75t_L g4023 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4023)
);

AND2x2_ASAP7_75t_L g4024 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4024)
);

NAND2xp5_ASAP7_75t_L g4025 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4025)
);

AND2x4_ASAP7_75t_L g4026 ( 
.A(n_2098),
.B(n_2221),
.Y(n_4026)
);

AOI21x1_ASAP7_75t_L g4027 ( 
.A1(n_1988),
.A2(n_2167),
.B(n_1903),
.Y(n_4027)
);

BUFx2_ASAP7_75t_SL g4028 ( 
.A(n_2009),
.Y(n_4028)
);

NAND2xp5_ASAP7_75t_SL g4029 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4029)
);

AOI21xp5_ASAP7_75t_L g4030 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4030)
);

OAI21xp5_ASAP7_75t_L g4031 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4031)
);

AO21x1_ASAP7_75t_L g4032 ( 
.A1(n_1988),
.A2(n_2145),
.B(n_2363),
.Y(n_4032)
);

O2A1O1Ixp33_ASAP7_75t_L g4033 ( 
.A1(n_3040),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4033)
);

AOI21xp5_ASAP7_75t_L g4034 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4034)
);

OAI22xp5_ASAP7_75t_L g4035 ( 
.A1(n_3040),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_4035)
);

AOI21xp5_ASAP7_75t_L g4036 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4036)
);

NOR2xp33_ASAP7_75t_L g4037 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4037)
);

AO21x1_ASAP7_75t_L g4038 ( 
.A1(n_1988),
.A2(n_2145),
.B(n_2363),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_L g4039 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4039)
);

OR2x2_ASAP7_75t_L g4040 ( 
.A(n_1988),
.B(n_2016),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_L g4041 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4041)
);

A2O1A1Ixp33_ASAP7_75t_L g4042 ( 
.A1(n_2737),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4042)
);

HB1xp67_ASAP7_75t_L g4043 ( 
.A(n_2144),
.Y(n_4043)
);

OAI21xp5_ASAP7_75t_L g4044 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4044)
);

AOI21xp5_ASAP7_75t_L g4045 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4045)
);

INVx2_ASAP7_75t_SL g4046 ( 
.A(n_2054),
.Y(n_4046)
);

NOR2xp33_ASAP7_75t_L g4047 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4047)
);

AOI22xp5_ASAP7_75t_L g4048 ( 
.A1(n_3053),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_4048)
);

AND2x2_ASAP7_75t_L g4049 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4049)
);

INVx2_ASAP7_75t_SL g4050 ( 
.A(n_2054),
.Y(n_4050)
);

INVx1_ASAP7_75t_SL g4051 ( 
.A(n_2144),
.Y(n_4051)
);

INVx2_ASAP7_75t_SL g4052 ( 
.A(n_2054),
.Y(n_4052)
);

AOI21x1_ASAP7_75t_L g4053 ( 
.A1(n_1988),
.A2(n_2167),
.B(n_1903),
.Y(n_4053)
);

O2A1O1Ixp5_ASAP7_75t_L g4054 ( 
.A1(n_2393),
.A2(n_788),
.B(n_807),
.C(n_673),
.Y(n_4054)
);

NAND2xp5_ASAP7_75t_L g4055 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4055)
);

OAI21xp5_ASAP7_75t_L g4056 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4056)
);

NAND2xp5_ASAP7_75t_L g4057 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4057)
);

INVx4_ASAP7_75t_L g4058 ( 
.A(n_2009),
.Y(n_4058)
);

BUFx6f_ASAP7_75t_L g4059 ( 
.A(n_2098),
.Y(n_4059)
);

NOR2xp33_ASAP7_75t_L g4060 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4060)
);

AOI21xp5_ASAP7_75t_L g4061 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4061)
);

NOR2xp33_ASAP7_75t_L g4062 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4062)
);

INVx1_ASAP7_75t_L g4063 ( 
.A(n_2232),
.Y(n_4063)
);

INVxp67_ASAP7_75t_L g4064 ( 
.A(n_2760),
.Y(n_4064)
);

NAND2xp5_ASAP7_75t_L g4065 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4065)
);

BUFx3_ASAP7_75t_L g4066 ( 
.A(n_2719),
.Y(n_4066)
);

OAI22xp5_ASAP7_75t_L g4067 ( 
.A1(n_3040),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_4067)
);

AND2x2_ASAP7_75t_L g4068 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4068)
);

NAND2xp5_ASAP7_75t_L g4069 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4069)
);

AOI21x1_ASAP7_75t_L g4070 ( 
.A1(n_1988),
.A2(n_2167),
.B(n_1903),
.Y(n_4070)
);

OAI22xp5_ASAP7_75t_L g4071 ( 
.A1(n_3040),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_4071)
);

BUFx6f_ASAP7_75t_L g4072 ( 
.A(n_2098),
.Y(n_4072)
);

NAND2xp5_ASAP7_75t_L g4073 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4073)
);

OAI22xp5_ASAP7_75t_L g4074 ( 
.A1(n_3040),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_4074)
);

OAI21xp5_ASAP7_75t_L g4075 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4075)
);

NAND2xp5_ASAP7_75t_SL g4076 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4076)
);

NOR2x1p5_ASAP7_75t_SL g4077 ( 
.A(n_2614),
.B(n_1272),
.Y(n_4077)
);

AOI21xp5_ASAP7_75t_L g4078 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4078)
);

OAI21xp5_ASAP7_75t_L g4079 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4079)
);

NOR2xp33_ASAP7_75t_L g4080 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4080)
);

NAND2xp5_ASAP7_75t_SL g4081 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4081)
);

OAI21xp5_ASAP7_75t_L g4082 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4082)
);

AOI21xp5_ASAP7_75t_L g4083 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4083)
);

AOI21xp5_ASAP7_75t_L g4084 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4084)
);

AO21x1_ASAP7_75t_L g4085 ( 
.A1(n_1988),
.A2(n_2145),
.B(n_2363),
.Y(n_4085)
);

OAI21xp5_ASAP7_75t_L g4086 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4086)
);

NAND2xp5_ASAP7_75t_L g4087 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4087)
);

NOR2xp33_ASAP7_75t_L g4088 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4088)
);

O2A1O1Ixp33_ASAP7_75t_SL g4089 ( 
.A1(n_2383),
.A2(n_1719),
.B(n_1866),
.C(n_1779),
.Y(n_4089)
);

AND2x2_ASAP7_75t_L g4090 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4090)
);

NAND2xp5_ASAP7_75t_L g4091 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4091)
);

NAND2xp5_ASAP7_75t_L g4092 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4092)
);

NAND2xp5_ASAP7_75t_L g4093 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4093)
);

OR2x2_ASAP7_75t_L g4094 ( 
.A(n_1988),
.B(n_2016),
.Y(n_4094)
);

AO21x1_ASAP7_75t_L g4095 ( 
.A1(n_1988),
.A2(n_2145),
.B(n_2363),
.Y(n_4095)
);

NAND2xp5_ASAP7_75t_L g4096 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_SL g4097 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4097)
);

BUFx6f_ASAP7_75t_L g4098 ( 
.A(n_2098),
.Y(n_4098)
);

O2A1O1Ixp5_ASAP7_75t_L g4099 ( 
.A1(n_2393),
.A2(n_788),
.B(n_807),
.C(n_673),
.Y(n_4099)
);

OAI21xp5_ASAP7_75t_L g4100 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_2232),
.Y(n_4101)
);

OAI21xp5_ASAP7_75t_L g4102 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4102)
);

AOI21xp5_ASAP7_75t_L g4103 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4103)
);

AOI21xp5_ASAP7_75t_L g4104 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4104)
);

AOI21xp5_ASAP7_75t_L g4105 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4105)
);

NOR2xp33_ASAP7_75t_L g4106 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4106)
);

NAND2xp5_ASAP7_75t_L g4107 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4107)
);

BUFx6f_ASAP7_75t_L g4108 ( 
.A(n_2098),
.Y(n_4108)
);

AOI21xp5_ASAP7_75t_L g4109 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4109)
);

AND2x4_ASAP7_75t_L g4110 ( 
.A(n_2098),
.B(n_2221),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_SL g4111 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4112)
);

A2O1A1Ixp33_ASAP7_75t_L g4113 ( 
.A1(n_2737),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4113)
);

AOI21xp5_ASAP7_75t_L g4114 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4114)
);

NAND2x1_ASAP7_75t_L g4115 ( 
.A(n_2081),
.B(n_2252),
.Y(n_4115)
);

NAND2xp5_ASAP7_75t_SL g4116 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4116)
);

OAI21xp5_ASAP7_75t_L g4117 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4117)
);

AOI21xp5_ASAP7_75t_L g4118 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4118)
);

AOI21xp5_ASAP7_75t_L g4119 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4119)
);

AOI21xp5_ASAP7_75t_L g4120 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4120)
);

AOI21xp5_ASAP7_75t_L g4121 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4121)
);

BUFx6f_ASAP7_75t_L g4122 ( 
.A(n_2098),
.Y(n_4122)
);

AOI21xp5_ASAP7_75t_L g4123 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4123)
);

BUFx3_ASAP7_75t_L g4124 ( 
.A(n_2719),
.Y(n_4124)
);

A2O1A1Ixp33_ASAP7_75t_L g4125 ( 
.A1(n_2737),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4125)
);

AOI21xp5_ASAP7_75t_L g4126 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4126)
);

NAND2xp5_ASAP7_75t_L g4127 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4127)
);

HB1xp67_ASAP7_75t_L g4128 ( 
.A(n_2144),
.Y(n_4128)
);

O2A1O1Ixp33_ASAP7_75t_L g4129 ( 
.A1(n_3040),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4129)
);

AOI21xp5_ASAP7_75t_L g4130 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4130)
);

OAI21xp5_ASAP7_75t_L g4131 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4131)
);

NAND2xp5_ASAP7_75t_L g4132 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_2232),
.Y(n_4133)
);

AOI21xp5_ASAP7_75t_L g4134 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4134)
);

NAND2x1_ASAP7_75t_L g4135 ( 
.A(n_2081),
.B(n_2252),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_L g4136 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4136)
);

INVx1_ASAP7_75t_L g4137 ( 
.A(n_2232),
.Y(n_4137)
);

AOI21xp5_ASAP7_75t_L g4138 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4138)
);

INVxp67_ASAP7_75t_L g4139 ( 
.A(n_2760),
.Y(n_4139)
);

NOR3xp33_ASAP7_75t_L g4140 ( 
.A(n_2829),
.B(n_788),
.C(n_673),
.Y(n_4140)
);

NOR2xp33_ASAP7_75t_L g4141 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4141)
);

BUFx2_ASAP7_75t_L g4142 ( 
.A(n_2760),
.Y(n_4142)
);

NAND2xp33_ASAP7_75t_L g4143 ( 
.A(n_2416),
.B(n_1066),
.Y(n_4143)
);

AOI21xp5_ASAP7_75t_L g4144 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4144)
);

NOR2xp33_ASAP7_75t_L g4145 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4145)
);

NOR2xp33_ASAP7_75t_L g4146 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4146)
);

AND2x4_ASAP7_75t_L g4147 ( 
.A(n_2098),
.B(n_2221),
.Y(n_4147)
);

NAND2xp5_ASAP7_75t_L g4148 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4148)
);

NAND2xp5_ASAP7_75t_L g4149 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4149)
);

NAND2xp5_ASAP7_75t_L g4150 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4150)
);

AOI21x1_ASAP7_75t_L g4151 ( 
.A1(n_1988),
.A2(n_2167),
.B(n_1903),
.Y(n_4151)
);

BUFx2_ASAP7_75t_L g4152 ( 
.A(n_2760),
.Y(n_4152)
);

BUFx2_ASAP7_75t_L g4153 ( 
.A(n_2760),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_SL g4154 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4154)
);

NAND2xp5_ASAP7_75t_SL g4155 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4155)
);

NOR2xp33_ASAP7_75t_L g4156 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4156)
);

OAI21xp5_ASAP7_75t_L g4157 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4157)
);

OAI22xp33_ASAP7_75t_L g4158 ( 
.A1(n_2390),
.A2(n_1085),
.B1(n_1089),
.B2(n_1081),
.Y(n_4158)
);

NAND2xp5_ASAP7_75t_SL g4159 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4159)
);

O2A1O1Ixp33_ASAP7_75t_L g4160 ( 
.A1(n_3040),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_L g4161 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4161)
);

AOI21xp5_ASAP7_75t_L g4162 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4162)
);

AND2x2_ASAP7_75t_L g4163 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4163)
);

OAI21xp5_ASAP7_75t_L g4164 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4164)
);

NAND2xp5_ASAP7_75t_L g4165 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4165)
);

O2A1O1Ixp33_ASAP7_75t_L g4166 ( 
.A1(n_3040),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4166)
);

AOI21xp5_ASAP7_75t_L g4167 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4167)
);

OAI22xp5_ASAP7_75t_L g4168 ( 
.A1(n_3040),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_4168)
);

AOI21xp5_ASAP7_75t_L g4169 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4169)
);

NAND2xp5_ASAP7_75t_L g4170 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4170)
);

AOI21xp5_ASAP7_75t_L g4171 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4171)
);

NAND2xp33_ASAP7_75t_L g4172 ( 
.A(n_2416),
.B(n_1066),
.Y(n_4172)
);

NAND2xp5_ASAP7_75t_L g4173 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4173)
);

NOR2xp33_ASAP7_75t_L g4174 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4174)
);

NAND2xp5_ASAP7_75t_SL g4175 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4175)
);

AOI21xp5_ASAP7_75t_L g4176 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4176)
);

NAND2xp5_ASAP7_75t_L g4177 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4177)
);

NAND2xp5_ASAP7_75t_L g4178 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_L g4179 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_L g4180 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4180)
);

NAND2x1_ASAP7_75t_L g4181 ( 
.A(n_2081),
.B(n_2252),
.Y(n_4181)
);

INVx1_ASAP7_75t_SL g4182 ( 
.A(n_2144),
.Y(n_4182)
);

NAND2xp5_ASAP7_75t_L g4183 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4183)
);

NOR2xp33_ASAP7_75t_L g4184 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4184)
);

NOR2xp33_ASAP7_75t_L g4185 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4185)
);

AND2x2_ASAP7_75t_L g4186 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4186)
);

OR2x6_ASAP7_75t_L g4187 ( 
.A(n_2167),
.B(n_2221),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_2232),
.Y(n_4188)
);

NAND3x1_ASAP7_75t_L g4189 ( 
.A(n_2362),
.B(n_2387),
.C(n_2373),
.Y(n_4189)
);

BUFx3_ASAP7_75t_L g4190 ( 
.A(n_2719),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_L g4191 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4191)
);

AOI21xp5_ASAP7_75t_L g4192 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4192)
);

AOI21xp5_ASAP7_75t_L g4193 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_2232),
.Y(n_4194)
);

AND2x2_ASAP7_75t_L g4195 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4195)
);

AO21x1_ASAP7_75t_L g4196 ( 
.A1(n_1988),
.A2(n_2145),
.B(n_2363),
.Y(n_4196)
);

AOI21xp5_ASAP7_75t_L g4197 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4197)
);

A2O1A1Ixp33_ASAP7_75t_L g4198 ( 
.A1(n_2737),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4198)
);

BUFx6f_ASAP7_75t_L g4199 ( 
.A(n_2098),
.Y(n_4199)
);

CKINVDCx5p33_ASAP7_75t_R g4200 ( 
.A(n_2328),
.Y(n_4200)
);

NAND2xp5_ASAP7_75t_L g4201 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4201)
);

AOI21x1_ASAP7_75t_L g4202 ( 
.A1(n_1988),
.A2(n_2167),
.B(n_1903),
.Y(n_4202)
);

OAI21xp5_ASAP7_75t_L g4203 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4203)
);

OAI21xp5_ASAP7_75t_L g4204 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4204)
);

NOR2xp67_ASAP7_75t_L g4205 ( 
.A(n_2009),
.B(n_2743),
.Y(n_4205)
);

AOI21x1_ASAP7_75t_L g4206 ( 
.A1(n_1988),
.A2(n_2167),
.B(n_1903),
.Y(n_4206)
);

AND2x2_ASAP7_75t_L g4207 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4207)
);

NOR3xp33_ASAP7_75t_L g4208 ( 
.A(n_2829),
.B(n_788),
.C(n_673),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_2232),
.Y(n_4209)
);

AOI21xp5_ASAP7_75t_L g4210 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4210)
);

NAND2xp5_ASAP7_75t_L g4211 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4211)
);

NAND2xp5_ASAP7_75t_L g4212 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_SL g4213 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4213)
);

NAND2xp5_ASAP7_75t_SL g4214 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4214)
);

NAND2xp5_ASAP7_75t_L g4215 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4215)
);

CKINVDCx5p33_ASAP7_75t_R g4216 ( 
.A(n_2328),
.Y(n_4216)
);

HB1xp67_ASAP7_75t_L g4217 ( 
.A(n_2144),
.Y(n_4217)
);

INVx3_ASAP7_75t_L g4218 ( 
.A(n_2081),
.Y(n_4218)
);

NAND2xp5_ASAP7_75t_SL g4219 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_L g4220 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4220)
);

NAND2xp5_ASAP7_75t_L g4221 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4221)
);

AND2x6_ASAP7_75t_L g4222 ( 
.A(n_2081),
.B(n_2252),
.Y(n_4222)
);

NAND2x1p5_ASAP7_75t_L g4223 ( 
.A(n_2098),
.B(n_2027),
.Y(n_4223)
);

AOI22xp33_ASAP7_75t_L g4224 ( 
.A1(n_1987),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_4224)
);

HB1xp67_ASAP7_75t_L g4225 ( 
.A(n_2144),
.Y(n_4225)
);

BUFx6f_ASAP7_75t_L g4226 ( 
.A(n_2098),
.Y(n_4226)
);

HB1xp67_ASAP7_75t_L g4227 ( 
.A(n_2144),
.Y(n_4227)
);

AOI21xp5_ASAP7_75t_L g4228 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_2232),
.Y(n_4229)
);

NAND2xp5_ASAP7_75t_L g4230 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4230)
);

OAI21xp5_ASAP7_75t_L g4231 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_L g4232 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4232)
);

AND2x2_ASAP7_75t_L g4233 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_2232),
.Y(n_4234)
);

AOI21x1_ASAP7_75t_L g4235 ( 
.A1(n_1988),
.A2(n_2167),
.B(n_1903),
.Y(n_4235)
);

BUFx12f_ASAP7_75t_L g4236 ( 
.A(n_2328),
.Y(n_4236)
);

NAND2xp5_ASAP7_75t_L g4237 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_2232),
.Y(n_4238)
);

AOI21xp5_ASAP7_75t_L g4239 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4239)
);

NAND2xp5_ASAP7_75t_L g4240 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4240)
);

NAND2xp5_ASAP7_75t_L g4241 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4241)
);

AOI21xp5_ASAP7_75t_L g4242 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4242)
);

O2A1O1Ixp33_ASAP7_75t_L g4243 ( 
.A1(n_3040),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4243)
);

HB1xp67_ASAP7_75t_L g4244 ( 
.A(n_2144),
.Y(n_4244)
);

AOI21x1_ASAP7_75t_L g4245 ( 
.A1(n_1988),
.A2(n_2167),
.B(n_1903),
.Y(n_4245)
);

INVx4_ASAP7_75t_L g4246 ( 
.A(n_2009),
.Y(n_4246)
);

NAND2xp5_ASAP7_75t_L g4247 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4247)
);

BUFx6f_ASAP7_75t_L g4248 ( 
.A(n_2098),
.Y(n_4248)
);

AOI21xp5_ASAP7_75t_L g4249 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4249)
);

NOR3xp33_ASAP7_75t_L g4250 ( 
.A(n_2829),
.B(n_788),
.C(n_673),
.Y(n_4250)
);

OAI321xp33_ASAP7_75t_L g4251 ( 
.A1(n_3040),
.A2(n_1090),
.A3(n_1067),
.B1(n_1101),
.B2(n_1087),
.C(n_1072),
.Y(n_4251)
);

AOI33xp33_ASAP7_75t_L g4252 ( 
.A1(n_2703),
.A2(n_1136),
.A3(n_1155),
.B1(n_1209),
.B2(n_1205),
.B3(n_1066),
.Y(n_4252)
);

AO21x1_ASAP7_75t_L g4253 ( 
.A1(n_1988),
.A2(n_2145),
.B(n_2363),
.Y(n_4253)
);

AND2x2_ASAP7_75t_L g4254 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4254)
);

A2O1A1Ixp33_ASAP7_75t_L g4255 ( 
.A1(n_2737),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4255)
);

NAND2xp5_ASAP7_75t_L g4256 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4256)
);

AOI21xp5_ASAP7_75t_L g4257 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4257)
);

NAND2xp5_ASAP7_75t_L g4258 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4258)
);

HB1xp67_ASAP7_75t_L g4259 ( 
.A(n_2144),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_2232),
.Y(n_4260)
);

NAND2xp5_ASAP7_75t_L g4261 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4261)
);

AOI21xp5_ASAP7_75t_L g4262 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4262)
);

NOR2xp33_ASAP7_75t_L g4263 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4263)
);

BUFx6f_ASAP7_75t_L g4264 ( 
.A(n_2098),
.Y(n_4264)
);

AOI21xp5_ASAP7_75t_L g4265 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4265)
);

NOR2xp33_ASAP7_75t_L g4266 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4266)
);

AOI21xp5_ASAP7_75t_L g4267 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4267)
);

A2O1A1Ixp33_ASAP7_75t_L g4268 ( 
.A1(n_2737),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4268)
);

AND2x2_ASAP7_75t_L g4269 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4269)
);

A2O1A1Ixp33_ASAP7_75t_L g4270 ( 
.A1(n_2737),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4270)
);

O2A1O1Ixp33_ASAP7_75t_SL g4271 ( 
.A1(n_2383),
.A2(n_1719),
.B(n_1866),
.C(n_1779),
.Y(n_4271)
);

BUFx3_ASAP7_75t_L g4272 ( 
.A(n_2719),
.Y(n_4272)
);

AOI21xp5_ASAP7_75t_L g4273 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_L g4274 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4274)
);

NOR2xp33_ASAP7_75t_L g4275 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4275)
);

NAND2xp5_ASAP7_75t_L g4276 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4276)
);

A2O1A1Ixp33_ASAP7_75t_L g4277 ( 
.A1(n_2737),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4277)
);

AOI21xp5_ASAP7_75t_L g4278 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_L g4279 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4279)
);

NAND2xp5_ASAP7_75t_SL g4280 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4280)
);

BUFx6f_ASAP7_75t_L g4281 ( 
.A(n_2098),
.Y(n_4281)
);

AOI21xp5_ASAP7_75t_L g4282 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4282)
);

NAND2xp5_ASAP7_75t_L g4283 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4283)
);

NAND2xp5_ASAP7_75t_L g4284 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4284)
);

NAND2xp5_ASAP7_75t_L g4285 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4285)
);

NOR2xp33_ASAP7_75t_L g4286 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4286)
);

AOI21xp5_ASAP7_75t_L g4287 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4287)
);

AOI21xp5_ASAP7_75t_L g4288 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4288)
);

AOI21xp5_ASAP7_75t_L g4289 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4289)
);

AOI22xp5_ASAP7_75t_L g4290 ( 
.A1(n_3053),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_4290)
);

OAI21xp33_ASAP7_75t_L g4291 ( 
.A1(n_2374),
.A2(n_1072),
.B(n_1067),
.Y(n_4291)
);

AOI21xp5_ASAP7_75t_L g4292 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4292)
);

NOR2xp33_ASAP7_75t_SL g4293 ( 
.A(n_3040),
.B(n_1067),
.Y(n_4293)
);

AOI22xp5_ASAP7_75t_L g4294 ( 
.A1(n_3053),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_4294)
);

OAI21xp5_ASAP7_75t_L g4295 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4295)
);

AND2x2_ASAP7_75t_L g4296 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4296)
);

NAND2xp33_ASAP7_75t_L g4297 ( 
.A(n_2416),
.B(n_1066),
.Y(n_4297)
);

INVxp67_ASAP7_75t_L g4298 ( 
.A(n_2760),
.Y(n_4298)
);

AOI21xp5_ASAP7_75t_L g4299 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4299)
);

BUFx3_ASAP7_75t_L g4300 ( 
.A(n_2719),
.Y(n_4300)
);

AOI22xp5_ASAP7_75t_L g4301 ( 
.A1(n_3053),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_4301)
);

NOR2xp33_ASAP7_75t_L g4302 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4302)
);

BUFx6f_ASAP7_75t_L g4303 ( 
.A(n_2098),
.Y(n_4303)
);

OR2x6_ASAP7_75t_L g4304 ( 
.A(n_2167),
.B(n_2221),
.Y(n_4304)
);

BUFx2_ASAP7_75t_L g4305 ( 
.A(n_2760),
.Y(n_4305)
);

AOI21xp5_ASAP7_75t_L g4306 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4306)
);

NOR2xp33_ASAP7_75t_L g4307 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4307)
);

NAND2xp5_ASAP7_75t_L g4308 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4308)
);

NOR3xp33_ASAP7_75t_L g4309 ( 
.A(n_2829),
.B(n_788),
.C(n_673),
.Y(n_4309)
);

AOI21xp5_ASAP7_75t_L g4310 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4310)
);

AOI22xp5_ASAP7_75t_L g4311 ( 
.A1(n_3053),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_4311)
);

HB1xp67_ASAP7_75t_L g4312 ( 
.A(n_2144),
.Y(n_4312)
);

A2O1A1Ixp33_ASAP7_75t_L g4313 ( 
.A1(n_2737),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4313)
);

OAI21xp33_ASAP7_75t_L g4314 ( 
.A1(n_2374),
.A2(n_1072),
.B(n_1067),
.Y(n_4314)
);

NAND2xp5_ASAP7_75t_SL g4315 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4315)
);

INVx4_ASAP7_75t_L g4316 ( 
.A(n_2009),
.Y(n_4316)
);

AOI21xp5_ASAP7_75t_L g4317 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4317)
);

AOI21xp5_ASAP7_75t_L g4318 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4318)
);

AOI21xp5_ASAP7_75t_L g4319 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4319)
);

NOR2xp33_ASAP7_75t_L g4320 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4320)
);

NAND2xp5_ASAP7_75t_SL g4321 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4321)
);

OAI22xp5_ASAP7_75t_L g4322 ( 
.A1(n_3040),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_4322)
);

OAI21xp5_ASAP7_75t_L g4323 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4323)
);

NAND2xp5_ASAP7_75t_L g4324 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4324)
);

O2A1O1Ixp33_ASAP7_75t_L g4325 ( 
.A1(n_3040),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4325)
);

NAND2xp5_ASAP7_75t_SL g4326 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4326)
);

NAND2xp5_ASAP7_75t_L g4327 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4327)
);

AOI21xp5_ASAP7_75t_L g4328 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4328)
);

O2A1O1Ixp33_ASAP7_75t_L g4329 ( 
.A1(n_3040),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4329)
);

BUFx3_ASAP7_75t_L g4330 ( 
.A(n_2719),
.Y(n_4330)
);

AOI21xp5_ASAP7_75t_L g4331 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4331)
);

NAND2xp5_ASAP7_75t_L g4332 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4332)
);

INVx3_ASAP7_75t_L g4333 ( 
.A(n_2081),
.Y(n_4333)
);

NAND2xp5_ASAP7_75t_L g4334 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4334)
);

NAND2xp5_ASAP7_75t_SL g4335 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4335)
);

NAND2xp5_ASAP7_75t_L g4336 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_2232),
.Y(n_4337)
);

NAND2xp5_ASAP7_75t_L g4338 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4338)
);

AOI21xp5_ASAP7_75t_L g4339 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_L g4340 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4340)
);

NAND2xp5_ASAP7_75t_SL g4341 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4341)
);

AOI21x1_ASAP7_75t_L g4342 ( 
.A1(n_1988),
.A2(n_2167),
.B(n_1903),
.Y(n_4342)
);

NAND2xp5_ASAP7_75t_L g4343 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4343)
);

OAI321xp33_ASAP7_75t_L g4344 ( 
.A1(n_3040),
.A2(n_1090),
.A3(n_1067),
.B1(n_1101),
.B2(n_1087),
.C(n_1072),
.Y(n_4344)
);

NOR2xp33_ASAP7_75t_L g4345 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4345)
);

NAND2xp5_ASAP7_75t_L g4346 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4346)
);

AOI21xp5_ASAP7_75t_L g4347 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4347)
);

AOI21xp5_ASAP7_75t_L g4348 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4348)
);

AND2x2_ASAP7_75t_L g4349 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4349)
);

O2A1O1Ixp33_ASAP7_75t_L g4350 ( 
.A1(n_3040),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4350)
);

NAND2xp5_ASAP7_75t_L g4351 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4351)
);

NAND2xp5_ASAP7_75t_L g4352 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4352)
);

AOI22xp33_ASAP7_75t_L g4353 ( 
.A1(n_1987),
.A2(n_1072),
.B1(n_1087),
.B2(n_1067),
.Y(n_4353)
);

NAND2xp5_ASAP7_75t_SL g4354 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4354)
);

AND2x2_ASAP7_75t_L g4355 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4355)
);

NAND2xp5_ASAP7_75t_SL g4356 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4356)
);

AOI22xp5_ASAP7_75t_L g4357 ( 
.A1(n_3053),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_4357)
);

AND2x2_ASAP7_75t_L g4358 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4358)
);

AOI21xp5_ASAP7_75t_L g4359 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4359)
);

BUFx4f_ASAP7_75t_L g4360 ( 
.A(n_2566),
.Y(n_4360)
);

BUFx4f_ASAP7_75t_L g4361 ( 
.A(n_2566),
.Y(n_4361)
);

BUFx3_ASAP7_75t_L g4362 ( 
.A(n_2719),
.Y(n_4362)
);

AOI21xp5_ASAP7_75t_L g4363 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4363)
);

OAI21xp5_ASAP7_75t_L g4364 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4364)
);

NAND2xp5_ASAP7_75t_L g4365 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4365)
);

BUFx3_ASAP7_75t_L g4366 ( 
.A(n_2719),
.Y(n_4366)
);

INVx3_ASAP7_75t_L g4367 ( 
.A(n_2081),
.Y(n_4367)
);

NAND2xp5_ASAP7_75t_L g4368 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4368)
);

AO21x1_ASAP7_75t_L g4369 ( 
.A1(n_1988),
.A2(n_2145),
.B(n_2363),
.Y(n_4369)
);

BUFx8_ASAP7_75t_L g4370 ( 
.A(n_2180),
.Y(n_4370)
);

NAND2xp5_ASAP7_75t_L g4371 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4371)
);

AOI21xp5_ASAP7_75t_L g4372 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4372)
);

OAI22xp5_ASAP7_75t_L g4373 ( 
.A1(n_3040),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_4373)
);

CKINVDCx5p33_ASAP7_75t_R g4374 ( 
.A(n_2328),
.Y(n_4374)
);

NAND2xp5_ASAP7_75t_L g4375 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4375)
);

AO21x1_ASAP7_75t_L g4376 ( 
.A1(n_1988),
.A2(n_2145),
.B(n_2363),
.Y(n_4376)
);

AND2x2_ASAP7_75t_L g4377 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_2232),
.Y(n_4378)
);

NAND2xp5_ASAP7_75t_SL g4379 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4379)
);

NAND2xp5_ASAP7_75t_L g4380 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4380)
);

NOR2xp33_ASAP7_75t_L g4381 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4381)
);

NAND2xp33_ASAP7_75t_L g4382 ( 
.A(n_2416),
.B(n_1066),
.Y(n_4382)
);

AO21x1_ASAP7_75t_L g4383 ( 
.A1(n_1988),
.A2(n_2145),
.B(n_2363),
.Y(n_4383)
);

AOI21xp5_ASAP7_75t_L g4384 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4384)
);

O2A1O1Ixp33_ASAP7_75t_L g4385 ( 
.A1(n_3040),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4385)
);

AND2x2_ASAP7_75t_L g4386 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4386)
);

AOI21xp5_ASAP7_75t_L g4387 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4387)
);

AND2x4_ASAP7_75t_L g4388 ( 
.A(n_2098),
.B(n_2221),
.Y(n_4388)
);

AOI21xp5_ASAP7_75t_L g4389 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4389)
);

AOI21xp5_ASAP7_75t_L g4390 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4390)
);

AOI21xp5_ASAP7_75t_L g4391 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_2232),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_2232),
.Y(n_4393)
);

HB1xp67_ASAP7_75t_L g4394 ( 
.A(n_2144),
.Y(n_4394)
);

NAND2xp5_ASAP7_75t_L g4395 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4395)
);

NAND2xp5_ASAP7_75t_L g4396 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_2232),
.Y(n_4397)
);

AO21x1_ASAP7_75t_L g4398 ( 
.A1(n_1988),
.A2(n_2145),
.B(n_2363),
.Y(n_4398)
);

NAND2xp5_ASAP7_75t_L g4399 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4399)
);

AOI21xp5_ASAP7_75t_L g4400 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4400)
);

NAND2xp5_ASAP7_75t_L g4401 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4401)
);

AOI21xp5_ASAP7_75t_L g4402 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4402)
);

AOI21xp33_ASAP7_75t_L g4403 ( 
.A1(n_2374),
.A2(n_1072),
.B(n_1067),
.Y(n_4403)
);

BUFx3_ASAP7_75t_L g4404 ( 
.A(n_2719),
.Y(n_4404)
);

NOR2xp33_ASAP7_75t_SL g4405 ( 
.A(n_3040),
.B(n_1067),
.Y(n_4405)
);

NOR2x1_ASAP7_75t_L g4406 ( 
.A(n_2145),
.B(n_2203),
.Y(n_4406)
);

NOR2xp33_ASAP7_75t_L g4407 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4407)
);

NAND2xp5_ASAP7_75t_L g4408 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4408)
);

AOI21xp5_ASAP7_75t_L g4409 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4409)
);

AOI21xp5_ASAP7_75t_L g4410 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4410)
);

NAND2xp5_ASAP7_75t_L g4411 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4411)
);

O2A1O1Ixp33_ASAP7_75t_L g4412 ( 
.A1(n_3040),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4412)
);

NOR2xp33_ASAP7_75t_L g4413 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4413)
);

OR2x6_ASAP7_75t_L g4414 ( 
.A(n_2167),
.B(n_2221),
.Y(n_4414)
);

AOI21xp5_ASAP7_75t_L g4415 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4415)
);

NOR3xp33_ASAP7_75t_L g4416 ( 
.A(n_2829),
.B(n_788),
.C(n_673),
.Y(n_4416)
);

BUFx2_ASAP7_75t_L g4417 ( 
.A(n_2760),
.Y(n_4417)
);

AOI21x1_ASAP7_75t_L g4418 ( 
.A1(n_1988),
.A2(n_2167),
.B(n_1903),
.Y(n_4418)
);

AND2x2_ASAP7_75t_L g4419 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4419)
);

INVxp67_ASAP7_75t_SL g4420 ( 
.A(n_2760),
.Y(n_4420)
);

NAND2xp5_ASAP7_75t_SL g4421 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4421)
);

NAND2xp5_ASAP7_75t_L g4422 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4422)
);

NAND2xp5_ASAP7_75t_L g4423 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4423)
);

NAND2xp5_ASAP7_75t_L g4424 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4424)
);

AOI21xp5_ASAP7_75t_L g4425 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4425)
);

AOI21xp5_ASAP7_75t_L g4426 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4426)
);

OAI22xp5_ASAP7_75t_L g4427 ( 
.A1(n_3040),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_4427)
);

INVx2_ASAP7_75t_SL g4428 ( 
.A(n_2054),
.Y(n_4428)
);

AOI21xp5_ASAP7_75t_L g4429 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4429)
);

AOI33xp33_ASAP7_75t_L g4430 ( 
.A1(n_2703),
.A2(n_1136),
.A3(n_1155),
.B1(n_1209),
.B2(n_1205),
.B3(n_1066),
.Y(n_4430)
);

NOR2xp67_ASAP7_75t_SL g4431 ( 
.A(n_2009),
.B(n_2743),
.Y(n_4431)
);

OAI21xp33_ASAP7_75t_L g4432 ( 
.A1(n_2374),
.A2(n_1072),
.B(n_1067),
.Y(n_4432)
);

OAI21xp5_ASAP7_75t_L g4433 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4433)
);

OAI22xp5_ASAP7_75t_L g4434 ( 
.A1(n_3040),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_4434)
);

AOI22xp5_ASAP7_75t_L g4435 ( 
.A1(n_3053),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_4435)
);

NAND2xp5_ASAP7_75t_L g4436 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4436)
);

NAND2xp5_ASAP7_75t_L g4437 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4437)
);

OAI22xp5_ASAP7_75t_L g4438 ( 
.A1(n_3040),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_4438)
);

NAND2xp5_ASAP7_75t_L g4439 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4439)
);

AOI22xp5_ASAP7_75t_L g4440 ( 
.A1(n_3053),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_4440)
);

NOR2xp33_ASAP7_75t_L g4441 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4441)
);

A2O1A1Ixp33_ASAP7_75t_L g4442 ( 
.A1(n_2737),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4442)
);

NAND2xp5_ASAP7_75t_L g4443 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4443)
);

HB1xp67_ASAP7_75t_L g4444 ( 
.A(n_2144),
.Y(n_4444)
);

INVx1_ASAP7_75t_L g4445 ( 
.A(n_2232),
.Y(n_4445)
);

AOI21xp5_ASAP7_75t_L g4446 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4446)
);

NAND2xp5_ASAP7_75t_L g4447 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4447)
);

AOI21xp5_ASAP7_75t_L g4448 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4448)
);

NAND2xp5_ASAP7_75t_L g4449 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4449)
);

OAI21xp5_ASAP7_75t_L g4450 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4450)
);

AOI21x1_ASAP7_75t_L g4451 ( 
.A1(n_1988),
.A2(n_2167),
.B(n_1903),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_SL g4452 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4452)
);

NAND2xp5_ASAP7_75t_L g4453 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4453)
);

BUFx2_ASAP7_75t_L g4454 ( 
.A(n_2760),
.Y(n_4454)
);

BUFx3_ASAP7_75t_L g4455 ( 
.A(n_2719),
.Y(n_4455)
);

AOI21xp5_ASAP7_75t_L g4456 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4456)
);

NAND2xp5_ASAP7_75t_L g4457 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4457)
);

AOI21xp5_ASAP7_75t_L g4458 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4458)
);

OAI21xp5_ASAP7_75t_L g4459 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4459)
);

NOR2xp33_ASAP7_75t_L g4460 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4460)
);

OAI21xp5_ASAP7_75t_L g4461 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4461)
);

XOR2x2_ASAP7_75t_L g4462 ( 
.A(n_3049),
.B(n_1993),
.Y(n_4462)
);

NOR2xp33_ASAP7_75t_L g4463 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4463)
);

CKINVDCx14_ASAP7_75t_R g4464 ( 
.A(n_2172),
.Y(n_4464)
);

OAI321xp33_ASAP7_75t_L g4465 ( 
.A1(n_3040),
.A2(n_1090),
.A3(n_1067),
.B1(n_1101),
.B2(n_1087),
.C(n_1072),
.Y(n_4465)
);

NAND2xp5_ASAP7_75t_SL g4466 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4466)
);

AND2x2_ASAP7_75t_L g4467 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4467)
);

BUFx12f_ASAP7_75t_L g4468 ( 
.A(n_2328),
.Y(n_4468)
);

O2A1O1Ixp33_ASAP7_75t_L g4469 ( 
.A1(n_3040),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4469)
);

AND2x2_ASAP7_75t_L g4470 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4470)
);

AND2x2_ASAP7_75t_L g4471 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4471)
);

AOI21xp5_ASAP7_75t_L g4472 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4472)
);

AOI21xp5_ASAP7_75t_L g4473 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4473)
);

OAI21xp5_ASAP7_75t_L g4474 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4474)
);

OAI22xp5_ASAP7_75t_L g4475 ( 
.A1(n_3040),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_4475)
);

AND2x2_ASAP7_75t_L g4476 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4476)
);

INVx1_ASAP7_75t_L g4477 ( 
.A(n_2232),
.Y(n_4477)
);

NOR3xp33_ASAP7_75t_L g4478 ( 
.A(n_2829),
.B(n_788),
.C(n_673),
.Y(n_4478)
);

NAND2xp5_ASAP7_75t_L g4479 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4479)
);

NAND2xp5_ASAP7_75t_L g4480 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4480)
);

OAI21xp5_ASAP7_75t_L g4481 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4481)
);

NOR2xp33_ASAP7_75t_L g4482 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4482)
);

AOI22xp5_ASAP7_75t_L g4483 ( 
.A1(n_3053),
.A2(n_1067),
.B1(n_1087),
.B2(n_1072),
.Y(n_4483)
);

INVxp67_ASAP7_75t_L g4484 ( 
.A(n_2760),
.Y(n_4484)
);

OAI321xp33_ASAP7_75t_L g4485 ( 
.A1(n_3040),
.A2(n_1090),
.A3(n_1067),
.B1(n_1101),
.B2(n_1087),
.C(n_1072),
.Y(n_4485)
);

NAND2xp5_ASAP7_75t_SL g4486 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4486)
);

NOR2xp33_ASAP7_75t_L g4487 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4487)
);

NOR2xp33_ASAP7_75t_L g4488 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4488)
);

INVx1_ASAP7_75t_L g4489 ( 
.A(n_2232),
.Y(n_4489)
);

AO21x1_ASAP7_75t_L g4490 ( 
.A1(n_1988),
.A2(n_2145),
.B(n_2363),
.Y(n_4490)
);

NOR2xp33_ASAP7_75t_L g4491 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4491)
);

AO21x1_ASAP7_75t_L g4492 ( 
.A1(n_1988),
.A2(n_2145),
.B(n_2363),
.Y(n_4492)
);

NOR2xp33_ASAP7_75t_L g4493 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4493)
);

HB1xp67_ASAP7_75t_L g4494 ( 
.A(n_2144),
.Y(n_4494)
);

AND2x2_ASAP7_75t_L g4495 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4495)
);

AOI21xp5_ASAP7_75t_L g4496 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4496)
);

INVx3_ASAP7_75t_L g4497 ( 
.A(n_2081),
.Y(n_4497)
);

AOI21xp5_ASAP7_75t_L g4498 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4498)
);

NAND2xp5_ASAP7_75t_L g4499 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4499)
);

AOI21xp5_ASAP7_75t_L g4500 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4500)
);

AOI21xp5_ASAP7_75t_L g4501 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4501)
);

BUFx6f_ASAP7_75t_L g4502 ( 
.A(n_2098),
.Y(n_4502)
);

INVx1_ASAP7_75t_L g4503 ( 
.A(n_2232),
.Y(n_4503)
);

O2A1O1Ixp33_ASAP7_75t_L g4504 ( 
.A1(n_3040),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4504)
);

AOI21xp5_ASAP7_75t_L g4505 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4505)
);

NOR2xp33_ASAP7_75t_L g4506 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4506)
);

NAND2xp5_ASAP7_75t_L g4507 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4507)
);

INVx1_ASAP7_75t_SL g4508 ( 
.A(n_2144),
.Y(n_4508)
);

NAND2xp5_ASAP7_75t_L g4509 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4509)
);

NAND2xp5_ASAP7_75t_L g4510 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4510)
);

OAI21xp5_ASAP7_75t_L g4511 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4511)
);

OAI21xp5_ASAP7_75t_L g4512 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4512)
);

HB1xp67_ASAP7_75t_L g4513 ( 
.A(n_2144),
.Y(n_4513)
);

OAI21xp33_ASAP7_75t_L g4514 ( 
.A1(n_2374),
.A2(n_1072),
.B(n_1067),
.Y(n_4514)
);

INVx1_ASAP7_75t_L g4515 ( 
.A(n_2232),
.Y(n_4515)
);

NAND2xp5_ASAP7_75t_SL g4516 ( 
.A(n_2374),
.B(n_1096),
.Y(n_4516)
);

O2A1O1Ixp33_ASAP7_75t_L g4517 ( 
.A1(n_3040),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4517)
);

NAND2xp5_ASAP7_75t_L g4518 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4518)
);

OAI21xp33_ASAP7_75t_L g4519 ( 
.A1(n_2374),
.A2(n_1072),
.B(n_1067),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_L g4520 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4520)
);

OAI21xp5_ASAP7_75t_L g4521 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4521)
);

NAND2xp5_ASAP7_75t_L g4522 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4522)
);

OAI21xp5_ASAP7_75t_L g4523 ( 
.A1(n_2393),
.A2(n_2829),
.B(n_2424),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_2232),
.Y(n_4524)
);

NAND2xp5_ASAP7_75t_L g4525 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4525)
);

AOI21xp5_ASAP7_75t_L g4526 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4526)
);

AOI21xp5_ASAP7_75t_L g4527 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4527)
);

CKINVDCx6p67_ASAP7_75t_R g4528 ( 
.A(n_2180),
.Y(n_4528)
);

NAND2xp5_ASAP7_75t_L g4529 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_L g4530 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4530)
);

AOI21x1_ASAP7_75t_L g4531 ( 
.A1(n_1988),
.A2(n_2167),
.B(n_1903),
.Y(n_4531)
);

NAND2xp5_ASAP7_75t_L g4532 ( 
.A(n_2135),
.B(n_2050),
.Y(n_4532)
);

BUFx6f_ASAP7_75t_L g4533 ( 
.A(n_2098),
.Y(n_4533)
);

O2A1O1Ixp33_ASAP7_75t_SL g4534 ( 
.A1(n_2383),
.A2(n_1719),
.B(n_1866),
.C(n_1779),
.Y(n_4534)
);

BUFx3_ASAP7_75t_L g4535 ( 
.A(n_2719),
.Y(n_4535)
);

A2O1A1Ixp33_ASAP7_75t_L g4536 ( 
.A1(n_2737),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4536)
);

INVx4_ASAP7_75t_L g4537 ( 
.A(n_2009),
.Y(n_4537)
);

O2A1O1Ixp33_ASAP7_75t_L g4538 ( 
.A1(n_3040),
.A2(n_1072),
.B(n_1087),
.C(n_1067),
.Y(n_4538)
);

INVx3_ASAP7_75t_L g4539 ( 
.A(n_2081),
.Y(n_4539)
);

AND2x2_ASAP7_75t_L g4540 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4540)
);

NAND2xp5_ASAP7_75t_L g4541 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4541)
);

BUFx6f_ASAP7_75t_L g4542 ( 
.A(n_2098),
.Y(n_4542)
);

AND2x2_ASAP7_75t_L g4543 ( 
.A(n_2549),
.B(n_2780),
.Y(n_4543)
);

AOI21xp5_ASAP7_75t_L g4544 ( 
.A1(n_2568),
.A2(n_2613),
.B(n_2586),
.Y(n_4544)
);

NOR2xp33_ASAP7_75t_L g4545 ( 
.A(n_2025),
.B(n_1067),
.Y(n_4545)
);

NAND2xp5_ASAP7_75t_L g4546 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4546)
);

INVxp67_ASAP7_75t_L g4547 ( 
.A(n_2760),
.Y(n_4547)
);

NAND2xp5_ASAP7_75t_L g4548 ( 
.A(n_2091),
.B(n_1067),
.Y(n_4548)
);

AOI21x1_ASAP7_75t_L g4549 ( 
.A1(n_1988),
.A2(n_2167),
.B(n_1903),
.Y(n_4549)
);

CKINVDCx20_ASAP7_75t_R g4550 ( 
.A(n_2480),
.Y(n_4550)
);

INVx2_ASAP7_75t_L g4551 ( 
.A(n_3694),
.Y(n_4551)
);

INVx1_ASAP7_75t_L g4552 ( 
.A(n_3694),
.Y(n_4552)
);

INVx1_ASAP7_75t_L g4553 ( 
.A(n_3563),
.Y(n_4553)
);

INVx2_ASAP7_75t_L g4554 ( 
.A(n_3564),
.Y(n_4554)
);

INVxp33_ASAP7_75t_L g4555 ( 
.A(n_3655),
.Y(n_4555)
);

NAND2xp5_ASAP7_75t_L g4556 ( 
.A(n_3170),
.B(n_3182),
.Y(n_4556)
);

HB1xp67_ASAP7_75t_L g4557 ( 
.A(n_3419),
.Y(n_4557)
);

CKINVDCx20_ASAP7_75t_R g4558 ( 
.A(n_3341),
.Y(n_4558)
);

INVx1_ASAP7_75t_L g4559 ( 
.A(n_3563),
.Y(n_4559)
);

AND2x4_ASAP7_75t_L g4560 ( 
.A(n_3541),
.B(n_3559),
.Y(n_4560)
);

INVx1_ASAP7_75t_L g4561 ( 
.A(n_3564),
.Y(n_4561)
);

AND3x1_ASAP7_75t_SL g4562 ( 
.A(n_3582),
.B(n_3415),
.C(n_4251),
.Y(n_4562)
);

BUFx12f_ASAP7_75t_L g4563 ( 
.A(n_3830),
.Y(n_4563)
);

AND2x4_ASAP7_75t_L g4564 ( 
.A(n_3541),
.B(n_3559),
.Y(n_4564)
);

INVx2_ASAP7_75t_L g4565 ( 
.A(n_3580),
.Y(n_4565)
);

AOI22xp33_ASAP7_75t_L g4566 ( 
.A1(n_3243),
.A2(n_3271),
.B1(n_3373),
.B2(n_3197),
.Y(n_4566)
);

INVx1_ASAP7_75t_L g4567 ( 
.A(n_3580),
.Y(n_4567)
);

BUFx6f_ASAP7_75t_L g4568 ( 
.A(n_3541),
.Y(n_4568)
);

BUFx3_ASAP7_75t_L g4569 ( 
.A(n_3541),
.Y(n_4569)
);

NAND2xp5_ASAP7_75t_L g4570 ( 
.A(n_3170),
.B(n_3182),
.Y(n_4570)
);

INVx2_ASAP7_75t_L g4571 ( 
.A(n_3705),
.Y(n_4571)
);

INVx2_ASAP7_75t_SL g4572 ( 
.A(n_3541),
.Y(n_4572)
);

HB1xp67_ASAP7_75t_L g4573 ( 
.A(n_3419),
.Y(n_4573)
);

INVx2_ASAP7_75t_L g4574 ( 
.A(n_3705),
.Y(n_4574)
);

HB1xp67_ASAP7_75t_L g4575 ( 
.A(n_3204),
.Y(n_4575)
);

NAND2x1p5_ASAP7_75t_L g4576 ( 
.A(n_4406),
.B(n_3195),
.Y(n_4576)
);

BUFx3_ASAP7_75t_L g4577 ( 
.A(n_3541),
.Y(n_4577)
);

CKINVDCx5p33_ASAP7_75t_R g4578 ( 
.A(n_3977),
.Y(n_4578)
);

OAI22xp5_ASAP7_75t_L g4579 ( 
.A1(n_3983),
.A2(n_4224),
.B1(n_4353),
.B2(n_4018),
.Y(n_4579)
);

INVx2_ASAP7_75t_SL g4580 ( 
.A(n_3559),
.Y(n_4580)
);

AND2x2_ASAP7_75t_L g4581 ( 
.A(n_3162),
.B(n_3165),
.Y(n_4581)
);

INVx1_ASAP7_75t_L g4582 ( 
.A(n_3204),
.Y(n_4582)
);

BUFx3_ASAP7_75t_L g4583 ( 
.A(n_3559),
.Y(n_4583)
);

BUFx3_ASAP7_75t_L g4584 ( 
.A(n_3561),
.Y(n_4584)
);

OAI21x1_ASAP7_75t_L g4585 ( 
.A1(n_3158),
.A2(n_3171),
.B(n_3167),
.Y(n_4585)
);

INVx2_ASAP7_75t_L g4586 ( 
.A(n_3450),
.Y(n_4586)
);

INVx1_ASAP7_75t_SL g4587 ( 
.A(n_3342),
.Y(n_4587)
);

NAND2xp5_ASAP7_75t_L g4588 ( 
.A(n_3170),
.B(n_3186),
.Y(n_4588)
);

NAND2xp5_ASAP7_75t_L g4589 ( 
.A(n_3186),
.B(n_3284),
.Y(n_4589)
);

HB1xp67_ASAP7_75t_L g4590 ( 
.A(n_3329),
.Y(n_4590)
);

INVx2_ASAP7_75t_L g4591 ( 
.A(n_3450),
.Y(n_4591)
);

NAND2xp5_ASAP7_75t_L g4592 ( 
.A(n_3284),
.B(n_3406),
.Y(n_4592)
);

NAND2xp5_ASAP7_75t_L g4593 ( 
.A(n_3410),
.B(n_3344),
.Y(n_4593)
);

A2O1A1Ixp33_ASAP7_75t_L g4594 ( 
.A1(n_3836),
.A2(n_3847),
.B(n_3949),
.C(n_3887),
.Y(n_4594)
);

BUFx4f_ASAP7_75t_SL g4595 ( 
.A(n_3337),
.Y(n_4595)
);

INVxp67_ASAP7_75t_L g4596 ( 
.A(n_3179),
.Y(n_4596)
);

HB1xp67_ASAP7_75t_L g4597 ( 
.A(n_3329),
.Y(n_4597)
);

NAND2xp5_ASAP7_75t_L g4598 ( 
.A(n_3344),
.B(n_3384),
.Y(n_4598)
);

NOR2xp33_ASAP7_75t_L g4599 ( 
.A(n_3954),
.B(n_4293),
.Y(n_4599)
);

NAND2xp5_ASAP7_75t_L g4600 ( 
.A(n_3384),
.B(n_3418),
.Y(n_4600)
);

BUFx2_ASAP7_75t_L g4601 ( 
.A(n_3875),
.Y(n_4601)
);

NAND2xp5_ASAP7_75t_L g4602 ( 
.A(n_3418),
.B(n_3312),
.Y(n_4602)
);

BUFx4f_ASAP7_75t_L g4603 ( 
.A(n_3498),
.Y(n_4603)
);

INVx2_ASAP7_75t_L g4604 ( 
.A(n_3473),
.Y(n_4604)
);

NAND2xp5_ASAP7_75t_L g4605 ( 
.A(n_3312),
.B(n_3164),
.Y(n_4605)
);

INVx2_ASAP7_75t_L g4606 ( 
.A(n_3473),
.Y(n_4606)
);

BUFx3_ASAP7_75t_L g4607 ( 
.A(n_3561),
.Y(n_4607)
);

INVx2_ASAP7_75t_L g4608 ( 
.A(n_3438),
.Y(n_4608)
);

NAND2xp5_ASAP7_75t_L g4609 ( 
.A(n_3164),
.B(n_3192),
.Y(n_4609)
);

INVx2_ASAP7_75t_L g4610 ( 
.A(n_3438),
.Y(n_4610)
);

NAND2xp5_ASAP7_75t_SL g4611 ( 
.A(n_3954),
.B(n_4293),
.Y(n_4611)
);

OR2x6_ASAP7_75t_L g4612 ( 
.A(n_3793),
.B(n_3799),
.Y(n_4612)
);

NAND2xp5_ASAP7_75t_L g4613 ( 
.A(n_3192),
.B(n_3196),
.Y(n_4613)
);

NAND2xp5_ASAP7_75t_L g4614 ( 
.A(n_3196),
.B(n_3218),
.Y(n_4614)
);

O2A1O1Ixp33_ASAP7_75t_L g4615 ( 
.A1(n_3807),
.A2(n_3890),
.B(n_3921),
.C(n_3839),
.Y(n_4615)
);

NAND2xp5_ASAP7_75t_L g4616 ( 
.A(n_3218),
.B(n_3219),
.Y(n_4616)
);

AND2x2_ASAP7_75t_L g4617 ( 
.A(n_3162),
.B(n_3165),
.Y(n_4617)
);

AOI221xp5_ASAP7_75t_L g4618 ( 
.A1(n_3807),
.A2(n_3890),
.B1(n_4035),
.B2(n_3921),
.C(n_3839),
.Y(n_4618)
);

OR2x2_ASAP7_75t_L g4619 ( 
.A(n_3224),
.B(n_3226),
.Y(n_4619)
);

INVxp67_ASAP7_75t_L g4620 ( 
.A(n_3179),
.Y(n_4620)
);

NAND2xp5_ASAP7_75t_L g4621 ( 
.A(n_3219),
.B(n_3223),
.Y(n_4621)
);

OR2x2_ASAP7_75t_L g4622 ( 
.A(n_3224),
.B(n_3226),
.Y(n_4622)
);

BUFx4f_ASAP7_75t_L g4623 ( 
.A(n_3498),
.Y(n_4623)
);

NOR2xp33_ASAP7_75t_SL g4624 ( 
.A(n_4431),
.B(n_4405),
.Y(n_4624)
);

BUFx2_ASAP7_75t_L g4625 ( 
.A(n_3875),
.Y(n_4625)
);

NAND2xp5_ASAP7_75t_L g4626 ( 
.A(n_3223),
.B(n_3521),
.Y(n_4626)
);

NAND2xp5_ASAP7_75t_SL g4627 ( 
.A(n_4405),
.B(n_3814),
.Y(n_4627)
);

NAND2xp5_ASAP7_75t_L g4628 ( 
.A(n_3521),
.B(n_3388),
.Y(n_4628)
);

INVx1_ASAP7_75t_SL g4629 ( 
.A(n_3342),
.Y(n_4629)
);

BUFx12f_ASAP7_75t_L g4630 ( 
.A(n_3830),
.Y(n_4630)
);

INVx2_ASAP7_75t_SL g4631 ( 
.A(n_3561),
.Y(n_4631)
);

AOI22xp5_ASAP7_75t_L g4632 ( 
.A1(n_4035),
.A2(n_4071),
.B1(n_4074),
.B2(n_4067),
.Y(n_4632)
);

CKINVDCx5p33_ASAP7_75t_R g4633 ( 
.A(n_3977),
.Y(n_4633)
);

AOI22xp5_ASAP7_75t_L g4634 ( 
.A1(n_4067),
.A2(n_4074),
.B1(n_4168),
.B2(n_4071),
.Y(n_4634)
);

HB1xp67_ASAP7_75t_L g4635 ( 
.A(n_3329),
.Y(n_4635)
);

NAND2xp5_ASAP7_75t_L g4636 ( 
.A(n_3521),
.B(n_3388),
.Y(n_4636)
);

NAND2xp5_ASAP7_75t_L g4637 ( 
.A(n_3322),
.B(n_3340),
.Y(n_4637)
);

NOR2xp33_ASAP7_75t_L g4638 ( 
.A(n_3814),
.B(n_3936),
.Y(n_4638)
);

OAI22xp5_ASAP7_75t_L g4639 ( 
.A1(n_3936),
.A2(n_3987),
.B1(n_4048),
.B2(n_3984),
.Y(n_4639)
);

AND2x4_ASAP7_75t_L g4640 ( 
.A(n_3568),
.B(n_3567),
.Y(n_4640)
);

AOI22xp33_ASAP7_75t_SL g4641 ( 
.A1(n_3290),
.A2(n_3313),
.B1(n_3315),
.B2(n_3308),
.Y(n_4641)
);

NAND2xp33_ASAP7_75t_R g4642 ( 
.A(n_3308),
.B(n_3329),
.Y(n_4642)
);

NAND2xp5_ASAP7_75t_L g4643 ( 
.A(n_3322),
.B(n_3340),
.Y(n_4643)
);

NAND2xp5_ASAP7_75t_L g4644 ( 
.A(n_3400),
.B(n_3350),
.Y(n_4644)
);

NAND2xp5_ASAP7_75t_L g4645 ( 
.A(n_3400),
.B(n_3350),
.Y(n_4645)
);

NAND2xp5_ASAP7_75t_L g4646 ( 
.A(n_3156),
.B(n_3176),
.Y(n_4646)
);

AND2x2_ASAP7_75t_L g4647 ( 
.A(n_3794),
.B(n_3812),
.Y(n_4647)
);

AOI22xp5_ASAP7_75t_L g4648 ( 
.A1(n_4168),
.A2(n_4373),
.B1(n_4427),
.B2(n_4322),
.Y(n_4648)
);

NAND2xp5_ASAP7_75t_L g4649 ( 
.A(n_3156),
.B(n_3176),
.Y(n_4649)
);

NAND2xp5_ASAP7_75t_L g4650 ( 
.A(n_3795),
.B(n_3796),
.Y(n_4650)
);

OR2x4_ASAP7_75t_L g4651 ( 
.A(n_4040),
.B(n_4094),
.Y(n_4651)
);

AOI22xp5_ASAP7_75t_L g4652 ( 
.A1(n_4322),
.A2(n_4427),
.B1(n_4434),
.B2(n_4373),
.Y(n_4652)
);

HB1xp67_ASAP7_75t_L g4653 ( 
.A(n_3817),
.Y(n_4653)
);

CKINVDCx5p33_ASAP7_75t_R g4654 ( 
.A(n_3776),
.Y(n_4654)
);

BUFx3_ASAP7_75t_L g4655 ( 
.A(n_3195),
.Y(n_4655)
);

NOR2xp33_ASAP7_75t_L g4656 ( 
.A(n_3984),
.B(n_3987),
.Y(n_4656)
);

BUFx12f_ASAP7_75t_L g4657 ( 
.A(n_3830),
.Y(n_4657)
);

BUFx6f_ASAP7_75t_L g4658 ( 
.A(n_3195),
.Y(n_4658)
);

INVx2_ASAP7_75t_SL g4659 ( 
.A(n_3195),
.Y(n_4659)
);

CKINVDCx16_ASAP7_75t_R g4660 ( 
.A(n_3513),
.Y(n_4660)
);

NAND2x1p5_ASAP7_75t_L g4661 ( 
.A(n_4406),
.B(n_3431),
.Y(n_4661)
);

NAND2xp5_ASAP7_75t_L g4662 ( 
.A(n_3795),
.B(n_3796),
.Y(n_4662)
);

NAND2xp5_ASAP7_75t_L g4663 ( 
.A(n_3797),
.B(n_3798),
.Y(n_4663)
);

HB1xp67_ASAP7_75t_L g4664 ( 
.A(n_3817),
.Y(n_4664)
);

AOI22xp5_ASAP7_75t_L g4665 ( 
.A1(n_4434),
.A2(n_4475),
.B1(n_4438),
.B2(n_4290),
.Y(n_4665)
);

BUFx12f_ASAP7_75t_L g4666 ( 
.A(n_3830),
.Y(n_4666)
);

AO22x1_ASAP7_75t_L g4667 ( 
.A1(n_3210),
.A2(n_3475),
.B1(n_3445),
.B2(n_3439),
.Y(n_4667)
);

HB1xp67_ASAP7_75t_L g4668 ( 
.A(n_3853),
.Y(n_4668)
);

AOI22xp5_ASAP7_75t_L g4669 ( 
.A1(n_4438),
.A2(n_4475),
.B1(n_4290),
.B2(n_4294),
.Y(n_4669)
);

INVx4_ASAP7_75t_L g4670 ( 
.A(n_3429),
.Y(n_4670)
);

AOI22xp5_ASAP7_75t_L g4671 ( 
.A1(n_4048),
.A2(n_4301),
.B1(n_4311),
.B2(n_4294),
.Y(n_4671)
);

INVx4_ASAP7_75t_L g4672 ( 
.A(n_3429),
.Y(n_4672)
);

BUFx2_ASAP7_75t_L g4673 ( 
.A(n_3875),
.Y(n_4673)
);

BUFx8_ASAP7_75t_L g4674 ( 
.A(n_3461),
.Y(n_4674)
);

AOI22xp5_ASAP7_75t_L g4675 ( 
.A1(n_4301),
.A2(n_4357),
.B1(n_4435),
.B2(n_4311),
.Y(n_4675)
);

NAND3xp33_ASAP7_75t_SL g4676 ( 
.A(n_3960),
.B(n_4129),
.C(n_4033),
.Y(n_4676)
);

NAND2xp5_ASAP7_75t_L g4677 ( 
.A(n_3797),
.B(n_3798),
.Y(n_4677)
);

CKINVDCx5p33_ASAP7_75t_R g4678 ( 
.A(n_3899),
.Y(n_4678)
);

BUFx2_ASAP7_75t_L g4679 ( 
.A(n_3875),
.Y(n_4679)
);

AND2x2_ASAP7_75t_L g4680 ( 
.A(n_3794),
.B(n_3812),
.Y(n_4680)
);

CKINVDCx5p33_ASAP7_75t_R g4681 ( 
.A(n_4200),
.Y(n_4681)
);

BUFx2_ASAP7_75t_L g4682 ( 
.A(n_3875),
.Y(n_4682)
);

NAND2xp5_ASAP7_75t_L g4683 ( 
.A(n_3800),
.B(n_3806),
.Y(n_4683)
);

NOR2x1_ASAP7_75t_L g4684 ( 
.A(n_3317),
.B(n_3365),
.Y(n_4684)
);

BUFx4f_ASAP7_75t_L g4685 ( 
.A(n_3498),
.Y(n_4685)
);

NAND2xp5_ASAP7_75t_L g4686 ( 
.A(n_3800),
.B(n_3806),
.Y(n_4686)
);

NAND2xp5_ASAP7_75t_L g4687 ( 
.A(n_3809),
.B(n_3822),
.Y(n_4687)
);

AOI22xp33_ASAP7_75t_L g4688 ( 
.A1(n_3243),
.A2(n_3271),
.B1(n_3333),
.B2(n_3318),
.Y(n_4688)
);

BUFx3_ASAP7_75t_L g4689 ( 
.A(n_3431),
.Y(n_4689)
);

BUFx3_ASAP7_75t_L g4690 ( 
.A(n_3431),
.Y(n_4690)
);

NOR2xp33_ASAP7_75t_L g4691 ( 
.A(n_4357),
.B(n_4435),
.Y(n_4691)
);

AOI221xp5_ASAP7_75t_L g4692 ( 
.A1(n_4160),
.A2(n_4243),
.B1(n_4329),
.B2(n_4325),
.C(n_4166),
.Y(n_4692)
);

NAND2xp5_ASAP7_75t_L g4693 ( 
.A(n_3809),
.B(n_3822),
.Y(n_4693)
);

A2O1A1Ixp33_ASAP7_75t_L g4694 ( 
.A1(n_4350),
.A2(n_4412),
.B(n_4469),
.C(n_4385),
.Y(n_4694)
);

BUFx6f_ASAP7_75t_L g4695 ( 
.A(n_3431),
.Y(n_4695)
);

BUFx6f_ASAP7_75t_L g4696 ( 
.A(n_3441),
.Y(n_4696)
);

NAND2xp5_ASAP7_75t_L g4697 ( 
.A(n_3828),
.B(n_3974),
.Y(n_4697)
);

NAND2xp5_ASAP7_75t_L g4698 ( 
.A(n_3828),
.B(n_3974),
.Y(n_4698)
);

AOI21xp5_ASAP7_75t_L g4699 ( 
.A1(n_3815),
.A2(n_3818),
.B(n_3816),
.Y(n_4699)
);

AND2x2_ASAP7_75t_L g4700 ( 
.A(n_3855),
.B(n_3894),
.Y(n_4700)
);

BUFx6f_ASAP7_75t_L g4701 ( 
.A(n_3441),
.Y(n_4701)
);

CKINVDCx5p33_ASAP7_75t_R g4702 ( 
.A(n_4216),
.Y(n_4702)
);

OR2x6_ASAP7_75t_L g4703 ( 
.A(n_3825),
.B(n_3826),
.Y(n_4703)
);

INVxp67_ASAP7_75t_SL g4704 ( 
.A(n_3217),
.Y(n_4704)
);

BUFx3_ASAP7_75t_L g4705 ( 
.A(n_3441),
.Y(n_4705)
);

NAND2xp5_ASAP7_75t_SL g4706 ( 
.A(n_4440),
.B(n_4483),
.Y(n_4706)
);

BUFx2_ASAP7_75t_L g4707 ( 
.A(n_3918),
.Y(n_4707)
);

NAND2xp5_ASAP7_75t_L g4708 ( 
.A(n_3978),
.B(n_3982),
.Y(n_4708)
);

HB1xp67_ASAP7_75t_L g4709 ( 
.A(n_3853),
.Y(n_4709)
);

NAND2xp5_ASAP7_75t_L g4710 ( 
.A(n_3978),
.B(n_3982),
.Y(n_4710)
);

NAND2xp5_ASAP7_75t_L g4711 ( 
.A(n_3991),
.B(n_4001),
.Y(n_4711)
);

OAI22xp5_ASAP7_75t_SL g4712 ( 
.A1(n_3257),
.A2(n_3300),
.B1(n_3163),
.B2(n_3191),
.Y(n_4712)
);

AND2x4_ASAP7_75t_L g4713 ( 
.A(n_3567),
.B(n_3918),
.Y(n_4713)
);

INVx1_ASAP7_75t_SL g4714 ( 
.A(n_3343),
.Y(n_4714)
);

AND2x2_ASAP7_75t_L g4715 ( 
.A(n_3896),
.B(n_3902),
.Y(n_4715)
);

HB1xp67_ASAP7_75t_L g4716 ( 
.A(n_3941),
.Y(n_4716)
);

BUFx12f_ASAP7_75t_L g4717 ( 
.A(n_4370),
.Y(n_4717)
);

INVx1_ASAP7_75t_SL g4718 ( 
.A(n_3343),
.Y(n_4718)
);

INVx5_ASAP7_75t_L g4719 ( 
.A(n_3918),
.Y(n_4719)
);

BUFx3_ASAP7_75t_L g4720 ( 
.A(n_3441),
.Y(n_4720)
);

NOR2xp33_ASAP7_75t_R g4721 ( 
.A(n_4464),
.B(n_3220),
.Y(n_4721)
);

NOR2xp33_ASAP7_75t_L g4722 ( 
.A(n_4440),
.B(n_4483),
.Y(n_4722)
);

NAND2xp5_ASAP7_75t_L g4723 ( 
.A(n_3991),
.B(n_4001),
.Y(n_4723)
);

INVx4_ASAP7_75t_L g4724 ( 
.A(n_3429),
.Y(n_4724)
);

NAND2xp5_ASAP7_75t_L g4725 ( 
.A(n_4011),
.B(n_4013),
.Y(n_4725)
);

OR2x6_ASAP7_75t_L g4726 ( 
.A(n_3843),
.B(n_3844),
.Y(n_4726)
);

AND3x1_ASAP7_75t_L g4727 ( 
.A(n_3354),
.B(n_3380),
.C(n_3358),
.Y(n_4727)
);

NAND2xp5_ASAP7_75t_SL g4728 ( 
.A(n_4251),
.B(n_4344),
.Y(n_4728)
);

BUFx2_ASAP7_75t_L g4729 ( 
.A(n_3918),
.Y(n_4729)
);

BUFx3_ASAP7_75t_L g4730 ( 
.A(n_3455),
.Y(n_4730)
);

BUFx6f_ASAP7_75t_L g4731 ( 
.A(n_3455),
.Y(n_4731)
);

NAND2x1p5_ASAP7_75t_L g4732 ( 
.A(n_3455),
.B(n_3833),
.Y(n_4732)
);

BUFx6f_ASAP7_75t_L g4733 ( 
.A(n_3455),
.Y(n_4733)
);

AND2x4_ASAP7_75t_L g4734 ( 
.A(n_3918),
.B(n_4187),
.Y(n_4734)
);

AND3x2_ASAP7_75t_SL g4735 ( 
.A(n_4344),
.B(n_4485),
.C(n_4465),
.Y(n_4735)
);

AND2x4_ASAP7_75t_SL g4736 ( 
.A(n_3202),
.B(n_3850),
.Y(n_4736)
);

NOR2xp33_ASAP7_75t_SL g4737 ( 
.A(n_4431),
.B(n_3513),
.Y(n_4737)
);

AND2x6_ASAP7_75t_SL g4738 ( 
.A(n_3785),
.B(n_3791),
.Y(n_4738)
);

INVx5_ASAP7_75t_L g4739 ( 
.A(n_4187),
.Y(n_4739)
);

AND2x2_ASAP7_75t_L g4740 ( 
.A(n_3896),
.B(n_3902),
.Y(n_4740)
);

A2O1A1Ixp33_ASAP7_75t_L g4741 ( 
.A1(n_4504),
.A2(n_4538),
.B(n_4517),
.C(n_3966),
.Y(n_4741)
);

AND2x2_ASAP7_75t_L g4742 ( 
.A(n_3919),
.B(n_3924),
.Y(n_4742)
);

NOR2xp67_ASAP7_75t_L g4743 ( 
.A(n_3332),
.B(n_3574),
.Y(n_4743)
);

NAND2xp5_ASAP7_75t_L g4744 ( 
.A(n_4011),
.B(n_4013),
.Y(n_4744)
);

BUFx2_ASAP7_75t_R g4745 ( 
.A(n_3402),
.Y(n_4745)
);

AND2x4_ASAP7_75t_L g4746 ( 
.A(n_4187),
.B(n_4304),
.Y(n_4746)
);

AOI21xp5_ASAP7_75t_L g4747 ( 
.A1(n_3845),
.A2(n_3864),
.B(n_3861),
.Y(n_4747)
);

NAND2xp5_ASAP7_75t_SL g4748 ( 
.A(n_4465),
.B(n_4485),
.Y(n_4748)
);

AND2x2_ASAP7_75t_L g4749 ( 
.A(n_3919),
.B(n_3924),
.Y(n_4749)
);

CKINVDCx5p33_ASAP7_75t_R g4750 ( 
.A(n_4374),
.Y(n_4750)
);

O2A1O1Ixp5_ASAP7_75t_L g4751 ( 
.A1(n_3803),
.A2(n_4099),
.B(n_4054),
.C(n_3871),
.Y(n_4751)
);

NAND2xp5_ASAP7_75t_SL g4752 ( 
.A(n_3309),
.B(n_3323),
.Y(n_4752)
);

NAND2xp5_ASAP7_75t_SL g4753 ( 
.A(n_3309),
.B(n_3323),
.Y(n_4753)
);

AOI22xp33_ASAP7_75t_L g4754 ( 
.A1(n_3413),
.A2(n_3428),
.B1(n_3228),
.B2(n_3279),
.Y(n_4754)
);

BUFx3_ASAP7_75t_L g4755 ( 
.A(n_3833),
.Y(n_4755)
);

NAND2xp5_ASAP7_75t_L g4756 ( 
.A(n_4023),
.B(n_4025),
.Y(n_4756)
);

NOR2xp33_ASAP7_75t_L g4757 ( 
.A(n_3209),
.B(n_3263),
.Y(n_4757)
);

AND2x2_ASAP7_75t_L g4758 ( 
.A(n_3956),
.B(n_3970),
.Y(n_4758)
);

AND2x4_ASAP7_75t_L g4759 ( 
.A(n_4187),
.B(n_4304),
.Y(n_4759)
);

AND2x4_ASAP7_75t_L g4760 ( 
.A(n_4187),
.B(n_4304),
.Y(n_4760)
);

NAND2xp5_ASAP7_75t_L g4761 ( 
.A(n_4023),
.B(n_4025),
.Y(n_4761)
);

NAND2xp5_ASAP7_75t_SL g4762 ( 
.A(n_3346),
.B(n_3362),
.Y(n_4762)
);

NAND2x1p5_ASAP7_75t_L g4763 ( 
.A(n_3833),
.B(n_3939),
.Y(n_4763)
);

BUFx6f_ASAP7_75t_L g4764 ( 
.A(n_3833),
.Y(n_4764)
);

BUFx2_ASAP7_75t_L g4765 ( 
.A(n_4304),
.Y(n_4765)
);

INVx5_ASAP7_75t_L g4766 ( 
.A(n_4304),
.Y(n_4766)
);

O2A1O1Ixp33_ASAP7_75t_L g4767 ( 
.A1(n_3237),
.A2(n_3294),
.B(n_3327),
.C(n_3255),
.Y(n_4767)
);

INVxp67_ASAP7_75t_SL g4768 ( 
.A(n_3217),
.Y(n_4768)
);

NAND2xp5_ASAP7_75t_L g4769 ( 
.A(n_4039),
.B(n_4041),
.Y(n_4769)
);

HB1xp67_ASAP7_75t_L g4770 ( 
.A(n_3941),
.Y(n_4770)
);

NAND2xp5_ASAP7_75t_L g4771 ( 
.A(n_4039),
.B(n_4041),
.Y(n_4771)
);

NAND2xp5_ASAP7_75t_L g4772 ( 
.A(n_4055),
.B(n_4057),
.Y(n_4772)
);

NOR2xp33_ASAP7_75t_L g4773 ( 
.A(n_3190),
.B(n_4158),
.Y(n_4773)
);

INVx1_ASAP7_75t_SL g4774 ( 
.A(n_3447),
.Y(n_4774)
);

NAND2xp5_ASAP7_75t_L g4775 ( 
.A(n_4055),
.B(n_4057),
.Y(n_4775)
);

NAND2xp5_ASAP7_75t_L g4776 ( 
.A(n_4065),
.B(n_4069),
.Y(n_4776)
);

BUFx3_ASAP7_75t_L g4777 ( 
.A(n_3939),
.Y(n_4777)
);

BUFx6f_ASAP7_75t_L g4778 ( 
.A(n_3939),
.Y(n_4778)
);

NOR2x1p5_ASAP7_75t_L g4779 ( 
.A(n_4040),
.B(n_4094),
.Y(n_4779)
);

OR2x2_ASAP7_75t_L g4780 ( 
.A(n_3956),
.B(n_3970),
.Y(n_4780)
);

BUFx3_ASAP7_75t_L g4781 ( 
.A(n_3939),
.Y(n_4781)
);

O2A1O1Ixp33_ASAP7_75t_L g4782 ( 
.A1(n_3363),
.A2(n_3371),
.B(n_3392),
.C(n_3389),
.Y(n_4782)
);

OAI22xp5_ASAP7_75t_L g4783 ( 
.A1(n_3820),
.A2(n_3876),
.B1(n_3882),
.B2(n_3846),
.Y(n_4783)
);

NAND3xp33_ASAP7_75t_L g4784 ( 
.A(n_3975),
.B(n_4140),
.C(n_3985),
.Y(n_4784)
);

AOI22xp5_ASAP7_75t_L g4785 ( 
.A1(n_3290),
.A2(n_3805),
.B1(n_3819),
.B2(n_3801),
.Y(n_4785)
);

NAND2xp5_ASAP7_75t_L g4786 ( 
.A(n_4065),
.B(n_4069),
.Y(n_4786)
);

NAND2xp5_ASAP7_75t_SL g4787 ( 
.A(n_3346),
.B(n_3362),
.Y(n_4787)
);

BUFx2_ASAP7_75t_L g4788 ( 
.A(n_4414),
.Y(n_4788)
);

CKINVDCx5p33_ASAP7_75t_R g4789 ( 
.A(n_3293),
.Y(n_4789)
);

NOR2xp33_ASAP7_75t_R g4790 ( 
.A(n_3434),
.B(n_3556),
.Y(n_4790)
);

AND2x4_ASAP7_75t_L g4791 ( 
.A(n_4414),
.B(n_3485),
.Y(n_4791)
);

NOR2xp33_ASAP7_75t_SL g4792 ( 
.A(n_3556),
.B(n_3429),
.Y(n_4792)
);

AOI22xp5_ASAP7_75t_L g4793 ( 
.A1(n_3838),
.A2(n_3904),
.B1(n_3920),
.B2(n_3891),
.Y(n_4793)
);

NAND2xp5_ASAP7_75t_L g4794 ( 
.A(n_4073),
.B(n_4087),
.Y(n_4794)
);

BUFx4f_ASAP7_75t_L g4795 ( 
.A(n_3461),
.Y(n_4795)
);

NAND2xp5_ASAP7_75t_SL g4796 ( 
.A(n_3379),
.B(n_3395),
.Y(n_4796)
);

BUFx6f_ASAP7_75t_L g4797 ( 
.A(n_4360),
.Y(n_4797)
);

AND2x4_ASAP7_75t_L g4798 ( 
.A(n_4414),
.B(n_3488),
.Y(n_4798)
);

NAND2xp5_ASAP7_75t_L g4799 ( 
.A(n_4073),
.B(n_4087),
.Y(n_4799)
);

BUFx6f_ASAP7_75t_L g4800 ( 
.A(n_4360),
.Y(n_4800)
);

AND3x2_ASAP7_75t_SL g4801 ( 
.A(n_3808),
.B(n_3925),
.C(n_3813),
.Y(n_4801)
);

NAND2xp5_ASAP7_75t_L g4802 ( 
.A(n_4091),
.B(n_4092),
.Y(n_4802)
);

INVxp67_ASAP7_75t_SL g4803 ( 
.A(n_3246),
.Y(n_4803)
);

BUFx4f_ASAP7_75t_L g4804 ( 
.A(n_3461),
.Y(n_4804)
);

NAND2xp5_ASAP7_75t_L g4805 ( 
.A(n_4091),
.B(n_4092),
.Y(n_4805)
);

INVx4_ASAP7_75t_L g4806 ( 
.A(n_3429),
.Y(n_4806)
);

NAND2xp5_ASAP7_75t_L g4807 ( 
.A(n_4093),
.B(n_4096),
.Y(n_4807)
);

NOR2xp33_ASAP7_75t_L g4808 ( 
.A(n_3824),
.B(n_3932),
.Y(n_4808)
);

NAND2xp5_ASAP7_75t_L g4809 ( 
.A(n_4093),
.B(n_4096),
.Y(n_4809)
);

NAND2xp5_ASAP7_75t_SL g4810 ( 
.A(n_3379),
.B(n_3395),
.Y(n_4810)
);

INVxp67_ASAP7_75t_L g4811 ( 
.A(n_4142),
.Y(n_4811)
);

O2A1O1Ixp33_ASAP7_75t_L g4812 ( 
.A1(n_3905),
.A2(n_3906),
.B(n_4113),
.C(n_4042),
.Y(n_4812)
);

BUFx2_ASAP7_75t_L g4813 ( 
.A(n_4414),
.Y(n_4813)
);

NOR2x1p5_ASAP7_75t_SL g4814 ( 
.A(n_3203),
.B(n_3239),
.Y(n_4814)
);

AOI22xp5_ASAP7_75t_L g4815 ( 
.A1(n_3945),
.A2(n_3952),
.B1(n_3992),
.B2(n_3946),
.Y(n_4815)
);

NAND2xp5_ASAP7_75t_L g4816 ( 
.A(n_4107),
.B(n_4177),
.Y(n_4816)
);

AND2x4_ASAP7_75t_L g4817 ( 
.A(n_3488),
.B(n_3671),
.Y(n_4817)
);

NAND2xp5_ASAP7_75t_L g4818 ( 
.A(n_4107),
.B(n_4177),
.Y(n_4818)
);

BUFx6f_ASAP7_75t_L g4819 ( 
.A(n_4360),
.Y(n_4819)
);

AOI22xp33_ASAP7_75t_SL g4820 ( 
.A1(n_3315),
.A2(n_3425),
.B1(n_3405),
.B2(n_3325),
.Y(n_4820)
);

BUFx2_ASAP7_75t_L g4821 ( 
.A(n_3581),
.Y(n_4821)
);

NAND2x1_ASAP7_75t_L g4822 ( 
.A(n_3202),
.B(n_3850),
.Y(n_4822)
);

NAND2xp5_ASAP7_75t_L g4823 ( 
.A(n_4178),
.B(n_4179),
.Y(n_4823)
);

INVxp67_ASAP7_75t_SL g4824 ( 
.A(n_3246),
.Y(n_4824)
);

CKINVDCx20_ASAP7_75t_R g4825 ( 
.A(n_4550),
.Y(n_4825)
);

NAND2xp5_ASAP7_75t_L g4826 ( 
.A(n_4178),
.B(n_4179),
.Y(n_4826)
);

NAND2xp5_ASAP7_75t_SL g4827 ( 
.A(n_3361),
.B(n_3377),
.Y(n_4827)
);

BUFx2_ASAP7_75t_L g4828 ( 
.A(n_3581),
.Y(n_4828)
);

NAND2xp5_ASAP7_75t_L g4829 ( 
.A(n_4183),
.B(n_4201),
.Y(n_4829)
);

BUFx4f_ASAP7_75t_SL g4830 ( 
.A(n_3337),
.Y(n_4830)
);

NOR2xp67_ASAP7_75t_L g4831 ( 
.A(n_3515),
.B(n_3486),
.Y(n_4831)
);

AND2x4_ASAP7_75t_L g4832 ( 
.A(n_3671),
.B(n_3202),
.Y(n_4832)
);

NAND2xp5_ASAP7_75t_L g4833 ( 
.A(n_4183),
.B(n_4201),
.Y(n_4833)
);

NAND2xp5_ASAP7_75t_L g4834 ( 
.A(n_4240),
.B(n_4241),
.Y(n_4834)
);

BUFx3_ASAP7_75t_L g4835 ( 
.A(n_4360),
.Y(n_4835)
);

AOI22xp33_ASAP7_75t_L g4836 ( 
.A1(n_3391),
.A2(n_3385),
.B1(n_3466),
.B2(n_3824),
.Y(n_4836)
);

NAND2xp5_ASAP7_75t_L g4837 ( 
.A(n_4240),
.B(n_4241),
.Y(n_4837)
);

INVxp33_ASAP7_75t_L g4838 ( 
.A(n_3572),
.Y(n_4838)
);

NAND2xp5_ASAP7_75t_L g4839 ( 
.A(n_4247),
.B(n_4256),
.Y(n_4839)
);

NAND2xp5_ASAP7_75t_L g4840 ( 
.A(n_4247),
.B(n_4256),
.Y(n_4840)
);

NAND2xp5_ASAP7_75t_L g4841 ( 
.A(n_4258),
.B(n_4261),
.Y(n_4841)
);

AOI22xp5_ASAP7_75t_L g4842 ( 
.A1(n_3995),
.A2(n_4037),
.B1(n_4060),
.B2(n_4047),
.Y(n_4842)
);

O2A1O1Ixp33_ASAP7_75t_L g4843 ( 
.A1(n_4125),
.A2(n_4198),
.B(n_4268),
.C(n_4255),
.Y(n_4843)
);

AOI22xp33_ASAP7_75t_L g4844 ( 
.A1(n_3391),
.A2(n_4012),
.B1(n_4291),
.B2(n_3932),
.Y(n_4844)
);

NAND2xp5_ASAP7_75t_L g4845 ( 
.A(n_4258),
.B(n_4261),
.Y(n_4845)
);

BUFx6f_ASAP7_75t_L g4846 ( 
.A(n_4361),
.Y(n_4846)
);

NAND2xp5_ASAP7_75t_SL g4847 ( 
.A(n_3274),
.B(n_3296),
.Y(n_4847)
);

BUFx2_ASAP7_75t_L g4848 ( 
.A(n_3979),
.Y(n_4848)
);

AND2x4_ASAP7_75t_L g4849 ( 
.A(n_3202),
.B(n_3850),
.Y(n_4849)
);

NAND2xp5_ASAP7_75t_L g4850 ( 
.A(n_4274),
.B(n_4276),
.Y(n_4850)
);

NAND2xp5_ASAP7_75t_L g4851 ( 
.A(n_4274),
.B(n_4276),
.Y(n_4851)
);

BUFx3_ASAP7_75t_L g4852 ( 
.A(n_4361),
.Y(n_4852)
);

AOI22xp5_ASAP7_75t_L g4853 ( 
.A1(n_4062),
.A2(n_4080),
.B1(n_4106),
.B2(n_4088),
.Y(n_4853)
);

BUFx6f_ASAP7_75t_L g4854 ( 
.A(n_4361),
.Y(n_4854)
);

NOR2xp33_ASAP7_75t_L g4855 ( 
.A(n_4012),
.B(n_4291),
.Y(n_4855)
);

BUFx8_ASAP7_75t_L g4856 ( 
.A(n_3461),
.Y(n_4856)
);

NOR2x1_ASAP7_75t_L g4857 ( 
.A(n_3365),
.B(n_3201),
.Y(n_4857)
);

AND2x4_ASAP7_75t_L g4858 ( 
.A(n_3850),
.B(n_3912),
.Y(n_4858)
);

OAI21xp5_ASAP7_75t_L g4859 ( 
.A1(n_3200),
.A2(n_3349),
.B(n_4270),
.Y(n_4859)
);

BUFx8_ASAP7_75t_SL g4860 ( 
.A(n_3337),
.Y(n_4860)
);

NAND2xp5_ASAP7_75t_L g4861 ( 
.A(n_4279),
.B(n_4283),
.Y(n_4861)
);

NOR2xp33_ASAP7_75t_L g4862 ( 
.A(n_4314),
.B(n_4432),
.Y(n_4862)
);

BUFx4f_ASAP7_75t_L g4863 ( 
.A(n_3461),
.Y(n_4863)
);

CKINVDCx20_ASAP7_75t_R g4864 ( 
.A(n_3759),
.Y(n_4864)
);

INVx3_ASAP7_75t_L g4865 ( 
.A(n_3668),
.Y(n_4865)
);

AND2x2_ASAP7_75t_L g4866 ( 
.A(n_3979),
.B(n_3980),
.Y(n_4866)
);

NAND2xp5_ASAP7_75t_L g4867 ( 
.A(n_4279),
.B(n_4283),
.Y(n_4867)
);

OR2x6_ASAP7_75t_L g4868 ( 
.A(n_3867),
.B(n_3870),
.Y(n_4868)
);

BUFx8_ASAP7_75t_SL g4869 ( 
.A(n_3293),
.Y(n_4869)
);

NOR2xp33_ASAP7_75t_L g4870 ( 
.A(n_4314),
.B(n_4432),
.Y(n_4870)
);

NAND2xp5_ASAP7_75t_L g4871 ( 
.A(n_4284),
.B(n_4285),
.Y(n_4871)
);

NOR2xp33_ASAP7_75t_L g4872 ( 
.A(n_4514),
.B(n_4519),
.Y(n_4872)
);

BUFx6f_ASAP7_75t_L g4873 ( 
.A(n_4361),
.Y(n_4873)
);

INVx3_ASAP7_75t_L g4874 ( 
.A(n_3668),
.Y(n_4874)
);

AOI221xp5_ASAP7_75t_L g4875 ( 
.A1(n_3368),
.A2(n_3420),
.B1(n_4403),
.B2(n_3427),
.C(n_4514),
.Y(n_4875)
);

BUFx12f_ASAP7_75t_L g4876 ( 
.A(n_4370),
.Y(n_4876)
);

AND2x2_ASAP7_75t_L g4877 ( 
.A(n_3980),
.B(n_4014),
.Y(n_4877)
);

AOI22xp5_ASAP7_75t_L g4878 ( 
.A1(n_4141),
.A2(n_4145),
.B1(n_4156),
.B2(n_4146),
.Y(n_4878)
);

AOI22xp5_ASAP7_75t_L g4879 ( 
.A1(n_4174),
.A2(n_4185),
.B1(n_4263),
.B2(n_4184),
.Y(n_4879)
);

NAND2xp5_ASAP7_75t_L g4880 ( 
.A(n_4284),
.B(n_4285),
.Y(n_4880)
);

BUFx2_ASAP7_75t_L g4881 ( 
.A(n_4014),
.Y(n_4881)
);

INVx5_ASAP7_75t_L g4882 ( 
.A(n_3668),
.Y(n_4882)
);

NAND2xp5_ASAP7_75t_L g4883 ( 
.A(n_4346),
.B(n_4351),
.Y(n_4883)
);

CKINVDCx5p33_ASAP7_75t_R g4884 ( 
.A(n_3293),
.Y(n_4884)
);

CKINVDCx11_ASAP7_75t_R g4885 ( 
.A(n_3402),
.Y(n_4885)
);

AND2x4_ASAP7_75t_L g4886 ( 
.A(n_3912),
.B(n_3951),
.Y(n_4886)
);

BUFx2_ASAP7_75t_L g4887 ( 
.A(n_4031),
.Y(n_4887)
);

OR2x2_ASAP7_75t_SL g4888 ( 
.A(n_4346),
.B(n_4351),
.Y(n_4888)
);

BUFx6f_ASAP7_75t_L g4889 ( 
.A(n_3231),
.Y(n_4889)
);

BUFx8_ASAP7_75t_L g4890 ( 
.A(n_3461),
.Y(n_4890)
);

AOI22xp33_ASAP7_75t_L g4891 ( 
.A1(n_4519),
.A2(n_3468),
.B1(n_4172),
.B2(n_4143),
.Y(n_4891)
);

NAND2xp5_ASAP7_75t_L g4892 ( 
.A(n_4352),
.B(n_4365),
.Y(n_4892)
);

INVxp67_ASAP7_75t_L g4893 ( 
.A(n_4142),
.Y(n_4893)
);

INVx2_ASAP7_75t_SL g4894 ( 
.A(n_3429),
.Y(n_4894)
);

AND2x4_ASAP7_75t_L g4895 ( 
.A(n_3912),
.B(n_3951),
.Y(n_4895)
);

INVx2_ASAP7_75t_L g4896 ( 
.A(n_3234),
.Y(n_4896)
);

AND2x4_ASAP7_75t_L g4897 ( 
.A(n_3912),
.B(n_3951),
.Y(n_4897)
);

NAND2xp5_ASAP7_75t_L g4898 ( 
.A(n_4352),
.B(n_4365),
.Y(n_4898)
);

NOR2xp33_ASAP7_75t_L g4899 ( 
.A(n_3393),
.B(n_3474),
.Y(n_4899)
);

AND2x2_ASAP7_75t_L g4900 ( 
.A(n_4031),
.B(n_4044),
.Y(n_4900)
);

A2O1A1Ixp33_ASAP7_75t_L g4901 ( 
.A1(n_4277),
.A2(n_4442),
.B(n_4536),
.C(n_4313),
.Y(n_4901)
);

AND2x4_ASAP7_75t_L g4902 ( 
.A(n_3951),
.B(n_4026),
.Y(n_4902)
);

INVx1_ASAP7_75t_L g4903 ( 
.A(n_3161),
.Y(n_4903)
);

BUFx2_ASAP7_75t_L g4904 ( 
.A(n_4044),
.Y(n_4904)
);

NAND2xp5_ASAP7_75t_L g4905 ( 
.A(n_4368),
.B(n_4371),
.Y(n_4905)
);

BUFx2_ASAP7_75t_L g4906 ( 
.A(n_4056),
.Y(n_4906)
);

OR2x2_ASAP7_75t_L g4907 ( 
.A(n_4056),
.B(n_4075),
.Y(n_4907)
);

NAND2xp5_ASAP7_75t_L g4908 ( 
.A(n_4368),
.B(n_4371),
.Y(n_4908)
);

INVx1_ASAP7_75t_L g4909 ( 
.A(n_3161),
.Y(n_4909)
);

AND3x1_ASAP7_75t_L g4910 ( 
.A(n_3347),
.B(n_3790),
.C(n_3435),
.Y(n_4910)
);

INVx1_ASAP7_75t_L g4911 ( 
.A(n_3168),
.Y(n_4911)
);

NAND2xp5_ASAP7_75t_L g4912 ( 
.A(n_4375),
.B(n_4380),
.Y(n_4912)
);

INVx1_ASAP7_75t_L g4913 ( 
.A(n_3168),
.Y(n_4913)
);

INVx2_ASAP7_75t_L g4914 ( 
.A(n_3234),
.Y(n_4914)
);

CKINVDCx5p33_ASAP7_75t_R g4915 ( 
.A(n_3923),
.Y(n_4915)
);

BUFx3_ASAP7_75t_L g4916 ( 
.A(n_3208),
.Y(n_4916)
);

HB1xp67_ASAP7_75t_L g4917 ( 
.A(n_3947),
.Y(n_4917)
);

INVx1_ASAP7_75t_L g4918 ( 
.A(n_3804),
.Y(n_4918)
);

NAND2xp5_ASAP7_75t_L g4919 ( 
.A(n_4375),
.B(n_4380),
.Y(n_4919)
);

BUFx3_ASAP7_75t_L g4920 ( 
.A(n_3208),
.Y(n_4920)
);

BUFx2_ASAP7_75t_L g4921 ( 
.A(n_4075),
.Y(n_4921)
);

OR2x2_ASAP7_75t_L g4922 ( 
.A(n_4079),
.B(n_4082),
.Y(n_4922)
);

INVx1_ASAP7_75t_L g4923 ( 
.A(n_3804),
.Y(n_4923)
);

CKINVDCx5p33_ASAP7_75t_R g4924 ( 
.A(n_3923),
.Y(n_4924)
);

NAND2xp5_ASAP7_75t_SL g4925 ( 
.A(n_3479),
.B(n_3808),
.Y(n_4925)
);

INVxp67_ASAP7_75t_L g4926 ( 
.A(n_4152),
.Y(n_4926)
);

NAND2xp5_ASAP7_75t_L g4927 ( 
.A(n_4395),
.B(n_4396),
.Y(n_4927)
);

AOI22xp33_ASAP7_75t_L g4928 ( 
.A1(n_3468),
.A2(n_4297),
.B1(n_4382),
.B2(n_3427),
.Y(n_4928)
);

NAND2xp5_ASAP7_75t_L g4929 ( 
.A(n_4395),
.B(n_4396),
.Y(n_4929)
);

BUFx3_ASAP7_75t_L g4930 ( 
.A(n_3208),
.Y(n_4930)
);

NOR2xp33_ASAP7_75t_R g4931 ( 
.A(n_3782),
.B(n_4370),
.Y(n_4931)
);

NAND2xp5_ASAP7_75t_L g4932 ( 
.A(n_4399),
.B(n_4401),
.Y(n_4932)
);

BUFx4f_ASAP7_75t_L g4933 ( 
.A(n_3481),
.Y(n_4933)
);

INVx1_ASAP7_75t_L g4934 ( 
.A(n_3827),
.Y(n_4934)
);

BUFx6f_ASAP7_75t_L g4935 ( 
.A(n_3231),
.Y(n_4935)
);

BUFx2_ASAP7_75t_L g4936 ( 
.A(n_4079),
.Y(n_4936)
);

NAND2xp5_ASAP7_75t_L g4937 ( 
.A(n_4399),
.B(n_4401),
.Y(n_4937)
);

AND2x4_ASAP7_75t_L g4938 ( 
.A(n_4026),
.B(n_4110),
.Y(n_4938)
);

NAND2xp5_ASAP7_75t_SL g4939 ( 
.A(n_3479),
.B(n_3808),
.Y(n_4939)
);

INVx2_ASAP7_75t_L g4940 ( 
.A(n_3234),
.Y(n_4940)
);

NOR2xp33_ASAP7_75t_L g4941 ( 
.A(n_3286),
.B(n_3222),
.Y(n_4941)
);

INVx2_ASAP7_75t_L g4942 ( 
.A(n_3236),
.Y(n_4942)
);

INVx1_ASAP7_75t_L g4943 ( 
.A(n_3827),
.Y(n_4943)
);

AOI22xp33_ASAP7_75t_L g4944 ( 
.A1(n_4403),
.A2(n_3425),
.B1(n_3405),
.B2(n_3475),
.Y(n_4944)
);

INVx1_ASAP7_75t_SL g4945 ( 
.A(n_3447),
.Y(n_4945)
);

BUFx6f_ASAP7_75t_L g4946 ( 
.A(n_3947),
.Y(n_4946)
);

NAND2xp5_ASAP7_75t_SL g4947 ( 
.A(n_3813),
.B(n_3925),
.Y(n_4947)
);

NAND2xp5_ASAP7_75t_L g4948 ( 
.A(n_4408),
.B(n_4411),
.Y(n_4948)
);

INVx4_ASAP7_75t_L g4949 ( 
.A(n_4026),
.Y(n_4949)
);

HB1xp67_ASAP7_75t_L g4950 ( 
.A(n_4019),
.Y(n_4950)
);

NOR2xp33_ASAP7_75t_L g4951 ( 
.A(n_3492),
.B(n_3435),
.Y(n_4951)
);

INVx2_ASAP7_75t_SL g4952 ( 
.A(n_3477),
.Y(n_4952)
);

AND2x2_ASAP7_75t_L g4953 ( 
.A(n_4082),
.B(n_4086),
.Y(n_4953)
);

AND2x2_ASAP7_75t_L g4954 ( 
.A(n_4086),
.B(n_4100),
.Y(n_4954)
);

BUFx2_ASAP7_75t_L g4955 ( 
.A(n_4100),
.Y(n_4955)
);

INVxp67_ASAP7_75t_SL g4956 ( 
.A(n_3871),
.Y(n_4956)
);

CKINVDCx5p33_ASAP7_75t_R g4957 ( 
.A(n_3923),
.Y(n_4957)
);

NAND2xp5_ASAP7_75t_L g4958 ( 
.A(n_4408),
.B(n_4411),
.Y(n_4958)
);

INVx1_ASAP7_75t_L g4959 ( 
.A(n_3835),
.Y(n_4959)
);

INVxp67_ASAP7_75t_SL g4960 ( 
.A(n_3898),
.Y(n_4960)
);

NAND2xp5_ASAP7_75t_L g4961 ( 
.A(n_4422),
.B(n_4423),
.Y(n_4961)
);

BUFx2_ASAP7_75t_L g4962 ( 
.A(n_4102),
.Y(n_4962)
);

CKINVDCx20_ASAP7_75t_R g4963 ( 
.A(n_4370),
.Y(n_4963)
);

AND2x2_ASAP7_75t_L g4964 ( 
.A(n_4102),
.B(n_4117),
.Y(n_4964)
);

NOR2xp33_ASAP7_75t_L g4965 ( 
.A(n_3840),
.B(n_3841),
.Y(n_4965)
);

AND2x2_ASAP7_75t_L g4966 ( 
.A(n_4117),
.B(n_4131),
.Y(n_4966)
);

INVx2_ASAP7_75t_SL g4967 ( 
.A(n_3477),
.Y(n_4967)
);

AND2x4_ASAP7_75t_L g4968 ( 
.A(n_4026),
.B(n_4110),
.Y(n_4968)
);

OR2x6_ASAP7_75t_L g4969 ( 
.A(n_3873),
.B(n_3881),
.Y(n_4969)
);

AND2x2_ASAP7_75t_L g4970 ( 
.A(n_4131),
.B(n_4157),
.Y(n_4970)
);

NOR2xp33_ASAP7_75t_R g4971 ( 
.A(n_3675),
.B(n_3570),
.Y(n_4971)
);

INVx1_ASAP7_75t_L g4972 ( 
.A(n_3835),
.Y(n_4972)
);

INVx1_ASAP7_75t_L g4973 ( 
.A(n_3848),
.Y(n_4973)
);

AND2x2_ASAP7_75t_L g4974 ( 
.A(n_4157),
.B(n_4164),
.Y(n_4974)
);

INVx1_ASAP7_75t_L g4975 ( 
.A(n_3848),
.Y(n_4975)
);

INVx1_ASAP7_75t_L g4976 ( 
.A(n_3854),
.Y(n_4976)
);

INVxp67_ASAP7_75t_L g4977 ( 
.A(n_4152),
.Y(n_4977)
);

NOR2xp67_ASAP7_75t_L g4978 ( 
.A(n_3352),
.B(n_3357),
.Y(n_4978)
);

INVx3_ASAP7_75t_L g4979 ( 
.A(n_4110),
.Y(n_4979)
);

INVx1_ASAP7_75t_L g4980 ( 
.A(n_3854),
.Y(n_4980)
);

INVx4_ASAP7_75t_L g4981 ( 
.A(n_4110),
.Y(n_4981)
);

NAND2xp5_ASAP7_75t_L g4982 ( 
.A(n_4422),
.B(n_4423),
.Y(n_4982)
);

NAND2xp5_ASAP7_75t_L g4983 ( 
.A(n_4424),
.B(n_4436),
.Y(n_4983)
);

NAND2xp5_ASAP7_75t_L g4984 ( 
.A(n_4424),
.B(n_4436),
.Y(n_4984)
);

AND2x2_ASAP7_75t_L g4985 ( 
.A(n_4164),
.B(n_4203),
.Y(n_4985)
);

OAI22xp5_ASAP7_75t_L g4986 ( 
.A1(n_4266),
.A2(n_4286),
.B1(n_4302),
.B2(n_4275),
.Y(n_4986)
);

INVx1_ASAP7_75t_L g4987 ( 
.A(n_3860),
.Y(n_4987)
);

NAND2xp5_ASAP7_75t_L g4988 ( 
.A(n_4437),
.B(n_4439),
.Y(n_4988)
);

INVx1_ASAP7_75t_SL g4989 ( 
.A(n_4153),
.Y(n_4989)
);

BUFx3_ASAP7_75t_L g4990 ( 
.A(n_3208),
.Y(n_4990)
);

INVx1_ASAP7_75t_L g4991 ( 
.A(n_3860),
.Y(n_4991)
);

A2O1A1Ixp33_ASAP7_75t_L g4992 ( 
.A1(n_4252),
.A2(n_4430),
.B(n_3306),
.C(n_3264),
.Y(n_4992)
);

INVx1_ASAP7_75t_L g4993 ( 
.A(n_3866),
.Y(n_4993)
);

AND2x4_ASAP7_75t_L g4994 ( 
.A(n_4147),
.B(n_4388),
.Y(n_4994)
);

NAND2x1p5_ASAP7_75t_L g4995 ( 
.A(n_4027),
.B(n_4151),
.Y(n_4995)
);

INVx3_ASAP7_75t_L g4996 ( 
.A(n_4147),
.Y(n_4996)
);

NAND2xp5_ASAP7_75t_L g4997 ( 
.A(n_4437),
.B(n_4439),
.Y(n_4997)
);

NOR2xp33_ASAP7_75t_L g4998 ( 
.A(n_3852),
.B(n_3857),
.Y(n_4998)
);

BUFx2_ASAP7_75t_L g4999 ( 
.A(n_4203),
.Y(n_4999)
);

OR2x6_ASAP7_75t_L g5000 ( 
.A(n_3900),
.B(n_3903),
.Y(n_5000)
);

NAND2xp5_ASAP7_75t_L g5001 ( 
.A(n_4443),
.B(n_4520),
.Y(n_5001)
);

NOR2xp67_ASAP7_75t_L g5002 ( 
.A(n_3381),
.B(n_3382),
.Y(n_5002)
);

INVx3_ASAP7_75t_SL g5003 ( 
.A(n_3606),
.Y(n_5003)
);

INVx1_ASAP7_75t_L g5004 ( 
.A(n_3866),
.Y(n_5004)
);

NOR2xp33_ASAP7_75t_L g5005 ( 
.A(n_3858),
.B(n_3863),
.Y(n_5005)
);

INVx1_ASAP7_75t_L g5006 ( 
.A(n_3869),
.Y(n_5006)
);

BUFx2_ASAP7_75t_L g5007 ( 
.A(n_4204),
.Y(n_5007)
);

INVx4_ASAP7_75t_L g5008 ( 
.A(n_4147),
.Y(n_5008)
);

CKINVDCx14_ASAP7_75t_R g5009 ( 
.A(n_3159),
.Y(n_5009)
);

AOI221x1_ASAP7_75t_L g5010 ( 
.A1(n_4208),
.A2(n_4416),
.B1(n_4478),
.B2(n_4309),
.C(n_4250),
.Y(n_5010)
);

INVx1_ASAP7_75t_L g5011 ( 
.A(n_3869),
.Y(n_5011)
);

CKINVDCx20_ASAP7_75t_R g5012 ( 
.A(n_3213),
.Y(n_5012)
);

CKINVDCx5p33_ASAP7_75t_R g5013 ( 
.A(n_4236),
.Y(n_5013)
);

AND2x2_ASAP7_75t_SL g5014 ( 
.A(n_3813),
.B(n_3925),
.Y(n_5014)
);

NAND2xp5_ASAP7_75t_L g5015 ( 
.A(n_4443),
.B(n_4520),
.Y(n_5015)
);

BUFx2_ASAP7_75t_L g5016 ( 
.A(n_4204),
.Y(n_5016)
);

NAND2xp5_ASAP7_75t_L g5017 ( 
.A(n_4522),
.B(n_4525),
.Y(n_5017)
);

AOI22xp33_ASAP7_75t_L g5018 ( 
.A1(n_3405),
.A2(n_3425),
.B1(n_3360),
.B2(n_3369),
.Y(n_5018)
);

INVx4_ASAP7_75t_L g5019 ( 
.A(n_4147),
.Y(n_5019)
);

BUFx6f_ASAP7_75t_L g5020 ( 
.A(n_4019),
.Y(n_5020)
);

NAND2xp5_ASAP7_75t_L g5021 ( 
.A(n_4522),
.B(n_4525),
.Y(n_5021)
);

CKINVDCx5p33_ASAP7_75t_R g5022 ( 
.A(n_4236),
.Y(n_5022)
);

NAND2xp5_ASAP7_75t_L g5023 ( 
.A(n_4529),
.B(n_4530),
.Y(n_5023)
);

AND2x4_ASAP7_75t_L g5024 ( 
.A(n_4388),
.B(n_3583),
.Y(n_5024)
);

CKINVDCx20_ASAP7_75t_R g5025 ( 
.A(n_3213),
.Y(n_5025)
);

INVx3_ASAP7_75t_L g5026 ( 
.A(n_4388),
.Y(n_5026)
);

NOR2xp33_ASAP7_75t_L g5027 ( 
.A(n_3872),
.B(n_3874),
.Y(n_5027)
);

NAND2xp5_ASAP7_75t_L g5028 ( 
.A(n_4529),
.B(n_4530),
.Y(n_5028)
);

HB1xp67_ASAP7_75t_L g5029 ( 
.A(n_4027),
.Y(n_5029)
);

BUFx6f_ASAP7_75t_L g5030 ( 
.A(n_4053),
.Y(n_5030)
);

INVxp67_ASAP7_75t_L g5031 ( 
.A(n_4153),
.Y(n_5031)
);

BUFx6f_ASAP7_75t_L g5032 ( 
.A(n_4053),
.Y(n_5032)
);

NAND2xp5_ASAP7_75t_L g5033 ( 
.A(n_4532),
.B(n_3173),
.Y(n_5033)
);

AND2x6_ASAP7_75t_L g5034 ( 
.A(n_4388),
.B(n_3481),
.Y(n_5034)
);

AND2x6_ASAP7_75t_L g5035 ( 
.A(n_3481),
.B(n_3242),
.Y(n_5035)
);

AND2x2_ASAP7_75t_L g5036 ( 
.A(n_4231),
.B(n_4295),
.Y(n_5036)
);

INVx1_ASAP7_75t_L g5037 ( 
.A(n_3879),
.Y(n_5037)
);

NOR2xp33_ASAP7_75t_L g5038 ( 
.A(n_3877),
.B(n_3878),
.Y(n_5038)
);

NAND2xp5_ASAP7_75t_SL g5039 ( 
.A(n_3898),
.B(n_3910),
.Y(n_5039)
);

A2O1A1Ixp33_ASAP7_75t_L g5040 ( 
.A1(n_3233),
.A2(n_3432),
.B(n_3198),
.C(n_3439),
.Y(n_5040)
);

NOR2xp33_ASAP7_75t_L g5041 ( 
.A(n_3880),
.B(n_3883),
.Y(n_5041)
);

NAND2xp5_ASAP7_75t_L g5042 ( 
.A(n_4532),
.B(n_3166),
.Y(n_5042)
);

NAND2xp5_ASAP7_75t_L g5043 ( 
.A(n_3169),
.B(n_3375),
.Y(n_5043)
);

AND3x1_ASAP7_75t_L g5044 ( 
.A(n_3347),
.B(n_3232),
.C(n_3570),
.Y(n_5044)
);

AND2x2_ASAP7_75t_L g5045 ( 
.A(n_4231),
.B(n_4295),
.Y(n_5045)
);

BUFx6f_ASAP7_75t_L g5046 ( 
.A(n_4070),
.Y(n_5046)
);

INVx1_ASAP7_75t_L g5047 ( 
.A(n_3879),
.Y(n_5047)
);

HB1xp67_ASAP7_75t_L g5048 ( 
.A(n_4070),
.Y(n_5048)
);

NOR2xp33_ASAP7_75t_L g5049 ( 
.A(n_3886),
.B(n_3888),
.Y(n_5049)
);

AND2x2_ASAP7_75t_L g5050 ( 
.A(n_4323),
.B(n_4364),
.Y(n_5050)
);

O2A1O1Ixp33_ASAP7_75t_L g5051 ( 
.A1(n_3849),
.A2(n_4271),
.B(n_4534),
.C(n_4089),
.Y(n_5051)
);

BUFx6f_ASAP7_75t_L g5052 ( 
.A(n_4151),
.Y(n_5052)
);

INVx1_ASAP7_75t_L g5053 ( 
.A(n_3915),
.Y(n_5053)
);

INVx1_ASAP7_75t_L g5054 ( 
.A(n_3915),
.Y(n_5054)
);

BUFx2_ASAP7_75t_L g5055 ( 
.A(n_4323),
.Y(n_5055)
);

HB1xp67_ASAP7_75t_L g5056 ( 
.A(n_4202),
.Y(n_5056)
);

CKINVDCx20_ASAP7_75t_R g5057 ( 
.A(n_3213),
.Y(n_5057)
);

INVx1_ASAP7_75t_L g5058 ( 
.A(n_3937),
.Y(n_5058)
);

INVx1_ASAP7_75t_L g5059 ( 
.A(n_3937),
.Y(n_5059)
);

INVx1_ASAP7_75t_L g5060 ( 
.A(n_3965),
.Y(n_5060)
);

INVx2_ASAP7_75t_SL g5061 ( 
.A(n_3493),
.Y(n_5061)
);

AOI221xp5_ASAP7_75t_L g5062 ( 
.A1(n_3432),
.A2(n_4345),
.B1(n_4381),
.B2(n_4320),
.C(n_4307),
.Y(n_5062)
);

INVx1_ASAP7_75t_L g5063 ( 
.A(n_3965),
.Y(n_5063)
);

INVx1_ASAP7_75t_L g5064 ( 
.A(n_3968),
.Y(n_5064)
);

BUFx3_ASAP7_75t_L g5065 ( 
.A(n_3968),
.Y(n_5065)
);

INVx4_ASAP7_75t_L g5066 ( 
.A(n_3481),
.Y(n_5066)
);

AND2x2_ASAP7_75t_L g5067 ( 
.A(n_4364),
.B(n_4433),
.Y(n_5067)
);

INVx1_ASAP7_75t_L g5068 ( 
.A(n_3973),
.Y(n_5068)
);

NAND2xp5_ASAP7_75t_L g5069 ( 
.A(n_3375),
.B(n_3277),
.Y(n_5069)
);

NAND2xp5_ASAP7_75t_L g5070 ( 
.A(n_3277),
.B(n_3355),
.Y(n_5070)
);

AOI22xp5_ASAP7_75t_L g5071 ( 
.A1(n_4407),
.A2(n_4413),
.B1(n_4460),
.B2(n_4441),
.Y(n_5071)
);

NAND2xp5_ASAP7_75t_L g5072 ( 
.A(n_3355),
.B(n_3497),
.Y(n_5072)
);

NAND2xp5_ASAP7_75t_L g5073 ( 
.A(n_3497),
.B(n_3530),
.Y(n_5073)
);

NAND2xp5_ASAP7_75t_SL g5074 ( 
.A(n_3910),
.B(n_4009),
.Y(n_5074)
);

BUFx6f_ASAP7_75t_L g5075 ( 
.A(n_4202),
.Y(n_5075)
);

NOR2xp33_ASAP7_75t_R g5076 ( 
.A(n_3654),
.B(n_3159),
.Y(n_5076)
);

NAND2xp5_ASAP7_75t_L g5077 ( 
.A(n_3530),
.B(n_3417),
.Y(n_5077)
);

OR2x6_ASAP7_75t_L g5078 ( 
.A(n_3907),
.B(n_3908),
.Y(n_5078)
);

AND2x2_ASAP7_75t_L g5079 ( 
.A(n_4433),
.B(n_4450),
.Y(n_5079)
);

NAND2xp5_ASAP7_75t_SL g5080 ( 
.A(n_4009),
.B(n_4032),
.Y(n_5080)
);

AND2x2_ASAP7_75t_SL g5081 ( 
.A(n_3180),
.B(n_3184),
.Y(n_5081)
);

INVx5_ASAP7_75t_L g5082 ( 
.A(n_4222),
.Y(n_5082)
);

INVx1_ASAP7_75t_L g5083 ( 
.A(n_3973),
.Y(n_5083)
);

NOR2xp33_ASAP7_75t_L g5084 ( 
.A(n_3892),
.B(n_3895),
.Y(n_5084)
);

BUFx2_ASAP7_75t_L g5085 ( 
.A(n_4450),
.Y(n_5085)
);

INVx1_ASAP7_75t_L g5086 ( 
.A(n_4000),
.Y(n_5086)
);

INVx1_ASAP7_75t_L g5087 ( 
.A(n_4000),
.Y(n_5087)
);

OAI21xp5_ASAP7_75t_L g5088 ( 
.A1(n_4189),
.A2(n_3215),
.B(n_3185),
.Y(n_5088)
);

NOR2xp33_ASAP7_75t_L g5089 ( 
.A(n_3897),
.B(n_3911),
.Y(n_5089)
);

CKINVDCx5p33_ASAP7_75t_R g5090 ( 
.A(n_4236),
.Y(n_5090)
);

INVx1_ASAP7_75t_L g5091 ( 
.A(n_4003),
.Y(n_5091)
);

NAND2xp5_ASAP7_75t_L g5092 ( 
.A(n_3440),
.B(n_3442),
.Y(n_5092)
);

NAND2xp5_ASAP7_75t_L g5093 ( 
.A(n_3448),
.B(n_3451),
.Y(n_5093)
);

NAND2xp5_ASAP7_75t_L g5094 ( 
.A(n_3452),
.B(n_3453),
.Y(n_5094)
);

AND2x2_ASAP7_75t_L g5095 ( 
.A(n_4459),
.B(n_4461),
.Y(n_5095)
);

BUFx2_ASAP7_75t_L g5096 ( 
.A(n_4459),
.Y(n_5096)
);

BUFx6f_ASAP7_75t_L g5097 ( 
.A(n_4206),
.Y(n_5097)
);

BUFx3_ASAP7_75t_L g5098 ( 
.A(n_4003),
.Y(n_5098)
);

BUFx12f_ASAP7_75t_L g5099 ( 
.A(n_3213),
.Y(n_5099)
);

NAND2xp5_ASAP7_75t_L g5100 ( 
.A(n_3462),
.B(n_3465),
.Y(n_5100)
);

NAND2xp5_ASAP7_75t_L g5101 ( 
.A(n_3470),
.B(n_3472),
.Y(n_5101)
);

INVx1_ASAP7_75t_L g5102 ( 
.A(n_4006),
.Y(n_5102)
);

BUFx4f_ASAP7_75t_L g5103 ( 
.A(n_3481),
.Y(n_5103)
);

INVx2_ASAP7_75t_SL g5104 ( 
.A(n_3493),
.Y(n_5104)
);

HB1xp67_ASAP7_75t_L g5105 ( 
.A(n_4206),
.Y(n_5105)
);

INVx2_ASAP7_75t_SL g5106 ( 
.A(n_3242),
.Y(n_5106)
);

BUFx3_ASAP7_75t_L g5107 ( 
.A(n_4006),
.Y(n_5107)
);

NAND2xp5_ASAP7_75t_L g5108 ( 
.A(n_3160),
.B(n_3509),
.Y(n_5108)
);

HB1xp67_ASAP7_75t_L g5109 ( 
.A(n_4235),
.Y(n_5109)
);

AND2x4_ASAP7_75t_L g5110 ( 
.A(n_4077),
.B(n_4461),
.Y(n_5110)
);

BUFx2_ASAP7_75t_R g5111 ( 
.A(n_3788),
.Y(n_5111)
);

OR2x6_ASAP7_75t_L g5112 ( 
.A(n_3909),
.B(n_3917),
.Y(n_5112)
);

NAND2xp5_ASAP7_75t_L g5113 ( 
.A(n_3509),
.B(n_3538),
.Y(n_5113)
);

NAND2xp5_ASAP7_75t_L g5114 ( 
.A(n_3538),
.B(n_3334),
.Y(n_5114)
);

HB1xp67_ASAP7_75t_L g5115 ( 
.A(n_4235),
.Y(n_5115)
);

INVx2_ASAP7_75t_L g5116 ( 
.A(n_3319),
.Y(n_5116)
);

NAND2xp5_ASAP7_75t_L g5117 ( 
.A(n_3372),
.B(n_3565),
.Y(n_5117)
);

INVx2_ASAP7_75t_L g5118 ( 
.A(n_3319),
.Y(n_5118)
);

NAND2xp5_ASAP7_75t_SL g5119 ( 
.A(n_4032),
.B(n_4038),
.Y(n_5119)
);

INVx4_ASAP7_75t_L g5120 ( 
.A(n_3481),
.Y(n_5120)
);

INVx3_ASAP7_75t_L g5121 ( 
.A(n_3353),
.Y(n_5121)
);

INVx2_ASAP7_75t_SL g5122 ( 
.A(n_3242),
.Y(n_5122)
);

AND3x1_ASAP7_75t_SL g5123 ( 
.A(n_3582),
.B(n_3415),
.C(n_4189),
.Y(n_5123)
);

INVx1_ASAP7_75t_L g5124 ( 
.A(n_4022),
.Y(n_5124)
);

INVx3_ASAP7_75t_L g5125 ( 
.A(n_3353),
.Y(n_5125)
);

INVx1_ASAP7_75t_L g5126 ( 
.A(n_4022),
.Y(n_5126)
);

AOI21xp5_ASAP7_75t_L g5127 ( 
.A1(n_3922),
.A2(n_3933),
.B(n_3930),
.Y(n_5127)
);

NAND2xp5_ASAP7_75t_SL g5128 ( 
.A(n_4038),
.B(n_4085),
.Y(n_5128)
);

A2O1A1Ixp33_ASAP7_75t_L g5129 ( 
.A1(n_3198),
.A2(n_3445),
.B(n_3459),
.C(n_3436),
.Y(n_5129)
);

BUFx6f_ASAP7_75t_L g5130 ( 
.A(n_4245),
.Y(n_5130)
);

INVxp67_ASAP7_75t_SL g5131 ( 
.A(n_4085),
.Y(n_5131)
);

NAND2xp5_ASAP7_75t_SL g5132 ( 
.A(n_4095),
.B(n_4196),
.Y(n_5132)
);

BUFx6f_ASAP7_75t_L g5133 ( 
.A(n_4245),
.Y(n_5133)
);

OR2x2_ASAP7_75t_L g5134 ( 
.A(n_4474),
.B(n_4481),
.Y(n_5134)
);

AND2x4_ASAP7_75t_L g5135 ( 
.A(n_4077),
.B(n_4474),
.Y(n_5135)
);

NAND2xp5_ASAP7_75t_L g5136 ( 
.A(n_3508),
.B(n_3519),
.Y(n_5136)
);

OAI21x1_ASAP7_75t_L g5137 ( 
.A1(n_3938),
.A2(n_4544),
.B(n_3944),
.Y(n_5137)
);

OAI221xp5_ASAP7_75t_L g5138 ( 
.A1(n_3811),
.A2(n_3851),
.B1(n_3868),
.B2(n_3837),
.C(n_3829),
.Y(n_5138)
);

NOR2x1_ASAP7_75t_L g5139 ( 
.A(n_3336),
.B(n_3338),
.Y(n_5139)
);

AND2x6_ASAP7_75t_L g5140 ( 
.A(n_3242),
.B(n_3823),
.Y(n_5140)
);

AOI22xp5_ASAP7_75t_L g5141 ( 
.A1(n_4463),
.A2(n_4487),
.B1(n_4488),
.B2(n_4482),
.Y(n_5141)
);

INVx2_ASAP7_75t_L g5142 ( 
.A(n_3351),
.Y(n_5142)
);

NAND2xp5_ASAP7_75t_SL g5143 ( 
.A(n_4095),
.B(n_4196),
.Y(n_5143)
);

INVx2_ASAP7_75t_L g5144 ( 
.A(n_3351),
.Y(n_5144)
);

INVxp67_ASAP7_75t_L g5145 ( 
.A(n_4305),
.Y(n_5145)
);

INVx1_ASAP7_75t_L g5146 ( 
.A(n_4063),
.Y(n_5146)
);

INVx2_ASAP7_75t_L g5147 ( 
.A(n_3351),
.Y(n_5147)
);

INVx1_ASAP7_75t_SL g5148 ( 
.A(n_4305),
.Y(n_5148)
);

NAND2xp5_ASAP7_75t_L g5149 ( 
.A(n_3550),
.B(n_3177),
.Y(n_5149)
);

CKINVDCx5p33_ASAP7_75t_R g5150 ( 
.A(n_4468),
.Y(n_5150)
);

AOI22xp33_ASAP7_75t_L g5151 ( 
.A1(n_3325),
.A2(n_3369),
.B1(n_3383),
.B2(n_3360),
.Y(n_5151)
);

INVx1_ASAP7_75t_L g5152 ( 
.A(n_4063),
.Y(n_5152)
);

INVx1_ASAP7_75t_L g5153 ( 
.A(n_4101),
.Y(n_5153)
);

BUFx12f_ASAP7_75t_L g5154 ( 
.A(n_3386),
.Y(n_5154)
);

INVx1_ASAP7_75t_L g5155 ( 
.A(n_4101),
.Y(n_5155)
);

INVx1_ASAP7_75t_L g5156 ( 
.A(n_4133),
.Y(n_5156)
);

NAND2xp5_ASAP7_75t_SL g5157 ( 
.A(n_4253),
.B(n_4369),
.Y(n_5157)
);

NAND2xp5_ASAP7_75t_L g5158 ( 
.A(n_3183),
.B(n_3188),
.Y(n_5158)
);

OR2x6_ASAP7_75t_L g5159 ( 
.A(n_3942),
.B(n_3948),
.Y(n_5159)
);

BUFx6f_ASAP7_75t_L g5160 ( 
.A(n_4342),
.Y(n_5160)
);

INVx4_ASAP7_75t_L g5161 ( 
.A(n_3935),
.Y(n_5161)
);

INVx2_ASAP7_75t_L g5162 ( 
.A(n_3387),
.Y(n_5162)
);

INVxp67_ASAP7_75t_L g5163 ( 
.A(n_4417),
.Y(n_5163)
);

AOI21xp5_ASAP7_75t_L g5164 ( 
.A1(n_3961),
.A2(n_3971),
.B(n_3964),
.Y(n_5164)
);

BUFx2_ASAP7_75t_L g5165 ( 
.A(n_4481),
.Y(n_5165)
);

INVx2_ASAP7_75t_SL g5166 ( 
.A(n_4533),
.Y(n_5166)
);

BUFx12f_ASAP7_75t_L g5167 ( 
.A(n_3386),
.Y(n_5167)
);

INVx2_ASAP7_75t_L g5168 ( 
.A(n_3387),
.Y(n_5168)
);

BUFx3_ASAP7_75t_L g5169 ( 
.A(n_4133),
.Y(n_5169)
);

NOR2xp33_ASAP7_75t_SL g5170 ( 
.A(n_3178),
.B(n_3245),
.Y(n_5170)
);

NAND2xp5_ASAP7_75t_L g5171 ( 
.A(n_3189),
.B(n_3207),
.Y(n_5171)
);

NAND2xp5_ASAP7_75t_L g5172 ( 
.A(n_3211),
.B(n_3216),
.Y(n_5172)
);

AND2x2_ASAP7_75t_L g5173 ( 
.A(n_4511),
.B(n_4512),
.Y(n_5173)
);

CKINVDCx5p33_ASAP7_75t_R g5174 ( 
.A(n_4468),
.Y(n_5174)
);

INVx1_ASAP7_75t_L g5175 ( 
.A(n_4137),
.Y(n_5175)
);

NAND2xp5_ASAP7_75t_L g5176 ( 
.A(n_3225),
.B(n_3229),
.Y(n_5176)
);

INVx1_ASAP7_75t_L g5177 ( 
.A(n_4137),
.Y(n_5177)
);

AND2x2_ASAP7_75t_L g5178 ( 
.A(n_4511),
.B(n_4512),
.Y(n_5178)
);

BUFx4f_ASAP7_75t_L g5179 ( 
.A(n_3242),
.Y(n_5179)
);

NAND2xp5_ASAP7_75t_SL g5180 ( 
.A(n_4253),
.B(n_4369),
.Y(n_5180)
);

INVx1_ASAP7_75t_L g5181 ( 
.A(n_4188),
.Y(n_5181)
);

NAND2xp5_ASAP7_75t_L g5182 ( 
.A(n_3241),
.B(n_3244),
.Y(n_5182)
);

NAND2xp5_ASAP7_75t_L g5183 ( 
.A(n_3247),
.B(n_3253),
.Y(n_5183)
);

AOI22xp5_ASAP7_75t_L g5184 ( 
.A1(n_4491),
.A2(n_4506),
.B1(n_4545),
.B2(n_4493),
.Y(n_5184)
);

NAND2xp5_ASAP7_75t_L g5185 ( 
.A(n_3260),
.B(n_3269),
.Y(n_5185)
);

NAND2xp5_ASAP7_75t_L g5186 ( 
.A(n_3272),
.B(n_3278),
.Y(n_5186)
);

NAND2xp5_ASAP7_75t_L g5187 ( 
.A(n_3280),
.B(n_3289),
.Y(n_5187)
);

BUFx3_ASAP7_75t_L g5188 ( 
.A(n_4188),
.Y(n_5188)
);

INVxp67_ASAP7_75t_SL g5189 ( 
.A(n_4376),
.Y(n_5189)
);

NAND2xp5_ASAP7_75t_L g5190 ( 
.A(n_3302),
.B(n_3528),
.Y(n_5190)
);

INVx1_ASAP7_75t_L g5191 ( 
.A(n_4194),
.Y(n_5191)
);

OAI21xp5_ASAP7_75t_L g5192 ( 
.A1(n_3175),
.A2(n_3928),
.B(n_3884),
.Y(n_5192)
);

BUFx6f_ASAP7_75t_SL g5193 ( 
.A(n_4542),
.Y(n_5193)
);

INVx1_ASAP7_75t_L g5194 ( 
.A(n_4194),
.Y(n_5194)
);

INVx4_ASAP7_75t_L g5195 ( 
.A(n_3242),
.Y(n_5195)
);

INVx1_ASAP7_75t_L g5196 ( 
.A(n_4209),
.Y(n_5196)
);

NAND2xp5_ASAP7_75t_L g5197 ( 
.A(n_3533),
.B(n_3545),
.Y(n_5197)
);

INVx3_ASAP7_75t_L g5198 ( 
.A(n_3206),
.Y(n_5198)
);

NAND2xp5_ASAP7_75t_SL g5199 ( 
.A(n_4376),
.B(n_4383),
.Y(n_5199)
);

NOR2xp33_ASAP7_75t_L g5200 ( 
.A(n_3913),
.B(n_3916),
.Y(n_5200)
);

CKINVDCx20_ASAP7_75t_R g5201 ( 
.A(n_3386),
.Y(n_5201)
);

AND2x4_ASAP7_75t_L g5202 ( 
.A(n_4521),
.B(n_4523),
.Y(n_5202)
);

AOI22xp33_ASAP7_75t_L g5203 ( 
.A1(n_3383),
.A2(n_3443),
.B1(n_3446),
.B2(n_3444),
.Y(n_5203)
);

OR2x2_ASAP7_75t_L g5204 ( 
.A(n_4521),
.B(n_4523),
.Y(n_5204)
);

BUFx6f_ASAP7_75t_L g5205 ( 
.A(n_4342),
.Y(n_5205)
);

AOI22xp5_ASAP7_75t_L g5206 ( 
.A1(n_3443),
.A2(n_3446),
.B1(n_3454),
.B2(n_3444),
.Y(n_5206)
);

INVx1_ASAP7_75t_L g5207 ( 
.A(n_4209),
.Y(n_5207)
);

AND2x2_ASAP7_75t_L g5208 ( 
.A(n_3157),
.B(n_3258),
.Y(n_5208)
);

AND2x2_ASAP7_75t_L g5209 ( 
.A(n_3157),
.B(n_3258),
.Y(n_5209)
);

NAND2xp5_ASAP7_75t_L g5210 ( 
.A(n_3547),
.B(n_3552),
.Y(n_5210)
);

NAND2xp5_ASAP7_75t_L g5211 ( 
.A(n_3553),
.B(n_3554),
.Y(n_5211)
);

OR2x6_ASAP7_75t_L g5212 ( 
.A(n_3989),
.B(n_3990),
.Y(n_5212)
);

NAND2xp5_ASAP7_75t_SL g5213 ( 
.A(n_4383),
.B(n_4398),
.Y(n_5213)
);

HB1xp67_ASAP7_75t_L g5214 ( 
.A(n_4418),
.Y(n_5214)
);

AND2x2_ASAP7_75t_SL g5215 ( 
.A(n_3180),
.B(n_3184),
.Y(n_5215)
);

INVx1_ASAP7_75t_L g5216 ( 
.A(n_4229),
.Y(n_5216)
);

INVxp67_ASAP7_75t_SL g5217 ( 
.A(n_4398),
.Y(n_5217)
);

AOI211xp5_ASAP7_75t_L g5218 ( 
.A1(n_3589),
.A2(n_3252),
.B(n_3464),
.C(n_3454),
.Y(n_5218)
);

INVx2_ASAP7_75t_SL g5219 ( 
.A(n_4533),
.Y(n_5219)
);

HB1xp67_ASAP7_75t_L g5220 ( 
.A(n_4418),
.Y(n_5220)
);

NAND2xp5_ASAP7_75t_L g5221 ( 
.A(n_3301),
.B(n_3544),
.Y(n_5221)
);

AOI221xp5_ASAP7_75t_L g5222 ( 
.A1(n_3464),
.A2(n_3927),
.B1(n_3943),
.B2(n_3940),
.C(n_3934),
.Y(n_5222)
);

AND2x4_ASAP7_75t_L g5223 ( 
.A(n_3496),
.B(n_3501),
.Y(n_5223)
);

NAND2xp5_ASAP7_75t_SL g5224 ( 
.A(n_4490),
.B(n_4492),
.Y(n_5224)
);

INVx3_ASAP7_75t_L g5225 ( 
.A(n_3206),
.Y(n_5225)
);

NAND2xp5_ASAP7_75t_L g5226 ( 
.A(n_3544),
.B(n_3394),
.Y(n_5226)
);

OR2x2_ASAP7_75t_L g5227 ( 
.A(n_3205),
.B(n_3212),
.Y(n_5227)
);

OAI22xp5_ASAP7_75t_SL g5228 ( 
.A1(n_3955),
.A2(n_3963),
.B1(n_3967),
.B2(n_3957),
.Y(n_5228)
);

AND2x2_ASAP7_75t_L g5229 ( 
.A(n_3276),
.B(n_3834),
.Y(n_5229)
);

INVx1_ASAP7_75t_L g5230 ( 
.A(n_4229),
.Y(n_5230)
);

INVx2_ASAP7_75t_SL g5231 ( 
.A(n_4542),
.Y(n_5231)
);

INVx1_ASAP7_75t_L g5232 ( 
.A(n_4234),
.Y(n_5232)
);

INVx5_ASAP7_75t_L g5233 ( 
.A(n_4222),
.Y(n_5233)
);

INVx3_ASAP7_75t_L g5234 ( 
.A(n_4222),
.Y(n_5234)
);

NAND2xp5_ASAP7_75t_L g5235 ( 
.A(n_3396),
.B(n_3397),
.Y(n_5235)
);

AND2x4_ASAP7_75t_L g5236 ( 
.A(n_3205),
.B(n_3212),
.Y(n_5236)
);

INVx3_ASAP7_75t_L g5237 ( 
.A(n_4222),
.Y(n_5237)
);

INVx1_ASAP7_75t_L g5238 ( 
.A(n_4234),
.Y(n_5238)
);

NOR2xp33_ASAP7_75t_L g5239 ( 
.A(n_3962),
.B(n_3972),
.Y(n_5239)
);

INVx2_ASAP7_75t_SL g5240 ( 
.A(n_3823),
.Y(n_5240)
);

NAND2x1p5_ASAP7_75t_L g5241 ( 
.A(n_4451),
.B(n_4531),
.Y(n_5241)
);

AND2x4_ASAP7_75t_L g5242 ( 
.A(n_3221),
.B(n_3303),
.Y(n_5242)
);

NAND2xp5_ASAP7_75t_L g5243 ( 
.A(n_3401),
.B(n_3404),
.Y(n_5243)
);

NOR2xp33_ASAP7_75t_L g5244 ( 
.A(n_4112),
.B(n_4127),
.Y(n_5244)
);

BUFx2_ASAP7_75t_L g5245 ( 
.A(n_4238),
.Y(n_5245)
);

A2O1A1Ixp33_ASAP7_75t_L g5246 ( 
.A1(n_3433),
.A2(n_3303),
.B(n_3305),
.C(n_3221),
.Y(n_5246)
);

NAND2xp5_ASAP7_75t_L g5247 ( 
.A(n_3480),
.B(n_3482),
.Y(n_5247)
);

AND2x2_ASAP7_75t_L g5248 ( 
.A(n_3276),
.B(n_3834),
.Y(n_5248)
);

NAND2xp5_ASAP7_75t_L g5249 ( 
.A(n_3480),
.B(n_3482),
.Y(n_5249)
);

NAND2xp5_ASAP7_75t_L g5250 ( 
.A(n_3490),
.B(n_3494),
.Y(n_5250)
);

NOR2xp33_ASAP7_75t_L g5251 ( 
.A(n_4132),
.B(n_4136),
.Y(n_5251)
);

NAND2xp5_ASAP7_75t_L g5252 ( 
.A(n_3490),
.B(n_3494),
.Y(n_5252)
);

INVx1_ASAP7_75t_L g5253 ( 
.A(n_4238),
.Y(n_5253)
);

AND2x4_ASAP7_75t_L g5254 ( 
.A(n_3305),
.B(n_3239),
.Y(n_5254)
);

BUFx3_ASAP7_75t_L g5255 ( 
.A(n_4260),
.Y(n_5255)
);

AND2x4_ASAP7_75t_L g5256 ( 
.A(n_3993),
.B(n_3994),
.Y(n_5256)
);

INVxp67_ASAP7_75t_SL g5257 ( 
.A(n_4490),
.Y(n_5257)
);

BUFx6f_ASAP7_75t_L g5258 ( 
.A(n_4451),
.Y(n_5258)
);

INVx2_ASAP7_75t_L g5259 ( 
.A(n_3463),
.Y(n_5259)
);

NAND2xp5_ASAP7_75t_SL g5260 ( 
.A(n_4492),
.B(n_3495),
.Y(n_5260)
);

NAND2xp5_ASAP7_75t_L g5261 ( 
.A(n_3503),
.B(n_3511),
.Y(n_5261)
);

OR2x2_ASAP7_75t_L g5262 ( 
.A(n_3339),
.B(n_3558),
.Y(n_5262)
);

AOI22xp33_ASAP7_75t_L g5263 ( 
.A1(n_3471),
.A2(n_4155),
.B1(n_4214),
.B2(n_4111),
.Y(n_5263)
);

INVx1_ASAP7_75t_SL g5264 ( 
.A(n_4417),
.Y(n_5264)
);

NAND2xp5_ASAP7_75t_L g5265 ( 
.A(n_3503),
.B(n_3511),
.Y(n_5265)
);

NAND2xp5_ASAP7_75t_L g5266 ( 
.A(n_3518),
.B(n_3523),
.Y(n_5266)
);

BUFx2_ASAP7_75t_L g5267 ( 
.A(n_4337),
.Y(n_5267)
);

BUFx2_ASAP7_75t_L g5268 ( 
.A(n_4337),
.Y(n_5268)
);

INVx2_ASAP7_75t_L g5269 ( 
.A(n_3463),
.Y(n_5269)
);

INVx2_ASAP7_75t_L g5270 ( 
.A(n_3476),
.Y(n_5270)
);

BUFx2_ASAP7_75t_L g5271 ( 
.A(n_4378),
.Y(n_5271)
);

AND2x4_ASAP7_75t_L g5272 ( 
.A(n_3998),
.B(n_3999),
.Y(n_5272)
);

HB1xp67_ASAP7_75t_L g5273 ( 
.A(n_4531),
.Y(n_5273)
);

INVx2_ASAP7_75t_L g5274 ( 
.A(n_3476),
.Y(n_5274)
);

NAND2xp5_ASAP7_75t_SL g5275 ( 
.A(n_3495),
.B(n_3555),
.Y(n_5275)
);

CKINVDCx6p67_ASAP7_75t_R g5276 ( 
.A(n_3181),
.Y(n_5276)
);

NAND2xp5_ASAP7_75t_L g5277 ( 
.A(n_3518),
.B(n_3523),
.Y(n_5277)
);

NAND2xp5_ASAP7_75t_L g5278 ( 
.A(n_3532),
.B(n_3534),
.Y(n_5278)
);

BUFx4f_ASAP7_75t_L g5279 ( 
.A(n_3823),
.Y(n_5279)
);

NAND2xp5_ASAP7_75t_L g5280 ( 
.A(n_3532),
.B(n_3534),
.Y(n_5280)
);

NAND2x1p5_ASAP7_75t_L g5281 ( 
.A(n_4549),
.B(n_4002),
.Y(n_5281)
);

NAND2xp5_ASAP7_75t_SL g5282 ( 
.A(n_3520),
.B(n_3433),
.Y(n_5282)
);

BUFx6f_ASAP7_75t_L g5283 ( 
.A(n_4549),
.Y(n_5283)
);

NAND2xp5_ASAP7_75t_L g5284 ( 
.A(n_3540),
.B(n_3542),
.Y(n_5284)
);

NOR2xp33_ASAP7_75t_L g5285 ( 
.A(n_4148),
.B(n_4149),
.Y(n_5285)
);

OR2x6_ASAP7_75t_L g5286 ( 
.A(n_4008),
.B(n_4010),
.Y(n_5286)
);

BUFx8_ASAP7_75t_L g5287 ( 
.A(n_3823),
.Y(n_5287)
);

NAND2xp5_ASAP7_75t_L g5288 ( 
.A(n_3540),
.B(n_3542),
.Y(n_5288)
);

NAND2xp5_ASAP7_75t_L g5289 ( 
.A(n_4150),
.B(n_4161),
.Y(n_5289)
);

INVx2_ASAP7_75t_L g5290 ( 
.A(n_3476),
.Y(n_5290)
);

INVx2_ASAP7_75t_L g5291 ( 
.A(n_3478),
.Y(n_5291)
);

HB1xp67_ASAP7_75t_L g5292 ( 
.A(n_4392),
.Y(n_5292)
);

NOR2xp33_ASAP7_75t_L g5293 ( 
.A(n_4165),
.B(n_4170),
.Y(n_5293)
);

NAND2xp5_ASAP7_75t_L g5294 ( 
.A(n_4173),
.B(n_4180),
.Y(n_5294)
);

NAND2xp5_ASAP7_75t_L g5295 ( 
.A(n_4191),
.B(n_4211),
.Y(n_5295)
);

BUFx12f_ASAP7_75t_L g5296 ( 
.A(n_3386),
.Y(n_5296)
);

BUFx4f_ASAP7_75t_L g5297 ( 
.A(n_3823),
.Y(n_5297)
);

NOR2xp33_ASAP7_75t_L g5298 ( 
.A(n_4212),
.B(n_4215),
.Y(n_5298)
);

NAND2x1p5_ASAP7_75t_L g5299 ( 
.A(n_4015),
.B(n_4016),
.Y(n_5299)
);

CKINVDCx5p33_ASAP7_75t_R g5300 ( 
.A(n_4468),
.Y(n_5300)
);

INVx4_ASAP7_75t_L g5301 ( 
.A(n_4533),
.Y(n_5301)
);

HB1xp67_ASAP7_75t_L g5302 ( 
.A(n_4393),
.Y(n_5302)
);

BUFx2_ASAP7_75t_L g5303 ( 
.A(n_4397),
.Y(n_5303)
);

AND2x2_ASAP7_75t_L g5304 ( 
.A(n_3859),
.B(n_3926),
.Y(n_5304)
);

AND2x2_ASAP7_75t_L g5305 ( 
.A(n_3859),
.B(n_3926),
.Y(n_5305)
);

INVx2_ASAP7_75t_L g5306 ( 
.A(n_3478),
.Y(n_5306)
);

CKINVDCx5p33_ASAP7_75t_R g5307 ( 
.A(n_3194),
.Y(n_5307)
);

NOR2xp67_ASAP7_75t_L g5308 ( 
.A(n_3414),
.B(n_3504),
.Y(n_5308)
);

INVx2_ASAP7_75t_L g5309 ( 
.A(n_3514),
.Y(n_5309)
);

INVx2_ASAP7_75t_SL g5310 ( 
.A(n_3823),
.Y(n_5310)
);

AND2x2_ASAP7_75t_L g5311 ( 
.A(n_3953),
.B(n_3959),
.Y(n_5311)
);

HB1xp67_ASAP7_75t_L g5312 ( 
.A(n_4445),
.Y(n_5312)
);

INVx2_ASAP7_75t_L g5313 ( 
.A(n_3514),
.Y(n_5313)
);

BUFx2_ASAP7_75t_L g5314 ( 
.A(n_4477),
.Y(n_5314)
);

NAND2xp5_ASAP7_75t_SL g5315 ( 
.A(n_3520),
.B(n_3931),
.Y(n_5315)
);

OR2x2_ASAP7_75t_SL g5316 ( 
.A(n_3460),
.B(n_3467),
.Y(n_5316)
);

BUFx2_ASAP7_75t_SL g5317 ( 
.A(n_3295),
.Y(n_5317)
);

INVx2_ASAP7_75t_L g5318 ( 
.A(n_3514),
.Y(n_5318)
);

NAND2xp5_ASAP7_75t_L g5319 ( 
.A(n_4220),
.B(n_4221),
.Y(n_5319)
);

INVx3_ASAP7_75t_L g5320 ( 
.A(n_4222),
.Y(n_5320)
);

INVxp67_ASAP7_75t_L g5321 ( 
.A(n_4454),
.Y(n_5321)
);

AOI22xp33_ASAP7_75t_L g5322 ( 
.A1(n_4341),
.A2(n_3981),
.B1(n_3997),
.B2(n_3958),
.Y(n_5322)
);

INVx2_ASAP7_75t_L g5323 ( 
.A(n_3539),
.Y(n_5323)
);

AND2x2_ASAP7_75t_L g5324 ( 
.A(n_3953),
.B(n_3959),
.Y(n_5324)
);

NOR2x1_ASAP7_75t_L g5325 ( 
.A(n_3591),
.B(n_3562),
.Y(n_5325)
);

NAND2xp5_ASAP7_75t_SL g5326 ( 
.A(n_4005),
.B(n_4007),
.Y(n_5326)
);

NAND2xp5_ASAP7_75t_L g5327 ( 
.A(n_4230),
.B(n_4232),
.Y(n_5327)
);

BUFx4f_ASAP7_75t_L g5328 ( 
.A(n_3865),
.Y(n_5328)
);

NAND2xp5_ASAP7_75t_SL g5329 ( 
.A(n_4017),
.B(n_4029),
.Y(n_5329)
);

CKINVDCx20_ASAP7_75t_R g5330 ( 
.A(n_3181),
.Y(n_5330)
);

NAND2xp5_ASAP7_75t_L g5331 ( 
.A(n_4237),
.B(n_4308),
.Y(n_5331)
);

AOI22xp5_ASAP7_75t_L g5332 ( 
.A1(n_3456),
.A2(n_3505),
.B1(n_3558),
.B2(n_4076),
.Y(n_5332)
);

A2O1A1Ixp33_ASAP7_75t_L g5333 ( 
.A1(n_4081),
.A2(n_4116),
.B(n_4154),
.C(n_4097),
.Y(n_5333)
);

A2O1A1Ixp33_ASAP7_75t_L g5334 ( 
.A1(n_4159),
.A2(n_4213),
.B(n_4219),
.C(n_4175),
.Y(n_5334)
);

BUFx6f_ASAP7_75t_L g5335 ( 
.A(n_4533),
.Y(n_5335)
);

BUFx2_ASAP7_75t_L g5336 ( 
.A(n_4489),
.Y(n_5336)
);

AOI22xp33_ASAP7_75t_L g5337 ( 
.A1(n_4326),
.A2(n_4486),
.B1(n_4354),
.B2(n_4315),
.Y(n_5337)
);

NAND2xp5_ASAP7_75t_SL g5338 ( 
.A(n_4280),
.B(n_4321),
.Y(n_5338)
);

NAND2xp5_ASAP7_75t_SL g5339 ( 
.A(n_4335),
.B(n_4356),
.Y(n_5339)
);

AOI21xp5_ASAP7_75t_L g5340 ( 
.A1(n_4030),
.A2(n_4036),
.B(n_4034),
.Y(n_5340)
);

NAND2xp5_ASAP7_75t_L g5341 ( 
.A(n_4324),
.B(n_4327),
.Y(n_5341)
);

INVx2_ASAP7_75t_SL g5342 ( 
.A(n_4533),
.Y(n_5342)
);

INVx3_ASAP7_75t_L g5343 ( 
.A(n_4222),
.Y(n_5343)
);

INVx6_ASAP7_75t_L g5344 ( 
.A(n_3230),
.Y(n_5344)
);

BUFx2_ASAP7_75t_L g5345 ( 
.A(n_4503),
.Y(n_5345)
);

AO221x1_ASAP7_75t_L g5346 ( 
.A1(n_3600),
.A2(n_4524),
.B1(n_4515),
.B2(n_3710),
.C(n_3711),
.Y(n_5346)
);

NAND2xp5_ASAP7_75t_L g5347 ( 
.A(n_4332),
.B(n_4334),
.Y(n_5347)
);

AND2x2_ASAP7_75t_L g5348 ( 
.A(n_4020),
.B(n_4024),
.Y(n_5348)
);

CKINVDCx5p33_ASAP7_75t_R g5349 ( 
.A(n_3194),
.Y(n_5349)
);

AO22x1_ASAP7_75t_L g5350 ( 
.A1(n_3600),
.A2(n_3562),
.B1(n_4024),
.B2(n_4020),
.Y(n_5350)
);

NAND2xp5_ASAP7_75t_L g5351 ( 
.A(n_4336),
.B(n_4338),
.Y(n_5351)
);

NAND2xp5_ASAP7_75t_L g5352 ( 
.A(n_4340),
.B(n_4343),
.Y(n_5352)
);

NAND2xp5_ASAP7_75t_L g5353 ( 
.A(n_4447),
.B(n_4449),
.Y(n_5353)
);

BUFx3_ASAP7_75t_L g5354 ( 
.A(n_4515),
.Y(n_5354)
);

OR2x6_ASAP7_75t_SL g5355 ( 
.A(n_3460),
.B(n_3467),
.Y(n_5355)
);

NAND2xp5_ASAP7_75t_L g5356 ( 
.A(n_4453),
.B(n_4457),
.Y(n_5356)
);

OR2x2_ASAP7_75t_L g5357 ( 
.A(n_3573),
.B(n_4045),
.Y(n_5357)
);

NAND2xp5_ASAP7_75t_SL g5358 ( 
.A(n_4379),
.B(n_4421),
.Y(n_5358)
);

BUFx2_ASAP7_75t_L g5359 ( 
.A(n_3557),
.Y(n_5359)
);

OAI22xp5_ASAP7_75t_L g5360 ( 
.A1(n_4479),
.A2(n_4499),
.B1(n_4507),
.B2(n_4480),
.Y(n_5360)
);

INVx1_ASAP7_75t_L g5361 ( 
.A(n_3560),
.Y(n_5361)
);

NAND2xp5_ASAP7_75t_SL g5362 ( 
.A(n_4452),
.B(n_4466),
.Y(n_5362)
);

INVx3_ASAP7_75t_L g5363 ( 
.A(n_4222),
.Y(n_5363)
);

HB1xp67_ASAP7_75t_L g5364 ( 
.A(n_4454),
.Y(n_5364)
);

BUFx6f_ASAP7_75t_L g5365 ( 
.A(n_4533),
.Y(n_5365)
);

INVx1_ASAP7_75t_L g5366 ( 
.A(n_3599),
.Y(n_5366)
);

INVx1_ASAP7_75t_L g5367 ( 
.A(n_3599),
.Y(n_5367)
);

AOI22xp33_ASAP7_75t_L g5368 ( 
.A1(n_4516),
.A2(n_4462),
.B1(n_4546),
.B2(n_4541),
.Y(n_5368)
);

OAI22xp5_ASAP7_75t_L g5369 ( 
.A1(n_4509),
.A2(n_4518),
.B1(n_4548),
.B2(n_4510),
.Y(n_5369)
);

NAND2xp5_ASAP7_75t_SL g5370 ( 
.A(n_3500),
.B(n_3586),
.Y(n_5370)
);

INVx1_ASAP7_75t_L g5371 ( 
.A(n_3620),
.Y(n_5371)
);

OR2x6_ASAP7_75t_L g5372 ( 
.A(n_4061),
.B(n_4078),
.Y(n_5372)
);

NAND2xp5_ASAP7_75t_L g5373 ( 
.A(n_3484),
.B(n_3235),
.Y(n_5373)
);

INVx5_ASAP7_75t_L g5374 ( 
.A(n_4502),
.Y(n_5374)
);

INVx1_ASAP7_75t_L g5375 ( 
.A(n_3620),
.Y(n_5375)
);

AND2x4_ASAP7_75t_L g5376 ( 
.A(n_4083),
.B(n_4084),
.Y(n_5376)
);

INVx1_ASAP7_75t_L g5377 ( 
.A(n_3620),
.Y(n_5377)
);

OAI22xp5_ASAP7_75t_L g5378 ( 
.A1(n_3524),
.A2(n_3249),
.B1(n_3250),
.B2(n_3248),
.Y(n_5378)
);

CKINVDCx5p33_ASAP7_75t_R g5379 ( 
.A(n_3330),
.Y(n_5379)
);

NAND2xp5_ASAP7_75t_SL g5380 ( 
.A(n_3596),
.B(n_3625),
.Y(n_5380)
);

NAND2xp5_ASAP7_75t_L g5381 ( 
.A(n_3261),
.B(n_3265),
.Y(n_5381)
);

BUFx6f_ASAP7_75t_L g5382 ( 
.A(n_4542),
.Y(n_5382)
);

NAND2xp5_ASAP7_75t_L g5383 ( 
.A(n_3266),
.B(n_3267),
.Y(n_5383)
);

NAND2xp5_ASAP7_75t_L g5384 ( 
.A(n_3268),
.B(n_3270),
.Y(n_5384)
);

NAND2xp5_ASAP7_75t_SL g5385 ( 
.A(n_3625),
.B(n_3524),
.Y(n_5385)
);

INVx1_ASAP7_75t_L g5386 ( 
.A(n_3661),
.Y(n_5386)
);

NOR2xp33_ASAP7_75t_L g5387 ( 
.A(n_3522),
.B(n_3506),
.Y(n_5387)
);

INVx1_ASAP7_75t_L g5388 ( 
.A(n_3661),
.Y(n_5388)
);

INVxp67_ASAP7_75t_SL g5389 ( 
.A(n_3298),
.Y(n_5389)
);

NAND2xp5_ASAP7_75t_L g5390 ( 
.A(n_3273),
.B(n_3281),
.Y(n_5390)
);

OR2x6_ASAP7_75t_L g5391 ( 
.A(n_4103),
.B(n_4104),
.Y(n_5391)
);

INVx1_ASAP7_75t_SL g5392 ( 
.A(n_3251),
.Y(n_5392)
);

INVx3_ASAP7_75t_L g5393 ( 
.A(n_3282),
.Y(n_5393)
);

NAND2xp5_ASAP7_75t_SL g5394 ( 
.A(n_3516),
.B(n_3605),
.Y(n_5394)
);

BUFx3_ASAP7_75t_L g5395 ( 
.A(n_3573),
.Y(n_5395)
);

INVx2_ASAP7_75t_SL g5396 ( 
.A(n_3865),
.Y(n_5396)
);

NAND2xp5_ASAP7_75t_L g5397 ( 
.A(n_3283),
.B(n_3288),
.Y(n_5397)
);

NAND2xp5_ASAP7_75t_SL g5398 ( 
.A(n_3579),
.B(n_3585),
.Y(n_5398)
);

NAND2xp5_ASAP7_75t_L g5399 ( 
.A(n_3292),
.B(n_3297),
.Y(n_5399)
);

INVx1_ASAP7_75t_L g5400 ( 
.A(n_3666),
.Y(n_5400)
);

HB1xp67_ASAP7_75t_L g5401 ( 
.A(n_3449),
.Y(n_5401)
);

AOI22xp33_ASAP7_75t_L g5402 ( 
.A1(n_4462),
.A2(n_3651),
.B1(n_3489),
.B2(n_4049),
.Y(n_5402)
);

AND2x2_ASAP7_75t_L g5403 ( 
.A(n_4049),
.B(n_4068),
.Y(n_5403)
);

HB1xp67_ASAP7_75t_L g5404 ( 
.A(n_4420),
.Y(n_5404)
);

INVx2_ASAP7_75t_L g5405 ( 
.A(n_3193),
.Y(n_5405)
);

NAND2x1p5_ASAP7_75t_L g5406 ( 
.A(n_4105),
.B(n_4109),
.Y(n_5406)
);

NOR2xp33_ASAP7_75t_L g5407 ( 
.A(n_3571),
.B(n_3672),
.Y(n_5407)
);

BUFx2_ASAP7_75t_L g5408 ( 
.A(n_3557),
.Y(n_5408)
);

NAND2xp5_ASAP7_75t_L g5409 ( 
.A(n_3299),
.B(n_3307),
.Y(n_5409)
);

INVxp67_ASAP7_75t_SL g5410 ( 
.A(n_3298),
.Y(n_5410)
);

NAND2xp5_ASAP7_75t_L g5411 ( 
.A(n_3310),
.B(n_3311),
.Y(n_5411)
);

INVx1_ASAP7_75t_L g5412 ( 
.A(n_3193),
.Y(n_5412)
);

BUFx2_ASAP7_75t_L g5413 ( 
.A(n_4068),
.Y(n_5413)
);

BUFx6f_ASAP7_75t_L g5414 ( 
.A(n_3865),
.Y(n_5414)
);

NAND2xp5_ASAP7_75t_SL g5415 ( 
.A(n_3588),
.B(n_3603),
.Y(n_5415)
);

BUFx6f_ASAP7_75t_L g5416 ( 
.A(n_3865),
.Y(n_5416)
);

HB1xp67_ASAP7_75t_L g5417 ( 
.A(n_3512),
.Y(n_5417)
);

INVxp67_ASAP7_75t_L g5418 ( 
.A(n_3703),
.Y(n_5418)
);

NAND2xp5_ASAP7_75t_L g5419 ( 
.A(n_3314),
.B(n_3316),
.Y(n_5419)
);

NAND2xp5_ASAP7_75t_SL g5420 ( 
.A(n_3690),
.B(n_3592),
.Y(n_5420)
);

INVx2_ASAP7_75t_L g5421 ( 
.A(n_3199),
.Y(n_5421)
);

HB1xp67_ASAP7_75t_L g5422 ( 
.A(n_3512),
.Y(n_5422)
);

HB1xp67_ASAP7_75t_L g5423 ( 
.A(n_3667),
.Y(n_5423)
);

BUFx6f_ASAP7_75t_L g5424 ( 
.A(n_3865),
.Y(n_5424)
);

CKINVDCx5p33_ASAP7_75t_R g5425 ( 
.A(n_3330),
.Y(n_5425)
);

INVx3_ASAP7_75t_SL g5426 ( 
.A(n_3230),
.Y(n_5426)
);

NAND2xp5_ASAP7_75t_L g5427 ( 
.A(n_3320),
.B(n_3326),
.Y(n_5427)
);

NAND2xp5_ASAP7_75t_L g5428 ( 
.A(n_3335),
.B(n_3345),
.Y(n_5428)
);

INVx2_ASAP7_75t_L g5429 ( 
.A(n_3214),
.Y(n_5429)
);

NAND2xp5_ASAP7_75t_L g5430 ( 
.A(n_3356),
.B(n_3359),
.Y(n_5430)
);

AOI22xp5_ASAP7_75t_L g5431 ( 
.A1(n_3610),
.A2(n_4090),
.B1(n_4186),
.B2(n_4163),
.Y(n_5431)
);

NAND2xp5_ASAP7_75t_SL g5432 ( 
.A(n_3690),
.B(n_3669),
.Y(n_5432)
);

NAND2xp5_ASAP7_75t_L g5433 ( 
.A(n_3366),
.B(n_3370),
.Y(n_5433)
);

AND2x4_ASAP7_75t_L g5434 ( 
.A(n_4114),
.B(n_4118),
.Y(n_5434)
);

INVx2_ASAP7_75t_L g5435 ( 
.A(n_3227),
.Y(n_5435)
);

NAND2xp5_ASAP7_75t_L g5436 ( 
.A(n_3374),
.B(n_3390),
.Y(n_5436)
);

INVx2_ASAP7_75t_L g5437 ( 
.A(n_3238),
.Y(n_5437)
);

NAND2xp5_ASAP7_75t_L g5438 ( 
.A(n_3399),
.B(n_3403),
.Y(n_5438)
);

AND2x2_ASAP7_75t_L g5439 ( 
.A(n_4090),
.B(n_4163),
.Y(n_5439)
);

BUFx6f_ASAP7_75t_L g5440 ( 
.A(n_3865),
.Y(n_5440)
);

NAND2xp5_ASAP7_75t_L g5441 ( 
.A(n_3407),
.B(n_3409),
.Y(n_5441)
);

INVx1_ASAP7_75t_SL g5442 ( 
.A(n_3251),
.Y(n_5442)
);

BUFx4f_ASAP7_75t_L g5443 ( 
.A(n_3929),
.Y(n_5443)
);

AND2x2_ASAP7_75t_L g5444 ( 
.A(n_4186),
.B(n_4195),
.Y(n_5444)
);

BUFx6f_ASAP7_75t_L g5445 ( 
.A(n_3929),
.Y(n_5445)
);

BUFx6f_ASAP7_75t_L g5446 ( 
.A(n_3929),
.Y(n_5446)
);

BUFx6f_ASAP7_75t_L g5447 ( 
.A(n_3929),
.Y(n_5447)
);

BUFx6f_ASAP7_75t_L g5448 ( 
.A(n_3929),
.Y(n_5448)
);

BUFx6f_ASAP7_75t_L g5449 ( 
.A(n_3929),
.Y(n_5449)
);

BUFx4f_ASAP7_75t_L g5450 ( 
.A(n_3935),
.Y(n_5450)
);

NOR2xp33_ASAP7_75t_L g5451 ( 
.A(n_3672),
.B(n_3531),
.Y(n_5451)
);

NAND2xp5_ASAP7_75t_L g5452 ( 
.A(n_3416),
.B(n_3422),
.Y(n_5452)
);

BUFx6f_ASAP7_75t_L g5453 ( 
.A(n_3935),
.Y(n_5453)
);

AND2x2_ASAP7_75t_L g5454 ( 
.A(n_4195),
.B(n_4207),
.Y(n_5454)
);

CKINVDCx5p33_ASAP7_75t_R g5455 ( 
.A(n_3616),
.Y(n_5455)
);

INVx2_ASAP7_75t_L g5456 ( 
.A(n_3240),
.Y(n_5456)
);

AND2x2_ASAP7_75t_L g5457 ( 
.A(n_4207),
.B(n_4233),
.Y(n_5457)
);

BUFx6f_ASAP7_75t_L g5458 ( 
.A(n_3935),
.Y(n_5458)
);

AND2x2_ASAP7_75t_L g5459 ( 
.A(n_4233),
.B(n_4254),
.Y(n_5459)
);

NAND2xp5_ASAP7_75t_L g5460 ( 
.A(n_3423),
.B(n_3424),
.Y(n_5460)
);

CKINVDCx5p33_ASAP7_75t_R g5461 ( 
.A(n_3616),
.Y(n_5461)
);

INVx2_ASAP7_75t_L g5462 ( 
.A(n_3254),
.Y(n_5462)
);

BUFx6f_ASAP7_75t_L g5463 ( 
.A(n_3935),
.Y(n_5463)
);

INVx2_ASAP7_75t_SL g5464 ( 
.A(n_3935),
.Y(n_5464)
);

NOR2x1_ASAP7_75t_L g5465 ( 
.A(n_4028),
.B(n_3230),
.Y(n_5465)
);

NAND2xp5_ASAP7_75t_SL g5466 ( 
.A(n_3669),
.B(n_3608),
.Y(n_5466)
);

INVx2_ASAP7_75t_L g5467 ( 
.A(n_3256),
.Y(n_5467)
);

BUFx3_ASAP7_75t_L g5468 ( 
.A(n_4254),
.Y(n_5468)
);

BUFx6f_ASAP7_75t_L g5469 ( 
.A(n_3950),
.Y(n_5469)
);

CKINVDCx5p33_ASAP7_75t_R g5470 ( 
.A(n_3856),
.Y(n_5470)
);

NAND2xp33_ASAP7_75t_L g5471 ( 
.A(n_3950),
.B(n_4059),
.Y(n_5471)
);

NAND2xp5_ASAP7_75t_SL g5472 ( 
.A(n_3601),
.B(n_3607),
.Y(n_5472)
);

AO22x1_ASAP7_75t_L g5473 ( 
.A1(n_4269),
.A2(n_4349),
.B1(n_4355),
.B2(n_4296),
.Y(n_5473)
);

BUFx2_ASAP7_75t_L g5474 ( 
.A(n_4269),
.Y(n_5474)
);

CKINVDCx16_ASAP7_75t_R g5475 ( 
.A(n_4296),
.Y(n_5475)
);

NAND2xp5_ASAP7_75t_L g5476 ( 
.A(n_3437),
.B(n_4349),
.Y(n_5476)
);

AOI22xp33_ASAP7_75t_L g5477 ( 
.A1(n_4355),
.A2(n_4358),
.B1(n_4386),
.B2(n_4377),
.Y(n_5477)
);

INVx2_ASAP7_75t_L g5478 ( 
.A(n_3259),
.Y(n_5478)
);

NAND2xp5_ASAP7_75t_L g5479 ( 
.A(n_4358),
.B(n_4377),
.Y(n_5479)
);

AND2x4_ASAP7_75t_L g5480 ( 
.A(n_4119),
.B(n_4120),
.Y(n_5480)
);

AOI22xp5_ASAP7_75t_L g5481 ( 
.A1(n_3610),
.A2(n_4386),
.B1(n_4467),
.B2(n_4419),
.Y(n_5481)
);

NAND2xp5_ASAP7_75t_L g5482 ( 
.A(n_4419),
.B(n_4467),
.Y(n_5482)
);

INVx4_ASAP7_75t_L g5483 ( 
.A(n_3950),
.Y(n_5483)
);

BUFx6f_ASAP7_75t_L g5484 ( 
.A(n_3950),
.Y(n_5484)
);

INVx4_ASAP7_75t_L g5485 ( 
.A(n_3950),
.Y(n_5485)
);

AOI22xp5_ASAP7_75t_L g5486 ( 
.A1(n_4470),
.A2(n_4471),
.B1(n_4495),
.B2(n_4476),
.Y(n_5486)
);

AND2x2_ASAP7_75t_L g5487 ( 
.A(n_4470),
.B(n_4471),
.Y(n_5487)
);

NAND2xp5_ASAP7_75t_L g5488 ( 
.A(n_4476),
.B(n_4495),
.Y(n_5488)
);

INVx2_ASAP7_75t_L g5489 ( 
.A(n_3275),
.Y(n_5489)
);

NAND2xp33_ASAP7_75t_SL g5490 ( 
.A(n_3696),
.B(n_3624),
.Y(n_5490)
);

INVx2_ASAP7_75t_L g5491 ( 
.A(n_3291),
.Y(n_5491)
);

INVx4_ASAP7_75t_L g5492 ( 
.A(n_3950),
.Y(n_5492)
);

HB1xp67_ASAP7_75t_L g5493 ( 
.A(n_3667),
.Y(n_5493)
);

NAND2x1p5_ASAP7_75t_L g5494 ( 
.A(n_4121),
.B(n_4123),
.Y(n_5494)
);

NOR2xp33_ASAP7_75t_R g5495 ( 
.A(n_3654),
.B(n_4528),
.Y(n_5495)
);

NAND2xp5_ASAP7_75t_L g5496 ( 
.A(n_4540),
.B(n_4543),
.Y(n_5496)
);

BUFx2_ASAP7_75t_L g5497 ( 
.A(n_4540),
.Y(n_5497)
);

NAND2xp5_ASAP7_75t_L g5498 ( 
.A(n_4543),
.B(n_3549),
.Y(n_5498)
);

INVx3_ASAP7_75t_SL g5499 ( 
.A(n_3230),
.Y(n_5499)
);

BUFx6f_ASAP7_75t_L g5500 ( 
.A(n_4059),
.Y(n_5500)
);

NOR2x1_ASAP7_75t_L g5501 ( 
.A(n_4028),
.B(n_3821),
.Y(n_5501)
);

BUFx3_ASAP7_75t_L g5502 ( 
.A(n_3893),
.Y(n_5502)
);

INVx2_ASAP7_75t_SL g5503 ( 
.A(n_4059),
.Y(n_5503)
);

BUFx2_ASAP7_75t_L g5504 ( 
.A(n_3684),
.Y(n_5504)
);

INVxp67_ASAP7_75t_L g5505 ( 
.A(n_3703),
.Y(n_5505)
);

NOR2xp33_ASAP7_75t_L g5506 ( 
.A(n_3551),
.B(n_3618),
.Y(n_5506)
);

BUFx2_ASAP7_75t_L g5507 ( 
.A(n_3684),
.Y(n_5507)
);

BUFx2_ASAP7_75t_SL g5508 ( 
.A(n_3295),
.Y(n_5508)
);

INVx2_ASAP7_75t_L g5509 ( 
.A(n_3321),
.Y(n_5509)
);

BUFx6f_ASAP7_75t_L g5510 ( 
.A(n_4059),
.Y(n_5510)
);

NAND2xp5_ASAP7_75t_SL g5511 ( 
.A(n_3601),
.B(n_3607),
.Y(n_5511)
);

AND2x4_ASAP7_75t_L g5512 ( 
.A(n_4126),
.B(n_4130),
.Y(n_5512)
);

INVx4_ASAP7_75t_L g5513 ( 
.A(n_4059),
.Y(n_5513)
);

NOR2xp33_ASAP7_75t_L g5514 ( 
.A(n_3618),
.B(n_3656),
.Y(n_5514)
);

INVx4_ASAP7_75t_L g5515 ( 
.A(n_4059),
.Y(n_5515)
);

NAND2xp5_ASAP7_75t_SL g5516 ( 
.A(n_3689),
.B(n_3613),
.Y(n_5516)
);

NAND2xp5_ASAP7_75t_L g5517 ( 
.A(n_3469),
.B(n_3502),
.Y(n_5517)
);

INVx2_ASAP7_75t_L g5518 ( 
.A(n_3324),
.Y(n_5518)
);

O2A1O1Ixp33_ASAP7_75t_L g5519 ( 
.A1(n_3710),
.A2(n_3662),
.B(n_3709),
.C(n_3659),
.Y(n_5519)
);

AND3x1_ASAP7_75t_SL g5520 ( 
.A(n_3328),
.B(n_3348),
.C(n_3331),
.Y(n_5520)
);

NAND2x2_ASAP7_75t_L g5521 ( 
.A(n_3304),
.B(n_3536),
.Y(n_5521)
);

INVx2_ASAP7_75t_L g5522 ( 
.A(n_3328),
.Y(n_5522)
);

AND2x6_ASAP7_75t_L g5523 ( 
.A(n_4072),
.B(n_4098),
.Y(n_5523)
);

INVx6_ASAP7_75t_L g5524 ( 
.A(n_3821),
.Y(n_5524)
);

OAI21xp5_ASAP7_75t_L g5525 ( 
.A1(n_4134),
.A2(n_4144),
.B(n_4138),
.Y(n_5525)
);

NOR2xp67_ASAP7_75t_L g5526 ( 
.A(n_3507),
.B(n_3617),
.Y(n_5526)
);

AOI22xp33_ASAP7_75t_L g5527 ( 
.A1(n_3656),
.A2(n_3619),
.B1(n_3566),
.B2(n_3502),
.Y(n_5527)
);

AND3x1_ASAP7_75t_SL g5528 ( 
.A(n_3331),
.B(n_3367),
.C(n_3348),
.Y(n_5528)
);

OAI22xp5_ASAP7_75t_SL g5529 ( 
.A1(n_3715),
.A2(n_3736),
.B1(n_3756),
.B2(n_3744),
.Y(n_5529)
);

BUFx2_ASAP7_75t_L g5530 ( 
.A(n_3693),
.Y(n_5530)
);

NAND2x1p5_ASAP7_75t_L g5531 ( 
.A(n_4162),
.B(n_4167),
.Y(n_5531)
);

INVxp67_ASAP7_75t_L g5532 ( 
.A(n_3703),
.Y(n_5532)
);

INVx4_ASAP7_75t_L g5533 ( 
.A(n_4072),
.Y(n_5533)
);

AND2x6_ASAP7_75t_L g5534 ( 
.A(n_4072),
.B(n_4098),
.Y(n_5534)
);

CKINVDCx5p33_ASAP7_75t_R g5535 ( 
.A(n_3856),
.Y(n_5535)
);

NAND2xp5_ASAP7_75t_SL g5536 ( 
.A(n_3609),
.B(n_3604),
.Y(n_5536)
);

NOR2xp33_ASAP7_75t_L g5537 ( 
.A(n_3469),
.B(n_3569),
.Y(n_5537)
);

INVx5_ASAP7_75t_L g5538 ( 
.A(n_4072),
.Y(n_5538)
);

HB1xp67_ASAP7_75t_L g5539 ( 
.A(n_3398),
.Y(n_5539)
);

BUFx6f_ASAP7_75t_L g5540 ( 
.A(n_4072),
.Y(n_5540)
);

NOR2xp33_ASAP7_75t_SL g5541 ( 
.A(n_3842),
.B(n_3996),
.Y(n_5541)
);

OR2x6_ASAP7_75t_L g5542 ( 
.A(n_4169),
.B(n_4171),
.Y(n_5542)
);

NOR2xp67_ASAP7_75t_L g5543 ( 
.A(n_3622),
.B(n_3626),
.Y(n_5543)
);

BUFx4f_ASAP7_75t_L g5544 ( 
.A(n_4072),
.Y(n_5544)
);

NAND2xp5_ASAP7_75t_L g5545 ( 
.A(n_3569),
.B(n_3693),
.Y(n_5545)
);

INVx1_ASAP7_75t_SL g5546 ( 
.A(n_3832),
.Y(n_5546)
);

NAND2xp5_ASAP7_75t_L g5547 ( 
.A(n_3412),
.B(n_3421),
.Y(n_5547)
);

INVxp67_ASAP7_75t_SL g5548 ( 
.A(n_4176),
.Y(n_5548)
);

NOR2xp33_ASAP7_75t_L g5549 ( 
.A(n_3680),
.B(n_3526),
.Y(n_5549)
);

BUFx6f_ASAP7_75t_L g5550 ( 
.A(n_4098),
.Y(n_5550)
);

NOR2xp33_ASAP7_75t_L g5551 ( 
.A(n_3680),
.B(n_3584),
.Y(n_5551)
);

NOR2xp33_ASAP7_75t_L g5552 ( 
.A(n_3624),
.B(n_3832),
.Y(n_5552)
);

BUFx6f_ASAP7_75t_L g5553 ( 
.A(n_4098),
.Y(n_5553)
);

INVx5_ASAP7_75t_L g5554 ( 
.A(n_4098),
.Y(n_5554)
);

AOI22xp5_ASAP7_75t_L g5555 ( 
.A1(n_3576),
.A2(n_3587),
.B1(n_3578),
.B2(n_3685),
.Y(n_5555)
);

CKINVDCx5p33_ASAP7_75t_R g5556 ( 
.A(n_4528),
.Y(n_5556)
);

NAND2xp5_ASAP7_75t_L g5557 ( 
.A(n_3426),
.B(n_3430),
.Y(n_5557)
);

AOI22xp33_ASAP7_75t_L g5558 ( 
.A1(n_3566),
.A2(n_3619),
.B1(n_3525),
.B2(n_3543),
.Y(n_5558)
);

NAND2xp5_ASAP7_75t_SL g5559 ( 
.A(n_3575),
.B(n_3636),
.Y(n_5559)
);

HB1xp67_ASAP7_75t_L g5560 ( 
.A(n_3426),
.Y(n_5560)
);

NAND2xp5_ASAP7_75t_L g5561 ( 
.A(n_3458),
.B(n_3483),
.Y(n_5561)
);

INVxp67_ASAP7_75t_L g5562 ( 
.A(n_3703),
.Y(n_5562)
);

NAND2xp5_ASAP7_75t_L g5563 ( 
.A(n_3499),
.B(n_3510),
.Y(n_5563)
);

INVxp67_ASAP7_75t_L g5564 ( 
.A(n_3597),
.Y(n_5564)
);

NAND2xp5_ASAP7_75t_L g5565 ( 
.A(n_3527),
.B(n_3546),
.Y(n_5565)
);

OR2x2_ASAP7_75t_L g5566 ( 
.A(n_4192),
.B(n_4193),
.Y(n_5566)
);

NAND2xp5_ASAP7_75t_L g5567 ( 
.A(n_3527),
.B(n_3546),
.Y(n_5567)
);

NAND2xp5_ASAP7_75t_L g5568 ( 
.A(n_3594),
.B(n_3611),
.Y(n_5568)
);

NOR2xp33_ASAP7_75t_L g5569 ( 
.A(n_3624),
.B(n_3901),
.Y(n_5569)
);

NAND2xp5_ASAP7_75t_L g5570 ( 
.A(n_3611),
.B(n_3623),
.Y(n_5570)
);

NAND2xp5_ASAP7_75t_SL g5571 ( 
.A(n_3624),
.B(n_3706),
.Y(n_5571)
);

NAND2xp5_ASAP7_75t_L g5572 ( 
.A(n_3548),
.B(n_3670),
.Y(n_5572)
);

BUFx2_ASAP7_75t_L g5573 ( 
.A(n_3629),
.Y(n_5573)
);

NAND2xp5_ASAP7_75t_L g5574 ( 
.A(n_3548),
.B(n_3670),
.Y(n_5574)
);

NAND2xp5_ASAP7_75t_L g5575 ( 
.A(n_3688),
.B(n_3597),
.Y(n_5575)
);

NAND2xp5_ASAP7_75t_SL g5576 ( 
.A(n_3624),
.B(n_4197),
.Y(n_5576)
);

INVx1_ASAP7_75t_L g5577 ( 
.A(n_3529),
.Y(n_5577)
);

INVx2_ASAP7_75t_L g5578 ( 
.A(n_3529),
.Y(n_5578)
);

INVx4_ASAP7_75t_L g5579 ( 
.A(n_4098),
.Y(n_5579)
);

INVx4_ASAP7_75t_L g5580 ( 
.A(n_4108),
.Y(n_5580)
);

NAND2xp5_ASAP7_75t_SL g5581 ( 
.A(n_3624),
.B(n_4210),
.Y(n_5581)
);

NAND2xp5_ASAP7_75t_L g5582 ( 
.A(n_3602),
.B(n_3612),
.Y(n_5582)
);

INVx1_ASAP7_75t_L g5583 ( 
.A(n_3491),
.Y(n_5583)
);

AND2x4_ASAP7_75t_L g5584 ( 
.A(n_4228),
.B(n_4239),
.Y(n_5584)
);

NAND2xp5_ASAP7_75t_L g5585 ( 
.A(n_3602),
.B(n_3612),
.Y(n_5585)
);

NAND2xp5_ASAP7_75t_L g5586 ( 
.A(n_3614),
.B(n_3621),
.Y(n_5586)
);

BUFx6f_ASAP7_75t_L g5587 ( 
.A(n_4108),
.Y(n_5587)
);

NAND2xp5_ASAP7_75t_L g5588 ( 
.A(n_3614),
.B(n_3621),
.Y(n_5588)
);

INVx3_ASAP7_75t_L g5589 ( 
.A(n_3282),
.Y(n_5589)
);

O2A1O1Ixp33_ASAP7_75t_L g5590 ( 
.A1(n_3653),
.A2(n_3711),
.B(n_3715),
.C(n_3590),
.Y(n_5590)
);

NAND2xp5_ASAP7_75t_SL g5591 ( 
.A(n_4242),
.B(n_4249),
.Y(n_5591)
);

INVx1_ASAP7_75t_L g5592 ( 
.A(n_3615),
.Y(n_5592)
);

AND2x4_ASAP7_75t_L g5593 ( 
.A(n_4257),
.B(n_4262),
.Y(n_5593)
);

INVx1_ASAP7_75t_L g5594 ( 
.A(n_3615),
.Y(n_5594)
);

BUFx6f_ASAP7_75t_L g5595 ( 
.A(n_4108),
.Y(n_5595)
);

NAND2xp5_ASAP7_75t_L g5596 ( 
.A(n_3627),
.B(n_3631),
.Y(n_5596)
);

AO221x1_ASAP7_75t_L g5597 ( 
.A1(n_3718),
.A2(n_4122),
.B1(n_4226),
.B2(n_4199),
.C(n_4108),
.Y(n_5597)
);

INVx1_ASAP7_75t_L g5598 ( 
.A(n_3649),
.Y(n_5598)
);

INVx1_ASAP7_75t_L g5599 ( 
.A(n_3649),
.Y(n_5599)
);

NAND2xp5_ASAP7_75t_L g5600 ( 
.A(n_3627),
.B(n_3631),
.Y(n_5600)
);

INVx6_ASAP7_75t_L g5601 ( 
.A(n_3821),
.Y(n_5601)
);

INVx1_ASAP7_75t_L g5602 ( 
.A(n_3635),
.Y(n_5602)
);

BUFx2_ASAP7_75t_L g5603 ( 
.A(n_3629),
.Y(n_5603)
);

AOI22xp33_ASAP7_75t_L g5604 ( 
.A1(n_3525),
.A2(n_3543),
.B1(n_3641),
.B2(n_3889),
.Y(n_5604)
);

BUFx6f_ASAP7_75t_L g5605 ( 
.A(n_4108),
.Y(n_5605)
);

NAND2xp5_ASAP7_75t_L g5606 ( 
.A(n_3635),
.B(n_3645),
.Y(n_5606)
);

INVx1_ASAP7_75t_L g5607 ( 
.A(n_3645),
.Y(n_5607)
);

HB1xp67_ASAP7_75t_L g5608 ( 
.A(n_4265),
.Y(n_5608)
);

NAND2x1p5_ASAP7_75t_L g5609 ( 
.A(n_4267),
.B(n_4273),
.Y(n_5609)
);

HB1xp67_ASAP7_75t_L g5610 ( 
.A(n_4278),
.Y(n_5610)
);

OR2x6_ASAP7_75t_L g5611 ( 
.A(n_4282),
.B(n_4287),
.Y(n_5611)
);

INVx1_ASAP7_75t_L g5612 ( 
.A(n_3646),
.Y(n_5612)
);

AND2x4_ASAP7_75t_L g5613 ( 
.A(n_4288),
.B(n_4289),
.Y(n_5613)
);

AOI22xp33_ASAP7_75t_L g5614 ( 
.A1(n_4043),
.A2(n_4217),
.B1(n_4225),
.B2(n_4128),
.Y(n_5614)
);

AND2x4_ASAP7_75t_L g5615 ( 
.A(n_4292),
.B(n_4299),
.Y(n_5615)
);

NAND2xp5_ASAP7_75t_L g5616 ( 
.A(n_3647),
.B(n_3648),
.Y(n_5616)
);

HB1xp67_ASAP7_75t_L g5617 ( 
.A(n_4306),
.Y(n_5617)
);

NAND2xp5_ASAP7_75t_L g5618 ( 
.A(n_3648),
.B(n_3657),
.Y(n_5618)
);

BUFx6f_ASAP7_75t_L g5619 ( 
.A(n_4108),
.Y(n_5619)
);

NAND2xp5_ASAP7_75t_L g5620 ( 
.A(n_3657),
.B(n_3663),
.Y(n_5620)
);

NAND2xp5_ASAP7_75t_SL g5621 ( 
.A(n_4310),
.B(n_4317),
.Y(n_5621)
);

NOR2xp33_ASAP7_75t_L g5622 ( 
.A(n_3901),
.B(n_4051),
.Y(n_5622)
);

INVx1_ASAP7_75t_L g5623 ( 
.A(n_3663),
.Y(n_5623)
);

CKINVDCx5p33_ASAP7_75t_R g5624 ( 
.A(n_3742),
.Y(n_5624)
);

INVx1_ASAP7_75t_L g5625 ( 
.A(n_3676),
.Y(n_5625)
);

NAND2xp5_ASAP7_75t_L g5626 ( 
.A(n_3637),
.B(n_4318),
.Y(n_5626)
);

BUFx12f_ASAP7_75t_L g5627 ( 
.A(n_4122),
.Y(n_5627)
);

CKINVDCx11_ASAP7_75t_R g5628 ( 
.A(n_3632),
.Y(n_5628)
);

AO22x1_ASAP7_75t_L g5629 ( 
.A1(n_3821),
.A2(n_3969),
.B1(n_3988),
.B2(n_3914),
.Y(n_5629)
);

NAND2xp5_ASAP7_75t_L g5630 ( 
.A(n_3637),
.B(n_4319),
.Y(n_5630)
);

NAND2xp5_ASAP7_75t_L g5631 ( 
.A(n_4328),
.B(n_4331),
.Y(n_5631)
);

AND2x2_ASAP7_75t_SL g5632 ( 
.A(n_3914),
.B(n_3969),
.Y(n_5632)
);

NAND2xp5_ASAP7_75t_SL g5633 ( 
.A(n_4339),
.B(n_4347),
.Y(n_5633)
);

INVx2_ASAP7_75t_SL g5634 ( 
.A(n_4122),
.Y(n_5634)
);

NAND2xp5_ASAP7_75t_L g5635 ( 
.A(n_4348),
.B(n_4359),
.Y(n_5635)
);

AND2x2_ASAP7_75t_L g5636 ( 
.A(n_4363),
.B(n_4372),
.Y(n_5636)
);

INVx2_ASAP7_75t_SL g5637 ( 
.A(n_4122),
.Y(n_5637)
);

INVx1_ASAP7_75t_L g5638 ( 
.A(n_4384),
.Y(n_5638)
);

AOI22xp5_ASAP7_75t_L g5639 ( 
.A1(n_3576),
.A2(n_3587),
.B1(n_3578),
.B2(n_3577),
.Y(n_5639)
);

AND2x2_ASAP7_75t_L g5640 ( 
.A(n_4387),
.B(n_4389),
.Y(n_5640)
);

BUFx6f_ASAP7_75t_L g5641 ( 
.A(n_4122),
.Y(n_5641)
);

NAND2xp5_ASAP7_75t_L g5642 ( 
.A(n_4390),
.B(n_4391),
.Y(n_5642)
);

INVx1_ASAP7_75t_L g5643 ( 
.A(n_4400),
.Y(n_5643)
);

INVx2_ASAP7_75t_SL g5644 ( 
.A(n_4122),
.Y(n_5644)
);

AND2x2_ASAP7_75t_L g5645 ( 
.A(n_4402),
.B(n_4409),
.Y(n_5645)
);

BUFx2_ASAP7_75t_L g5646 ( 
.A(n_3262),
.Y(n_5646)
);

NAND2xp5_ASAP7_75t_SL g5647 ( 
.A(n_4410),
.B(n_4415),
.Y(n_5647)
);

AOI22x1_ASAP7_75t_L g5648 ( 
.A1(n_4425),
.A2(n_4429),
.B1(n_4446),
.B2(n_4426),
.Y(n_5648)
);

INVx1_ASAP7_75t_L g5649 ( 
.A(n_4448),
.Y(n_5649)
);

AOI21xp5_ASAP7_75t_L g5650 ( 
.A1(n_4456),
.A2(n_4472),
.B(n_4458),
.Y(n_5650)
);

HB1xp67_ASAP7_75t_L g5651 ( 
.A(n_4473),
.Y(n_5651)
);

AND2x4_ASAP7_75t_SL g5652 ( 
.A(n_4199),
.B(n_4226),
.Y(n_5652)
);

AND2x4_ASAP7_75t_L g5653 ( 
.A(n_4496),
.B(n_4498),
.Y(n_5653)
);

BUFx2_ASAP7_75t_L g5654 ( 
.A(n_3633),
.Y(n_5654)
);

NAND2xp5_ASAP7_75t_SL g5655 ( 
.A(n_4500),
.B(n_4501),
.Y(n_5655)
);

NAND2xp5_ASAP7_75t_SL g5656 ( 
.A(n_4505),
.B(n_4526),
.Y(n_5656)
);

INVx1_ASAP7_75t_L g5657 ( 
.A(n_4527),
.Y(n_5657)
);

AND2x2_ASAP7_75t_L g5658 ( 
.A(n_3652),
.B(n_3681),
.Y(n_5658)
);

NAND2xp5_ASAP7_75t_L g5659 ( 
.A(n_3639),
.B(n_3652),
.Y(n_5659)
);

INVx4_ASAP7_75t_L g5660 ( 
.A(n_4199),
.Y(n_5660)
);

NAND2xp5_ASAP7_75t_L g5661 ( 
.A(n_3639),
.B(n_3681),
.Y(n_5661)
);

NAND2xp5_ASAP7_75t_L g5662 ( 
.A(n_3673),
.B(n_3683),
.Y(n_5662)
);

NAND2xp5_ASAP7_75t_L g5663 ( 
.A(n_3673),
.B(n_3683),
.Y(n_5663)
);

NAND2xp5_ASAP7_75t_L g5664 ( 
.A(n_3687),
.B(n_3692),
.Y(n_5664)
);

OR2x2_ASAP7_75t_L g5665 ( 
.A(n_4051),
.B(n_4182),
.Y(n_5665)
);

NOR2xp33_ASAP7_75t_SL g5666 ( 
.A(n_3842),
.B(n_3996),
.Y(n_5666)
);

OR2x2_ASAP7_75t_L g5667 ( 
.A(n_4182),
.B(n_4508),
.Y(n_5667)
);

BUFx2_ASAP7_75t_L g5668 ( 
.A(n_3633),
.Y(n_5668)
);

NAND2xp5_ASAP7_75t_L g5669 ( 
.A(n_3692),
.B(n_3697),
.Y(n_5669)
);

NAND2xp5_ASAP7_75t_L g5670 ( 
.A(n_3697),
.B(n_3698),
.Y(n_5670)
);

BUFx8_ASAP7_75t_L g5671 ( 
.A(n_4199),
.Y(n_5671)
);

HB1xp67_ASAP7_75t_L g5672 ( 
.A(n_3628),
.Y(n_5672)
);

BUFx6f_ASAP7_75t_L g5673 ( 
.A(n_4199),
.Y(n_5673)
);

NAND2xp5_ASAP7_75t_L g5674 ( 
.A(n_3701),
.B(n_3702),
.Y(n_5674)
);

INVx1_ASAP7_75t_L g5675 ( 
.A(n_3701),
.Y(n_5675)
);

NAND2xp5_ASAP7_75t_L g5676 ( 
.A(n_3702),
.B(n_3642),
.Y(n_5676)
);

INVx1_ASAP7_75t_L g5677 ( 
.A(n_3674),
.Y(n_5677)
);

BUFx6f_ASAP7_75t_L g5678 ( 
.A(n_4199),
.Y(n_5678)
);

INVx1_ASAP7_75t_L g5679 ( 
.A(n_3678),
.Y(n_5679)
);

INVx1_ASAP7_75t_SL g5680 ( 
.A(n_4508),
.Y(n_5680)
);

A2O1A1Ixp33_ASAP7_75t_L g5681 ( 
.A1(n_3630),
.A2(n_3640),
.B(n_3644),
.C(n_3650),
.Y(n_5681)
);

OR2x6_ASAP7_75t_L g5682 ( 
.A(n_4223),
.B(n_3914),
.Y(n_5682)
);

NAND2xp5_ASAP7_75t_L g5683 ( 
.A(n_3642),
.B(n_3643),
.Y(n_5683)
);

NAND2xp5_ASAP7_75t_L g5684 ( 
.A(n_3643),
.B(n_3660),
.Y(n_5684)
);

INVx1_ASAP7_75t_L g5685 ( 
.A(n_3691),
.Y(n_5685)
);

INVx1_ASAP7_75t_L g5686 ( 
.A(n_3638),
.Y(n_5686)
);

INVx2_ASAP7_75t_SL g5687 ( 
.A(n_4226),
.Y(n_5687)
);

INVx1_ASAP7_75t_L g5688 ( 
.A(n_3658),
.Y(n_5688)
);

CKINVDCx8_ASAP7_75t_R g5689 ( 
.A(n_4226),
.Y(n_5689)
);

OAI21xp5_ASAP7_75t_L g5690 ( 
.A1(n_3665),
.A2(n_3679),
.B(n_3677),
.Y(n_5690)
);

INVx1_ASAP7_75t_L g5691 ( 
.A(n_3695),
.Y(n_5691)
);

NAND2xp5_ASAP7_75t_L g5692 ( 
.A(n_3660),
.B(n_3700),
.Y(n_5692)
);

NAND2xp5_ASAP7_75t_L g5693 ( 
.A(n_3598),
.B(n_3634),
.Y(n_5693)
);

AOI22xp33_ASAP7_75t_L g5694 ( 
.A1(n_4227),
.A2(n_4244),
.B1(n_4259),
.B2(n_4513),
.Y(n_5694)
);

INVx1_ASAP7_75t_L g5695 ( 
.A(n_4218),
.Y(n_5695)
);

INVx1_ASAP7_75t_L g5696 ( 
.A(n_4218),
.Y(n_5696)
);

HB1xp67_ASAP7_75t_L g5697 ( 
.A(n_3628),
.Y(n_5697)
);

INVx1_ASAP7_75t_L g5698 ( 
.A(n_4218),
.Y(n_5698)
);

INVx3_ASAP7_75t_SL g5699 ( 
.A(n_3914),
.Y(n_5699)
);

NOR2xp67_ASAP7_75t_L g5700 ( 
.A(n_3969),
.B(n_3988),
.Y(n_5700)
);

NAND2xp5_ASAP7_75t_L g5701 ( 
.A(n_3598),
.B(n_4333),
.Y(n_5701)
);

NOR2xp33_ASAP7_75t_L g5702 ( 
.A(n_3686),
.B(n_3457),
.Y(n_5702)
);

BUFx4f_ASAP7_75t_L g5703 ( 
.A(n_4226),
.Y(n_5703)
);

NAND2xp5_ASAP7_75t_L g5704 ( 
.A(n_3598),
.B(n_4333),
.Y(n_5704)
);

NAND2xp5_ASAP7_75t_L g5705 ( 
.A(n_3598),
.B(n_4367),
.Y(n_5705)
);

AOI22xp33_ASAP7_75t_L g5706 ( 
.A1(n_4312),
.A2(n_4494),
.B1(n_4444),
.B2(n_4394),
.Y(n_5706)
);

BUFx6f_ASAP7_75t_L g5707 ( 
.A(n_4226),
.Y(n_5707)
);

NAND2xp5_ASAP7_75t_SL g5708 ( 
.A(n_3727),
.B(n_3708),
.Y(n_5708)
);

NAND2xp5_ASAP7_75t_L g5709 ( 
.A(n_4497),
.B(n_4539),
.Y(n_5709)
);

NOR2xp33_ASAP7_75t_L g5710 ( 
.A(n_3457),
.B(n_3708),
.Y(n_5710)
);

BUFx6f_ASAP7_75t_L g5711 ( 
.A(n_4248),
.Y(n_5711)
);

AOI22x1_ASAP7_75t_L g5712 ( 
.A1(n_3969),
.A2(n_4246),
.B1(n_4058),
.B2(n_3988),
.Y(n_5712)
);

NAND2xp5_ASAP7_75t_L g5713 ( 
.A(n_4539),
.B(n_3174),
.Y(n_5713)
);

AND2x2_ASAP7_75t_L g5714 ( 
.A(n_3595),
.B(n_3716),
.Y(n_5714)
);

INVx1_ASAP7_75t_L g5715 ( 
.A(n_3810),
.Y(n_5715)
);

BUFx6f_ASAP7_75t_L g5716 ( 
.A(n_4248),
.Y(n_5716)
);

BUFx6f_ASAP7_75t_L g5717 ( 
.A(n_4248),
.Y(n_5717)
);

INVx2_ASAP7_75t_L g5718 ( 
.A(n_3810),
.Y(n_5718)
);

BUFx3_ASAP7_75t_L g5719 ( 
.A(n_4248),
.Y(n_5719)
);

INVx2_ASAP7_75t_SL g5720 ( 
.A(n_4248),
.Y(n_5720)
);

INVx1_ASAP7_75t_L g5721 ( 
.A(n_4115),
.Y(n_5721)
);

CKINVDCx5p33_ASAP7_75t_R g5722 ( 
.A(n_3742),
.Y(n_5722)
);

INVx1_ASAP7_75t_L g5723 ( 
.A(n_4135),
.Y(n_5723)
);

NAND2xp5_ASAP7_75t_L g5724 ( 
.A(n_3187),
.B(n_3287),
.Y(n_5724)
);

INVx3_ASAP7_75t_L g5725 ( 
.A(n_3282),
.Y(n_5725)
);

BUFx3_ASAP7_75t_L g5726 ( 
.A(n_4248),
.Y(n_5726)
);

AOI22x1_ASAP7_75t_L g5727 ( 
.A1(n_3988),
.A2(n_4316),
.B1(n_4246),
.B2(n_4058),
.Y(n_5727)
);

INVx1_ASAP7_75t_L g5728 ( 
.A(n_4181),
.Y(n_5728)
);

INVx1_ASAP7_75t_L g5729 ( 
.A(n_3704),
.Y(n_5729)
);

AND2x4_ASAP7_75t_L g5730 ( 
.A(n_3282),
.B(n_3378),
.Y(n_5730)
);

INVx2_ASAP7_75t_L g5731 ( 
.A(n_3282),
.Y(n_5731)
);

NOR2xp33_ASAP7_75t_L g5732 ( 
.A(n_3721),
.B(n_3831),
.Y(n_5732)
);

AOI22xp5_ASAP7_75t_L g5733 ( 
.A1(n_3788),
.A2(n_3789),
.B1(n_3593),
.B2(n_3595),
.Y(n_5733)
);

AOI22xp33_ASAP7_75t_L g5734 ( 
.A1(n_3736),
.A2(n_3756),
.B1(n_3789),
.B2(n_3593),
.Y(n_5734)
);

INVx1_ASAP7_75t_L g5735 ( 
.A(n_4264),
.Y(n_5735)
);

BUFx3_ASAP7_75t_L g5736 ( 
.A(n_4264),
.Y(n_5736)
);

BUFx2_ASAP7_75t_L g5737 ( 
.A(n_3862),
.Y(n_5737)
);

NOR2xp33_ASAP7_75t_L g5738 ( 
.A(n_3721),
.B(n_4064),
.Y(n_5738)
);

NAND2xp5_ASAP7_75t_L g5739 ( 
.A(n_4139),
.B(n_4298),
.Y(n_5739)
);

HB1xp67_ASAP7_75t_L g5740 ( 
.A(n_4484),
.Y(n_5740)
);

INVx2_ASAP7_75t_L g5741 ( 
.A(n_3282),
.Y(n_5741)
);

AND2x4_ASAP7_75t_L g5742 ( 
.A(n_3378),
.B(n_3408),
.Y(n_5742)
);

AND2x2_ASAP7_75t_L g5743 ( 
.A(n_3595),
.B(n_3716),
.Y(n_5743)
);

NAND2xp5_ASAP7_75t_L g5744 ( 
.A(n_4547),
.B(n_3595),
.Y(n_5744)
);

OR2x2_ASAP7_75t_L g5745 ( 
.A(n_3718),
.B(n_4264),
.Y(n_5745)
);

NOR2xp33_ASAP7_75t_L g5746 ( 
.A(n_3792),
.B(n_3720),
.Y(n_5746)
);

NAND2xp5_ASAP7_75t_L g5747 ( 
.A(n_3720),
.B(n_3593),
.Y(n_5747)
);

NAND2xp5_ASAP7_75t_L g5748 ( 
.A(n_3593),
.B(n_4264),
.Y(n_5748)
);

NAND2xp5_ASAP7_75t_SL g5749 ( 
.A(n_3727),
.B(n_4264),
.Y(n_5749)
);

NOR2xp33_ASAP7_75t_L g5750 ( 
.A(n_3792),
.B(n_3743),
.Y(n_5750)
);

BUFx12f_ASAP7_75t_L g5751 ( 
.A(n_4264),
.Y(n_5751)
);

INVx1_ASAP7_75t_L g5752 ( 
.A(n_4281),
.Y(n_5752)
);

NAND2xp5_ASAP7_75t_L g5753 ( 
.A(n_4281),
.B(n_4303),
.Y(n_5753)
);

NAND2xp5_ASAP7_75t_L g5754 ( 
.A(n_4281),
.B(n_4303),
.Y(n_5754)
);

INVx1_ASAP7_75t_L g5755 ( 
.A(n_4281),
.Y(n_5755)
);

INVx2_ASAP7_75t_L g5756 ( 
.A(n_3378),
.Y(n_5756)
);

INVx1_ASAP7_75t_L g5757 ( 
.A(n_4281),
.Y(n_5757)
);

INVx1_ASAP7_75t_L g5758 ( 
.A(n_4281),
.Y(n_5758)
);

NAND2xp5_ASAP7_75t_L g5759 ( 
.A(n_4303),
.B(n_4502),
.Y(n_5759)
);

INVx1_ASAP7_75t_L g5760 ( 
.A(n_4303),
.Y(n_5760)
);

INVx1_ASAP7_75t_L g5761 ( 
.A(n_4303),
.Y(n_5761)
);

NOR2x1_ASAP7_75t_L g5762 ( 
.A(n_4058),
.B(n_4246),
.Y(n_5762)
);

BUFx2_ASAP7_75t_L g5763 ( 
.A(n_4303),
.Y(n_5763)
);

INVx2_ASAP7_75t_L g5764 ( 
.A(n_4896),
.Y(n_5764)
);

NAND2xp5_ASAP7_75t_SL g5765 ( 
.A(n_5014),
.B(n_4502),
.Y(n_5765)
);

AND2x2_ASAP7_75t_SL g5766 ( 
.A(n_5014),
.B(n_4058),
.Y(n_5766)
);

OAI22xp5_ASAP7_75t_L g5767 ( 
.A1(n_4785),
.A2(n_3744),
.B1(n_3787),
.B2(n_3707),
.Y(n_5767)
);

INVx4_ASAP7_75t_L g5768 ( 
.A(n_5082),
.Y(n_5768)
);

OAI22xp33_ASAP7_75t_L g5769 ( 
.A1(n_4671),
.A2(n_3713),
.B1(n_3712),
.B2(n_4316),
.Y(n_5769)
);

OAI22xp5_ASAP7_75t_L g5770 ( 
.A1(n_4785),
.A2(n_3744),
.B1(n_3729),
.B2(n_4205),
.Y(n_5770)
);

INVx4_ASAP7_75t_L g5771 ( 
.A(n_5082),
.Y(n_5771)
);

NAND2xp5_ASAP7_75t_L g5772 ( 
.A(n_5113),
.B(n_3753),
.Y(n_5772)
);

INVx2_ASAP7_75t_L g5773 ( 
.A(n_4896),
.Y(n_5773)
);

OAI22xp5_ASAP7_75t_SL g5774 ( 
.A1(n_4712),
.A2(n_3769),
.B1(n_3729),
.B2(n_3767),
.Y(n_5774)
);

AOI21xp5_ASAP7_75t_L g5775 ( 
.A1(n_5398),
.A2(n_5093),
.B(n_5092),
.Y(n_5775)
);

NAND2xp5_ASAP7_75t_L g5776 ( 
.A(n_4613),
.B(n_3719),
.Y(n_5776)
);

INVx1_ASAP7_75t_L g5777 ( 
.A(n_5412),
.Y(n_5777)
);

OAI21xp5_ASAP7_75t_L g5778 ( 
.A1(n_4594),
.A2(n_3802),
.B(n_3487),
.Y(n_5778)
);

CKINVDCx5p33_ASAP7_75t_R g5779 ( 
.A(n_4558),
.Y(n_5779)
);

BUFx6f_ASAP7_75t_L g5780 ( 
.A(n_4658),
.Y(n_5780)
);

INVx1_ASAP7_75t_L g5781 ( 
.A(n_5412),
.Y(n_5781)
);

NAND2xp5_ASAP7_75t_SL g5782 ( 
.A(n_5014),
.B(n_4502),
.Y(n_5782)
);

AOI22xp5_ASAP7_75t_L g5783 ( 
.A1(n_4579),
.A2(n_4757),
.B1(n_4712),
.B2(n_4773),
.Y(n_5783)
);

BUFx6f_ASAP7_75t_L g5784 ( 
.A(n_4658),
.Y(n_5784)
);

INVx1_ASAP7_75t_L g5785 ( 
.A(n_5412),
.Y(n_5785)
);

AOI21xp5_ASAP7_75t_L g5786 ( 
.A1(n_5398),
.A2(n_3802),
.B(n_3411),
.Y(n_5786)
);

O2A1O1Ixp33_ASAP7_75t_L g5787 ( 
.A1(n_4594),
.A2(n_3733),
.B(n_3664),
.C(n_3682),
.Y(n_5787)
);

AOI22xp5_ASAP7_75t_L g5788 ( 
.A1(n_4579),
.A2(n_3761),
.B1(n_3758),
.B2(n_3517),
.Y(n_5788)
);

NAND2xp5_ASAP7_75t_L g5789 ( 
.A(n_4592),
.B(n_3725),
.Y(n_5789)
);

NOR2xp33_ASAP7_75t_L g5790 ( 
.A(n_4899),
.B(n_3378),
.Y(n_5790)
);

INVx2_ASAP7_75t_SL g5791 ( 
.A(n_4916),
.Y(n_5791)
);

AOI21xp5_ASAP7_75t_L g5792 ( 
.A1(n_5092),
.A2(n_4205),
.B(n_3376),
.Y(n_5792)
);

O2A1O1Ixp33_ASAP7_75t_L g5793 ( 
.A1(n_4694),
.A2(n_3767),
.B(n_3748),
.C(n_3752),
.Y(n_5793)
);

AOI21xp5_ASAP7_75t_L g5794 ( 
.A1(n_5093),
.A2(n_3411),
.B(n_3376),
.Y(n_5794)
);

NOR2xp33_ASAP7_75t_L g5795 ( 
.A(n_4899),
.B(n_4757),
.Y(n_5795)
);

BUFx2_ASAP7_75t_L g5796 ( 
.A(n_4979),
.Y(n_5796)
);

AOI221xp5_ASAP7_75t_L g5797 ( 
.A1(n_4639),
.A2(n_4618),
.B1(n_4692),
.B2(n_4667),
.C(n_4566),
.Y(n_5797)
);

INVx2_ASAP7_75t_L g5798 ( 
.A(n_4896),
.Y(n_5798)
);

NAND2xp5_ASAP7_75t_L g5799 ( 
.A(n_4646),
.B(n_3734),
.Y(n_5799)
);

HB1xp67_ASAP7_75t_L g5800 ( 
.A(n_4557),
.Y(n_5800)
);

NOR2xp33_ASAP7_75t_R g5801 ( 
.A(n_4558),
.B(n_3632),
.Y(n_5801)
);

NAND2xp5_ASAP7_75t_L g5802 ( 
.A(n_4649),
.B(n_3734),
.Y(n_5802)
);

OAI22xp5_ASAP7_75t_L g5803 ( 
.A1(n_4688),
.A2(n_3487),
.B1(n_3774),
.B2(n_3784),
.Y(n_5803)
);

BUFx3_ASAP7_75t_L g5804 ( 
.A(n_5502),
.Y(n_5804)
);

O2A1O1Ixp33_ASAP7_75t_L g5805 ( 
.A1(n_4694),
.A2(n_3752),
.B(n_3738),
.C(n_3730),
.Y(n_5805)
);

INVx4_ASAP7_75t_L g5806 ( 
.A(n_5082),
.Y(n_5806)
);

OAI21xp5_ASAP7_75t_L g5807 ( 
.A1(n_4741),
.A2(n_3738),
.B(n_3741),
.Y(n_5807)
);

OR2x2_ASAP7_75t_L g5808 ( 
.A(n_5357),
.B(n_3735),
.Y(n_5808)
);

INVx2_ASAP7_75t_L g5809 ( 
.A(n_4896),
.Y(n_5809)
);

A2O1A1Ixp33_ASAP7_75t_L g5810 ( 
.A1(n_5519),
.A2(n_3717),
.B(n_3731),
.C(n_3723),
.Y(n_5810)
);

OR2x6_ASAP7_75t_L g5811 ( 
.A(n_4734),
.B(n_4746),
.Y(n_5811)
);

INVx4_ASAP7_75t_L g5812 ( 
.A(n_5082),
.Y(n_5812)
);

INVx1_ASAP7_75t_SL g5813 ( 
.A(n_5392),
.Y(n_5813)
);

BUFx6f_ASAP7_75t_L g5814 ( 
.A(n_4658),
.Y(n_5814)
);

INVx1_ASAP7_75t_SL g5815 ( 
.A(n_5392),
.Y(n_5815)
);

INVx4_ASAP7_75t_L g5816 ( 
.A(n_5082),
.Y(n_5816)
);

CKINVDCx20_ASAP7_75t_R g5817 ( 
.A(n_4864),
.Y(n_5817)
);

NAND2xp5_ASAP7_75t_L g5818 ( 
.A(n_4649),
.B(n_3735),
.Y(n_5818)
);

AOI21xp5_ASAP7_75t_L g5819 ( 
.A1(n_5094),
.A2(n_5101),
.B(n_5100),
.Y(n_5819)
);

AOI22xp33_ASAP7_75t_L g5820 ( 
.A1(n_4688),
.A2(n_3761),
.B1(n_3747),
.B2(n_3714),
.Y(n_5820)
);

AND2x4_ASAP7_75t_L g5821 ( 
.A(n_4832),
.B(n_3378),
.Y(n_5821)
);

INVx4_ASAP7_75t_L g5822 ( 
.A(n_5082),
.Y(n_5822)
);

AOI21xp5_ASAP7_75t_L g5823 ( 
.A1(n_5094),
.A2(n_4537),
.B(n_4246),
.Y(n_5823)
);

BUFx2_ASAP7_75t_L g5824 ( 
.A(n_4979),
.Y(n_5824)
);

CKINVDCx5p33_ASAP7_75t_R g5825 ( 
.A(n_4678),
.Y(n_5825)
);

NOR2xp33_ASAP7_75t_SL g5826 ( 
.A(n_4792),
.B(n_4316),
.Y(n_5826)
);

BUFx6f_ASAP7_75t_L g5827 ( 
.A(n_4658),
.Y(n_5827)
);

OAI22xp5_ASAP7_75t_L g5828 ( 
.A1(n_4641),
.A2(n_3774),
.B1(n_4537),
.B2(n_4316),
.Y(n_5828)
);

AOI21xp5_ASAP7_75t_L g5829 ( 
.A1(n_5100),
.A2(n_4537),
.B(n_4542),
.Y(n_5829)
);

OR2x2_ASAP7_75t_L g5830 ( 
.A(n_5357),
.B(n_3735),
.Y(n_5830)
);

BUFx3_ASAP7_75t_L g5831 ( 
.A(n_5502),
.Y(n_5831)
);

AOI22xp33_ASAP7_75t_L g5832 ( 
.A1(n_4827),
.A2(n_3747),
.B1(n_3535),
.B2(n_3517),
.Y(n_5832)
);

INVx2_ASAP7_75t_L g5833 ( 
.A(n_4914),
.Y(n_5833)
);

INVx3_ASAP7_75t_SL g5834 ( 
.A(n_5394),
.Y(n_5834)
);

NAND2xp5_ASAP7_75t_L g5835 ( 
.A(n_4650),
.B(n_3768),
.Y(n_5835)
);

O2A1O1Ixp33_ASAP7_75t_L g5836 ( 
.A1(n_4741),
.A2(n_3770),
.B(n_3775),
.C(n_3783),
.Y(n_5836)
);

AOI22xp5_ASAP7_75t_L g5837 ( 
.A1(n_4773),
.A2(n_3517),
.B1(n_3537),
.B2(n_3535),
.Y(n_5837)
);

NOR3xp33_ASAP7_75t_L g5838 ( 
.A(n_4676),
.B(n_4537),
.C(n_3764),
.Y(n_5838)
);

AOI22xp33_ASAP7_75t_L g5839 ( 
.A1(n_4827),
.A2(n_3537),
.B1(n_3535),
.B2(n_3517),
.Y(n_5839)
);

INVxp67_ASAP7_75t_L g5840 ( 
.A(n_4557),
.Y(n_5840)
);

BUFx8_ASAP7_75t_SL g5841 ( 
.A(n_4578),
.Y(n_5841)
);

AOI21xp5_ASAP7_75t_L g5842 ( 
.A1(n_5101),
.A2(n_4542),
.B(n_4502),
.Y(n_5842)
);

CKINVDCx5p33_ASAP7_75t_R g5843 ( 
.A(n_4678),
.Y(n_5843)
);

NOR2xp33_ASAP7_75t_L g5844 ( 
.A(n_4941),
.B(n_5221),
.Y(n_5844)
);

BUFx2_ASAP7_75t_L g5845 ( 
.A(n_4979),
.Y(n_5845)
);

AND2x2_ASAP7_75t_L g5846 ( 
.A(n_4581),
.B(n_3768),
.Y(n_5846)
);

NAND2xp5_ASAP7_75t_L g5847 ( 
.A(n_4650),
.B(n_3768),
.Y(n_5847)
);

AOI21xp5_ASAP7_75t_L g5848 ( 
.A1(n_4699),
.A2(n_4542),
.B(n_4502),
.Y(n_5848)
);

O2A1O1Ixp33_ASAP7_75t_L g5849 ( 
.A1(n_4676),
.A2(n_3783),
.B(n_3745),
.C(n_3751),
.Y(n_5849)
);

NAND2xp5_ASAP7_75t_SL g5850 ( 
.A(n_5014),
.B(n_3408),
.Y(n_5850)
);

OAI22xp5_ASAP7_75t_L g5851 ( 
.A1(n_4641),
.A2(n_3537),
.B1(n_3535),
.B2(n_3304),
.Y(n_5851)
);

INVx2_ASAP7_75t_SL g5852 ( 
.A(n_4916),
.Y(n_5852)
);

OR2x2_ASAP7_75t_L g5853 ( 
.A(n_5357),
.B(n_3771),
.Y(n_5853)
);

INVx2_ASAP7_75t_L g5854 ( 
.A(n_4914),
.Y(n_5854)
);

O2A1O1Ixp5_ASAP7_75t_L g5855 ( 
.A1(n_4728),
.A2(n_3537),
.B(n_3757),
.C(n_3750),
.Y(n_5855)
);

INVxp67_ASAP7_75t_SL g5856 ( 
.A(n_4553),
.Y(n_5856)
);

A2O1A1Ixp33_ASAP7_75t_L g5857 ( 
.A1(n_5519),
.A2(n_3364),
.B(n_4455),
.C(n_3304),
.Y(n_5857)
);

BUFx2_ASAP7_75t_L g5858 ( 
.A(n_4979),
.Y(n_5858)
);

NOR2xp33_ASAP7_75t_SL g5859 ( 
.A(n_4792),
.B(n_3696),
.Y(n_5859)
);

INVx5_ASAP7_75t_L g5860 ( 
.A(n_4946),
.Y(n_5860)
);

OAI22x1_ASAP7_75t_L g5861 ( 
.A1(n_5039),
.A2(n_3750),
.B1(n_3757),
.B2(n_3771),
.Y(n_5861)
);

CKINVDCx16_ASAP7_75t_R g5862 ( 
.A(n_5076),
.Y(n_5862)
);

INVx2_ASAP7_75t_L g5863 ( 
.A(n_4914),
.Y(n_5863)
);

BUFx6f_ASAP7_75t_L g5864 ( 
.A(n_4658),
.Y(n_5864)
);

BUFx6f_ASAP7_75t_L g5865 ( 
.A(n_4658),
.Y(n_5865)
);

INVx2_ASAP7_75t_L g5866 ( 
.A(n_4914),
.Y(n_5866)
);

NOR2xp33_ASAP7_75t_L g5867 ( 
.A(n_4941),
.B(n_3408),
.Y(n_5867)
);

INVx3_ASAP7_75t_L g5868 ( 
.A(n_4713),
.Y(n_5868)
);

INVx3_ASAP7_75t_L g5869 ( 
.A(n_4713),
.Y(n_5869)
);

AOI21xp5_ASAP7_75t_L g5870 ( 
.A1(n_4699),
.A2(n_3408),
.B(n_3364),
.Y(n_5870)
);

O2A1O1Ixp33_ASAP7_75t_L g5871 ( 
.A1(n_4728),
.A2(n_3765),
.B(n_3754),
.C(n_3781),
.Y(n_5871)
);

NOR2xp33_ASAP7_75t_SL g5872 ( 
.A(n_5111),
.B(n_3696),
.Y(n_5872)
);

BUFx12f_ASAP7_75t_L g5873 ( 
.A(n_4578),
.Y(n_5873)
);

HB1xp67_ASAP7_75t_L g5874 ( 
.A(n_4573),
.Y(n_5874)
);

O2A1O1Ixp33_ASAP7_75t_L g5875 ( 
.A1(n_4748),
.A2(n_3772),
.B(n_3746),
.C(n_3781),
.Y(n_5875)
);

INVx2_ASAP7_75t_SL g5876 ( 
.A(n_4916),
.Y(n_5876)
);

AOI22xp33_ASAP7_75t_L g5877 ( 
.A1(n_5062),
.A2(n_3762),
.B1(n_3740),
.B2(n_3408),
.Y(n_5877)
);

NAND2xp5_ASAP7_75t_L g5878 ( 
.A(n_4662),
.B(n_3732),
.Y(n_5878)
);

OAI21xp5_ASAP7_75t_L g5879 ( 
.A1(n_4692),
.A2(n_3777),
.B(n_3766),
.Y(n_5879)
);

NAND2xp5_ASAP7_75t_SL g5880 ( 
.A(n_4566),
.B(n_5332),
.Y(n_5880)
);

OAI22xp5_ASAP7_75t_L g5881 ( 
.A1(n_5018),
.A2(n_4535),
.B1(n_4455),
.B2(n_4004),
.Y(n_5881)
);

INVx2_ASAP7_75t_L g5882 ( 
.A(n_4940),
.Y(n_5882)
);

AOI21xp5_ASAP7_75t_L g5883 ( 
.A1(n_4747),
.A2(n_3364),
.B(n_3763),
.Y(n_5883)
);

HB1xp67_ASAP7_75t_L g5884 ( 
.A(n_4573),
.Y(n_5884)
);

OAI22xp33_ASAP7_75t_L g5885 ( 
.A1(n_4671),
.A2(n_3696),
.B1(n_4455),
.B2(n_3536),
.Y(n_5885)
);

BUFx8_ASAP7_75t_L g5886 ( 
.A(n_5193),
.Y(n_5886)
);

AND2x2_ASAP7_75t_L g5887 ( 
.A(n_4581),
.B(n_4617),
.Y(n_5887)
);

OAI22xp5_ASAP7_75t_L g5888 ( 
.A1(n_5018),
.A2(n_4535),
.B1(n_4404),
.B2(n_3536),
.Y(n_5888)
);

INVx5_ASAP7_75t_L g5889 ( 
.A(n_4946),
.Y(n_5889)
);

AO22x1_ASAP7_75t_L g5890 ( 
.A1(n_4857),
.A2(n_4535),
.B1(n_4404),
.B2(n_3699),
.Y(n_5890)
);

HB1xp67_ASAP7_75t_L g5891 ( 
.A(n_5404),
.Y(n_5891)
);

BUFx3_ASAP7_75t_L g5892 ( 
.A(n_5502),
.Y(n_5892)
);

NAND3xp33_ASAP7_75t_L g5893 ( 
.A(n_4754),
.B(n_3722),
.C(n_3739),
.Y(n_5893)
);

AND2x2_ASAP7_75t_L g5894 ( 
.A(n_4581),
.B(n_3724),
.Y(n_5894)
);

NAND2x1_ASAP7_75t_L g5895 ( 
.A(n_5597),
.B(n_3732),
.Y(n_5895)
);

OAI22xp33_ASAP7_75t_L g5896 ( 
.A1(n_4675),
.A2(n_4004),
.B1(n_4404),
.B2(n_3699),
.Y(n_5896)
);

AND2x4_ASAP7_75t_L g5897 ( 
.A(n_4832),
.B(n_4366),
.Y(n_5897)
);

OAI22xp5_ASAP7_75t_L g5898 ( 
.A1(n_4754),
.A2(n_4004),
.B1(n_4366),
.B2(n_3699),
.Y(n_5898)
);

NAND2xp5_ASAP7_75t_L g5899 ( 
.A(n_4662),
.B(n_3732),
.Y(n_5899)
);

INVx2_ASAP7_75t_L g5900 ( 
.A(n_4940),
.Y(n_5900)
);

OR2x2_ASAP7_75t_L g5901 ( 
.A(n_5359),
.B(n_3779),
.Y(n_5901)
);

INVx3_ASAP7_75t_L g5902 ( 
.A(n_4713),
.Y(n_5902)
);

INVx2_ASAP7_75t_L g5903 ( 
.A(n_4940),
.Y(n_5903)
);

INVx4_ASAP7_75t_L g5904 ( 
.A(n_5082),
.Y(n_5904)
);

INVx2_ASAP7_75t_L g5905 ( 
.A(n_4940),
.Y(n_5905)
);

OAI22xp5_ASAP7_75t_L g5906 ( 
.A1(n_4820),
.A2(n_4066),
.B1(n_4366),
.B2(n_4362),
.Y(n_5906)
);

HB1xp67_ASAP7_75t_L g5907 ( 
.A(n_5404),
.Y(n_5907)
);

OR2x6_ASAP7_75t_L g5908 ( 
.A(n_4734),
.B(n_4066),
.Y(n_5908)
);

AOI22xp5_ASAP7_75t_L g5909 ( 
.A1(n_4638),
.A2(n_4656),
.B1(n_4722),
.B2(n_4691),
.Y(n_5909)
);

NOR2x1_ASAP7_75t_L g5910 ( 
.A(n_4684),
.B(n_4066),
.Y(n_5910)
);

AOI21xp5_ASAP7_75t_L g5911 ( 
.A1(n_4747),
.A2(n_5164),
.B(n_5127),
.Y(n_5911)
);

AOI21xp5_ASAP7_75t_L g5912 ( 
.A1(n_5127),
.A2(n_3763),
.B(n_3780),
.Y(n_5912)
);

O2A1O1Ixp33_ASAP7_75t_L g5913 ( 
.A1(n_4748),
.A2(n_3778),
.B(n_3779),
.C(n_3780),
.Y(n_5913)
);

AOI21x1_ASAP7_75t_L g5914 ( 
.A1(n_5275),
.A2(n_3773),
.B(n_3755),
.Y(n_5914)
);

O2A1O1Ixp33_ASAP7_75t_SL g5915 ( 
.A1(n_5040),
.A2(n_3773),
.B(n_3778),
.C(n_3772),
.Y(n_5915)
);

AND2x2_ASAP7_75t_L g5916 ( 
.A(n_4617),
.B(n_3724),
.Y(n_5916)
);

OR2x6_ASAP7_75t_L g5917 ( 
.A(n_4734),
.B(n_4362),
.Y(n_5917)
);

AOI21xp5_ASAP7_75t_L g5918 ( 
.A1(n_5164),
.A2(n_3763),
.B(n_3755),
.Y(n_5918)
);

INVxp67_ASAP7_75t_SL g5919 ( 
.A(n_4553),
.Y(n_5919)
);

INVx4_ASAP7_75t_L g5920 ( 
.A(n_5082),
.Y(n_5920)
);

NOR2xp33_ASAP7_75t_L g5921 ( 
.A(n_5221),
.B(n_3732),
.Y(n_5921)
);

INVx2_ASAP7_75t_L g5922 ( 
.A(n_4942),
.Y(n_5922)
);

O2A1O1Ixp33_ASAP7_75t_L g5923 ( 
.A1(n_4706),
.A2(n_3754),
.B(n_3726),
.C(n_3749),
.Y(n_5923)
);

AOI21xp33_ASAP7_75t_L g5924 ( 
.A1(n_4767),
.A2(n_3749),
.B(n_3726),
.Y(n_5924)
);

AOI22xp33_ASAP7_75t_L g5925 ( 
.A1(n_5062),
.A2(n_3762),
.B1(n_3740),
.B2(n_4190),
.Y(n_5925)
);

NOR2xp33_ASAP7_75t_L g5926 ( 
.A(n_4706),
.B(n_3746),
.Y(n_5926)
);

NAND2xp5_ASAP7_75t_L g5927 ( 
.A(n_4663),
.B(n_4677),
.Y(n_5927)
);

AOI21xp5_ASAP7_75t_L g5928 ( 
.A1(n_5340),
.A2(n_3763),
.B(n_3739),
.Y(n_5928)
);

OAI22xp5_ASAP7_75t_L g5929 ( 
.A1(n_4820),
.A2(n_4362),
.B1(n_4330),
.B2(n_4300),
.Y(n_5929)
);

BUFx3_ASAP7_75t_L g5930 ( 
.A(n_5502),
.Y(n_5930)
);

INVxp33_ASAP7_75t_SL g5931 ( 
.A(n_4633),
.Y(n_5931)
);

NAND2xp5_ASAP7_75t_L g5932 ( 
.A(n_4663),
.B(n_3763),
.Y(n_5932)
);

INVx2_ASAP7_75t_SL g5933 ( 
.A(n_4916),
.Y(n_5933)
);

INVx4_ASAP7_75t_L g5934 ( 
.A(n_5082),
.Y(n_5934)
);

NOR2x1_ASAP7_75t_L g5935 ( 
.A(n_4684),
.B(n_4330),
.Y(n_5935)
);

AND2x2_ASAP7_75t_L g5936 ( 
.A(n_4617),
.B(n_3763),
.Y(n_5936)
);

INVx4_ASAP7_75t_L g5937 ( 
.A(n_5233),
.Y(n_5937)
);

BUFx6f_ASAP7_75t_L g5938 ( 
.A(n_4658),
.Y(n_5938)
);

O2A1O1Ixp5_ASAP7_75t_SL g5939 ( 
.A1(n_5275),
.A2(n_3737),
.B(n_3786),
.C(n_3986),
.Y(n_5939)
);

INVx3_ASAP7_75t_L g5940 ( 
.A(n_4713),
.Y(n_5940)
);

AOI21xp5_ASAP7_75t_L g5941 ( 
.A1(n_5340),
.A2(n_3737),
.B(n_3285),
.Y(n_5941)
);

A2O1A1Ixp33_ASAP7_75t_SL g5942 ( 
.A1(n_4859),
.A2(n_4599),
.B(n_4656),
.C(n_4638),
.Y(n_5942)
);

NAND2xp5_ASAP7_75t_L g5943 ( 
.A(n_4677),
.B(n_4683),
.Y(n_5943)
);

O2A1O1Ixp5_ASAP7_75t_SL g5944 ( 
.A1(n_5260),
.A2(n_3172),
.B(n_3285),
.C(n_4428),
.Y(n_5944)
);

AND2x2_ASAP7_75t_L g5945 ( 
.A(n_4647),
.B(n_3172),
.Y(n_5945)
);

AND2x2_ASAP7_75t_L g5946 ( 
.A(n_4647),
.B(n_4046),
.Y(n_5946)
);

AND2x2_ASAP7_75t_L g5947 ( 
.A(n_4647),
.B(n_4046),
.Y(n_5947)
);

INVx8_ASAP7_75t_L g5948 ( 
.A(n_5035),
.Y(n_5948)
);

AOI21xp5_ASAP7_75t_L g5949 ( 
.A1(n_5650),
.A2(n_4050),
.B(n_4052),
.Y(n_5949)
);

NAND2xp5_ASAP7_75t_L g5950 ( 
.A(n_4683),
.B(n_4050),
.Y(n_5950)
);

INVx5_ASAP7_75t_L g5951 ( 
.A(n_4946),
.Y(n_5951)
);

O2A1O1Ixp33_ASAP7_75t_L g5952 ( 
.A1(n_4639),
.A2(n_4330),
.B(n_4300),
.C(n_4272),
.Y(n_5952)
);

AOI22xp33_ASAP7_75t_SL g5953 ( 
.A1(n_4691),
.A2(n_4300),
.B1(n_4272),
.B2(n_4190),
.Y(n_5953)
);

AOI22xp33_ASAP7_75t_L g5954 ( 
.A1(n_4722),
.A2(n_3740),
.B1(n_3762),
.B2(n_4272),
.Y(n_5954)
);

O2A1O1Ixp5_ASAP7_75t_L g5955 ( 
.A1(n_4667),
.A2(n_5260),
.B(n_5074),
.C(n_5080),
.Y(n_5955)
);

O2A1O1Ixp33_ASAP7_75t_SL g5956 ( 
.A1(n_5040),
.A2(n_3986),
.B(n_4052),
.C(n_4021),
.Y(n_5956)
);

NAND2x1_ASAP7_75t_L g5957 ( 
.A(n_5597),
.B(n_3976),
.Y(n_5957)
);

NAND2xp5_ASAP7_75t_L g5958 ( 
.A(n_4686),
.B(n_3976),
.Y(n_5958)
);

AND2x2_ASAP7_75t_L g5959 ( 
.A(n_4680),
.B(n_3885),
.Y(n_5959)
);

AND2x4_ASAP7_75t_L g5960 ( 
.A(n_4832),
.B(n_4190),
.Y(n_5960)
);

NOR2xp33_ASAP7_75t_L g5961 ( 
.A(n_5149),
.B(n_4124),
.Y(n_5961)
);

INVxp67_ASAP7_75t_L g5962 ( 
.A(n_5746),
.Y(n_5962)
);

O2A1O1Ixp5_ASAP7_75t_SL g5963 ( 
.A1(n_5039),
.A2(n_3885),
.B(n_4021),
.C(n_4428),
.Y(n_5963)
);

INVx4_ASAP7_75t_L g5964 ( 
.A(n_5233),
.Y(n_5964)
);

BUFx6f_ASAP7_75t_L g5965 ( 
.A(n_4658),
.Y(n_5965)
);

AOI21xp5_ASAP7_75t_L g5966 ( 
.A1(n_5650),
.A2(n_4124),
.B(n_3760),
.Y(n_5966)
);

NAND2xp5_ASAP7_75t_SL g5967 ( 
.A(n_5332),
.B(n_3760),
.Y(n_5967)
);

OA21x2_ASAP7_75t_L g5968 ( 
.A1(n_5010),
.A2(n_3740),
.B(n_3762),
.Y(n_5968)
);

INVx1_ASAP7_75t_SL g5969 ( 
.A(n_5442),
.Y(n_5969)
);

NAND2xp5_ASAP7_75t_L g5970 ( 
.A(n_4686),
.B(n_4124),
.Y(n_5970)
);

INVx1_ASAP7_75t_SL g5971 ( 
.A(n_5442),
.Y(n_5971)
);

INVx3_ASAP7_75t_L g5972 ( 
.A(n_4713),
.Y(n_5972)
);

BUFx12f_ASAP7_75t_L g5973 ( 
.A(n_4633),
.Y(n_5973)
);

OAI21x1_ASAP7_75t_SL g5974 ( 
.A1(n_5590),
.A2(n_3728),
.B(n_4859),
.Y(n_5974)
);

NOR3xp33_ASAP7_75t_L g5975 ( 
.A(n_5138),
.B(n_4667),
.C(n_4847),
.Y(n_5975)
);

OR2x2_ASAP7_75t_L g5976 ( 
.A(n_5359),
.B(n_5408),
.Y(n_5976)
);

NOR2xp33_ASAP7_75t_L g5977 ( 
.A(n_5149),
.B(n_5451),
.Y(n_5977)
);

INVx6_ASAP7_75t_L g5978 ( 
.A(n_4674),
.Y(n_5978)
);

BUFx2_ASAP7_75t_L g5979 ( 
.A(n_4979),
.Y(n_5979)
);

AND2x4_ASAP7_75t_L g5980 ( 
.A(n_4832),
.B(n_4734),
.Y(n_5980)
);

AOI222xp33_ASAP7_75t_L g5981 ( 
.A1(n_4618),
.A2(n_5368),
.B1(n_5514),
.B2(n_4986),
.C1(n_5203),
.C2(n_5151),
.Y(n_5981)
);

A2O1A1Ixp33_ASAP7_75t_SL g5982 ( 
.A1(n_4599),
.A2(n_5746),
.B(n_5138),
.C(n_5218),
.Y(n_5982)
);

NAND2xp5_ASAP7_75t_L g5983 ( 
.A(n_4687),
.B(n_4693),
.Y(n_5983)
);

NAND2xp5_ASAP7_75t_SL g5984 ( 
.A(n_5218),
.B(n_4857),
.Y(n_5984)
);

NOR2xp33_ASAP7_75t_L g5985 ( 
.A(n_5451),
.B(n_5370),
.Y(n_5985)
);

OR2x2_ASAP7_75t_L g5986 ( 
.A(n_5359),
.B(n_5408),
.Y(n_5986)
);

A2O1A1Ixp33_ASAP7_75t_L g5987 ( 
.A1(n_5051),
.A2(n_4782),
.B(n_4767),
.C(n_4675),
.Y(n_5987)
);

AOI22xp5_ASAP7_75t_L g5988 ( 
.A1(n_5514),
.A2(n_4727),
.B1(n_5170),
.B2(n_4669),
.Y(n_5988)
);

HB1xp67_ASAP7_75t_L g5989 ( 
.A(n_4575),
.Y(n_5989)
);

O2A1O1Ixp33_ASAP7_75t_L g5990 ( 
.A1(n_4901),
.A2(n_4627),
.B(n_4847),
.C(n_5333),
.Y(n_5990)
);

NAND2xp5_ASAP7_75t_L g5991 ( 
.A(n_4687),
.B(n_4693),
.Y(n_5991)
);

NAND2xp5_ASAP7_75t_L g5992 ( 
.A(n_4697),
.B(n_4698),
.Y(n_5992)
);

NAND2x1p5_ASAP7_75t_L g5993 ( 
.A(n_4719),
.B(n_4739),
.Y(n_5993)
);

INVx4_ASAP7_75t_L g5994 ( 
.A(n_5233),
.Y(n_5994)
);

NAND2x1p5_ASAP7_75t_L g5995 ( 
.A(n_4719),
.B(n_4739),
.Y(n_5995)
);

INVx2_ASAP7_75t_SL g5996 ( 
.A(n_4920),
.Y(n_5996)
);

A2O1A1Ixp33_ASAP7_75t_SL g5997 ( 
.A1(n_5192),
.A2(n_5088),
.B(n_4812),
.C(n_4843),
.Y(n_5997)
);

AOI21xp5_ASAP7_75t_L g5998 ( 
.A1(n_5415),
.A2(n_5525),
.B(n_5591),
.Y(n_5998)
);

O2A1O1Ixp33_ASAP7_75t_L g5999 ( 
.A1(n_4901),
.A2(n_4627),
.B(n_5334),
.C(n_5333),
.Y(n_5999)
);

AOI21xp5_ASAP7_75t_L g6000 ( 
.A1(n_5415),
.A2(n_5525),
.B(n_5591),
.Y(n_6000)
);

AOI22xp33_ASAP7_75t_L g6001 ( 
.A1(n_4753),
.A2(n_4752),
.B1(n_4669),
.B2(n_4605),
.Y(n_6001)
);

OAI22xp5_ASAP7_75t_L g6002 ( 
.A1(n_5368),
.A2(n_4665),
.B1(n_5203),
.B2(n_5151),
.Y(n_6002)
);

CKINVDCx8_ASAP7_75t_R g6003 ( 
.A(n_4660),
.Y(n_6003)
);

NOR2xp33_ASAP7_75t_L g6004 ( 
.A(n_5370),
.B(n_5073),
.Y(n_6004)
);

INVx1_ASAP7_75t_SL g6005 ( 
.A(n_5546),
.Y(n_6005)
);

NAND2xp5_ASAP7_75t_SL g6006 ( 
.A(n_4782),
.B(n_4727),
.Y(n_6006)
);

NAND2xp5_ASAP7_75t_L g6007 ( 
.A(n_4697),
.B(n_4698),
.Y(n_6007)
);

OR2x2_ASAP7_75t_L g6008 ( 
.A(n_5408),
.B(n_4590),
.Y(n_6008)
);

INVxp67_ASAP7_75t_L g6009 ( 
.A(n_5539),
.Y(n_6009)
);

NAND2xp5_ASAP7_75t_SL g6010 ( 
.A(n_5077),
.B(n_5334),
.Y(n_6010)
);

BUFx4_ASAP7_75t_SL g6011 ( 
.A(n_4864),
.Y(n_6011)
);

INVx2_ASAP7_75t_SL g6012 ( 
.A(n_4920),
.Y(n_6012)
);

INVx1_ASAP7_75t_SL g6013 ( 
.A(n_5546),
.Y(n_6013)
);

INVx1_ASAP7_75t_SL g6014 ( 
.A(n_5680),
.Y(n_6014)
);

NAND2xp5_ASAP7_75t_L g6015 ( 
.A(n_4708),
.B(n_4710),
.Y(n_6015)
);

INVx3_ASAP7_75t_L g6016 ( 
.A(n_4791),
.Y(n_6016)
);

O2A1O1Ixp5_ASAP7_75t_SL g6017 ( 
.A1(n_5074),
.A2(n_5119),
.B(n_5128),
.C(n_5080),
.Y(n_6017)
);

INVxp67_ASAP7_75t_L g6018 ( 
.A(n_5539),
.Y(n_6018)
);

BUFx4f_ASAP7_75t_L g6019 ( 
.A(n_4732),
.Y(n_6019)
);

NOR2xp33_ASAP7_75t_L g6020 ( 
.A(n_5073),
.B(n_5228),
.Y(n_6020)
);

AOI21xp5_ASAP7_75t_L g6021 ( 
.A1(n_5621),
.A2(n_5647),
.B(n_5633),
.Y(n_6021)
);

NAND2xp5_ASAP7_75t_L g6022 ( 
.A(n_4708),
.B(n_4710),
.Y(n_6022)
);

NOR2xp67_ASAP7_75t_SL g6023 ( 
.A(n_4563),
.B(n_4630),
.Y(n_6023)
);

A2O1A1Ixp33_ASAP7_75t_L g6024 ( 
.A1(n_5051),
.A2(n_4615),
.B(n_4939),
.C(n_4925),
.Y(n_6024)
);

AOI21xp5_ASAP7_75t_L g6025 ( 
.A1(n_5621),
.A2(n_5647),
.B(n_5633),
.Y(n_6025)
);

BUFx2_ASAP7_75t_L g6026 ( 
.A(n_4996),
.Y(n_6026)
);

AOI21xp5_ASAP7_75t_L g6027 ( 
.A1(n_5655),
.A2(n_5656),
.B(n_5210),
.Y(n_6027)
);

INVx5_ASAP7_75t_L g6028 ( 
.A(n_4946),
.Y(n_6028)
);

BUFx12f_ASAP7_75t_L g6029 ( 
.A(n_4885),
.Y(n_6029)
);

AND2x6_ASAP7_75t_L g6030 ( 
.A(n_4695),
.B(n_4696),
.Y(n_6030)
);

OAI22xp5_ASAP7_75t_L g6031 ( 
.A1(n_4665),
.A2(n_4634),
.B1(n_4648),
.B2(n_4632),
.Y(n_6031)
);

NAND2x1p5_ASAP7_75t_L g6032 ( 
.A(n_4719),
.B(n_4739),
.Y(n_6032)
);

A2O1A1Ixp33_ASAP7_75t_SL g6033 ( 
.A1(n_5192),
.A2(n_5088),
.B(n_4812),
.C(n_4843),
.Y(n_6033)
);

CKINVDCx5p33_ASAP7_75t_R g6034 ( 
.A(n_4681),
.Y(n_6034)
);

A2O1A1Ixp33_ASAP7_75t_L g6035 ( 
.A1(n_4615),
.A2(n_4939),
.B(n_4925),
.C(n_5129),
.Y(n_6035)
);

INVx5_ASAP7_75t_L g6036 ( 
.A(n_4946),
.Y(n_6036)
);

CKINVDCx5p33_ASAP7_75t_R g6037 ( 
.A(n_4681),
.Y(n_6037)
);

BUFx2_ASAP7_75t_L g6038 ( 
.A(n_4996),
.Y(n_6038)
);

BUFx12f_ASAP7_75t_L g6039 ( 
.A(n_4885),
.Y(n_6039)
);

O2A1O1Ixp33_ASAP7_75t_L g6040 ( 
.A1(n_4783),
.A2(n_4753),
.B(n_4752),
.C(n_4611),
.Y(n_6040)
);

OAI22xp5_ASAP7_75t_L g6041 ( 
.A1(n_4632),
.A2(n_4648),
.B1(n_4652),
.B2(n_4634),
.Y(n_6041)
);

NOR2xp33_ASAP7_75t_L g6042 ( 
.A(n_5228),
.B(n_5373),
.Y(n_6042)
);

INVx5_ASAP7_75t_L g6043 ( 
.A(n_4946),
.Y(n_6043)
);

NOR2xp33_ASAP7_75t_L g6044 ( 
.A(n_5373),
.B(n_5072),
.Y(n_6044)
);

INVxp67_ASAP7_75t_L g6045 ( 
.A(n_5560),
.Y(n_6045)
);

O2A1O1Ixp33_ASAP7_75t_L g6046 ( 
.A1(n_4783),
.A2(n_4611),
.B(n_4992),
.C(n_4986),
.Y(n_6046)
);

AND2x4_ASAP7_75t_L g6047 ( 
.A(n_4734),
.B(n_4746),
.Y(n_6047)
);

OAI21xp33_ASAP7_75t_L g6048 ( 
.A1(n_4891),
.A2(n_4928),
.B(n_5170),
.Y(n_6048)
);

OR2x2_ASAP7_75t_L g6049 ( 
.A(n_4590),
.B(n_4597),
.Y(n_6049)
);

INVx5_ASAP7_75t_L g6050 ( 
.A(n_4946),
.Y(n_6050)
);

NAND2xp5_ASAP7_75t_L g6051 ( 
.A(n_4711),
.B(n_4723),
.Y(n_6051)
);

AND2x4_ASAP7_75t_L g6052 ( 
.A(n_4734),
.B(n_4746),
.Y(n_6052)
);

BUFx2_ASAP7_75t_L g6053 ( 
.A(n_4996),
.Y(n_6053)
);

A2O1A1Ixp33_ASAP7_75t_SL g6054 ( 
.A1(n_4808),
.A2(n_4855),
.B(n_4870),
.C(n_4862),
.Y(n_6054)
);

AOI22xp5_ASAP7_75t_L g6055 ( 
.A1(n_4605),
.A2(n_4652),
.B1(n_4910),
.B2(n_4951),
.Y(n_6055)
);

O2A1O1Ixp33_ASAP7_75t_L g6056 ( 
.A1(n_4992),
.A2(n_5129),
.B(n_5329),
.C(n_5326),
.Y(n_6056)
);

O2A1O1Ixp5_ASAP7_75t_SL g6057 ( 
.A1(n_5119),
.A2(n_5132),
.B(n_5143),
.C(n_5128),
.Y(n_6057)
);

AOI21xp5_ASAP7_75t_L g6058 ( 
.A1(n_5655),
.A2(n_5656),
.B(n_5210),
.Y(n_6058)
);

INVx1_ASAP7_75t_SL g6059 ( 
.A(n_5680),
.Y(n_6059)
);

OAI21x1_ASAP7_75t_L g6060 ( 
.A1(n_4585),
.A2(n_5137),
.B(n_5648),
.Y(n_6060)
);

NOR2xp33_ASAP7_75t_L g6061 ( 
.A(n_5072),
.B(n_5114),
.Y(n_6061)
);

AND2x4_ASAP7_75t_L g6062 ( 
.A(n_4746),
.B(n_4759),
.Y(n_6062)
);

CKINVDCx6p67_ASAP7_75t_R g6063 ( 
.A(n_4563),
.Y(n_6063)
);

NAND2xp5_ASAP7_75t_L g6064 ( 
.A(n_4711),
.B(n_4723),
.Y(n_6064)
);

BUFx2_ASAP7_75t_L g6065 ( 
.A(n_4996),
.Y(n_6065)
);

O2A1O1Ixp33_ASAP7_75t_L g6066 ( 
.A1(n_5326),
.A2(n_5338),
.B(n_5339),
.C(n_5329),
.Y(n_6066)
);

NAND2xp5_ASAP7_75t_L g6067 ( 
.A(n_4725),
.B(n_4744),
.Y(n_6067)
);

AOI22xp5_ASAP7_75t_L g6068 ( 
.A1(n_4910),
.A2(n_4951),
.B1(n_5402),
.B2(n_5206),
.Y(n_6068)
);

A2O1A1Ixp33_ASAP7_75t_L g6069 ( 
.A1(n_5206),
.A2(n_5246),
.B(n_4947),
.C(n_4960),
.Y(n_6069)
);

OAI22xp5_ASAP7_75t_SL g6070 ( 
.A1(n_5402),
.A2(n_4793),
.B1(n_4842),
.B2(n_4815),
.Y(n_6070)
);

OAI22xp5_ASAP7_75t_L g6071 ( 
.A1(n_4793),
.A2(n_4815),
.B1(n_4853),
.B2(n_4842),
.Y(n_6071)
);

NAND2xp5_ASAP7_75t_L g6072 ( 
.A(n_4725),
.B(n_4744),
.Y(n_6072)
);

NOR2xp67_ASAP7_75t_L g6073 ( 
.A(n_4784),
.B(n_5583),
.Y(n_6073)
);

INVx4_ASAP7_75t_L g6074 ( 
.A(n_5233),
.Y(n_6074)
);

OAI22xp5_ASAP7_75t_L g6075 ( 
.A1(n_4853),
.A2(n_4879),
.B1(n_5071),
.B2(n_4878),
.Y(n_6075)
);

AND2x4_ASAP7_75t_L g6076 ( 
.A(n_4746),
.B(n_4759),
.Y(n_6076)
);

NOR2xp33_ASAP7_75t_L g6077 ( 
.A(n_5114),
.B(n_5387),
.Y(n_6077)
);

O2A1O1Ixp33_ASAP7_75t_L g6078 ( 
.A1(n_5338),
.A2(n_5358),
.B(n_5362),
.C(n_5339),
.Y(n_6078)
);

NOR2x1_ASAP7_75t_L g6079 ( 
.A(n_5394),
.B(n_4784),
.Y(n_6079)
);

BUFx12f_ASAP7_75t_L g6080 ( 
.A(n_5307),
.Y(n_6080)
);

AOI222xp33_ASAP7_75t_L g6081 ( 
.A1(n_5472),
.A2(n_5511),
.B1(n_5222),
.B2(n_4928),
.C1(n_4891),
.C2(n_4836),
.Y(n_6081)
);

INVx3_ASAP7_75t_SL g6082 ( 
.A(n_5536),
.Y(n_6082)
);

AND2x4_ASAP7_75t_L g6083 ( 
.A(n_4746),
.B(n_4759),
.Y(n_6083)
);

INVxp67_ASAP7_75t_SL g6084 ( 
.A(n_4553),
.Y(n_6084)
);

CKINVDCx5p33_ASAP7_75t_R g6085 ( 
.A(n_4702),
.Y(n_6085)
);

BUFx2_ASAP7_75t_L g6086 ( 
.A(n_4996),
.Y(n_6086)
);

BUFx12f_ASAP7_75t_L g6087 ( 
.A(n_5307),
.Y(n_6087)
);

AOI21xp5_ASAP7_75t_L g6088 ( 
.A1(n_5197),
.A2(n_5211),
.B(n_5548),
.Y(n_6088)
);

INVx5_ASAP7_75t_L g6089 ( 
.A(n_4946),
.Y(n_6089)
);

AOI222xp33_ASAP7_75t_L g6090 ( 
.A1(n_5472),
.A2(n_5511),
.B1(n_5222),
.B2(n_4836),
.C1(n_4609),
.C2(n_4602),
.Y(n_6090)
);

OAI22xp5_ASAP7_75t_L g6091 ( 
.A1(n_4878),
.A2(n_4879),
.B1(n_5141),
.B2(n_5071),
.Y(n_6091)
);

AOI22xp5_ASAP7_75t_L g6092 ( 
.A1(n_5387),
.A2(n_5184),
.B1(n_5141),
.B2(n_4808),
.Y(n_6092)
);

NAND2xp5_ASAP7_75t_L g6093 ( 
.A(n_4756),
.B(n_4761),
.Y(n_6093)
);

NOR2xp33_ASAP7_75t_L g6094 ( 
.A(n_5590),
.B(n_5033),
.Y(n_6094)
);

NAND2xp5_ASAP7_75t_L g6095 ( 
.A(n_4756),
.B(n_4761),
.Y(n_6095)
);

INVx3_ASAP7_75t_L g6096 ( 
.A(n_4798),
.Y(n_6096)
);

O2A1O1Ixp33_ASAP7_75t_L g6097 ( 
.A1(n_5358),
.A2(n_5362),
.B(n_5378),
.C(n_5246),
.Y(n_6097)
);

AOI21x1_ASAP7_75t_L g6098 ( 
.A1(n_4831),
.A2(n_4743),
.B(n_5308),
.Y(n_6098)
);

NAND2xp5_ASAP7_75t_SL g6099 ( 
.A(n_5077),
.B(n_5322),
.Y(n_6099)
);

A2O1A1Ixp33_ASAP7_75t_L g6100 ( 
.A1(n_4947),
.A2(n_4956),
.B(n_5131),
.C(n_4960),
.Y(n_6100)
);

AOI21xp5_ASAP7_75t_L g6101 ( 
.A1(n_5197),
.A2(n_5211),
.B(n_5548),
.Y(n_6101)
);

OAI21x1_ASAP7_75t_L g6102 ( 
.A1(n_4585),
.A2(n_5137),
.B(n_5648),
.Y(n_6102)
);

NAND2xp5_ASAP7_75t_SL g6103 ( 
.A(n_5322),
.B(n_5337),
.Y(n_6103)
);

OAI22x1_ASAP7_75t_L g6104 ( 
.A1(n_5132),
.A2(n_5157),
.B1(n_5180),
.B2(n_5143),
.Y(n_6104)
);

OAI22xp5_ASAP7_75t_L g6105 ( 
.A1(n_5184),
.A2(n_4944),
.B1(n_5136),
.B2(n_5263),
.Y(n_6105)
);

INVx3_ASAP7_75t_L g6106 ( 
.A(n_4798),
.Y(n_6106)
);

AOI21xp5_ASAP7_75t_L g6107 ( 
.A1(n_5389),
.A2(n_5410),
.B(n_4703),
.Y(n_6107)
);

AND2x4_ASAP7_75t_L g6108 ( 
.A(n_4759),
.B(n_4760),
.Y(n_6108)
);

BUFx8_ASAP7_75t_L g6109 ( 
.A(n_5193),
.Y(n_6109)
);

O2A1O1Ixp33_ASAP7_75t_L g6110 ( 
.A1(n_5378),
.A2(n_5282),
.B(n_5385),
.C(n_5380),
.Y(n_6110)
);

BUFx2_ASAP7_75t_SL g6111 ( 
.A(n_5689),
.Y(n_6111)
);

BUFx8_ASAP7_75t_SL g6112 ( 
.A(n_4860),
.Y(n_6112)
);

AOI21x1_ASAP7_75t_L g6113 ( 
.A1(n_4831),
.A2(n_4743),
.B(n_5308),
.Y(n_6113)
);

INVx4_ASAP7_75t_L g6114 ( 
.A(n_5233),
.Y(n_6114)
);

OAI22xp5_ASAP7_75t_L g6115 ( 
.A1(n_4944),
.A2(n_5136),
.B1(n_5263),
.B2(n_5355),
.Y(n_6115)
);

NAND2xp5_ASAP7_75t_L g6116 ( 
.A(n_4769),
.B(n_4771),
.Y(n_6116)
);

A2O1A1Ixp33_ASAP7_75t_L g6117 ( 
.A1(n_4956),
.A2(n_5189),
.B(n_5217),
.C(n_5131),
.Y(n_6117)
);

INVx4_ASAP7_75t_L g6118 ( 
.A(n_5233),
.Y(n_6118)
);

INVx2_ASAP7_75t_SL g6119 ( 
.A(n_4920),
.Y(n_6119)
);

NOR2xp33_ASAP7_75t_L g6120 ( 
.A(n_5033),
.B(n_5506),
.Y(n_6120)
);

INVx4_ASAP7_75t_L g6121 ( 
.A(n_5233),
.Y(n_6121)
);

NAND2xp33_ASAP7_75t_L g6122 ( 
.A(n_5076),
.B(n_5495),
.Y(n_6122)
);

INVx4_ASAP7_75t_L g6123 ( 
.A(n_5233),
.Y(n_6123)
);

BUFx2_ASAP7_75t_SL g6124 ( 
.A(n_5689),
.Y(n_6124)
);

AOI21x1_ASAP7_75t_L g6125 ( 
.A1(n_5629),
.A2(n_5526),
.B(n_5536),
.Y(n_6125)
);

BUFx6f_ASAP7_75t_SL g6126 ( 
.A(n_5632),
.Y(n_6126)
);

NAND2xp5_ASAP7_75t_L g6127 ( 
.A(n_4769),
.B(n_4771),
.Y(n_6127)
);

AND2x2_ASAP7_75t_L g6128 ( 
.A(n_4700),
.B(n_4715),
.Y(n_6128)
);

OR2x6_ASAP7_75t_SL g6129 ( 
.A(n_4801),
.B(n_5262),
.Y(n_6129)
);

AOI21xp5_ASAP7_75t_L g6130 ( 
.A1(n_5389),
.A2(n_5410),
.B(n_4703),
.Y(n_6130)
);

OAI22xp33_ASAP7_75t_L g6131 ( 
.A1(n_4602),
.A2(n_5555),
.B1(n_4598),
.B2(n_4600),
.Y(n_6131)
);

NOR2xp67_ASAP7_75t_L g6132 ( 
.A(n_5583),
.B(n_5198),
.Y(n_6132)
);

BUFx2_ASAP7_75t_L g6133 ( 
.A(n_5026),
.Y(n_6133)
);

AND2x4_ASAP7_75t_L g6134 ( 
.A(n_4759),
.B(n_4760),
.Y(n_6134)
);

NOR2xp67_ASAP7_75t_L g6135 ( 
.A(n_5583),
.B(n_5198),
.Y(n_6135)
);

NAND2xp5_ASAP7_75t_L g6136 ( 
.A(n_4772),
.B(n_4775),
.Y(n_6136)
);

INVxp67_ASAP7_75t_SL g6137 ( 
.A(n_4559),
.Y(n_6137)
);

AOI22xp33_ASAP7_75t_L g6138 ( 
.A1(n_4598),
.A2(n_4600),
.B1(n_4862),
.B2(n_4855),
.Y(n_6138)
);

NAND2xp5_ASAP7_75t_L g6139 ( 
.A(n_4772),
.B(n_4775),
.Y(n_6139)
);

INVx4_ASAP7_75t_L g6140 ( 
.A(n_5233),
.Y(n_6140)
);

BUFx2_ASAP7_75t_L g6141 ( 
.A(n_5026),
.Y(n_6141)
);

OR2x2_ASAP7_75t_L g6142 ( 
.A(n_4597),
.B(n_4635),
.Y(n_6142)
);

O2A1O1Ixp33_ASAP7_75t_L g6143 ( 
.A1(n_5282),
.A2(n_5385),
.B(n_5380),
.C(n_5315),
.Y(n_6143)
);

NOR2xp33_ASAP7_75t_R g6144 ( 
.A(n_5349),
.B(n_5379),
.Y(n_6144)
);

NAND2xp5_ASAP7_75t_L g6145 ( 
.A(n_4776),
.B(n_4786),
.Y(n_6145)
);

AOI21xp5_ASAP7_75t_L g6146 ( 
.A1(n_4612),
.A2(n_4726),
.B(n_4703),
.Y(n_6146)
);

CKINVDCx6p67_ASAP7_75t_R g6147 ( 
.A(n_4563),
.Y(n_6147)
);

NOR2xp67_ASAP7_75t_L g6148 ( 
.A(n_5198),
.B(n_5225),
.Y(n_6148)
);

BUFx2_ASAP7_75t_L g6149 ( 
.A(n_5026),
.Y(n_6149)
);

BUFx2_ASAP7_75t_L g6150 ( 
.A(n_5026),
.Y(n_6150)
);

NAND2xp5_ASAP7_75t_L g6151 ( 
.A(n_4776),
.B(n_4786),
.Y(n_6151)
);

OAI22xp5_ASAP7_75t_L g6152 ( 
.A1(n_5355),
.A2(n_4844),
.B1(n_5527),
.B2(n_5337),
.Y(n_6152)
);

AND2x4_ASAP7_75t_L g6153 ( 
.A(n_4760),
.B(n_4640),
.Y(n_6153)
);

AOI21xp5_ASAP7_75t_L g6154 ( 
.A1(n_4612),
.A2(n_4726),
.B(n_4703),
.Y(n_6154)
);

INVx5_ASAP7_75t_L g6155 ( 
.A(n_4946),
.Y(n_6155)
);

NOR2xp33_ASAP7_75t_L g6156 ( 
.A(n_5506),
.B(n_4609),
.Y(n_6156)
);

AOI21xp5_ASAP7_75t_L g6157 ( 
.A1(n_4612),
.A2(n_4726),
.B(n_4703),
.Y(n_6157)
);

AOI22xp33_ASAP7_75t_L g6158 ( 
.A1(n_4870),
.A2(n_4872),
.B1(n_5346),
.B2(n_5549),
.Y(n_6158)
);

BUFx12f_ASAP7_75t_L g6159 ( 
.A(n_5349),
.Y(n_6159)
);

INVx1_ASAP7_75t_L g6160 ( 
.A(n_5405),
.Y(n_6160)
);

OAI22xp5_ASAP7_75t_L g6161 ( 
.A1(n_5355),
.A2(n_4844),
.B1(n_5527),
.B2(n_5044),
.Y(n_6161)
);

NOR2xp33_ASAP7_75t_R g6162 ( 
.A(n_5379),
.B(n_5425),
.Y(n_6162)
);

AOI21xp5_ASAP7_75t_L g6163 ( 
.A1(n_4612),
.A2(n_4726),
.B(n_4703),
.Y(n_6163)
);

INVxp67_ASAP7_75t_L g6164 ( 
.A(n_5560),
.Y(n_6164)
);

INVxp67_ASAP7_75t_L g6165 ( 
.A(n_5364),
.Y(n_6165)
);

INVx1_ASAP7_75t_L g6166 ( 
.A(n_5405),
.Y(n_6166)
);

AND2x4_ASAP7_75t_L g6167 ( 
.A(n_4760),
.B(n_4640),
.Y(n_6167)
);

INVx1_ASAP7_75t_L g6168 ( 
.A(n_5405),
.Y(n_6168)
);

O2A1O1Ixp5_ASAP7_75t_SL g6169 ( 
.A1(n_5157),
.A2(n_5199),
.B(n_5213),
.C(n_5180),
.Y(n_6169)
);

AND2x4_ASAP7_75t_L g6170 ( 
.A(n_4760),
.B(n_4640),
.Y(n_6170)
);

INVx4_ASAP7_75t_L g6171 ( 
.A(n_4696),
.Y(n_6171)
);

NAND2xp5_ASAP7_75t_L g6172 ( 
.A(n_4794),
.B(n_4799),
.Y(n_6172)
);

INVx1_ASAP7_75t_L g6173 ( 
.A(n_5405),
.Y(n_6173)
);

AOI22xp33_ASAP7_75t_SL g6174 ( 
.A1(n_5346),
.A2(n_5081),
.B1(n_5215),
.B2(n_4801),
.Y(n_6174)
);

INVx1_ASAP7_75t_L g6175 ( 
.A(n_5421),
.Y(n_6175)
);

BUFx8_ASAP7_75t_SL g6176 ( 
.A(n_4860),
.Y(n_6176)
);

A2O1A1Ixp33_ASAP7_75t_L g6177 ( 
.A1(n_5189),
.A2(n_5257),
.B(n_5217),
.C(n_5213),
.Y(n_6177)
);

O2A1O1Ixp33_ASAP7_75t_L g6178 ( 
.A1(n_5315),
.A2(n_5420),
.B(n_4593),
.C(n_5224),
.Y(n_6178)
);

INVx1_ASAP7_75t_L g6179 ( 
.A(n_5421),
.Y(n_6179)
);

OR2x2_ASAP7_75t_L g6180 ( 
.A(n_4635),
.B(n_4821),
.Y(n_6180)
);

O2A1O1Ixp33_ASAP7_75t_L g6181 ( 
.A1(n_5420),
.A2(n_4593),
.B(n_5224),
.C(n_5199),
.Y(n_6181)
);

A2O1A1Ixp33_ASAP7_75t_L g6182 ( 
.A1(n_5257),
.A2(n_5407),
.B(n_4801),
.C(n_4872),
.Y(n_6182)
);

NAND2x2_ASAP7_75t_L g6183 ( 
.A(n_4779),
.B(n_4655),
.Y(n_6183)
);

AO32x1_ASAP7_75t_L g6184 ( 
.A1(n_4700),
.A2(n_4715),
.A3(n_4749),
.B1(n_4742),
.B2(n_4740),
.Y(n_6184)
);

AOI22xp5_ASAP7_75t_SL g6185 ( 
.A1(n_4801),
.A2(n_5350),
.B1(n_5473),
.B2(n_5236),
.Y(n_6185)
);

CKINVDCx5p33_ASAP7_75t_R g6186 ( 
.A(n_4702),
.Y(n_6186)
);

INVx1_ASAP7_75t_L g6187 ( 
.A(n_5421),
.Y(n_6187)
);

OR2x6_ASAP7_75t_L g6188 ( 
.A(n_4822),
.B(n_4601),
.Y(n_6188)
);

NAND2xp5_ASAP7_75t_L g6189 ( 
.A(n_4794),
.B(n_4799),
.Y(n_6189)
);

CKINVDCx5p33_ASAP7_75t_R g6190 ( 
.A(n_4750),
.Y(n_6190)
);

NOR2xp33_ASAP7_75t_L g6191 ( 
.A(n_5407),
.B(n_5108),
.Y(n_6191)
);

NAND2xp5_ASAP7_75t_L g6192 ( 
.A(n_4802),
.B(n_4805),
.Y(n_6192)
);

INVx1_ASAP7_75t_L g6193 ( 
.A(n_5421),
.Y(n_6193)
);

NAND2xp5_ASAP7_75t_L g6194 ( 
.A(n_4802),
.B(n_4805),
.Y(n_6194)
);

A2O1A1Ixp33_ASAP7_75t_L g6195 ( 
.A1(n_4801),
.A2(n_4875),
.B(n_5559),
.C(n_4704),
.Y(n_6195)
);

AOI22xp33_ASAP7_75t_SL g6196 ( 
.A1(n_5346),
.A2(n_5081),
.B1(n_5215),
.B2(n_5236),
.Y(n_6196)
);

AOI21xp5_ASAP7_75t_L g6197 ( 
.A1(n_4612),
.A2(n_4726),
.B(n_4703),
.Y(n_6197)
);

AOI21xp5_ASAP7_75t_L g6198 ( 
.A1(n_4612),
.A2(n_4868),
.B(n_4726),
.Y(n_6198)
);

AOI22x1_ASAP7_75t_L g6199 ( 
.A1(n_4704),
.A2(n_4803),
.B1(n_4824),
.B2(n_4768),
.Y(n_6199)
);

O2A1O1Ixp5_ASAP7_75t_SL g6200 ( 
.A1(n_5516),
.A2(n_5577),
.B(n_5466),
.C(n_5708),
.Y(n_6200)
);

HB1xp67_ASAP7_75t_L g6201 ( 
.A(n_4554),
.Y(n_6201)
);

NAND2xp5_ASAP7_75t_L g6202 ( 
.A(n_4807),
.B(n_4809),
.Y(n_6202)
);

OAI222xp33_ASAP7_75t_L g6203 ( 
.A1(n_4762),
.A2(n_4796),
.B1(n_4810),
.B2(n_4787),
.C1(n_4589),
.C2(n_5555),
.Y(n_6203)
);

AOI21x1_ASAP7_75t_L g6204 ( 
.A1(n_5629),
.A2(n_5526),
.B(n_5516),
.Y(n_6204)
);

NOR2xp67_ASAP7_75t_L g6205 ( 
.A(n_5198),
.B(n_5225),
.Y(n_6205)
);

BUFx2_ASAP7_75t_L g6206 ( 
.A(n_5026),
.Y(n_6206)
);

NAND2xp5_ASAP7_75t_L g6207 ( 
.A(n_4807),
.B(n_4809),
.Y(n_6207)
);

NOR2xp33_ASAP7_75t_L g6208 ( 
.A(n_5108),
.B(n_4816),
.Y(n_6208)
);

BUFx2_ASAP7_75t_L g6209 ( 
.A(n_4930),
.Y(n_6209)
);

BUFx2_ASAP7_75t_L g6210 ( 
.A(n_4990),
.Y(n_6210)
);

CKINVDCx20_ASAP7_75t_R g6211 ( 
.A(n_4825),
.Y(n_6211)
);

OR2x2_ASAP7_75t_L g6212 ( 
.A(n_4821),
.B(n_4828),
.Y(n_6212)
);

AND2x2_ASAP7_75t_L g6213 ( 
.A(n_4715),
.B(n_4740),
.Y(n_6213)
);

AND2x2_ASAP7_75t_L g6214 ( 
.A(n_4740),
.B(n_4742),
.Y(n_6214)
);

AOI21xp5_ASAP7_75t_L g6215 ( 
.A1(n_4612),
.A2(n_4868),
.B(n_4726),
.Y(n_6215)
);

AOI21xp5_ASAP7_75t_L g6216 ( 
.A1(n_4868),
.A2(n_5000),
.B(n_4969),
.Y(n_6216)
);

AND2x2_ASAP7_75t_L g6217 ( 
.A(n_4742),
.B(n_4749),
.Y(n_6217)
);

INVx1_ASAP7_75t_L g6218 ( 
.A(n_5429),
.Y(n_6218)
);

INVx1_ASAP7_75t_L g6219 ( 
.A(n_5429),
.Y(n_6219)
);

INVx1_ASAP7_75t_L g6220 ( 
.A(n_5429),
.Y(n_6220)
);

NAND2xp5_ASAP7_75t_SL g6221 ( 
.A(n_4875),
.B(n_5044),
.Y(n_6221)
);

INVx1_ASAP7_75t_L g6222 ( 
.A(n_5429),
.Y(n_6222)
);

INVx1_ASAP7_75t_L g6223 ( 
.A(n_5435),
.Y(n_6223)
);

NAND2xp5_ASAP7_75t_L g6224 ( 
.A(n_4816),
.B(n_4818),
.Y(n_6224)
);

OAI221xp5_ASAP7_75t_L g6225 ( 
.A1(n_5559),
.A2(n_4796),
.B1(n_4810),
.B2(n_4787),
.C(n_4762),
.Y(n_6225)
);

O2A1O1Ixp5_ASAP7_75t_SL g6226 ( 
.A1(n_5577),
.A2(n_5466),
.B(n_5708),
.C(n_4567),
.Y(n_6226)
);

A2O1A1Ixp33_ASAP7_75t_L g6227 ( 
.A1(n_4768),
.A2(n_4803),
.B(n_4824),
.C(n_5325),
.Y(n_6227)
);

INVx1_ASAP7_75t_SL g6228 ( 
.A(n_5665),
.Y(n_6228)
);

NAND2xp5_ASAP7_75t_SL g6229 ( 
.A(n_4624),
.B(n_5117),
.Y(n_6229)
);

OA21x2_ASAP7_75t_L g6230 ( 
.A1(n_5010),
.A2(n_4751),
.B(n_4585),
.Y(n_6230)
);

NAND2xp5_ASAP7_75t_SL g6231 ( 
.A(n_4624),
.B(n_5117),
.Y(n_6231)
);

INVxp67_ASAP7_75t_L g6232 ( 
.A(n_5364),
.Y(n_6232)
);

AOI22x1_ASAP7_75t_L g6233 ( 
.A1(n_4735),
.A2(n_4660),
.B1(n_4661),
.B2(n_4576),
.Y(n_6233)
);

A2O1A1Ixp33_ASAP7_75t_L g6234 ( 
.A1(n_5325),
.A2(n_5139),
.B(n_5242),
.C(n_5236),
.Y(n_6234)
);

INVx1_ASAP7_75t_L g6235 ( 
.A(n_5435),
.Y(n_6235)
);

BUFx2_ASAP7_75t_L g6236 ( 
.A(n_4828),
.Y(n_6236)
);

AOI21x1_ASAP7_75t_SL g6237 ( 
.A1(n_4735),
.A2(n_4758),
.B(n_4749),
.Y(n_6237)
);

NOR2xp33_ASAP7_75t_SL g6238 ( 
.A(n_5111),
.B(n_4737),
.Y(n_6238)
);

INVx1_ASAP7_75t_L g6239 ( 
.A(n_5435),
.Y(n_6239)
);

NOR2xp33_ASAP7_75t_L g6240 ( 
.A(n_4818),
.B(n_4823),
.Y(n_6240)
);

BUFx8_ASAP7_75t_L g6241 ( 
.A(n_5193),
.Y(n_6241)
);

NAND2xp5_ASAP7_75t_L g6242 ( 
.A(n_4823),
.B(n_4826),
.Y(n_6242)
);

AND2x2_ASAP7_75t_L g6243 ( 
.A(n_4758),
.B(n_4866),
.Y(n_6243)
);

AND2x2_ASAP7_75t_L g6244 ( 
.A(n_4758),
.B(n_4866),
.Y(n_6244)
);

A2O1A1Ixp33_ASAP7_75t_L g6245 ( 
.A1(n_5139),
.A2(n_5236),
.B(n_5242),
.C(n_5190),
.Y(n_6245)
);

HB1xp67_ASAP7_75t_L g6246 ( 
.A(n_4554),
.Y(n_6246)
);

OAI22xp5_ASAP7_75t_L g6247 ( 
.A1(n_4965),
.A2(n_5005),
.B1(n_5027),
.B2(n_4998),
.Y(n_6247)
);

AOI222xp33_ASAP7_75t_L g6248 ( 
.A1(n_5360),
.A2(n_5369),
.B1(n_5027),
.B2(n_4965),
.C1(n_5038),
.C2(n_5005),
.Y(n_6248)
);

INVx5_ASAP7_75t_L g6249 ( 
.A(n_5020),
.Y(n_6249)
);

NAND2xp5_ASAP7_75t_L g6250 ( 
.A(n_4826),
.B(n_4829),
.Y(n_6250)
);

INVx1_ASAP7_75t_L g6251 ( 
.A(n_5435),
.Y(n_6251)
);

AND2x2_ASAP7_75t_L g6252 ( 
.A(n_4866),
.B(n_4877),
.Y(n_6252)
);

INVx1_ASAP7_75t_L g6253 ( 
.A(n_5437),
.Y(n_6253)
);

AOI22xp5_ASAP7_75t_L g6254 ( 
.A1(n_5549),
.A2(n_5551),
.B1(n_5369),
.B2(n_5360),
.Y(n_6254)
);

AOI21x1_ASAP7_75t_L g6255 ( 
.A1(n_5629),
.A2(n_5010),
.B(n_5749),
.Y(n_6255)
);

A2O1A1Ixp33_ASAP7_75t_L g6256 ( 
.A1(n_5236),
.A2(n_5242),
.B(n_5190),
.C(n_5432),
.Y(n_6256)
);

AOI21xp5_ASAP7_75t_L g6257 ( 
.A1(n_4868),
.A2(n_5000),
.B(n_4969),
.Y(n_6257)
);

NOR2xp33_ASAP7_75t_L g6258 ( 
.A(n_4829),
.B(n_4833),
.Y(n_6258)
);

BUFx2_ASAP7_75t_L g6259 ( 
.A(n_4849),
.Y(n_6259)
);

AOI222xp33_ASAP7_75t_L g6260 ( 
.A1(n_4998),
.A2(n_5084),
.B1(n_5038),
.B2(n_5089),
.C1(n_5049),
.C2(n_5041),
.Y(n_6260)
);

NAND2xp5_ASAP7_75t_L g6261 ( 
.A(n_4833),
.B(n_4834),
.Y(n_6261)
);

BUFx2_ASAP7_75t_L g6262 ( 
.A(n_4849),
.Y(n_6262)
);

NAND2xp5_ASAP7_75t_L g6263 ( 
.A(n_4834),
.B(n_4837),
.Y(n_6263)
);

AND2x4_ASAP7_75t_L g6264 ( 
.A(n_4849),
.B(n_4858),
.Y(n_6264)
);

NAND2x1p5_ASAP7_75t_L g6265 ( 
.A(n_4719),
.B(n_4739),
.Y(n_6265)
);

INVx1_ASAP7_75t_SL g6266 ( 
.A(n_5665),
.Y(n_6266)
);

AND2x2_ASAP7_75t_L g6267 ( 
.A(n_4877),
.B(n_4900),
.Y(n_6267)
);

AOI21xp5_ASAP7_75t_L g6268 ( 
.A1(n_4868),
.A2(n_5000),
.B(n_4969),
.Y(n_6268)
);

INVx1_ASAP7_75t_L g6269 ( 
.A(n_5437),
.Y(n_6269)
);

INVxp67_ASAP7_75t_L g6270 ( 
.A(n_5423),
.Y(n_6270)
);

INVx2_ASAP7_75t_SL g6271 ( 
.A(n_4736),
.Y(n_6271)
);

AOI21xp5_ASAP7_75t_L g6272 ( 
.A1(n_4868),
.A2(n_5000),
.B(n_4969),
.Y(n_6272)
);

NAND2xp5_ASAP7_75t_L g6273 ( 
.A(n_4837),
.B(n_4839),
.Y(n_6273)
);

O2A1O1Ixp33_ASAP7_75t_L g6274 ( 
.A1(n_5432),
.A2(n_4643),
.B(n_4637),
.C(n_5226),
.Y(n_6274)
);

INVxp67_ASAP7_75t_L g6275 ( 
.A(n_5423),
.Y(n_6275)
);

INVx2_ASAP7_75t_SL g6276 ( 
.A(n_4736),
.Y(n_6276)
);

INVxp67_ASAP7_75t_L g6277 ( 
.A(n_5493),
.Y(n_6277)
);

INVx4_ASAP7_75t_L g6278 ( 
.A(n_4701),
.Y(n_6278)
);

AOI21xp5_ASAP7_75t_L g6279 ( 
.A1(n_4868),
.A2(n_5000),
.B(n_4969),
.Y(n_6279)
);

INVx1_ASAP7_75t_L g6280 ( 
.A(n_5437),
.Y(n_6280)
);

INVx1_ASAP7_75t_SL g6281 ( 
.A(n_5665),
.Y(n_6281)
);

INVx2_ASAP7_75t_SL g6282 ( 
.A(n_4736),
.Y(n_6282)
);

INVx3_ASAP7_75t_L g6283 ( 
.A(n_4560),
.Y(n_6283)
);

NAND2xp5_ASAP7_75t_L g6284 ( 
.A(n_4839),
.B(n_4840),
.Y(n_6284)
);

INVx2_ASAP7_75t_SL g6285 ( 
.A(n_4736),
.Y(n_6285)
);

NOR2xp33_ASAP7_75t_L g6286 ( 
.A(n_4840),
.B(n_4841),
.Y(n_6286)
);

AOI22xp33_ASAP7_75t_L g6287 ( 
.A1(n_5551),
.A2(n_4643),
.B1(n_4637),
.B2(n_5215),
.Y(n_6287)
);

INVx3_ASAP7_75t_L g6288 ( 
.A(n_4560),
.Y(n_6288)
);

NAND2xp5_ASAP7_75t_L g6289 ( 
.A(n_4841),
.B(n_4845),
.Y(n_6289)
);

INVx4_ASAP7_75t_L g6290 ( 
.A(n_4701),
.Y(n_6290)
);

BUFx2_ASAP7_75t_L g6291 ( 
.A(n_4849),
.Y(n_6291)
);

NOR2xp33_ASAP7_75t_L g6292 ( 
.A(n_4845),
.B(n_4850),
.Y(n_6292)
);

AOI21xp5_ASAP7_75t_L g6293 ( 
.A1(n_4969),
.A2(n_5078),
.B(n_5000),
.Y(n_6293)
);

AOI22xp33_ASAP7_75t_L g6294 ( 
.A1(n_5081),
.A2(n_5215),
.B1(n_5049),
.B2(n_5084),
.Y(n_6294)
);

AOI21xp5_ASAP7_75t_L g6295 ( 
.A1(n_4969),
.A2(n_5078),
.B(n_5000),
.Y(n_6295)
);

AOI21xp5_ASAP7_75t_L g6296 ( 
.A1(n_5078),
.A2(n_5159),
.B(n_5112),
.Y(n_6296)
);

O2A1O1Ixp5_ASAP7_75t_L g6297 ( 
.A1(n_4751),
.A2(n_5350),
.B(n_5202),
.C(n_5571),
.Y(n_6297)
);

INVx1_ASAP7_75t_L g6298 ( 
.A(n_5437),
.Y(n_6298)
);

OR2x6_ASAP7_75t_L g6299 ( 
.A(n_4822),
.B(n_4601),
.Y(n_6299)
);

A2O1A1Ixp33_ASAP7_75t_L g6300 ( 
.A1(n_5236),
.A2(n_5242),
.B(n_5171),
.C(n_5172),
.Y(n_6300)
);

AOI21xp5_ASAP7_75t_L g6301 ( 
.A1(n_5078),
.A2(n_5159),
.B(n_5112),
.Y(n_6301)
);

NAND2xp5_ASAP7_75t_L g6302 ( 
.A(n_4850),
.B(n_4851),
.Y(n_6302)
);

INVx2_ASAP7_75t_SL g6303 ( 
.A(n_4822),
.Y(n_6303)
);

NOR2xp33_ASAP7_75t_L g6304 ( 
.A(n_4851),
.B(n_4861),
.Y(n_6304)
);

INVx1_ASAP7_75t_L g6305 ( 
.A(n_5456),
.Y(n_6305)
);

NAND2xp5_ASAP7_75t_L g6306 ( 
.A(n_4861),
.B(n_4867),
.Y(n_6306)
);

HB1xp67_ASAP7_75t_L g6307 ( 
.A(n_4554),
.Y(n_6307)
);

NAND2xp5_ASAP7_75t_SL g6308 ( 
.A(n_4660),
.B(n_4737),
.Y(n_6308)
);

AOI21xp5_ASAP7_75t_L g6309 ( 
.A1(n_5078),
.A2(n_5159),
.B(n_5112),
.Y(n_6309)
);

INVx4_ASAP7_75t_L g6310 ( 
.A(n_4731),
.Y(n_6310)
);

AND2x4_ASAP7_75t_L g6311 ( 
.A(n_4849),
.B(n_4858),
.Y(n_6311)
);

AND2x4_ASAP7_75t_SL g6312 ( 
.A(n_4731),
.B(n_4733),
.Y(n_6312)
);

INVx1_ASAP7_75t_L g6313 ( 
.A(n_5456),
.Y(n_6313)
);

INVx3_ASAP7_75t_L g6314 ( 
.A(n_4560),
.Y(n_6314)
);

NAND2x2_ASAP7_75t_L g6315 ( 
.A(n_4779),
.B(n_4655),
.Y(n_6315)
);

A2O1A1Ixp33_ASAP7_75t_L g6316 ( 
.A1(n_5242),
.A2(n_5171),
.B(n_5172),
.C(n_5158),
.Y(n_6316)
);

BUFx2_ASAP7_75t_L g6317 ( 
.A(n_4849),
.Y(n_6317)
);

NOR2xp33_ASAP7_75t_L g6318 ( 
.A(n_4867),
.B(n_4871),
.Y(n_6318)
);

AND2x2_ASAP7_75t_L g6319 ( 
.A(n_4877),
.B(n_4900),
.Y(n_6319)
);

AOI21xp33_ASAP7_75t_L g6320 ( 
.A1(n_4780),
.A2(n_4922),
.B(n_4907),
.Y(n_6320)
);

NAND2xp5_ASAP7_75t_L g6321 ( 
.A(n_4871),
.B(n_4880),
.Y(n_6321)
);

INVx1_ASAP7_75t_L g6322 ( 
.A(n_5456),
.Y(n_6322)
);

OAI21x1_ASAP7_75t_SL g6323 ( 
.A1(n_5226),
.A2(n_5733),
.B(n_5545),
.Y(n_6323)
);

BUFx10_ASAP7_75t_L g6324 ( 
.A(n_5193),
.Y(n_6324)
);

INVx1_ASAP7_75t_L g6325 ( 
.A(n_5456),
.Y(n_6325)
);

CKINVDCx20_ASAP7_75t_R g6326 ( 
.A(n_4825),
.Y(n_6326)
);

INVx1_ASAP7_75t_L g6327 ( 
.A(n_5462),
.Y(n_6327)
);

INVxp67_ASAP7_75t_L g6328 ( 
.A(n_5493),
.Y(n_6328)
);

NAND2xp5_ASAP7_75t_L g6329 ( 
.A(n_4880),
.B(n_4883),
.Y(n_6329)
);

OAI22xp5_ASAP7_75t_L g6330 ( 
.A1(n_5041),
.A2(n_5089),
.B1(n_5239),
.B2(n_5200),
.Y(n_6330)
);

INVx1_ASAP7_75t_L g6331 ( 
.A(n_5462),
.Y(n_6331)
);

HB1xp67_ASAP7_75t_L g6332 ( 
.A(n_4554),
.Y(n_6332)
);

INVx5_ASAP7_75t_L g6333 ( 
.A(n_5020),
.Y(n_6333)
);

O2A1O1Ixp5_ASAP7_75t_SL g6334 ( 
.A1(n_5577),
.A2(n_4567),
.B(n_4561),
.C(n_5417),
.Y(n_6334)
);

INVx1_ASAP7_75t_L g6335 ( 
.A(n_5462),
.Y(n_6335)
);

BUFx2_ASAP7_75t_SL g6336 ( 
.A(n_5689),
.Y(n_6336)
);

A2O1A1Ixp33_ASAP7_75t_SL g6337 ( 
.A1(n_5710),
.A2(n_5239),
.B(n_5244),
.C(n_5200),
.Y(n_6337)
);

NAND2xp5_ASAP7_75t_L g6338 ( 
.A(n_4883),
.B(n_4892),
.Y(n_6338)
);

NOR2xp33_ASAP7_75t_L g6339 ( 
.A(n_4892),
.B(n_4898),
.Y(n_6339)
);

NAND2xp5_ASAP7_75t_L g6340 ( 
.A(n_4898),
.B(n_4905),
.Y(n_6340)
);

AOI21xp5_ASAP7_75t_L g6341 ( 
.A1(n_5078),
.A2(n_5159),
.B(n_5112),
.Y(n_6341)
);

HB1xp67_ASAP7_75t_L g6342 ( 
.A(n_4565),
.Y(n_6342)
);

NOR2x1_ASAP7_75t_SL g6343 ( 
.A(n_5682),
.B(n_5749),
.Y(n_6343)
);

A2O1A1Ixp33_ASAP7_75t_L g6344 ( 
.A1(n_5242),
.A2(n_5176),
.B(n_5182),
.C(n_5158),
.Y(n_6344)
);

INVx1_ASAP7_75t_L g6345 ( 
.A(n_5462),
.Y(n_6345)
);

INVx1_ASAP7_75t_L g6346 ( 
.A(n_5467),
.Y(n_6346)
);

AND2x2_ASAP7_75t_L g6347 ( 
.A(n_4953),
.B(n_4954),
.Y(n_6347)
);

INVx2_ASAP7_75t_L g6348 ( 
.A(n_5116),
.Y(n_6348)
);

NAND2xp5_ASAP7_75t_SL g6349 ( 
.A(n_5081),
.B(n_4978),
.Y(n_6349)
);

AND2x2_ASAP7_75t_L g6350 ( 
.A(n_4953),
.B(n_4954),
.Y(n_6350)
);

INVx2_ASAP7_75t_L g6351 ( 
.A(n_5116),
.Y(n_6351)
);

O2A1O1Ixp5_ASAP7_75t_L g6352 ( 
.A1(n_5350),
.A2(n_5202),
.B(n_5571),
.C(n_5576),
.Y(n_6352)
);

NOR3xp33_ASAP7_75t_L g6353 ( 
.A(n_5750),
.B(n_5710),
.C(n_5383),
.Y(n_6353)
);

NOR2x1_ASAP7_75t_L g6354 ( 
.A(n_4978),
.B(n_5002),
.Y(n_6354)
);

CKINVDCx20_ASAP7_75t_R g6355 ( 
.A(n_4869),
.Y(n_6355)
);

INVx1_ASAP7_75t_L g6356 ( 
.A(n_5467),
.Y(n_6356)
);

INVx4_ASAP7_75t_SL g6357 ( 
.A(n_5034),
.Y(n_6357)
);

INVx1_ASAP7_75t_L g6358 ( 
.A(n_5467),
.Y(n_6358)
);

NAND2xp5_ASAP7_75t_L g6359 ( 
.A(n_4905),
.B(n_4908),
.Y(n_6359)
);

INVx1_ASAP7_75t_L g6360 ( 
.A(n_5467),
.Y(n_6360)
);

AND2x4_ASAP7_75t_L g6361 ( 
.A(n_4858),
.B(n_4886),
.Y(n_6361)
);

INVx1_ASAP7_75t_L g6362 ( 
.A(n_5478),
.Y(n_6362)
);

AOI21xp5_ASAP7_75t_L g6363 ( 
.A1(n_5078),
.A2(n_5159),
.B(n_5112),
.Y(n_6363)
);

AND2x4_ASAP7_75t_L g6364 ( 
.A(n_4858),
.B(n_4886),
.Y(n_6364)
);

NOR2x1_ASAP7_75t_L g6365 ( 
.A(n_5002),
.B(n_5235),
.Y(n_6365)
);

HB1xp67_ASAP7_75t_L g6366 ( 
.A(n_4565),
.Y(n_6366)
);

INVx2_ASAP7_75t_L g6367 ( 
.A(n_5116),
.Y(n_6367)
);

HB1xp67_ASAP7_75t_L g6368 ( 
.A(n_4565),
.Y(n_6368)
);

INVxp67_ASAP7_75t_L g6369 ( 
.A(n_5401),
.Y(n_6369)
);

CKINVDCx8_ASAP7_75t_R g6370 ( 
.A(n_5374),
.Y(n_6370)
);

INVx1_ASAP7_75t_L g6371 ( 
.A(n_5478),
.Y(n_6371)
);

INVx1_ASAP7_75t_SL g6372 ( 
.A(n_5667),
.Y(n_6372)
);

AOI21xp5_ASAP7_75t_L g6373 ( 
.A1(n_5112),
.A2(n_5212),
.B(n_5159),
.Y(n_6373)
);

AND2x4_ASAP7_75t_L g6374 ( 
.A(n_4858),
.B(n_4886),
.Y(n_6374)
);

INVx1_ASAP7_75t_L g6375 ( 
.A(n_5478),
.Y(n_6375)
);

BUFx2_ASAP7_75t_SL g6376 ( 
.A(n_5193),
.Y(n_6376)
);

INVx1_ASAP7_75t_L g6377 ( 
.A(n_5478),
.Y(n_6377)
);

OAI22xp5_ASAP7_75t_SL g6378 ( 
.A1(n_5529),
.A2(n_5722),
.B1(n_5624),
.B2(n_5003),
.Y(n_6378)
);

INVx2_ASAP7_75t_SL g6379 ( 
.A(n_4882),
.Y(n_6379)
);

HAxp5_ASAP7_75t_L g6380 ( 
.A(n_4735),
.B(n_4779),
.CON(n_6380),
.SN(n_6380)
);

AND2x2_ASAP7_75t_L g6381 ( 
.A(n_4954),
.B(n_4964),
.Y(n_6381)
);

INVx2_ASAP7_75t_L g6382 ( 
.A(n_5116),
.Y(n_6382)
);

INVx3_ASAP7_75t_L g6383 ( 
.A(n_4560),
.Y(n_6383)
);

AND2x4_ASAP7_75t_L g6384 ( 
.A(n_4858),
.B(n_4886),
.Y(n_6384)
);

AOI21xp5_ASAP7_75t_L g6385 ( 
.A1(n_5112),
.A2(n_5212),
.B(n_5159),
.Y(n_6385)
);

OR2x2_ASAP7_75t_L g6386 ( 
.A(n_4848),
.B(n_4881),
.Y(n_6386)
);

INVx1_ASAP7_75t_L g6387 ( 
.A(n_5489),
.Y(n_6387)
);

AND3x1_ASAP7_75t_SL g6388 ( 
.A(n_4735),
.B(n_4745),
.C(n_5003),
.Y(n_6388)
);

INVxp67_ASAP7_75t_SL g6389 ( 
.A(n_4559),
.Y(n_6389)
);

NAND2xp5_ASAP7_75t_L g6390 ( 
.A(n_4908),
.B(n_4912),
.Y(n_6390)
);

AOI22xp5_ASAP7_75t_L g6391 ( 
.A1(n_5639),
.A2(n_5244),
.B1(n_5285),
.B2(n_5251),
.Y(n_6391)
);

OAI21xp5_ASAP7_75t_L g6392 ( 
.A1(n_5681),
.A2(n_4645),
.B(n_4644),
.Y(n_6392)
);

INVx3_ASAP7_75t_L g6393 ( 
.A(n_4560),
.Y(n_6393)
);

INVx1_ASAP7_75t_SL g6394 ( 
.A(n_5667),
.Y(n_6394)
);

OAI22xp5_ASAP7_75t_L g6395 ( 
.A1(n_5251),
.A2(n_5293),
.B1(n_5298),
.B2(n_5285),
.Y(n_6395)
);

INVx3_ASAP7_75t_SL g6396 ( 
.A(n_5632),
.Y(n_6396)
);

NAND2xp5_ASAP7_75t_L g6397 ( 
.A(n_4912),
.B(n_4919),
.Y(n_6397)
);

AOI21x1_ASAP7_75t_L g6398 ( 
.A1(n_4653),
.A2(n_4668),
.B(n_4664),
.Y(n_6398)
);

AND2x4_ASAP7_75t_L g6399 ( 
.A(n_4886),
.B(n_4895),
.Y(n_6399)
);

INVx1_ASAP7_75t_L g6400 ( 
.A(n_5489),
.Y(n_6400)
);

CKINVDCx16_ASAP7_75t_R g6401 ( 
.A(n_5495),
.Y(n_6401)
);

BUFx2_ASAP7_75t_L g6402 ( 
.A(n_4886),
.Y(n_6402)
);

AOI21xp5_ASAP7_75t_L g6403 ( 
.A1(n_5212),
.A2(n_5372),
.B(n_5286),
.Y(n_6403)
);

NAND2xp5_ASAP7_75t_L g6404 ( 
.A(n_4919),
.B(n_4927),
.Y(n_6404)
);

OAI22xp5_ASAP7_75t_L g6405 ( 
.A1(n_5293),
.A2(n_5298),
.B1(n_5294),
.B2(n_5295),
.Y(n_6405)
);

NOR2xp33_ASAP7_75t_L g6406 ( 
.A(n_4927),
.B(n_4929),
.Y(n_6406)
);

BUFx2_ASAP7_75t_L g6407 ( 
.A(n_4895),
.Y(n_6407)
);

NAND2xp5_ASAP7_75t_SL g6408 ( 
.A(n_5235),
.B(n_5243),
.Y(n_6408)
);

INVx5_ASAP7_75t_L g6409 ( 
.A(n_5020),
.Y(n_6409)
);

INVx3_ASAP7_75t_L g6410 ( 
.A(n_4560),
.Y(n_6410)
);

AOI22xp5_ASAP7_75t_L g6411 ( 
.A1(n_5639),
.A2(n_5529),
.B1(n_5042),
.B2(n_5750),
.Y(n_6411)
);

AND2x2_ASAP7_75t_L g6412 ( 
.A(n_4964),
.B(n_4966),
.Y(n_6412)
);

AOI21xp5_ASAP7_75t_L g6413 ( 
.A1(n_5212),
.A2(n_5372),
.B(n_5286),
.Y(n_6413)
);

O2A1O1Ixp33_ASAP7_75t_L g6414 ( 
.A1(n_5381),
.A2(n_5384),
.B(n_5390),
.C(n_5383),
.Y(n_6414)
);

INVx1_ASAP7_75t_L g6415 ( 
.A(n_5489),
.Y(n_6415)
);

AND2x4_ASAP7_75t_L g6416 ( 
.A(n_4895),
.B(n_4897),
.Y(n_6416)
);

INVx1_ASAP7_75t_L g6417 ( 
.A(n_5489),
.Y(n_6417)
);

OAI22xp5_ASAP7_75t_L g6418 ( 
.A1(n_5289),
.A2(n_5295),
.B1(n_5319),
.B2(n_5294),
.Y(n_6418)
);

INVx2_ASAP7_75t_L g6419 ( 
.A(n_5118),
.Y(n_6419)
);

INVx2_ASAP7_75t_SL g6420 ( 
.A(n_4882),
.Y(n_6420)
);

AND2x4_ASAP7_75t_L g6421 ( 
.A(n_4895),
.B(n_4897),
.Y(n_6421)
);

OAI22xp5_ASAP7_75t_L g6422 ( 
.A1(n_5289),
.A2(n_5319),
.B1(n_5331),
.B2(n_5327),
.Y(n_6422)
);

INVx1_ASAP7_75t_L g6423 ( 
.A(n_5491),
.Y(n_6423)
);

AOI22xp5_ASAP7_75t_L g6424 ( 
.A1(n_5042),
.A2(n_4929),
.B1(n_4937),
.B2(n_4932),
.Y(n_6424)
);

NAND2xp5_ASAP7_75t_L g6425 ( 
.A(n_4932),
.B(n_4937),
.Y(n_6425)
);

NOR2xp33_ASAP7_75t_L g6426 ( 
.A(n_4948),
.B(n_4958),
.Y(n_6426)
);

A2O1A1Ixp33_ASAP7_75t_L g6427 ( 
.A1(n_5176),
.A2(n_5183),
.B(n_5185),
.C(n_5182),
.Y(n_6427)
);

OAI22xp5_ASAP7_75t_L g6428 ( 
.A1(n_5327),
.A2(n_5331),
.B1(n_5347),
.B2(n_5341),
.Y(n_6428)
);

AOI22xp5_ASAP7_75t_L g6429 ( 
.A1(n_4948),
.A2(n_4958),
.B1(n_4982),
.B2(n_4961),
.Y(n_6429)
);

INVx2_ASAP7_75t_L g6430 ( 
.A(n_5118),
.Y(n_6430)
);

INVx3_ASAP7_75t_L g6431 ( 
.A(n_4564),
.Y(n_6431)
);

INVxp33_ASAP7_75t_SL g6432 ( 
.A(n_4654),
.Y(n_6432)
);

NAND2xp5_ASAP7_75t_L g6433 ( 
.A(n_4961),
.B(n_4982),
.Y(n_6433)
);

INVx1_ASAP7_75t_L g6434 ( 
.A(n_5491),
.Y(n_6434)
);

AND2x4_ASAP7_75t_L g6435 ( 
.A(n_4895),
.B(n_4897),
.Y(n_6435)
);

A2O1A1Ixp33_ASAP7_75t_L g6436 ( 
.A1(n_5183),
.A2(n_5186),
.B(n_5187),
.C(n_5185),
.Y(n_6436)
);

INVx1_ASAP7_75t_L g6437 ( 
.A(n_5491),
.Y(n_6437)
);

INVx1_ASAP7_75t_L g6438 ( 
.A(n_5491),
.Y(n_6438)
);

INVx2_ASAP7_75t_L g6439 ( 
.A(n_5118),
.Y(n_6439)
);

BUFx2_ASAP7_75t_L g6440 ( 
.A(n_4895),
.Y(n_6440)
);

INVx3_ASAP7_75t_L g6441 ( 
.A(n_4564),
.Y(n_6441)
);

INVx5_ASAP7_75t_L g6442 ( 
.A(n_5020),
.Y(n_6442)
);

OAI21x1_ASAP7_75t_SL g6443 ( 
.A1(n_5733),
.A2(n_5545),
.B(n_4659),
.Y(n_6443)
);

AOI21xp5_ASAP7_75t_L g6444 ( 
.A1(n_5212),
.A2(n_5372),
.B(n_5286),
.Y(n_6444)
);

INVx2_ASAP7_75t_L g6445 ( 
.A(n_5118),
.Y(n_6445)
);

BUFx2_ASAP7_75t_L g6446 ( 
.A(n_4897),
.Y(n_6446)
);

INVx3_ASAP7_75t_L g6447 ( 
.A(n_4564),
.Y(n_6447)
);

AOI21xp5_ASAP7_75t_L g6448 ( 
.A1(n_5212),
.A2(n_5372),
.B(n_5286),
.Y(n_6448)
);

NOR2xp33_ASAP7_75t_R g6449 ( 
.A(n_5425),
.B(n_5455),
.Y(n_6449)
);

NAND2xp5_ASAP7_75t_L g6450 ( 
.A(n_4983),
.B(n_4984),
.Y(n_6450)
);

A2O1A1Ixp33_ASAP7_75t_L g6451 ( 
.A1(n_5186),
.A2(n_5187),
.B(n_5530),
.C(n_5227),
.Y(n_6451)
);

NAND2xp5_ASAP7_75t_L g6452 ( 
.A(n_4983),
.B(n_4984),
.Y(n_6452)
);

CKINVDCx20_ASAP7_75t_R g6453 ( 
.A(n_4869),
.Y(n_6453)
);

NAND2xp5_ASAP7_75t_L g6454 ( 
.A(n_4988),
.B(n_4997),
.Y(n_6454)
);

BUFx2_ASAP7_75t_L g6455 ( 
.A(n_4897),
.Y(n_6455)
);

INVx2_ASAP7_75t_L g6456 ( 
.A(n_5142),
.Y(n_6456)
);

O2A1O1Ixp33_ASAP7_75t_L g6457 ( 
.A1(n_5381),
.A2(n_5390),
.B(n_5397),
.C(n_5384),
.Y(n_6457)
);

INVx1_ASAP7_75t_SL g6458 ( 
.A(n_5667),
.Y(n_6458)
);

INVx1_ASAP7_75t_L g6459 ( 
.A(n_5509),
.Y(n_6459)
);

NAND2x2_ASAP7_75t_L g6460 ( 
.A(n_4655),
.B(n_4689),
.Y(n_6460)
);

OR2x6_ASAP7_75t_L g6461 ( 
.A(n_4601),
.B(n_4625),
.Y(n_6461)
);

BUFx8_ASAP7_75t_L g6462 ( 
.A(n_5099),
.Y(n_6462)
);

INVxp67_ASAP7_75t_L g6463 ( 
.A(n_5401),
.Y(n_6463)
);

INVx2_ASAP7_75t_L g6464 ( 
.A(n_5142),
.Y(n_6464)
);

NAND2xp5_ASAP7_75t_L g6465 ( 
.A(n_4988),
.B(n_4997),
.Y(n_6465)
);

INVx1_ASAP7_75t_L g6466 ( 
.A(n_5509),
.Y(n_6466)
);

INVx1_ASAP7_75t_L g6467 ( 
.A(n_5509),
.Y(n_6467)
);

INVx1_ASAP7_75t_L g6468 ( 
.A(n_5509),
.Y(n_6468)
);

OR2x6_ASAP7_75t_L g6469 ( 
.A(n_4625),
.B(n_4673),
.Y(n_6469)
);

O2A1O1Ixp33_ASAP7_75t_L g6470 ( 
.A1(n_5397),
.A2(n_5409),
.B(n_5411),
.C(n_5399),
.Y(n_6470)
);

OR2x2_ASAP7_75t_L g6471 ( 
.A(n_4848),
.B(n_4881),
.Y(n_6471)
);

INVx3_ASAP7_75t_L g6472 ( 
.A(n_4564),
.Y(n_6472)
);

INVx2_ASAP7_75t_L g6473 ( 
.A(n_5142),
.Y(n_6473)
);

INVx2_ASAP7_75t_SL g6474 ( 
.A(n_4882),
.Y(n_6474)
);

NAND2xp5_ASAP7_75t_L g6475 ( 
.A(n_5001),
.B(n_5015),
.Y(n_6475)
);

INVx1_ASAP7_75t_L g6476 ( 
.A(n_5518),
.Y(n_6476)
);

AOI21xp5_ASAP7_75t_L g6477 ( 
.A1(n_5212),
.A2(n_5372),
.B(n_5286),
.Y(n_6477)
);

INVx2_ASAP7_75t_SL g6478 ( 
.A(n_4882),
.Y(n_6478)
);

INVx1_ASAP7_75t_L g6479 ( 
.A(n_5518),
.Y(n_6479)
);

BUFx12f_ASAP7_75t_L g6480 ( 
.A(n_5455),
.Y(n_6480)
);

AOI21x1_ASAP7_75t_L g6481 ( 
.A1(n_4653),
.A2(n_4668),
.B(n_4664),
.Y(n_6481)
);

CKINVDCx11_ASAP7_75t_R g6482 ( 
.A(n_4563),
.Y(n_6482)
);

INVx1_ASAP7_75t_L g6483 ( 
.A(n_5518),
.Y(n_6483)
);

INVx1_ASAP7_75t_L g6484 ( 
.A(n_5518),
.Y(n_6484)
);

AOI22xp33_ASAP7_75t_L g6485 ( 
.A1(n_4589),
.A2(n_4555),
.B1(n_5227),
.B2(n_5341),
.Y(n_6485)
);

INVx2_ASAP7_75t_SL g6486 ( 
.A(n_4882),
.Y(n_6486)
);

BUFx12f_ASAP7_75t_L g6487 ( 
.A(n_5461),
.Y(n_6487)
);

NAND2xp5_ASAP7_75t_L g6488 ( 
.A(n_5001),
.B(n_5015),
.Y(n_6488)
);

O2A1O1Ixp33_ASAP7_75t_L g6489 ( 
.A1(n_5399),
.A2(n_5411),
.B(n_5419),
.C(n_5409),
.Y(n_6489)
);

INVx1_ASAP7_75t_L g6490 ( 
.A(n_5522),
.Y(n_6490)
);

HB1xp67_ASAP7_75t_L g6491 ( 
.A(n_4565),
.Y(n_6491)
);

HB1xp67_ASAP7_75t_L g6492 ( 
.A(n_4561),
.Y(n_6492)
);

NOR2xp33_ASAP7_75t_L g6493 ( 
.A(n_5017),
.B(n_5021),
.Y(n_6493)
);

INVx1_ASAP7_75t_L g6494 ( 
.A(n_5522),
.Y(n_6494)
);

NOR2xp33_ASAP7_75t_L g6495 ( 
.A(n_5017),
.B(n_5021),
.Y(n_6495)
);

AOI21x1_ASAP7_75t_L g6496 ( 
.A1(n_4709),
.A2(n_4770),
.B(n_4716),
.Y(n_6496)
);

AOI21xp5_ASAP7_75t_L g6497 ( 
.A1(n_5286),
.A2(n_5391),
.B(n_5372),
.Y(n_6497)
);

NOR2xp33_ASAP7_75t_L g6498 ( 
.A(n_5023),
.B(n_5028),
.Y(n_6498)
);

INVx2_ASAP7_75t_L g6499 ( 
.A(n_5142),
.Y(n_6499)
);

AOI21xp5_ASAP7_75t_L g6500 ( 
.A1(n_5286),
.A2(n_5391),
.B(n_5372),
.Y(n_6500)
);

A2O1A1Ixp33_ASAP7_75t_SL g6501 ( 
.A1(n_5690),
.A2(n_5738),
.B(n_5732),
.C(n_5643),
.Y(n_6501)
);

AND2x2_ASAP7_75t_SL g6502 ( 
.A(n_5475),
.B(n_4625),
.Y(n_6502)
);

AOI22xp5_ASAP7_75t_L g6503 ( 
.A1(n_5023),
.A2(n_5028),
.B1(n_5351),
.B2(n_5347),
.Y(n_6503)
);

OAI21xp33_ASAP7_75t_L g6504 ( 
.A1(n_4644),
.A2(n_4645),
.B(n_5227),
.Y(n_6504)
);

NAND2xp5_ASAP7_75t_L g6505 ( 
.A(n_4614),
.B(n_5564),
.Y(n_6505)
);

HB1xp67_ASAP7_75t_L g6506 ( 
.A(n_4561),
.Y(n_6506)
);

AND2x2_ASAP7_75t_L g6507 ( 
.A(n_4970),
.B(n_4974),
.Y(n_6507)
);

A2O1A1Ixp33_ASAP7_75t_L g6508 ( 
.A1(n_5530),
.A2(n_5262),
.B(n_4735),
.C(n_5573),
.Y(n_6508)
);

A2O1A1Ixp33_ASAP7_75t_SL g6509 ( 
.A1(n_5690),
.A2(n_5738),
.B(n_5732),
.C(n_5643),
.Y(n_6509)
);

A2O1A1Ixp33_ASAP7_75t_L g6510 ( 
.A1(n_5530),
.A2(n_5262),
.B(n_5603),
.C(n_5573),
.Y(n_6510)
);

O2A1O1Ixp5_ASAP7_75t_SL g6511 ( 
.A1(n_4567),
.A2(n_5422),
.B(n_5417),
.C(n_4559),
.Y(n_6511)
);

INVx2_ASAP7_75t_L g6512 ( 
.A(n_5144),
.Y(n_6512)
);

O2A1O1Ixp33_ASAP7_75t_L g6513 ( 
.A1(n_5419),
.A2(n_5428),
.B(n_5430),
.C(n_5427),
.Y(n_6513)
);

O2A1O1Ixp33_ASAP7_75t_L g6514 ( 
.A1(n_5427),
.A2(n_5430),
.B(n_5433),
.C(n_5428),
.Y(n_6514)
);

OR2x2_ASAP7_75t_L g6515 ( 
.A(n_4848),
.B(n_4881),
.Y(n_6515)
);

NOR2xp67_ASAP7_75t_L g6516 ( 
.A(n_5198),
.B(n_5225),
.Y(n_6516)
);

AOI21xp5_ASAP7_75t_L g6517 ( 
.A1(n_5391),
.A2(n_5611),
.B(n_5542),
.Y(n_6517)
);

INVx2_ASAP7_75t_L g6518 ( 
.A(n_5144),
.Y(n_6518)
);

HB1xp67_ASAP7_75t_L g6519 ( 
.A(n_4552),
.Y(n_6519)
);

AOI21xp5_ASAP7_75t_L g6520 ( 
.A1(n_5391),
.A2(n_5611),
.B(n_5542),
.Y(n_6520)
);

BUFx2_ASAP7_75t_L g6521 ( 
.A(n_4902),
.Y(n_6521)
);

NAND2xp5_ASAP7_75t_L g6522 ( 
.A(n_4614),
.B(n_5564),
.Y(n_6522)
);

INVx2_ASAP7_75t_L g6523 ( 
.A(n_5144),
.Y(n_6523)
);

AOI21xp5_ASAP7_75t_L g6524 ( 
.A1(n_5391),
.A2(n_5611),
.B(n_5542),
.Y(n_6524)
);

INVx3_ASAP7_75t_L g6525 ( 
.A(n_4564),
.Y(n_6525)
);

OAI21xp5_ASAP7_75t_L g6526 ( 
.A1(n_5681),
.A2(n_5243),
.B(n_5543),
.Y(n_6526)
);

AOI21xp5_ASAP7_75t_L g6527 ( 
.A1(n_5391),
.A2(n_5611),
.B(n_5542),
.Y(n_6527)
);

NAND2xp5_ASAP7_75t_L g6528 ( 
.A(n_4556),
.B(n_4570),
.Y(n_6528)
);

AOI21xp5_ASAP7_75t_L g6529 ( 
.A1(n_5391),
.A2(n_5611),
.B(n_5542),
.Y(n_6529)
);

A2O1A1Ixp33_ASAP7_75t_L g6530 ( 
.A1(n_5573),
.A2(n_5603),
.B(n_5254),
.C(n_5679),
.Y(n_6530)
);

OR2x2_ASAP7_75t_L g6531 ( 
.A(n_4887),
.B(n_4904),
.Y(n_6531)
);

INVx5_ASAP7_75t_L g6532 ( 
.A(n_5020),
.Y(n_6532)
);

NAND2xp5_ASAP7_75t_L g6533 ( 
.A(n_4556),
.B(n_4570),
.Y(n_6533)
);

AOI222xp33_ASAP7_75t_L g6534 ( 
.A1(n_5351),
.A2(n_5353),
.B1(n_5356),
.B2(n_5352),
.C1(n_5537),
.C2(n_5517),
.Y(n_6534)
);

OR2x6_ASAP7_75t_L g6535 ( 
.A(n_4673),
.B(n_4679),
.Y(n_6535)
);

AOI21xp5_ASAP7_75t_L g6536 ( 
.A1(n_5542),
.A2(n_5611),
.B(n_5631),
.Y(n_6536)
);

AOI21xp33_ASAP7_75t_L g6537 ( 
.A1(n_4780),
.A2(n_4922),
.B(n_4907),
.Y(n_6537)
);

BUFx2_ASAP7_75t_L g6538 ( 
.A(n_4902),
.Y(n_6538)
);

AOI21x1_ASAP7_75t_L g6539 ( 
.A1(n_4709),
.A2(n_4770),
.B(n_4716),
.Y(n_6539)
);

AOI22xp5_ASAP7_75t_L g6540 ( 
.A1(n_5352),
.A2(n_5353),
.B1(n_5356),
.B2(n_5734),
.Y(n_6540)
);

INVx2_ASAP7_75t_L g6541 ( 
.A(n_5144),
.Y(n_6541)
);

O2A1O1Ixp33_ASAP7_75t_L g6542 ( 
.A1(n_5433),
.A2(n_5438),
.B(n_5441),
.C(n_5436),
.Y(n_6542)
);

AOI21xp5_ASAP7_75t_L g6543 ( 
.A1(n_5542),
.A2(n_5611),
.B(n_5631),
.Y(n_6543)
);

HB1xp67_ASAP7_75t_L g6544 ( 
.A(n_4552),
.Y(n_6544)
);

INVx3_ASAP7_75t_L g6545 ( 
.A(n_4564),
.Y(n_6545)
);

INVx5_ASAP7_75t_L g6546 ( 
.A(n_5020),
.Y(n_6546)
);

INVx2_ASAP7_75t_L g6547 ( 
.A(n_5147),
.Y(n_6547)
);

AND2x2_ASAP7_75t_L g6548 ( 
.A(n_4970),
.B(n_4974),
.Y(n_6548)
);

AND2x2_ASAP7_75t_L g6549 ( 
.A(n_4974),
.B(n_4985),
.Y(n_6549)
);

CKINVDCx5p33_ASAP7_75t_R g6550 ( 
.A(n_4750),
.Y(n_6550)
);

OAI22xp5_ASAP7_75t_L g6551 ( 
.A1(n_5316),
.A2(n_5438),
.B1(n_5441),
.B2(n_5436),
.Y(n_6551)
);

A2O1A1Ixp33_ASAP7_75t_L g6552 ( 
.A1(n_5603),
.A2(n_5254),
.B(n_5679),
.C(n_5677),
.Y(n_6552)
);

INVx2_ASAP7_75t_SL g6553 ( 
.A(n_4882),
.Y(n_6553)
);

AOI22xp33_ASAP7_75t_SL g6554 ( 
.A1(n_5597),
.A2(n_5475),
.B1(n_4790),
.B2(n_4904),
.Y(n_6554)
);

OR2x6_ASAP7_75t_L g6555 ( 
.A(n_4673),
.B(n_4679),
.Y(n_6555)
);

OAI22xp5_ASAP7_75t_L g6556 ( 
.A1(n_5316),
.A2(n_5460),
.B1(n_5452),
.B2(n_5247),
.Y(n_6556)
);

OR2x2_ASAP7_75t_L g6557 ( 
.A(n_4887),
.B(n_4904),
.Y(n_6557)
);

NAND2xp5_ASAP7_75t_L g6558 ( 
.A(n_4588),
.B(n_5602),
.Y(n_6558)
);

NAND2xp5_ASAP7_75t_L g6559 ( 
.A(n_4588),
.B(n_5602),
.Y(n_6559)
);

BUFx2_ASAP7_75t_L g6560 ( 
.A(n_4902),
.Y(n_6560)
);

AOI21xp5_ASAP7_75t_L g6561 ( 
.A1(n_5635),
.A2(n_5642),
.B(n_5648),
.Y(n_6561)
);

AOI22xp33_ASAP7_75t_L g6562 ( 
.A1(n_4555),
.A2(n_5043),
.B1(n_5537),
.B2(n_4838),
.Y(n_6562)
);

AOI22xp33_ASAP7_75t_L g6563 ( 
.A1(n_5043),
.A2(n_4838),
.B1(n_5003),
.B2(n_5476),
.Y(n_6563)
);

NOR2xp33_ASAP7_75t_L g6564 ( 
.A(n_4888),
.B(n_4626),
.Y(n_6564)
);

HB1xp67_ASAP7_75t_L g6565 ( 
.A(n_4552),
.Y(n_6565)
);

AOI221xp5_ASAP7_75t_L g6566 ( 
.A1(n_5452),
.A2(n_5460),
.B1(n_5250),
.B2(n_5252),
.C(n_5249),
.Y(n_6566)
);

A2O1A1Ixp33_ASAP7_75t_L g6567 ( 
.A1(n_5254),
.A2(n_5679),
.B(n_5685),
.C(n_5677),
.Y(n_6567)
);

NAND2xp5_ASAP7_75t_L g6568 ( 
.A(n_5602),
.B(n_5607),
.Y(n_6568)
);

HAxp5_ASAP7_75t_L g6569 ( 
.A(n_5316),
.B(n_4888),
.CON(n_6569),
.SN(n_6569)
);

NAND2xp5_ASAP7_75t_L g6570 ( 
.A(n_5607),
.B(n_5612),
.Y(n_6570)
);

OAI222xp33_ASAP7_75t_L g6571 ( 
.A1(n_5431),
.A2(n_5481),
.B1(n_4619),
.B2(n_4622),
.C1(n_5486),
.C2(n_5477),
.Y(n_6571)
);

INVx4_ASAP7_75t_L g6572 ( 
.A(n_4764),
.Y(n_6572)
);

NAND3xp33_ASAP7_75t_SL g6573 ( 
.A(n_4790),
.B(n_4721),
.C(n_4971),
.Y(n_6573)
);

AOI22xp5_ASAP7_75t_L g6574 ( 
.A1(n_5734),
.A2(n_5702),
.B1(n_4562),
.B2(n_5476),
.Y(n_6574)
);

OAI22xp5_ASAP7_75t_SL g6575 ( 
.A1(n_5624),
.A2(n_5722),
.B1(n_5003),
.B2(n_5025),
.Y(n_6575)
);

O2A1O1Ixp33_ASAP7_75t_L g6576 ( 
.A1(n_5247),
.A2(n_5250),
.B(n_5252),
.C(n_5249),
.Y(n_6576)
);

AOI21xp5_ASAP7_75t_L g6577 ( 
.A1(n_5635),
.A2(n_5642),
.B(n_5406),
.Y(n_6577)
);

INVxp67_ASAP7_75t_L g6578 ( 
.A(n_5654),
.Y(n_6578)
);

AOI21xp5_ASAP7_75t_L g6579 ( 
.A1(n_5299),
.A2(n_5494),
.B(n_5406),
.Y(n_6579)
);

AOI21xp5_ASAP7_75t_L g6580 ( 
.A1(n_5299),
.A2(n_5494),
.B(n_5406),
.Y(n_6580)
);

INVx2_ASAP7_75t_SL g6581 ( 
.A(n_4882),
.Y(n_6581)
);

AOI22xp5_ASAP7_75t_L g6582 ( 
.A1(n_5702),
.A2(n_4562),
.B1(n_5481),
.B2(n_5431),
.Y(n_6582)
);

CKINVDCx14_ASAP7_75t_R g6583 ( 
.A(n_5009),
.Y(n_6583)
);

INVxp67_ASAP7_75t_L g6584 ( 
.A(n_5654),
.Y(n_6584)
);

BUFx6f_ASAP7_75t_SL g6585 ( 
.A(n_5632),
.Y(n_6585)
);

OR2x2_ASAP7_75t_L g6586 ( 
.A(n_4887),
.B(n_4906),
.Y(n_6586)
);

INVxp67_ASAP7_75t_L g6587 ( 
.A(n_5654),
.Y(n_6587)
);

AOI222xp33_ASAP7_75t_L g6588 ( 
.A1(n_5517),
.A2(n_4595),
.B1(n_4830),
.B2(n_5265),
.C1(n_5266),
.C2(n_5261),
.Y(n_6588)
);

AOI221xp5_ASAP7_75t_L g6589 ( 
.A1(n_5261),
.A2(n_5277),
.B1(n_5278),
.B2(n_5266),
.C(n_5265),
.Y(n_6589)
);

NAND2xp5_ASAP7_75t_SL g6590 ( 
.A(n_5683),
.B(n_5684),
.Y(n_6590)
);

A2O1A1Ixp33_ASAP7_75t_L g6591 ( 
.A1(n_5254),
.A2(n_5685),
.B(n_5677),
.C(n_4739),
.Y(n_6591)
);

NOR2xp33_ASAP7_75t_L g6592 ( 
.A(n_4888),
.B(n_4626),
.Y(n_6592)
);

CKINVDCx14_ASAP7_75t_R g6593 ( 
.A(n_5009),
.Y(n_6593)
);

NAND3xp33_ASAP7_75t_L g6594 ( 
.A(n_5614),
.B(n_5706),
.C(n_5694),
.Y(n_6594)
);

CKINVDCx5p33_ASAP7_75t_R g6595 ( 
.A(n_4654),
.Y(n_6595)
);

BUFx2_ASAP7_75t_L g6596 ( 
.A(n_4938),
.Y(n_6596)
);

CKINVDCx5p33_ASAP7_75t_R g6597 ( 
.A(n_5461),
.Y(n_6597)
);

HB1xp67_ASAP7_75t_L g6598 ( 
.A(n_4551),
.Y(n_6598)
);

NOR2xp33_ASAP7_75t_L g6599 ( 
.A(n_5069),
.B(n_5498),
.Y(n_6599)
);

OR2x6_ASAP7_75t_L g6600 ( 
.A(n_4679),
.B(n_4682),
.Y(n_6600)
);

AO22x1_ASAP7_75t_L g6601 ( 
.A1(n_5035),
.A2(n_5523),
.B1(n_5534),
.B2(n_5140),
.Y(n_6601)
);

NAND2xp5_ASAP7_75t_SL g6602 ( 
.A(n_5683),
.B(n_5684),
.Y(n_6602)
);

AND2x2_ASAP7_75t_L g6603 ( 
.A(n_4985),
.B(n_5036),
.Y(n_6603)
);

OR2x6_ASAP7_75t_L g6604 ( 
.A(n_4682),
.B(n_4707),
.Y(n_6604)
);

NOR2xp33_ASAP7_75t_L g6605 ( 
.A(n_5069),
.B(n_5498),
.Y(n_6605)
);

INVx4_ASAP7_75t_L g6606 ( 
.A(n_4764),
.Y(n_6606)
);

NOR2xp33_ASAP7_75t_L g6607 ( 
.A(n_5070),
.B(n_4616),
.Y(n_6607)
);

INVx4_ASAP7_75t_L g6608 ( 
.A(n_4764),
.Y(n_6608)
);

NOR2x1_ASAP7_75t_SL g6609 ( 
.A(n_5682),
.B(n_5317),
.Y(n_6609)
);

NAND2xp5_ASAP7_75t_SL g6610 ( 
.A(n_4616),
.B(n_4621),
.Y(n_6610)
);

O2A1O1Ixp33_ASAP7_75t_L g6611 ( 
.A1(n_5277),
.A2(n_5280),
.B(n_5284),
.C(n_5278),
.Y(n_6611)
);

NAND2xp5_ASAP7_75t_SL g6612 ( 
.A(n_4621),
.B(n_5692),
.Y(n_6612)
);

NAND2xp5_ASAP7_75t_SL g6613 ( 
.A(n_5692),
.B(n_4628),
.Y(n_6613)
);

AOI21x1_ASAP7_75t_SL g6614 ( 
.A1(n_4985),
.A2(n_5045),
.B(n_5036),
.Y(n_6614)
);

A2O1A1Ixp33_ASAP7_75t_L g6615 ( 
.A1(n_5254),
.A2(n_5685),
.B(n_4739),
.C(n_4766),
.Y(n_6615)
);

BUFx2_ASAP7_75t_L g6616 ( 
.A(n_4968),
.Y(n_6616)
);

HB1xp67_ASAP7_75t_L g6617 ( 
.A(n_4551),
.Y(n_6617)
);

A2O1A1Ixp33_ASAP7_75t_L g6618 ( 
.A1(n_5254),
.A2(n_4739),
.B(n_4766),
.C(n_4719),
.Y(n_6618)
);

INVx1_ASAP7_75t_L g6619 ( 
.A(n_5361),
.Y(n_6619)
);

INVx1_ASAP7_75t_L g6620 ( 
.A(n_5361),
.Y(n_6620)
);

AND2x4_ASAP7_75t_L g6621 ( 
.A(n_4968),
.B(n_4994),
.Y(n_6621)
);

OR2x6_ASAP7_75t_L g6622 ( 
.A(n_4682),
.B(n_4707),
.Y(n_6622)
);

A2O1A1Ixp33_ASAP7_75t_L g6623 ( 
.A1(n_4719),
.A2(n_4766),
.B(n_4739),
.C(n_4906),
.Y(n_6623)
);

INVx1_ASAP7_75t_L g6624 ( 
.A(n_5361),
.Y(n_6624)
);

INVx1_ASAP7_75t_L g6625 ( 
.A(n_5366),
.Y(n_6625)
);

OR2x6_ASAP7_75t_L g6626 ( 
.A(n_4707),
.B(n_4729),
.Y(n_6626)
);

AND2x2_ASAP7_75t_L g6627 ( 
.A(n_5036),
.B(n_5045),
.Y(n_6627)
);

OR2x6_ASAP7_75t_L g6628 ( 
.A(n_4729),
.B(n_4765),
.Y(n_6628)
);

INVx4_ASAP7_75t_L g6629 ( 
.A(n_4764),
.Y(n_6629)
);

AOI22xp33_ASAP7_75t_L g6630 ( 
.A1(n_5622),
.A2(n_5694),
.B1(n_5706),
.B2(n_5614),
.Y(n_6630)
);

AND2x2_ASAP7_75t_L g6631 ( 
.A(n_5045),
.B(n_5050),
.Y(n_6631)
);

BUFx2_ASAP7_75t_L g6632 ( 
.A(n_4968),
.Y(n_6632)
);

BUFx12f_ASAP7_75t_L g6633 ( 
.A(n_5470),
.Y(n_6633)
);

NAND2xp5_ASAP7_75t_L g6634 ( 
.A(n_5623),
.B(n_5676),
.Y(n_6634)
);

INVx2_ASAP7_75t_L g6635 ( 
.A(n_5162),
.Y(n_6635)
);

INVx1_ASAP7_75t_L g6636 ( 
.A(n_5366),
.Y(n_6636)
);

AOI22xp33_ASAP7_75t_SL g6637 ( 
.A1(n_5475),
.A2(n_4921),
.B1(n_4936),
.B2(n_4906),
.Y(n_6637)
);

A2O1A1Ixp33_ASAP7_75t_L g6638 ( 
.A1(n_4719),
.A2(n_4766),
.B(n_4739),
.C(n_4921),
.Y(n_6638)
);

NAND2xp5_ASAP7_75t_L g6639 ( 
.A(n_5623),
.B(n_5676),
.Y(n_6639)
);

CKINVDCx11_ASAP7_75t_R g6640 ( 
.A(n_4630),
.Y(n_6640)
);

HB1xp67_ASAP7_75t_L g6641 ( 
.A(n_4551),
.Y(n_6641)
);

NAND2xp5_ASAP7_75t_SL g6642 ( 
.A(n_4628),
.B(n_4636),
.Y(n_6642)
);

NOR2xp67_ASAP7_75t_L g6643 ( 
.A(n_5225),
.B(n_4949),
.Y(n_6643)
);

CKINVDCx11_ASAP7_75t_R g6644 ( 
.A(n_4630),
.Y(n_6644)
);

AOI21x1_ASAP7_75t_L g6645 ( 
.A1(n_4917),
.A2(n_5029),
.B(n_4950),
.Y(n_6645)
);

NAND2xp5_ASAP7_75t_L g6646 ( 
.A(n_4619),
.B(n_4622),
.Y(n_6646)
);

O2A1O1Ixp33_ASAP7_75t_L g6647 ( 
.A1(n_5280),
.A2(n_5284),
.B(n_5288),
.C(n_4636),
.Y(n_6647)
);

AND2x2_ASAP7_75t_L g6648 ( 
.A(n_5050),
.B(n_5067),
.Y(n_6648)
);

AOI22xp5_ASAP7_75t_L g6649 ( 
.A1(n_5604),
.A2(n_5622),
.B1(n_5288),
.B2(n_5693),
.Y(n_6649)
);

NOR2x1_ASAP7_75t_L g6650 ( 
.A(n_5715),
.B(n_5721),
.Y(n_6650)
);

INVx1_ASAP7_75t_L g6651 ( 
.A(n_5366),
.Y(n_6651)
);

INVx1_ASAP7_75t_L g6652 ( 
.A(n_5367),
.Y(n_6652)
);

AO22x1_ASAP7_75t_L g6653 ( 
.A1(n_5035),
.A2(n_5523),
.B1(n_5534),
.B2(n_5140),
.Y(n_6653)
);

AND2x4_ASAP7_75t_L g6654 ( 
.A(n_4994),
.B(n_4719),
.Y(n_6654)
);

AOI22xp5_ASAP7_75t_L g6655 ( 
.A1(n_5604),
.A2(n_5693),
.B1(n_5666),
.B2(n_5541),
.Y(n_6655)
);

NAND2xp5_ASAP7_75t_L g6656 ( 
.A(n_4619),
.B(n_4622),
.Y(n_6656)
);

AND2x2_ASAP7_75t_L g6657 ( 
.A(n_5050),
.B(n_5067),
.Y(n_6657)
);

NAND2x1p5_ASAP7_75t_L g6658 ( 
.A(n_4719),
.B(n_4766),
.Y(n_6658)
);

NOR2xp33_ASAP7_75t_L g6659 ( 
.A(n_5070),
.B(n_5479),
.Y(n_6659)
);

INVx1_ASAP7_75t_L g6660 ( 
.A(n_5367),
.Y(n_6660)
);

INVx2_ASAP7_75t_L g6661 ( 
.A(n_5168),
.Y(n_6661)
);

INVx1_ASAP7_75t_L g6662 ( 
.A(n_5367),
.Y(n_6662)
);

NOR2xp33_ASAP7_75t_L g6663 ( 
.A(n_5479),
.B(n_5482),
.Y(n_6663)
);

OAI22xp5_ASAP7_75t_L g6664 ( 
.A1(n_5558),
.A2(n_5477),
.B1(n_5486),
.B2(n_4651),
.Y(n_6664)
);

O2A1O1Ixp33_ASAP7_75t_L g6665 ( 
.A1(n_4780),
.A2(n_4922),
.B(n_5134),
.C(n_4907),
.Y(n_6665)
);

BUFx2_ASAP7_75t_L g6666 ( 
.A(n_4994),
.Y(n_6666)
);

INVx1_ASAP7_75t_L g6667 ( 
.A(n_5371),
.Y(n_6667)
);

INVx1_ASAP7_75t_L g6668 ( 
.A(n_5371),
.Y(n_6668)
);

O2A1O1Ixp5_ASAP7_75t_L g6669 ( 
.A1(n_5202),
.A2(n_5581),
.B(n_5576),
.C(n_5079),
.Y(n_6669)
);

NOR2xp33_ASAP7_75t_L g6670 ( 
.A(n_5482),
.B(n_5488),
.Y(n_6670)
);

INVx1_ASAP7_75t_L g6671 ( 
.A(n_5371),
.Y(n_6671)
);

INVx2_ASAP7_75t_L g6672 ( 
.A(n_5168),
.Y(n_6672)
);

AOI21xp5_ASAP7_75t_L g6673 ( 
.A1(n_5299),
.A2(n_5494),
.B(n_5406),
.Y(n_6673)
);

AOI21xp5_ASAP7_75t_L g6674 ( 
.A1(n_5299),
.A2(n_5494),
.B(n_5406),
.Y(n_6674)
);

OAI22xp5_ASAP7_75t_L g6675 ( 
.A1(n_5558),
.A2(n_4651),
.B1(n_4629),
.B2(n_4587),
.Y(n_6675)
);

O2A1O1Ixp5_ASAP7_75t_L g6676 ( 
.A1(n_5202),
.A2(n_5581),
.B(n_5079),
.C(n_5095),
.Y(n_6676)
);

BUFx12f_ASAP7_75t_L g6677 ( 
.A(n_5470),
.Y(n_6677)
);

AND2x4_ASAP7_75t_L g6678 ( 
.A(n_4994),
.B(n_4766),
.Y(n_6678)
);

O2A1O1Ixp33_ASAP7_75t_L g6679 ( 
.A1(n_5134),
.A2(n_5204),
.B(n_5740),
.C(n_5739),
.Y(n_6679)
);

INVx1_ASAP7_75t_L g6680 ( 
.A(n_5375),
.Y(n_6680)
);

NOR2xp67_ASAP7_75t_L g6681 ( 
.A(n_5225),
.B(n_4949),
.Y(n_6681)
);

INVx4_ASAP7_75t_L g6682 ( 
.A(n_4778),
.Y(n_6682)
);

INVx3_ASAP7_75t_SL g6683 ( 
.A(n_5632),
.Y(n_6683)
);

AOI21xp5_ASAP7_75t_L g6684 ( 
.A1(n_5299),
.A2(n_5531),
.B(n_5494),
.Y(n_6684)
);

OAI22xp5_ASAP7_75t_SL g6685 ( 
.A1(n_5012),
.A2(n_5057),
.B1(n_5201),
.B2(n_5025),
.Y(n_6685)
);

BUFx8_ASAP7_75t_L g6686 ( 
.A(n_5099),
.Y(n_6686)
);

AND2x4_ASAP7_75t_L g6687 ( 
.A(n_4994),
.B(n_4766),
.Y(n_6687)
);

O2A1O1Ixp33_ASAP7_75t_L g6688 ( 
.A1(n_5134),
.A2(n_5204),
.B(n_5740),
.C(n_5739),
.Y(n_6688)
);

AND2x2_ASAP7_75t_L g6689 ( 
.A(n_5067),
.B(n_5079),
.Y(n_6689)
);

NOR2xp33_ASAP7_75t_L g6690 ( 
.A(n_5488),
.B(n_5496),
.Y(n_6690)
);

BUFx4f_ASAP7_75t_SL g6691 ( 
.A(n_4630),
.Y(n_6691)
);

BUFx2_ASAP7_75t_L g6692 ( 
.A(n_4994),
.Y(n_6692)
);

INVx1_ASAP7_75t_L g6693 ( 
.A(n_5375),
.Y(n_6693)
);

INVx1_ASAP7_75t_SL g6694 ( 
.A(n_4989),
.Y(n_6694)
);

AOI21xp5_ASAP7_75t_L g6695 ( 
.A1(n_5531),
.A2(n_5609),
.B(n_5608),
.Y(n_6695)
);

NAND2xp5_ASAP7_75t_L g6696 ( 
.A(n_5675),
.B(n_5582),
.Y(n_6696)
);

HB1xp67_ASAP7_75t_L g6697 ( 
.A(n_4582),
.Y(n_6697)
);

NAND2x1p5_ASAP7_75t_L g6698 ( 
.A(n_4766),
.B(n_4670),
.Y(n_6698)
);

AOI22xp33_ASAP7_75t_L g6699 ( 
.A1(n_5099),
.A2(n_5154),
.B1(n_5296),
.B2(n_5167),
.Y(n_6699)
);

INVx1_ASAP7_75t_L g6700 ( 
.A(n_5375),
.Y(n_6700)
);

INVx2_ASAP7_75t_SL g6701 ( 
.A(n_5718),
.Y(n_6701)
);

NAND2xp5_ASAP7_75t_L g6702 ( 
.A(n_5675),
.B(n_5582),
.Y(n_6702)
);

CKINVDCx8_ASAP7_75t_R g6703 ( 
.A(n_5374),
.Y(n_6703)
);

NAND2xp5_ASAP7_75t_L g6704 ( 
.A(n_5675),
.B(n_5585),
.Y(n_6704)
);

INVx1_ASAP7_75t_L g6705 ( 
.A(n_5377),
.Y(n_6705)
);

INVx6_ASAP7_75t_L g6706 ( 
.A(n_4674),
.Y(n_6706)
);

AOI21xp5_ASAP7_75t_L g6707 ( 
.A1(n_5531),
.A2(n_5609),
.B(n_5608),
.Y(n_6707)
);

INVx5_ASAP7_75t_L g6708 ( 
.A(n_5020),
.Y(n_6708)
);

OR2x2_ASAP7_75t_L g6709 ( 
.A(n_4921),
.B(n_4936),
.Y(n_6709)
);

INVx1_ASAP7_75t_L g6710 ( 
.A(n_5377),
.Y(n_6710)
);

A2O1A1Ixp33_ASAP7_75t_L g6711 ( 
.A1(n_4766),
.A2(n_4955),
.B(n_4962),
.C(n_4936),
.Y(n_6711)
);

INVx1_ASAP7_75t_L g6712 ( 
.A(n_5377),
.Y(n_6712)
);

A2O1A1Ixp33_ASAP7_75t_L g6713 ( 
.A1(n_4955),
.A2(n_4999),
.B(n_5007),
.C(n_4962),
.Y(n_6713)
);

NAND2xp5_ASAP7_75t_SL g6714 ( 
.A(n_5659),
.B(n_5661),
.Y(n_6714)
);

OR2x6_ASAP7_75t_L g6715 ( 
.A(n_4729),
.B(n_4765),
.Y(n_6715)
);

NAND2xp5_ASAP7_75t_L g6716 ( 
.A(n_5585),
.B(n_5586),
.Y(n_6716)
);

A2O1A1Ixp33_ASAP7_75t_L g6717 ( 
.A1(n_4955),
.A2(n_4999),
.B(n_5007),
.C(n_4962),
.Y(n_6717)
);

NAND2xp5_ASAP7_75t_L g6718 ( 
.A(n_5586),
.B(n_5588),
.Y(n_6718)
);

HB1xp67_ASAP7_75t_L g6719 ( 
.A(n_4582),
.Y(n_6719)
);

AND2x4_ASAP7_75t_L g6720 ( 
.A(n_4949),
.B(n_4981),
.Y(n_6720)
);

NAND2xp5_ASAP7_75t_L g6721 ( 
.A(n_5588),
.B(n_5596),
.Y(n_6721)
);

AND2x2_ASAP7_75t_L g6722 ( 
.A(n_5095),
.B(n_5173),
.Y(n_6722)
);

OA21x2_ASAP7_75t_L g6723 ( 
.A1(n_4585),
.A2(n_5137),
.B(n_5578),
.Y(n_6723)
);

AND2x2_ASAP7_75t_L g6724 ( 
.A(n_5095),
.B(n_5173),
.Y(n_6724)
);

O2A1O1Ixp33_ASAP7_75t_L g6725 ( 
.A1(n_5204),
.A2(n_5724),
.B(n_5007),
.C(n_5016),
.Y(n_6725)
);

NAND2xp5_ASAP7_75t_L g6726 ( 
.A(n_5596),
.B(n_5600),
.Y(n_6726)
);

INVx1_ASAP7_75t_L g6727 ( 
.A(n_5386),
.Y(n_6727)
);

NAND2xp5_ASAP7_75t_L g6728 ( 
.A(n_5600),
.B(n_5606),
.Y(n_6728)
);

AOI22xp33_ASAP7_75t_L g6729 ( 
.A1(n_5099),
.A2(n_5167),
.B1(n_5296),
.B2(n_5154),
.Y(n_6729)
);

BUFx12f_ASAP7_75t_L g6730 ( 
.A(n_5535),
.Y(n_6730)
);

CKINVDCx5p33_ASAP7_75t_R g6731 ( 
.A(n_5535),
.Y(n_6731)
);

AOI22xp5_ASAP7_75t_L g6732 ( 
.A1(n_5541),
.A2(n_5666),
.B1(n_5552),
.B2(n_5569),
.Y(n_6732)
);

NAND2x1p5_ASAP7_75t_L g6733 ( 
.A(n_4670),
.B(n_4672),
.Y(n_6733)
);

A2O1A1Ixp33_ASAP7_75t_L g6734 ( 
.A1(n_4999),
.A2(n_5055),
.B(n_5085),
.C(n_5016),
.Y(n_6734)
);

INVx1_ASAP7_75t_SL g6735 ( 
.A(n_4989),
.Y(n_6735)
);

NAND2xp5_ASAP7_75t_SL g6736 ( 
.A(n_5659),
.B(n_5661),
.Y(n_6736)
);

A2O1A1Ixp33_ASAP7_75t_L g6737 ( 
.A1(n_5016),
.A2(n_5085),
.B(n_5096),
.C(n_5055),
.Y(n_6737)
);

NAND2xp5_ASAP7_75t_L g6738 ( 
.A(n_5606),
.B(n_5616),
.Y(n_6738)
);

NAND2xp5_ASAP7_75t_L g6739 ( 
.A(n_5616),
.B(n_5618),
.Y(n_6739)
);

AOI21xp5_ASAP7_75t_L g6740 ( 
.A1(n_5609),
.A2(n_5617),
.B(n_5610),
.Y(n_6740)
);

HB1xp67_ASAP7_75t_L g6741 ( 
.A(n_4582),
.Y(n_6741)
);

INVx4_ASAP7_75t_L g6742 ( 
.A(n_4778),
.Y(n_6742)
);

INVx1_ASAP7_75t_L g6743 ( 
.A(n_5386),
.Y(n_6743)
);

AOI21xp5_ASAP7_75t_L g6744 ( 
.A1(n_5610),
.A2(n_5651),
.B(n_5617),
.Y(n_6744)
);

OAI21x1_ASAP7_75t_L g6745 ( 
.A1(n_5137),
.A2(n_5281),
.B(n_5241),
.Y(n_6745)
);

NAND2xp5_ASAP7_75t_L g6746 ( 
.A(n_5618),
.B(n_5620),
.Y(n_6746)
);

NAND2x1p5_ASAP7_75t_L g6747 ( 
.A(n_4670),
.B(n_4672),
.Y(n_6747)
);

HB1xp67_ASAP7_75t_L g6748 ( 
.A(n_5626),
.Y(n_6748)
);

AOI22xp33_ASAP7_75t_L g6749 ( 
.A1(n_5154),
.A2(n_5296),
.B1(n_5167),
.B2(n_5178),
.Y(n_6749)
);

NOR2xp33_ASAP7_75t_L g6750 ( 
.A(n_5496),
.B(n_5395),
.Y(n_6750)
);

BUFx2_ASAP7_75t_L g6751 ( 
.A(n_5395),
.Y(n_6751)
);

INVx1_ASAP7_75t_L g6752 ( 
.A(n_5386),
.Y(n_6752)
);

NAND2xp5_ASAP7_75t_L g6753 ( 
.A(n_5620),
.B(n_5592),
.Y(n_6753)
);

AND2x2_ASAP7_75t_L g6754 ( 
.A(n_5173),
.B(n_5178),
.Y(n_6754)
);

AOI22xp5_ASAP7_75t_L g6755 ( 
.A1(n_5552),
.A2(n_5569),
.B1(n_4642),
.B2(n_5744),
.Y(n_6755)
);

BUFx2_ASAP7_75t_L g6756 ( 
.A(n_5395),
.Y(n_6756)
);

NOR2xp33_ASAP7_75t_L g6757 ( 
.A(n_5395),
.B(n_4651),
.Y(n_6757)
);

NOR2xp67_ASAP7_75t_L g6758 ( 
.A(n_4949),
.B(n_4981),
.Y(n_6758)
);

NAND2xp5_ASAP7_75t_SL g6759 ( 
.A(n_5543),
.B(n_4971),
.Y(n_6759)
);

BUFx8_ASAP7_75t_L g6760 ( 
.A(n_5154),
.Y(n_6760)
);

NOR2xp33_ASAP7_75t_L g6761 ( 
.A(n_4651),
.B(n_5208),
.Y(n_6761)
);

INVx1_ASAP7_75t_L g6762 ( 
.A(n_5388),
.Y(n_6762)
);

OA22x2_ASAP7_75t_L g6763 ( 
.A1(n_5148),
.A2(n_5264),
.B1(n_5474),
.B2(n_5413),
.Y(n_6763)
);

OAI22xp5_ASAP7_75t_SL g6764 ( 
.A1(n_5012),
.A2(n_5201),
.B1(n_5057),
.B2(n_4963),
.Y(n_6764)
);

OR2x6_ASAP7_75t_L g6765 ( 
.A(n_4765),
.B(n_4788),
.Y(n_6765)
);

AOI21x1_ASAP7_75t_L g6766 ( 
.A1(n_4917),
.A2(n_5029),
.B(n_4950),
.Y(n_6766)
);

AOI21xp5_ASAP7_75t_L g6767 ( 
.A1(n_5651),
.A2(n_5272),
.B(n_5256),
.Y(n_6767)
);

CKINVDCx11_ASAP7_75t_R g6768 ( 
.A(n_4657),
.Y(n_6768)
);

INVx1_ASAP7_75t_L g6769 ( 
.A(n_5388),
.Y(n_6769)
);

NAND2xp5_ASAP7_75t_L g6770 ( 
.A(n_5592),
.B(n_5594),
.Y(n_6770)
);

INVx5_ASAP7_75t_L g6771 ( 
.A(n_5020),
.Y(n_6771)
);

A2O1A1Ixp33_ASAP7_75t_SL g6772 ( 
.A1(n_5638),
.A2(n_5649),
.B(n_5657),
.C(n_5643),
.Y(n_6772)
);

A2O1A1Ixp33_ASAP7_75t_L g6773 ( 
.A1(n_5055),
.A2(n_5096),
.B(n_5165),
.C(n_5085),
.Y(n_6773)
);

NAND2xp5_ASAP7_75t_L g6774 ( 
.A(n_5592),
.B(n_5594),
.Y(n_6774)
);

OR2x6_ASAP7_75t_L g6775 ( 
.A(n_4788),
.B(n_4813),
.Y(n_6775)
);

INVx5_ASAP7_75t_L g6776 ( 
.A(n_5020),
.Y(n_6776)
);

NAND2xp5_ASAP7_75t_L g6777 ( 
.A(n_5594),
.B(n_5598),
.Y(n_6777)
);

OAI22xp33_ASAP7_75t_L g6778 ( 
.A1(n_4642),
.A2(n_4651),
.B1(n_5296),
.B2(n_5167),
.Y(n_6778)
);

AOI21xp5_ASAP7_75t_L g6779 ( 
.A1(n_5256),
.A2(n_5376),
.B(n_5272),
.Y(n_6779)
);

AOI21xp5_ASAP7_75t_L g6780 ( 
.A1(n_5256),
.A2(n_5376),
.B(n_5272),
.Y(n_6780)
);

A2O1A1Ixp33_ASAP7_75t_L g6781 ( 
.A1(n_5096),
.A2(n_5165),
.B(n_5202),
.C(n_5490),
.Y(n_6781)
);

O2A1O1Ixp5_ASAP7_75t_SL g6782 ( 
.A1(n_5422),
.A2(n_5649),
.B(n_5657),
.C(n_5638),
.Y(n_6782)
);

INVx6_ASAP7_75t_L g6783 ( 
.A(n_4674),
.Y(n_6783)
);

BUFx4f_ASAP7_75t_SL g6784 ( 
.A(n_4657),
.Y(n_6784)
);

AOI22xp33_ASAP7_75t_L g6785 ( 
.A1(n_5165),
.A2(n_4666),
.B1(n_4717),
.B2(n_4657),
.Y(n_6785)
);

INVx1_ASAP7_75t_L g6786 ( 
.A(n_5388),
.Y(n_6786)
);

AOI21xp5_ASAP7_75t_L g6787 ( 
.A1(n_5256),
.A2(n_5376),
.B(n_5272),
.Y(n_6787)
);

AND2x2_ASAP7_75t_L g6788 ( 
.A(n_4788),
.B(n_4813),
.Y(n_6788)
);

AOI21xp5_ASAP7_75t_L g6789 ( 
.A1(n_5256),
.A2(n_5376),
.B(n_5272),
.Y(n_6789)
);

INVx1_ASAP7_75t_L g6790 ( 
.A(n_5400),
.Y(n_6790)
);

INVx4_ASAP7_75t_L g6791 ( 
.A(n_4797),
.Y(n_6791)
);

OR2x6_ASAP7_75t_L g6792 ( 
.A(n_4813),
.B(n_4981),
.Y(n_6792)
);

AOI21xp5_ASAP7_75t_L g6793 ( 
.A1(n_5256),
.A2(n_5376),
.B(n_5272),
.Y(n_6793)
);

OR2x6_ASAP7_75t_L g6794 ( 
.A(n_4981),
.B(n_5008),
.Y(n_6794)
);

O2A1O1Ixp33_ASAP7_75t_L g6795 ( 
.A1(n_5724),
.A2(n_4629),
.B(n_4714),
.C(n_4587),
.Y(n_6795)
);

AOI22xp33_ASAP7_75t_L g6796 ( 
.A1(n_4657),
.A2(n_4717),
.B1(n_4876),
.B2(n_4666),
.Y(n_6796)
);

NAND2xp5_ASAP7_75t_SL g6797 ( 
.A(n_5504),
.B(n_5507),
.Y(n_6797)
);

NAND2xp5_ASAP7_75t_L g6798 ( 
.A(n_5598),
.B(n_5599),
.Y(n_6798)
);

OR2x6_ASAP7_75t_L g6799 ( 
.A(n_5008),
.B(n_5019),
.Y(n_6799)
);

INVx1_ASAP7_75t_L g6800 ( 
.A(n_5400),
.Y(n_6800)
);

BUFx2_ASAP7_75t_SL g6801 ( 
.A(n_5374),
.Y(n_6801)
);

INVx5_ASAP7_75t_L g6802 ( 
.A(n_5030),
.Y(n_6802)
);

AOI21xp33_ASAP7_75t_L g6803 ( 
.A1(n_5626),
.A2(n_5630),
.B(n_5566),
.Y(n_6803)
);

INVxp33_ASAP7_75t_SL g6804 ( 
.A(n_4789),
.Y(n_6804)
);

OAI21x1_ASAP7_75t_L g6805 ( 
.A1(n_5281),
.A2(n_5241),
.B(n_4995),
.Y(n_6805)
);

NOR2xp33_ASAP7_75t_L g6806 ( 
.A(n_5208),
.B(n_5209),
.Y(n_6806)
);

NAND2xp5_ASAP7_75t_SL g6807 ( 
.A(n_5504),
.B(n_5507),
.Y(n_6807)
);

AND2x2_ASAP7_75t_L g6808 ( 
.A(n_5636),
.B(n_5640),
.Y(n_6808)
);

CKINVDCx16_ASAP7_75t_R g6809 ( 
.A(n_4666),
.Y(n_6809)
);

AOI21x1_ASAP7_75t_L g6810 ( 
.A1(n_5048),
.A2(n_5105),
.B(n_5056),
.Y(n_6810)
);

AOI21x1_ASAP7_75t_L g6811 ( 
.A1(n_5048),
.A2(n_5105),
.B(n_5056),
.Y(n_6811)
);

NAND2xp5_ASAP7_75t_SL g6812 ( 
.A(n_5504),
.B(n_5507),
.Y(n_6812)
);

BUFx8_ASAP7_75t_SL g6813 ( 
.A(n_4666),
.Y(n_6813)
);

NOR2xp33_ASAP7_75t_L g6814 ( 
.A(n_5208),
.B(n_5209),
.Y(n_6814)
);

NAND2xp5_ASAP7_75t_L g6815 ( 
.A(n_5599),
.B(n_5625),
.Y(n_6815)
);

OAI21xp33_ASAP7_75t_SL g6816 ( 
.A1(n_4952),
.A2(n_5061),
.B(n_4967),
.Y(n_6816)
);

OAI22xp5_ASAP7_75t_L g6817 ( 
.A1(n_4714),
.A2(n_4774),
.B1(n_4945),
.B2(n_4718),
.Y(n_6817)
);

INVxp67_ASAP7_75t_SL g6818 ( 
.A(n_4571),
.Y(n_6818)
);

CKINVDCx8_ASAP7_75t_R g6819 ( 
.A(n_5374),
.Y(n_6819)
);

INVx1_ASAP7_75t_SL g6820 ( 
.A(n_5148),
.Y(n_6820)
);

AOI22xp33_ASAP7_75t_SL g6821 ( 
.A1(n_4576),
.A2(n_4661),
.B1(n_4876),
.B2(n_4717),
.Y(n_6821)
);

NOR2xp33_ASAP7_75t_L g6822 ( 
.A(n_5209),
.B(n_5229),
.Y(n_6822)
);

O2A1O1Ixp33_ASAP7_75t_L g6823 ( 
.A1(n_4718),
.A2(n_4945),
.B(n_4774),
.C(n_5630),
.Y(n_6823)
);

NOR2xp33_ASAP7_75t_L g6824 ( 
.A(n_5229),
.B(n_5248),
.Y(n_6824)
);

O2A1O1Ixp5_ASAP7_75t_SL g6825 ( 
.A1(n_5638),
.A2(n_5657),
.B(n_5649),
.C(n_5125),
.Y(n_6825)
);

INVx3_ASAP7_75t_L g6826 ( 
.A(n_5008),
.Y(n_6826)
);

INVx1_ASAP7_75t_SL g6827 ( 
.A(n_5264),
.Y(n_6827)
);

OAI22xp5_ASAP7_75t_L g6828 ( 
.A1(n_4745),
.A2(n_4620),
.B1(n_4811),
.B2(n_4596),
.Y(n_6828)
);

NAND2x1_ASAP7_75t_L g6829 ( 
.A(n_5035),
.B(n_5140),
.Y(n_6829)
);

AOI22xp33_ASAP7_75t_L g6830 ( 
.A1(n_4717),
.A2(n_4876),
.B1(n_5737),
.B2(n_4595),
.Y(n_6830)
);

CKINVDCx20_ASAP7_75t_R g6831 ( 
.A(n_4963),
.Y(n_6831)
);

INVx1_ASAP7_75t_SL g6832 ( 
.A(n_5668),
.Y(n_6832)
);

AND2x4_ASAP7_75t_L g6833 ( 
.A(n_5008),
.B(n_5019),
.Y(n_6833)
);

AOI21x1_ASAP7_75t_L g6834 ( 
.A1(n_5109),
.A2(n_5214),
.B(n_5115),
.Y(n_6834)
);

OAI22xp5_ASAP7_75t_L g6835 ( 
.A1(n_4596),
.A2(n_4811),
.B1(n_4893),
.B2(n_4620),
.Y(n_6835)
);

AOI22xp5_ASAP7_75t_L g6836 ( 
.A1(n_5744),
.A2(n_5123),
.B1(n_4876),
.B2(n_5330),
.Y(n_6836)
);

AND2x2_ASAP7_75t_L g6837 ( 
.A(n_5636),
.B(n_5640),
.Y(n_6837)
);

NAND2xp5_ASAP7_75t_R g6838 ( 
.A(n_4659),
.B(n_5636),
.Y(n_6838)
);

NAND2xp5_ASAP7_75t_SL g6839 ( 
.A(n_4576),
.B(n_4661),
.Y(n_6839)
);

OAI22xp5_ASAP7_75t_L g6840 ( 
.A1(n_4893),
.A2(n_4977),
.B1(n_5031),
.B2(n_4926),
.Y(n_6840)
);

INVx1_ASAP7_75t_SL g6841 ( 
.A(n_5668),
.Y(n_6841)
);

OAI22xp5_ASAP7_75t_L g6842 ( 
.A1(n_4926),
.A2(n_5031),
.B1(n_5145),
.B2(n_4977),
.Y(n_6842)
);

INVx5_ASAP7_75t_L g6843 ( 
.A(n_5030),
.Y(n_6843)
);

AOI22xp5_ASAP7_75t_L g6844 ( 
.A1(n_5123),
.A2(n_5330),
.B1(n_5248),
.B2(n_5304),
.Y(n_6844)
);

OAI22xp33_ASAP7_75t_L g6845 ( 
.A1(n_4576),
.A2(n_4661),
.B1(n_4830),
.B2(n_5745),
.Y(n_6845)
);

AOI22xp5_ASAP7_75t_L g6846 ( 
.A1(n_5229),
.A2(n_5304),
.B1(n_5305),
.B2(n_5248),
.Y(n_6846)
);

HB1xp67_ASAP7_75t_L g6847 ( 
.A(n_5292),
.Y(n_6847)
);

NOR2xp67_ASAP7_75t_L g6848 ( 
.A(n_5019),
.B(n_5121),
.Y(n_6848)
);

INVx3_ASAP7_75t_L g6849 ( 
.A(n_5019),
.Y(n_6849)
);

OAI22xp33_ASAP7_75t_L g6850 ( 
.A1(n_4576),
.A2(n_4661),
.B1(n_5745),
.B2(n_5521),
.Y(n_6850)
);

BUFx12f_ASAP7_75t_L g6851 ( 
.A(n_5628),
.Y(n_6851)
);

NOR2xp33_ASAP7_75t_L g6852 ( 
.A(n_5304),
.B(n_5305),
.Y(n_6852)
);

AO22x1_ASAP7_75t_L g6853 ( 
.A1(n_5035),
.A2(n_5523),
.B1(n_5534),
.B2(n_5140),
.Y(n_6853)
);

A2O1A1Ixp33_ASAP7_75t_L g6854 ( 
.A1(n_5490),
.A2(n_5471),
.B(n_4623),
.C(n_4685),
.Y(n_6854)
);

AND2x2_ASAP7_75t_L g6855 ( 
.A(n_5640),
.B(n_5645),
.Y(n_6855)
);

AOI21xp5_ASAP7_75t_L g6856 ( 
.A1(n_5376),
.A2(n_5480),
.B(n_5434),
.Y(n_6856)
);

OAI22xp5_ASAP7_75t_L g6857 ( 
.A1(n_5145),
.A2(n_5321),
.B1(n_5163),
.B2(n_5098),
.Y(n_6857)
);

INVx6_ASAP7_75t_L g6858 ( 
.A(n_4674),
.Y(n_6858)
);

A2O1A1Ixp33_ASAP7_75t_L g6859 ( 
.A1(n_5471),
.A2(n_4623),
.B(n_4685),
.C(n_4603),
.Y(n_6859)
);

AND2x2_ASAP7_75t_L g6860 ( 
.A(n_5645),
.B(n_4608),
.Y(n_6860)
);

BUFx12f_ASAP7_75t_L g6861 ( 
.A(n_5628),
.Y(n_6861)
);

INVx5_ASAP7_75t_L g6862 ( 
.A(n_5030),
.Y(n_6862)
);

AND2x2_ASAP7_75t_L g6863 ( 
.A(n_5645),
.B(n_4608),
.Y(n_6863)
);

AOI22xp33_ASAP7_75t_L g6864 ( 
.A1(n_5737),
.A2(n_5668),
.B1(n_4721),
.B2(n_5658),
.Y(n_6864)
);

NOR2xp67_ASAP7_75t_SL g6865 ( 
.A(n_4789),
.B(n_4884),
.Y(n_6865)
);

OAI22xp5_ASAP7_75t_L g6866 ( 
.A1(n_5163),
.A2(n_5321),
.B1(n_5098),
.B2(n_5107),
.Y(n_6866)
);

INVxp67_ASAP7_75t_L g6867 ( 
.A(n_5672),
.Y(n_6867)
);

CKINVDCx8_ASAP7_75t_R g6868 ( 
.A(n_5374),
.Y(n_6868)
);

AOI21x1_ASAP7_75t_L g6869 ( 
.A1(n_5109),
.A2(n_5214),
.B(n_5115),
.Y(n_6869)
);

O2A1O1Ixp33_ASAP7_75t_L g6870 ( 
.A1(n_5672),
.A2(n_5697),
.B(n_5713),
.C(n_5737),
.Y(n_6870)
);

AOI21xp5_ASAP7_75t_L g6871 ( 
.A1(n_5434),
.A2(n_5512),
.B(n_5480),
.Y(n_6871)
);

INVx4_ASAP7_75t_L g6872 ( 
.A(n_4800),
.Y(n_6872)
);

BUFx8_ASAP7_75t_L g6873 ( 
.A(n_4800),
.Y(n_6873)
);

OAI21xp5_ASAP7_75t_L g6874 ( 
.A1(n_5566),
.A2(n_5747),
.B(n_5688),
.Y(n_6874)
);

AOI21xp5_ASAP7_75t_L g6875 ( 
.A1(n_5434),
.A2(n_5512),
.B(n_5480),
.Y(n_6875)
);

A2O1A1Ixp33_ASAP7_75t_L g6876 ( 
.A1(n_4603),
.A2(n_4685),
.B(n_4623),
.C(n_5223),
.Y(n_6876)
);

CKINVDCx8_ASAP7_75t_R g6877 ( 
.A(n_5374),
.Y(n_6877)
);

CKINVDCx5p33_ASAP7_75t_R g6878 ( 
.A(n_5556),
.Y(n_6878)
);

NOR2x1_ASAP7_75t_SL g6879 ( 
.A(n_5682),
.B(n_5317),
.Y(n_6879)
);

NOR2xp33_ASAP7_75t_L g6880 ( 
.A(n_5305),
.B(n_5311),
.Y(n_6880)
);

AOI21xp5_ASAP7_75t_L g6881 ( 
.A1(n_5434),
.A2(n_5512),
.B(n_5480),
.Y(n_6881)
);

OAI22xp5_ASAP7_75t_L g6882 ( 
.A1(n_5065),
.A2(n_5107),
.B1(n_5169),
.B2(n_5098),
.Y(n_6882)
);

INVx5_ASAP7_75t_L g6883 ( 
.A(n_5030),
.Y(n_6883)
);

NOR2xp67_ASAP7_75t_L g6884 ( 
.A(n_5121),
.B(n_5125),
.Y(n_6884)
);

INVx1_ASAP7_75t_SL g6885 ( 
.A(n_5646),
.Y(n_6885)
);

AOI21xp5_ASAP7_75t_L g6886 ( 
.A1(n_5434),
.A2(n_5512),
.B(n_5480),
.Y(n_6886)
);

BUFx3_ASAP7_75t_L g6887 ( 
.A(n_5034),
.Y(n_6887)
);

AOI21xp5_ASAP7_75t_L g6888 ( 
.A1(n_5434),
.A2(n_5512),
.B(n_5480),
.Y(n_6888)
);

OAI21xp5_ASAP7_75t_L g6889 ( 
.A1(n_5566),
.A2(n_5747),
.B(n_5688),
.Y(n_6889)
);

BUFx8_ASAP7_75t_L g6890 ( 
.A(n_4819),
.Y(n_6890)
);

AO22x1_ASAP7_75t_L g6891 ( 
.A1(n_5035),
.A2(n_5523),
.B1(n_5534),
.B2(n_5140),
.Y(n_6891)
);

AOI21xp5_ASAP7_75t_L g6892 ( 
.A1(n_5512),
.A2(n_5593),
.B(n_5584),
.Y(n_6892)
);

CKINVDCx20_ASAP7_75t_R g6893 ( 
.A(n_5556),
.Y(n_6893)
);

NOR2xp33_ASAP7_75t_L g6894 ( 
.A(n_5311),
.B(n_5324),
.Y(n_6894)
);

INVx3_ASAP7_75t_L g6895 ( 
.A(n_5024),
.Y(n_6895)
);

OAI21xp5_ASAP7_75t_L g6896 ( 
.A1(n_5686),
.A2(n_5691),
.B(n_5688),
.Y(n_6896)
);

O2A1O1Ixp5_ASAP7_75t_L g6897 ( 
.A1(n_5110),
.A2(n_5135),
.B(n_5223),
.C(n_5473),
.Y(n_6897)
);

INVx3_ASAP7_75t_L g6898 ( 
.A(n_5024),
.Y(n_6898)
);

AO21x2_ASAP7_75t_L g6899 ( 
.A1(n_5578),
.A2(n_4610),
.B(n_4591),
.Y(n_6899)
);

CKINVDCx5p33_ASAP7_75t_R g6900 ( 
.A(n_5276),
.Y(n_6900)
);

A2O1A1Ixp33_ASAP7_75t_L g6901 ( 
.A1(n_4603),
.A2(n_4685),
.B(n_4623),
.C(n_5223),
.Y(n_6901)
);

OR2x6_ASAP7_75t_L g6902 ( 
.A(n_4732),
.B(n_4763),
.Y(n_6902)
);

NAND2xp5_ASAP7_75t_SL g6903 ( 
.A(n_5223),
.B(n_4603),
.Y(n_6903)
);

AND2x2_ASAP7_75t_L g6904 ( 
.A(n_4586),
.B(n_4591),
.Y(n_6904)
);

INVx3_ASAP7_75t_L g6905 ( 
.A(n_5024),
.Y(n_6905)
);

BUFx6f_ASAP7_75t_L g6906 ( 
.A(n_4819),
.Y(n_6906)
);

AND2x2_ASAP7_75t_L g6907 ( 
.A(n_6808),
.B(n_6837),
.Y(n_6907)
);

INVx1_ASAP7_75t_L g6908 ( 
.A(n_5777),
.Y(n_6908)
);

OAI21xp33_ASAP7_75t_L g6909 ( 
.A1(n_5880),
.A2(n_4931),
.B(n_5065),
.Y(n_6909)
);

OAI22xp5_ASAP7_75t_L g6910 ( 
.A1(n_5987),
.A2(n_5745),
.B1(n_5474),
.B2(n_5497),
.Y(n_6910)
);

INVx1_ASAP7_75t_SL g6911 ( 
.A(n_6180),
.Y(n_6911)
);

AND2x2_ASAP7_75t_L g6912 ( 
.A(n_6808),
.B(n_4586),
.Y(n_6912)
);

INVx5_ASAP7_75t_L g6913 ( 
.A(n_6030),
.Y(n_6913)
);

INVx3_ASAP7_75t_L g6914 ( 
.A(n_6016),
.Y(n_6914)
);

INVx2_ASAP7_75t_SL g6915 ( 
.A(n_6654),
.Y(n_6915)
);

BUFx6f_ASAP7_75t_L g6916 ( 
.A(n_5860),
.Y(n_6916)
);

AOI21xp5_ASAP7_75t_L g6917 ( 
.A1(n_5911),
.A2(n_5593),
.B(n_5584),
.Y(n_6917)
);

OAI21x1_ASAP7_75t_L g6918 ( 
.A1(n_6060),
.A2(n_5241),
.B(n_4995),
.Y(n_6918)
);

INVx2_ASAP7_75t_SL g6919 ( 
.A(n_6654),
.Y(n_6919)
);

INVx3_ASAP7_75t_SL g6920 ( 
.A(n_5834),
.Y(n_6920)
);

NOR2xp33_ASAP7_75t_SL g6921 ( 
.A(n_6195),
.B(n_5374),
.Y(n_6921)
);

AND2x4_ASAP7_75t_L g6922 ( 
.A(n_6047),
.B(n_5110),
.Y(n_6922)
);

INVx1_ASAP7_75t_L g6923 ( 
.A(n_5777),
.Y(n_6923)
);

INVx5_ASAP7_75t_L g6924 ( 
.A(n_6030),
.Y(n_6924)
);

O2A1O1Ixp5_ASAP7_75t_L g6925 ( 
.A1(n_6221),
.A2(n_5473),
.B(n_5223),
.C(n_5135),
.Y(n_6925)
);

BUFx3_ASAP7_75t_L g6926 ( 
.A(n_6829),
.Y(n_6926)
);

INVx2_ASAP7_75t_SL g6927 ( 
.A(n_6654),
.Y(n_6927)
);

AOI21xp5_ASAP7_75t_L g6928 ( 
.A1(n_5911),
.A2(n_5593),
.B(n_5584),
.Y(n_6928)
);

NAND2xp5_ASAP7_75t_SL g6929 ( 
.A(n_5975),
.B(n_5110),
.Y(n_6929)
);

BUFx3_ASAP7_75t_L g6930 ( 
.A(n_6829),
.Y(n_6930)
);

INVx2_ASAP7_75t_L g6931 ( 
.A(n_5764),
.Y(n_6931)
);

NOR2xp33_ASAP7_75t_L g6932 ( 
.A(n_5985),
.B(n_5311),
.Y(n_6932)
);

INVx2_ASAP7_75t_SL g6933 ( 
.A(n_6654),
.Y(n_6933)
);

NAND2xp33_ASAP7_75t_L g6934 ( 
.A(n_5975),
.B(n_4931),
.Y(n_6934)
);

INVx2_ASAP7_75t_SL g6935 ( 
.A(n_6654),
.Y(n_6935)
);

AND2x2_ASAP7_75t_L g6936 ( 
.A(n_6808),
.B(n_4586),
.Y(n_6936)
);

INVx3_ASAP7_75t_L g6937 ( 
.A(n_6016),
.Y(n_6937)
);

AND2x4_ASAP7_75t_L g6938 ( 
.A(n_6047),
.B(n_5135),
.Y(n_6938)
);

AOI22xp33_ASAP7_75t_L g6939 ( 
.A1(n_5880),
.A2(n_5348),
.B1(n_5403),
.B2(n_5324),
.Y(n_6939)
);

BUFx6f_ASAP7_75t_L g6940 ( 
.A(n_5860),
.Y(n_6940)
);

INVx2_ASAP7_75t_L g6941 ( 
.A(n_5764),
.Y(n_6941)
);

INVx1_ASAP7_75t_L g6942 ( 
.A(n_5781),
.Y(n_6942)
);

AOI22xp5_ASAP7_75t_L g6943 ( 
.A1(n_6070),
.A2(n_5324),
.B1(n_5403),
.B2(n_5348),
.Y(n_6943)
);

INVx1_ASAP7_75t_L g6944 ( 
.A(n_5781),
.Y(n_6944)
);

AND2x4_ASAP7_75t_L g6945 ( 
.A(n_6047),
.B(n_5110),
.Y(n_6945)
);

OR2x6_ASAP7_75t_L g6946 ( 
.A(n_5993),
.B(n_5584),
.Y(n_6946)
);

AND3x1_ASAP7_75t_SL g6947 ( 
.A(n_5797),
.B(n_5276),
.C(n_4738),
.Y(n_6947)
);

AND2x4_ASAP7_75t_L g6948 ( 
.A(n_6047),
.B(n_5110),
.Y(n_6948)
);

BUFx6f_ASAP7_75t_L g6949 ( 
.A(n_5860),
.Y(n_6949)
);

INVx3_ASAP7_75t_L g6950 ( 
.A(n_6016),
.Y(n_6950)
);

CKINVDCx20_ASAP7_75t_R g6951 ( 
.A(n_5817),
.Y(n_6951)
);

AOI22xp33_ASAP7_75t_L g6952 ( 
.A1(n_6070),
.A2(n_5403),
.B1(n_5439),
.B2(n_5348),
.Y(n_6952)
);

INVx2_ASAP7_75t_L g6953 ( 
.A(n_5764),
.Y(n_6953)
);

INVx1_ASAP7_75t_L g6954 ( 
.A(n_5785),
.Y(n_6954)
);

NAND2xp5_ASAP7_75t_L g6955 ( 
.A(n_6748),
.B(n_5223),
.Y(n_6955)
);

INVxp67_ASAP7_75t_L g6956 ( 
.A(n_6748),
.Y(n_6956)
);

INVx3_ASAP7_75t_L g6957 ( 
.A(n_6016),
.Y(n_6957)
);

OAI22xp33_ASAP7_75t_L g6958 ( 
.A1(n_5783),
.A2(n_5474),
.B1(n_5497),
.B2(n_5413),
.Y(n_6958)
);

NAND2xp5_ASAP7_75t_L g6959 ( 
.A(n_6647),
.B(n_6208),
.Y(n_6959)
);

BUFx6f_ASAP7_75t_L g6960 ( 
.A(n_5860),
.Y(n_6960)
);

BUFx3_ASAP7_75t_L g6961 ( 
.A(n_5948),
.Y(n_6961)
);

INVx2_ASAP7_75t_L g6962 ( 
.A(n_5773),
.Y(n_6962)
);

BUFx3_ASAP7_75t_L g6963 ( 
.A(n_5948),
.Y(n_6963)
);

OR2x2_ASAP7_75t_L g6964 ( 
.A(n_6049),
.B(n_6142),
.Y(n_6964)
);

INVxp67_ASAP7_75t_SL g6965 ( 
.A(n_6598),
.Y(n_6965)
);

AO32x1_ASAP7_75t_L g6966 ( 
.A1(n_6031),
.A2(n_4952),
.A3(n_5104),
.B1(n_5061),
.B2(n_4967),
.Y(n_6966)
);

NOR2xp33_ASAP7_75t_L g6967 ( 
.A(n_5985),
.B(n_5439),
.Y(n_6967)
);

NAND2xp5_ASAP7_75t_L g6968 ( 
.A(n_6647),
.B(n_5110),
.Y(n_6968)
);

OAI22xp33_ASAP7_75t_L g6969 ( 
.A1(n_5783),
.A2(n_5497),
.B1(n_5413),
.B2(n_5521),
.Y(n_6969)
);

AOI22xp5_ASAP7_75t_L g6970 ( 
.A1(n_6002),
.A2(n_5439),
.B1(n_5454),
.B2(n_5444),
.Y(n_6970)
);

AOI22xp33_ASAP7_75t_L g6971 ( 
.A1(n_5797),
.A2(n_5454),
.B1(n_5457),
.B2(n_5444),
.Y(n_6971)
);

AOI22x1_ASAP7_75t_L g6972 ( 
.A1(n_6081),
.A2(n_5508),
.B1(n_5317),
.B2(n_4670),
.Y(n_6972)
);

BUFx6f_ASAP7_75t_L g6973 ( 
.A(n_5860),
.Y(n_6973)
);

INVx2_ASAP7_75t_SL g6974 ( 
.A(n_6678),
.Y(n_6974)
);

INVx2_ASAP7_75t_L g6975 ( 
.A(n_5773),
.Y(n_6975)
);

AOI21xp5_ASAP7_75t_L g6976 ( 
.A1(n_5998),
.A2(n_5593),
.B(n_5584),
.Y(n_6976)
);

INVx5_ASAP7_75t_L g6977 ( 
.A(n_6030),
.Y(n_6977)
);

OAI21xp5_ASAP7_75t_L g6978 ( 
.A1(n_5999),
.A2(n_5593),
.B(n_5584),
.Y(n_6978)
);

BUFx3_ASAP7_75t_L g6979 ( 
.A(n_5948),
.Y(n_6979)
);

INVx2_ASAP7_75t_L g6980 ( 
.A(n_5773),
.Y(n_6980)
);

BUFx6f_ASAP7_75t_L g6981 ( 
.A(n_5860),
.Y(n_6981)
);

NAND2xp5_ASAP7_75t_SL g6982 ( 
.A(n_6195),
.B(n_5135),
.Y(n_6982)
);

INVx2_ASAP7_75t_L g6983 ( 
.A(n_5798),
.Y(n_6983)
);

BUFx2_ASAP7_75t_L g6984 ( 
.A(n_6188),
.Y(n_6984)
);

NOR2xp33_ASAP7_75t_L g6985 ( 
.A(n_6006),
.B(n_5444),
.Y(n_6985)
);

INVx1_ASAP7_75t_SL g6986 ( 
.A(n_6180),
.Y(n_6986)
);

AOI21xp5_ASAP7_75t_L g6987 ( 
.A1(n_5998),
.A2(n_5613),
.B(n_5593),
.Y(n_6987)
);

INVx2_ASAP7_75t_L g6988 ( 
.A(n_5798),
.Y(n_6988)
);

NAND2xp5_ASAP7_75t_L g6989 ( 
.A(n_6208),
.B(n_5819),
.Y(n_6989)
);

AND2x2_ASAP7_75t_SL g6990 ( 
.A(n_5766),
.B(n_5613),
.Y(n_6990)
);

AND2x4_ASAP7_75t_L g6991 ( 
.A(n_6047),
.B(n_5135),
.Y(n_6991)
);

NAND2xp5_ASAP7_75t_L g6992 ( 
.A(n_5819),
.B(n_6061),
.Y(n_6992)
);

NOR2xp33_ASAP7_75t_L g6993 ( 
.A(n_6006),
.B(n_5454),
.Y(n_6993)
);

INVx5_ASAP7_75t_L g6994 ( 
.A(n_6030),
.Y(n_6994)
);

AOI21x1_ASAP7_75t_L g6995 ( 
.A1(n_6255),
.A2(n_5273),
.B(n_5220),
.Y(n_6995)
);

AND2x4_ASAP7_75t_L g6996 ( 
.A(n_6052),
.B(n_5135),
.Y(n_6996)
);

AND2x2_ASAP7_75t_L g6997 ( 
.A(n_6837),
.B(n_4604),
.Y(n_6997)
);

AOI22xp33_ASAP7_75t_L g6998 ( 
.A1(n_6002),
.A2(n_5459),
.B1(n_5487),
.B2(n_5457),
.Y(n_6998)
);

INVx4_ASAP7_75t_L g6999 ( 
.A(n_6902),
.Y(n_6999)
);

CKINVDCx5p33_ASAP7_75t_R g7000 ( 
.A(n_6011),
.Y(n_7000)
);

INVx2_ASAP7_75t_L g7001 ( 
.A(n_5798),
.Y(n_7001)
);

NAND2xp5_ASAP7_75t_SL g7002 ( 
.A(n_6097),
.B(n_5024),
.Y(n_7002)
);

INVx4_ASAP7_75t_L g7003 ( 
.A(n_6902),
.Y(n_7003)
);

OAI22xp5_ASAP7_75t_SL g7004 ( 
.A1(n_6174),
.A2(n_4915),
.B1(n_4924),
.B2(n_4884),
.Y(n_7004)
);

AOI22xp33_ASAP7_75t_L g7005 ( 
.A1(n_5981),
.A2(n_5459),
.B1(n_5487),
.B2(n_5457),
.Y(n_7005)
);

INVx2_ASAP7_75t_L g7006 ( 
.A(n_5809),
.Y(n_7006)
);

AOI21xp5_ASAP7_75t_L g7007 ( 
.A1(n_6000),
.A2(n_5615),
.B(n_5613),
.Y(n_7007)
);

AND2x2_ASAP7_75t_L g7008 ( 
.A(n_6837),
.B(n_6855),
.Y(n_7008)
);

BUFx12f_ASAP7_75t_L g7009 ( 
.A(n_6851),
.Y(n_7009)
);

BUFx3_ASAP7_75t_L g7010 ( 
.A(n_5948),
.Y(n_7010)
);

NOR2xp33_ASAP7_75t_L g7011 ( 
.A(n_6094),
.B(n_5459),
.Y(n_7011)
);

OAI21xp33_ASAP7_75t_L g7012 ( 
.A1(n_5981),
.A2(n_5098),
.B(n_5065),
.Y(n_7012)
);

CKINVDCx6p67_ASAP7_75t_R g7013 ( 
.A(n_5834),
.Y(n_7013)
);

BUFx6f_ASAP7_75t_L g7014 ( 
.A(n_5860),
.Y(n_7014)
);

INVx2_ASAP7_75t_L g7015 ( 
.A(n_5809),
.Y(n_7015)
);

AOI21xp33_ASAP7_75t_SL g7016 ( 
.A1(n_5999),
.A2(n_4924),
.B(n_4915),
.Y(n_7016)
);

AOI221xp5_ASAP7_75t_L g7017 ( 
.A1(n_6071),
.A2(n_5574),
.B1(n_5572),
.B2(n_5658),
.C(n_5268),
.Y(n_7017)
);

BUFx6f_ASAP7_75t_L g7018 ( 
.A(n_5860),
.Y(n_7018)
);

OR2x6_ASAP7_75t_L g7019 ( 
.A(n_5993),
.B(n_5613),
.Y(n_7019)
);

BUFx6f_ASAP7_75t_L g7020 ( 
.A(n_5889),
.Y(n_7020)
);

NOR3xp33_ASAP7_75t_L g7021 ( 
.A(n_5990),
.B(n_5759),
.C(n_5754),
.Y(n_7021)
);

NOR2xp33_ASAP7_75t_L g7022 ( 
.A(n_6094),
.B(n_6042),
.Y(n_7022)
);

O2A1O1Ixp5_ASAP7_75t_L g7023 ( 
.A1(n_6221),
.A2(n_4623),
.B(n_4685),
.C(n_4603),
.Y(n_7023)
);

AOI21xp5_ASAP7_75t_L g7024 ( 
.A1(n_6000),
.A2(n_5615),
.B(n_5613),
.Y(n_7024)
);

OAI22xp5_ASAP7_75t_L g7025 ( 
.A1(n_5987),
.A2(n_5107),
.B1(n_5169),
.B2(n_5065),
.Y(n_7025)
);

NOR2xp33_ASAP7_75t_L g7026 ( 
.A(n_6042),
.B(n_5487),
.Y(n_7026)
);

NAND2xp5_ASAP7_75t_L g7027 ( 
.A(n_6061),
.B(n_5259),
.Y(n_7027)
);

AND2x4_ASAP7_75t_L g7028 ( 
.A(n_6052),
.B(n_5024),
.Y(n_7028)
);

AND2x4_ASAP7_75t_L g7029 ( 
.A(n_6052),
.B(n_5024),
.Y(n_7029)
);

INVx1_ASAP7_75t_SL g7030 ( 
.A(n_6008),
.Y(n_7030)
);

BUFx3_ASAP7_75t_L g7031 ( 
.A(n_5948),
.Y(n_7031)
);

AOI21xp33_ASAP7_75t_L g7032 ( 
.A1(n_6081),
.A2(n_5615),
.B(n_5613),
.Y(n_7032)
);

CKINVDCx5p33_ASAP7_75t_R g7033 ( 
.A(n_6011),
.Y(n_7033)
);

AOI21xp5_ASAP7_75t_L g7034 ( 
.A1(n_6088),
.A2(n_5653),
.B(n_5615),
.Y(n_7034)
);

A2O1A1Ixp33_ASAP7_75t_SL g7035 ( 
.A1(n_5990),
.A2(n_5589),
.B(n_5393),
.C(n_5725),
.Y(n_7035)
);

INVx1_ASAP7_75t_SL g7036 ( 
.A(n_6008),
.Y(n_7036)
);

NAND2xp5_ASAP7_75t_L g7037 ( 
.A(n_5962),
.B(n_6044),
.Y(n_7037)
);

NAND2xp5_ASAP7_75t_L g7038 ( 
.A(n_5962),
.B(n_5259),
.Y(n_7038)
);

AND2x2_ASAP7_75t_L g7039 ( 
.A(n_6855),
.B(n_4604),
.Y(n_7039)
);

INVx4_ASAP7_75t_L g7040 ( 
.A(n_6902),
.Y(n_7040)
);

INVx2_ASAP7_75t_SL g7041 ( 
.A(n_6678),
.Y(n_7041)
);

INVx2_ASAP7_75t_L g7042 ( 
.A(n_5809),
.Y(n_7042)
);

INVx6_ASAP7_75t_L g7043 ( 
.A(n_6460),
.Y(n_7043)
);

BUFx4f_ASAP7_75t_L g7044 ( 
.A(n_5766),
.Y(n_7044)
);

INVx4_ASAP7_75t_L g7045 ( 
.A(n_6902),
.Y(n_7045)
);

INVx4_ASAP7_75t_L g7046 ( 
.A(n_6902),
.Y(n_7046)
);

CKINVDCx8_ASAP7_75t_R g7047 ( 
.A(n_6111),
.Y(n_7047)
);

BUFx4f_ASAP7_75t_SL g7048 ( 
.A(n_5873),
.Y(n_7048)
);

BUFx2_ASAP7_75t_L g7049 ( 
.A(n_6188),
.Y(n_7049)
);

BUFx6f_ASAP7_75t_L g7050 ( 
.A(n_5889),
.Y(n_7050)
);

BUFx4f_ASAP7_75t_L g7051 ( 
.A(n_5766),
.Y(n_7051)
);

AOI21xp33_ASAP7_75t_L g7052 ( 
.A1(n_5997),
.A2(n_6033),
.B(n_6110),
.Y(n_7052)
);

INVxp67_ASAP7_75t_L g7053 ( 
.A(n_5800),
.Y(n_7053)
);

INVx2_ASAP7_75t_L g7054 ( 
.A(n_5833),
.Y(n_7054)
);

INVx1_ASAP7_75t_SL g7055 ( 
.A(n_6142),
.Y(n_7055)
);

AND2x2_ASAP7_75t_L g7056 ( 
.A(n_6855),
.B(n_4606),
.Y(n_7056)
);

AOI22xp5_ASAP7_75t_L g7057 ( 
.A1(n_6048),
.A2(n_5658),
.B1(n_5468),
.B2(n_5034),
.Y(n_7057)
);

INVx2_ASAP7_75t_SL g7058 ( 
.A(n_6678),
.Y(n_7058)
);

NOR2xp33_ASAP7_75t_L g7059 ( 
.A(n_5977),
.B(n_5468),
.Y(n_7059)
);

INVx3_ASAP7_75t_SL g7060 ( 
.A(n_5834),
.Y(n_7060)
);

INVx2_ASAP7_75t_L g7061 ( 
.A(n_5833),
.Y(n_7061)
);

AOI22xp33_ASAP7_75t_L g7062 ( 
.A1(n_6048),
.A2(n_5653),
.B1(n_5615),
.B2(n_5169),
.Y(n_7062)
);

OR2x6_ASAP7_75t_L g7063 ( 
.A(n_5993),
.B(n_5615),
.Y(n_7063)
);

A2O1A1Ixp33_ASAP7_75t_L g7064 ( 
.A1(n_6110),
.A2(n_5703),
.B(n_5450),
.C(n_4804),
.Y(n_7064)
);

BUFx6f_ASAP7_75t_L g7065 ( 
.A(n_5889),
.Y(n_7065)
);

NAND2xp5_ASAP7_75t_SL g7066 ( 
.A(n_6097),
.B(n_5335),
.Y(n_7066)
);

HB1xp67_ASAP7_75t_L g7067 ( 
.A(n_5800),
.Y(n_7067)
);

INVx2_ASAP7_75t_L g7068 ( 
.A(n_5833),
.Y(n_7068)
);

BUFx2_ASAP7_75t_L g7069 ( 
.A(n_6188),
.Y(n_7069)
);

NAND2xp5_ASAP7_75t_L g7070 ( 
.A(n_6044),
.B(n_5269),
.Y(n_7070)
);

AOI22xp33_ASAP7_75t_L g7071 ( 
.A1(n_6071),
.A2(n_6091),
.B1(n_6075),
.B2(n_6103),
.Y(n_7071)
);

INVx2_ASAP7_75t_L g7072 ( 
.A(n_5854),
.Y(n_7072)
);

NAND2xp5_ASAP7_75t_L g7073 ( 
.A(n_6613),
.B(n_6590),
.Y(n_7073)
);

BUFx2_ASAP7_75t_L g7074 ( 
.A(n_6188),
.Y(n_7074)
);

AOI22xp5_ASAP7_75t_L g7075 ( 
.A1(n_6103),
.A2(n_5468),
.B1(n_5034),
.B2(n_5418),
.Y(n_7075)
);

INVx2_ASAP7_75t_L g7076 ( 
.A(n_5854),
.Y(n_7076)
);

INVx2_ASAP7_75t_SL g7077 ( 
.A(n_6678),
.Y(n_7077)
);

AND2x2_ASAP7_75t_L g7078 ( 
.A(n_6860),
.B(n_6863),
.Y(n_7078)
);

BUFx8_ASAP7_75t_L g7079 ( 
.A(n_6126),
.Y(n_7079)
);

AOI21xp5_ASAP7_75t_L g7080 ( 
.A1(n_6088),
.A2(n_5653),
.B(n_5281),
.Y(n_7080)
);

BUFx2_ASAP7_75t_L g7081 ( 
.A(n_6188),
.Y(n_7081)
);

AOI21xp5_ASAP7_75t_L g7082 ( 
.A1(n_6101),
.A2(n_5653),
.B(n_5281),
.Y(n_7082)
);

INVx2_ASAP7_75t_L g7083 ( 
.A(n_5854),
.Y(n_7083)
);

NAND2xp5_ASAP7_75t_L g7084 ( 
.A(n_6613),
.B(n_6590),
.Y(n_7084)
);

NAND2xp5_ASAP7_75t_L g7085 ( 
.A(n_6602),
.B(n_5269),
.Y(n_7085)
);

AOI21xp5_ASAP7_75t_L g7086 ( 
.A1(n_6101),
.A2(n_5653),
.B(n_5281),
.Y(n_7086)
);

HB1xp67_ASAP7_75t_L g7087 ( 
.A(n_5874),
.Y(n_7087)
);

OAI221xp5_ASAP7_75t_L g7088 ( 
.A1(n_5997),
.A2(n_4763),
.B1(n_4732),
.B2(n_5521),
.C(n_5505),
.Y(n_7088)
);

NAND2xp5_ASAP7_75t_L g7089 ( 
.A(n_6602),
.B(n_5269),
.Y(n_7089)
);

AOI21xp5_ASAP7_75t_L g7090 ( 
.A1(n_6579),
.A2(n_6673),
.B(n_6580),
.Y(n_7090)
);

AOI22xp33_ASAP7_75t_L g7091 ( 
.A1(n_6075),
.A2(n_5169),
.B1(n_5188),
.B2(n_5107),
.Y(n_7091)
);

OAI221xp5_ASAP7_75t_L g7092 ( 
.A1(n_6033),
.A2(n_6046),
.B1(n_6040),
.B2(n_6091),
.C(n_6092),
.Y(n_7092)
);

NAND2xp5_ASAP7_75t_L g7093 ( 
.A(n_6534),
.B(n_5269),
.Y(n_7093)
);

INVx2_ASAP7_75t_L g7094 ( 
.A(n_5863),
.Y(n_7094)
);

AO32x2_ASAP7_75t_L g7095 ( 
.A1(n_6835),
.A2(n_6842),
.A3(n_6840),
.B1(n_6556),
.B2(n_6551),
.Y(n_7095)
);

AO21x2_ASAP7_75t_L g7096 ( 
.A1(n_6107),
.A2(n_4574),
.B(n_4571),
.Y(n_7096)
);

INVx2_ASAP7_75t_L g7097 ( 
.A(n_5863),
.Y(n_7097)
);

AOI22xp5_ASAP7_75t_L g7098 ( 
.A1(n_5909),
.A2(n_5468),
.B1(n_5034),
.B2(n_5418),
.Y(n_7098)
);

NAND2xp5_ASAP7_75t_L g7099 ( 
.A(n_6534),
.B(n_5270),
.Y(n_7099)
);

AOI21xp5_ASAP7_75t_L g7100 ( 
.A1(n_6579),
.A2(n_5241),
.B(n_4995),
.Y(n_7100)
);

BUFx6f_ASAP7_75t_L g7101 ( 
.A(n_5889),
.Y(n_7101)
);

INVx1_ASAP7_75t_SL g7102 ( 
.A(n_5834),
.Y(n_7102)
);

OAI22xp5_ASAP7_75t_L g7103 ( 
.A1(n_6174),
.A2(n_5255),
.B1(n_5354),
.B2(n_5188),
.Y(n_7103)
);

HB1xp67_ASAP7_75t_L g7104 ( 
.A(n_5874),
.Y(n_7104)
);

CKINVDCx5p33_ASAP7_75t_R g7105 ( 
.A(n_5841),
.Y(n_7105)
);

INVx2_ASAP7_75t_L g7106 ( 
.A(n_5863),
.Y(n_7106)
);

HAxp5_ASAP7_75t_L g7107 ( 
.A(n_6090),
.B(n_4738),
.CON(n_7107),
.SN(n_7107)
);

BUFx2_ASAP7_75t_L g7108 ( 
.A(n_6188),
.Y(n_7108)
);

OR2x6_ASAP7_75t_L g7109 ( 
.A(n_5993),
.B(n_5682),
.Y(n_7109)
);

INVx2_ASAP7_75t_L g7110 ( 
.A(n_5866),
.Y(n_7110)
);

NAND2xp5_ASAP7_75t_L g7111 ( 
.A(n_6427),
.B(n_5270),
.Y(n_7111)
);

BUFx2_ASAP7_75t_L g7112 ( 
.A(n_6299),
.Y(n_7112)
);

OAI22xp33_ASAP7_75t_L g7113 ( 
.A1(n_6068),
.A2(n_5521),
.B1(n_4846),
.B2(n_4854),
.Y(n_7113)
);

INVx2_ASAP7_75t_SL g7114 ( 
.A(n_6678),
.Y(n_7114)
);

INVx1_ASAP7_75t_SL g7115 ( 
.A(n_6885),
.Y(n_7115)
);

NAND2xp5_ASAP7_75t_SL g7116 ( 
.A(n_6040),
.B(n_5335),
.Y(n_7116)
);

BUFx2_ASAP7_75t_L g7117 ( 
.A(n_6299),
.Y(n_7117)
);

AOI22xp5_ASAP7_75t_L g7118 ( 
.A1(n_5909),
.A2(n_5034),
.B1(n_5532),
.B2(n_5505),
.Y(n_7118)
);

INVx2_ASAP7_75t_L g7119 ( 
.A(n_5866),
.Y(n_7119)
);

AND2x4_ASAP7_75t_L g7120 ( 
.A(n_6062),
.B(n_4817),
.Y(n_7120)
);

BUFx8_ASAP7_75t_L g7121 ( 
.A(n_6126),
.Y(n_7121)
);

INVx2_ASAP7_75t_L g7122 ( 
.A(n_5866),
.Y(n_7122)
);

NAND2xp5_ASAP7_75t_L g7123 ( 
.A(n_6427),
.B(n_5270),
.Y(n_7123)
);

OR2x2_ASAP7_75t_L g7124 ( 
.A(n_5976),
.B(n_5986),
.Y(n_7124)
);

NAND2x1p5_ASAP7_75t_L g7125 ( 
.A(n_5889),
.B(n_4670),
.Y(n_7125)
);

NAND2xp5_ASAP7_75t_L g7126 ( 
.A(n_6436),
.B(n_5270),
.Y(n_7126)
);

OAI22xp5_ASAP7_75t_L g7127 ( 
.A1(n_6068),
.A2(n_5255),
.B1(n_5354),
.B2(n_5188),
.Y(n_7127)
);

BUFx8_ASAP7_75t_L g7128 ( 
.A(n_6126),
.Y(n_7128)
);

CKINVDCx5p33_ASAP7_75t_R g7129 ( 
.A(n_5841),
.Y(n_7129)
);

NAND2xp5_ASAP7_75t_L g7130 ( 
.A(n_6436),
.B(n_5274),
.Y(n_7130)
);

INVx2_ASAP7_75t_L g7131 ( 
.A(n_5882),
.Y(n_7131)
);

INVx2_ASAP7_75t_SL g7132 ( 
.A(n_6687),
.Y(n_7132)
);

AND2x4_ASAP7_75t_L g7133 ( 
.A(n_6062),
.B(n_6076),
.Y(n_7133)
);

AO21x2_ASAP7_75t_L g7134 ( 
.A1(n_6107),
.A2(n_6130),
.B(n_6117),
.Y(n_7134)
);

BUFx12f_ASAP7_75t_L g7135 ( 
.A(n_6851),
.Y(n_7135)
);

NOR2xp33_ASAP7_75t_SL g7136 ( 
.A(n_5859),
.B(n_5374),
.Y(n_7136)
);

NAND2xp33_ASAP7_75t_L g7137 ( 
.A(n_6069),
.B(n_4957),
.Y(n_7137)
);

AOI22xp5_ASAP7_75t_L g7138 ( 
.A1(n_6105),
.A2(n_5034),
.B1(n_5562),
.B2(n_5532),
.Y(n_7138)
);

CKINVDCx5p33_ASAP7_75t_R g7139 ( 
.A(n_6112),
.Y(n_7139)
);

O2A1O1Ixp5_ASAP7_75t_SL g7140 ( 
.A1(n_6010),
.A2(n_5125),
.B(n_5121),
.C(n_5686),
.Y(n_7140)
);

BUFx12f_ASAP7_75t_L g7141 ( 
.A(n_6851),
.Y(n_7141)
);

AOI22xp33_ASAP7_75t_SL g7142 ( 
.A1(n_6185),
.A2(n_4935),
.B1(n_4889),
.B2(n_4689),
.Y(n_7142)
);

BUFx3_ASAP7_75t_L g7143 ( 
.A(n_6030),
.Y(n_7143)
);

HB1xp67_ASAP7_75t_L g7144 ( 
.A(n_5884),
.Y(n_7144)
);

INVx2_ASAP7_75t_L g7145 ( 
.A(n_5882),
.Y(n_7145)
);

OAI21xp33_ASAP7_75t_L g7146 ( 
.A1(n_6090),
.A2(n_5255),
.B(n_5188),
.Y(n_7146)
);

INVx2_ASAP7_75t_L g7147 ( 
.A(n_5882),
.Y(n_7147)
);

INVx2_ASAP7_75t_L g7148 ( 
.A(n_5900),
.Y(n_7148)
);

HB1xp67_ASAP7_75t_L g7149 ( 
.A(n_5884),
.Y(n_7149)
);

AND2x4_ASAP7_75t_L g7150 ( 
.A(n_6062),
.B(n_4817),
.Y(n_7150)
);

AOI22xp5_ASAP7_75t_L g7151 ( 
.A1(n_6105),
.A2(n_5034),
.B1(n_5562),
.B2(n_4689),
.Y(n_7151)
);

HB1xp67_ASAP7_75t_L g7152 ( 
.A(n_6201),
.Y(n_7152)
);

BUFx3_ASAP7_75t_L g7153 ( 
.A(n_6030),
.Y(n_7153)
);

INVx2_ASAP7_75t_L g7154 ( 
.A(n_5900),
.Y(n_7154)
);

OAI22xp5_ASAP7_75t_L g7155 ( 
.A1(n_6129),
.A2(n_5255),
.B1(n_5354),
.B2(n_5314),
.Y(n_7155)
);

NAND2xp5_ASAP7_75t_SL g7156 ( 
.A(n_6182),
.B(n_5335),
.Y(n_7156)
);

BUFx2_ASAP7_75t_L g7157 ( 
.A(n_6299),
.Y(n_7157)
);

INVx2_ASAP7_75t_L g7158 ( 
.A(n_5900),
.Y(n_7158)
);

INVx2_ASAP7_75t_L g7159 ( 
.A(n_5903),
.Y(n_7159)
);

BUFx2_ASAP7_75t_L g7160 ( 
.A(n_6299),
.Y(n_7160)
);

AOI21xp5_ASAP7_75t_L g7161 ( 
.A1(n_6580),
.A2(n_6674),
.B(n_6673),
.Y(n_7161)
);

AOI21xp5_ASAP7_75t_L g7162 ( 
.A1(n_6674),
.A2(n_5241),
.B(n_4995),
.Y(n_7162)
);

BUFx2_ASAP7_75t_L g7163 ( 
.A(n_6299),
.Y(n_7163)
);

AOI21xp5_ASAP7_75t_L g7164 ( 
.A1(n_6684),
.A2(n_4995),
.B(n_5686),
.Y(n_7164)
);

BUFx2_ASAP7_75t_L g7165 ( 
.A(n_6299),
.Y(n_7165)
);

INVxp67_ASAP7_75t_SL g7166 ( 
.A(n_6598),
.Y(n_7166)
);

INVx2_ASAP7_75t_SL g7167 ( 
.A(n_6687),
.Y(n_7167)
);

NAND3xp33_ASAP7_75t_L g7168 ( 
.A(n_6046),
.B(n_5691),
.C(n_5697),
.Y(n_7168)
);

AOI21xp33_ASAP7_75t_L g7169 ( 
.A1(n_6054),
.A2(n_5691),
.B(n_5729),
.Y(n_7169)
);

INVx2_ASAP7_75t_SL g7170 ( 
.A(n_6687),
.Y(n_7170)
);

CKINVDCx5p33_ASAP7_75t_R g7171 ( 
.A(n_6112),
.Y(n_7171)
);

A2O1A1Ixp33_ASAP7_75t_L g7172 ( 
.A1(n_6056),
.A2(n_5544),
.B(n_5279),
.C(n_4804),
.Y(n_7172)
);

AOI222xp33_ASAP7_75t_L g7173 ( 
.A1(n_6031),
.A2(n_5090),
.B1(n_5013),
.B2(n_5150),
.C1(n_5022),
.C2(n_4957),
.Y(n_7173)
);

AOI21xp5_ASAP7_75t_L g7174 ( 
.A1(n_6684),
.A2(n_5032),
.B(n_5030),
.Y(n_7174)
);

AOI21xp5_ASAP7_75t_L g7175 ( 
.A1(n_6561),
.A2(n_5032),
.B(n_5030),
.Y(n_7175)
);

INVx8_ASAP7_75t_L g7176 ( 
.A(n_6902),
.Y(n_7176)
);

HB1xp67_ASAP7_75t_L g7177 ( 
.A(n_6201),
.Y(n_7177)
);

INVx1_ASAP7_75t_SL g7178 ( 
.A(n_6885),
.Y(n_7178)
);

INVx2_ASAP7_75t_SL g7179 ( 
.A(n_6687),
.Y(n_7179)
);

OA21x2_ASAP7_75t_L g7180 ( 
.A1(n_6060),
.A2(n_4574),
.B(n_4571),
.Y(n_7180)
);

BUFx2_ASAP7_75t_L g7181 ( 
.A(n_6816),
.Y(n_7181)
);

OAI21xp5_ASAP7_75t_L g7182 ( 
.A1(n_5955),
.A2(n_5729),
.B(n_5762),
.Y(n_7182)
);

INVx2_ASAP7_75t_SL g7183 ( 
.A(n_6687),
.Y(n_7183)
);

INVx2_ASAP7_75t_L g7184 ( 
.A(n_5903),
.Y(n_7184)
);

NAND2xp5_ASAP7_75t_SL g7185 ( 
.A(n_6182),
.B(n_5335),
.Y(n_7185)
);

AND2x4_ASAP7_75t_L g7186 ( 
.A(n_6076),
.B(n_4817),
.Y(n_7186)
);

AOI22xp5_ASAP7_75t_L g7187 ( 
.A1(n_5795),
.A2(n_5034),
.B1(n_4689),
.B2(n_4690),
.Y(n_7187)
);

HB1xp67_ASAP7_75t_L g7188 ( 
.A(n_6246),
.Y(n_7188)
);

AOI22xp33_ASAP7_75t_L g7189 ( 
.A1(n_6248),
.A2(n_5354),
.B1(n_4846),
.B2(n_4854),
.Y(n_7189)
);

NOR2xp33_ASAP7_75t_L g7190 ( 
.A(n_5977),
.B(n_5572),
.Y(n_7190)
);

AOI21xp5_ASAP7_75t_L g7191 ( 
.A1(n_6561),
.A2(n_5032),
.B(n_5030),
.Y(n_7191)
);

INVx2_ASAP7_75t_L g7192 ( 
.A(n_5903),
.Y(n_7192)
);

NAND2xp5_ASAP7_75t_L g7193 ( 
.A(n_6504),
.B(n_5290),
.Y(n_7193)
);

BUFx8_ASAP7_75t_SL g7194 ( 
.A(n_6176),
.Y(n_7194)
);

OAI21x1_ASAP7_75t_L g7195 ( 
.A1(n_6060),
.A2(n_5125),
.B(n_5121),
.Y(n_7195)
);

BUFx2_ASAP7_75t_L g7196 ( 
.A(n_6816),
.Y(n_7196)
);

AOI21xp5_ASAP7_75t_L g7197 ( 
.A1(n_6536),
.A2(n_5032),
.B(n_5030),
.Y(n_7197)
);

AND2x4_ASAP7_75t_L g7198 ( 
.A(n_6076),
.B(n_4817),
.Y(n_7198)
);

NAND2x1p5_ASAP7_75t_L g7199 ( 
.A(n_5951),
.B(n_4670),
.Y(n_7199)
);

AOI22xp33_ASAP7_75t_L g7200 ( 
.A1(n_6248),
.A2(n_4846),
.B1(n_4854),
.B2(n_4819),
.Y(n_7200)
);

HB1xp67_ASAP7_75t_L g7201 ( 
.A(n_6246),
.Y(n_7201)
);

NAND2xp5_ASAP7_75t_L g7202 ( 
.A(n_6504),
.B(n_5290),
.Y(n_7202)
);

OAI21xp5_ASAP7_75t_L g7203 ( 
.A1(n_5955),
.A2(n_5729),
.B(n_5762),
.Y(n_7203)
);

AOI22xp5_ASAP7_75t_L g7204 ( 
.A1(n_5795),
.A2(n_4705),
.B1(n_4720),
.B2(n_4655),
.Y(n_7204)
);

CKINVDCx5p33_ASAP7_75t_R g7205 ( 
.A(n_6176),
.Y(n_7205)
);

NOR2xp33_ASAP7_75t_L g7206 ( 
.A(n_6004),
.B(n_5574),
.Y(n_7206)
);

AND2x4_ASAP7_75t_L g7207 ( 
.A(n_6076),
.B(n_6083),
.Y(n_7207)
);

NAND2xp5_ASAP7_75t_L g7208 ( 
.A(n_6612),
.B(n_5290),
.Y(n_7208)
);

O2A1O1Ixp33_ASAP7_75t_L g7209 ( 
.A1(n_6337),
.A2(n_5713),
.B(n_5754),
.C(n_5753),
.Y(n_7209)
);

BUFx6f_ASAP7_75t_L g7210 ( 
.A(n_5951),
.Y(n_7210)
);

CKINVDCx5p33_ASAP7_75t_R g7211 ( 
.A(n_5817),
.Y(n_7211)
);

NOR2xp33_ASAP7_75t_L g7212 ( 
.A(n_6004),
.B(n_5714),
.Y(n_7212)
);

BUFx2_ASAP7_75t_L g7213 ( 
.A(n_6461),
.Y(n_7213)
);

HB1xp67_ASAP7_75t_L g7214 ( 
.A(n_6307),
.Y(n_7214)
);

INVx2_ASAP7_75t_L g7215 ( 
.A(n_5905),
.Y(n_7215)
);

OR2x6_ASAP7_75t_L g7216 ( 
.A(n_5995),
.B(n_5682),
.Y(n_7216)
);

AOI22xp33_ASAP7_75t_L g7217 ( 
.A1(n_6020),
.A2(n_6001),
.B1(n_6041),
.B2(n_6092),
.Y(n_7217)
);

BUFx6f_ASAP7_75t_L g7218 ( 
.A(n_5951),
.Y(n_7218)
);

CKINVDCx16_ASAP7_75t_R g7219 ( 
.A(n_6129),
.Y(n_7219)
);

INVx1_ASAP7_75t_SL g7220 ( 
.A(n_6386),
.Y(n_7220)
);

CKINVDCx5p33_ASAP7_75t_R g7221 ( 
.A(n_6144),
.Y(n_7221)
);

INVx2_ASAP7_75t_L g7222 ( 
.A(n_5905),
.Y(n_7222)
);

NAND2x1p5_ASAP7_75t_L g7223 ( 
.A(n_5951),
.B(n_4672),
.Y(n_7223)
);

INVx2_ASAP7_75t_L g7224 ( 
.A(n_5905),
.Y(n_7224)
);

AOI21xp5_ASAP7_75t_L g7225 ( 
.A1(n_6536),
.A2(n_5046),
.B(n_5032),
.Y(n_7225)
);

INVx2_ASAP7_75t_L g7226 ( 
.A(n_5922),
.Y(n_7226)
);

AOI21xp5_ASAP7_75t_L g7227 ( 
.A1(n_6543),
.A2(n_5046),
.B(n_5032),
.Y(n_7227)
);

OAI22xp33_ASAP7_75t_L g7228 ( 
.A1(n_5988),
.A2(n_4846),
.B1(n_4854),
.B2(n_4819),
.Y(n_7228)
);

NAND2xp5_ASAP7_75t_L g7229 ( 
.A(n_6612),
.B(n_5291),
.Y(n_7229)
);

INVx2_ASAP7_75t_L g7230 ( 
.A(n_5922),
.Y(n_7230)
);

NAND2xp5_ASAP7_75t_SL g7231 ( 
.A(n_6254),
.B(n_5335),
.Y(n_7231)
);

AOI21xp5_ASAP7_75t_L g7232 ( 
.A1(n_6543),
.A2(n_5046),
.B(n_5032),
.Y(n_7232)
);

AOI21xp5_ASAP7_75t_L g7233 ( 
.A1(n_6272),
.A2(n_5046),
.B(n_5032),
.Y(n_7233)
);

INVx1_ASAP7_75t_SL g7234 ( 
.A(n_6386),
.Y(n_7234)
);

AOI21xp5_ASAP7_75t_L g7235 ( 
.A1(n_6272),
.A2(n_5046),
.B(n_5032),
.Y(n_7235)
);

AOI22xp33_ASAP7_75t_SL g7236 ( 
.A1(n_6185),
.A2(n_4935),
.B1(n_4889),
.B2(n_4705),
.Y(n_7236)
);

AND2x6_ASAP7_75t_L g7237 ( 
.A(n_5821),
.B(n_4819),
.Y(n_7237)
);

BUFx2_ASAP7_75t_L g7238 ( 
.A(n_6461),
.Y(n_7238)
);

AOI21xp5_ASAP7_75t_L g7239 ( 
.A1(n_6198),
.A2(n_5052),
.B(n_5046),
.Y(n_7239)
);

AND2x6_ASAP7_75t_L g7240 ( 
.A(n_5821),
.B(n_4846),
.Y(n_7240)
);

OAI22xp5_ASAP7_75t_L g7241 ( 
.A1(n_6129),
.A2(n_5267),
.B1(n_5268),
.B2(n_5245),
.Y(n_7241)
);

A2O1A1Ixp33_ASAP7_75t_L g7242 ( 
.A1(n_6056),
.A2(n_5328),
.B(n_4863),
.C(n_4804),
.Y(n_7242)
);

AOI21xp33_ASAP7_75t_L g7243 ( 
.A1(n_6054),
.A2(n_4967),
.B(n_4952),
.Y(n_7243)
);

BUFx12f_ASAP7_75t_L g7244 ( 
.A(n_6861),
.Y(n_7244)
);

BUFx10_ASAP7_75t_L g7245 ( 
.A(n_6126),
.Y(n_7245)
);

BUFx8_ASAP7_75t_L g7246 ( 
.A(n_6126),
.Y(n_7246)
);

BUFx8_ASAP7_75t_L g7247 ( 
.A(n_6585),
.Y(n_7247)
);

BUFx10_ASAP7_75t_L g7248 ( 
.A(n_6585),
.Y(n_7248)
);

AOI21xp33_ASAP7_75t_L g7249 ( 
.A1(n_5942),
.A2(n_5104),
.B(n_5061),
.Y(n_7249)
);

NAND2xp5_ASAP7_75t_SL g7250 ( 
.A(n_6254),
.B(n_5335),
.Y(n_7250)
);

BUFx4_ASAP7_75t_SL g7251 ( 
.A(n_6355),
.Y(n_7251)
);

CKINVDCx5p33_ASAP7_75t_R g7252 ( 
.A(n_6144),
.Y(n_7252)
);

BUFx2_ASAP7_75t_L g7253 ( 
.A(n_6461),
.Y(n_7253)
);

INVx1_ASAP7_75t_SL g7254 ( 
.A(n_6386),
.Y(n_7254)
);

CKINVDCx20_ASAP7_75t_R g7255 ( 
.A(n_6211),
.Y(n_7255)
);

NOR2xp33_ASAP7_75t_L g7256 ( 
.A(n_6191),
.B(n_5714),
.Y(n_7256)
);

AOI21xp5_ASAP7_75t_L g7257 ( 
.A1(n_6198),
.A2(n_5052),
.B(n_5046),
.Y(n_7257)
);

INVx4_ASAP7_75t_L g7258 ( 
.A(n_6019),
.Y(n_7258)
);

NAND2x1p5_ASAP7_75t_L g7259 ( 
.A(n_5951),
.B(n_4672),
.Y(n_7259)
);

HB1xp67_ASAP7_75t_L g7260 ( 
.A(n_6307),
.Y(n_7260)
);

O2A1O1Ixp33_ASAP7_75t_L g7261 ( 
.A1(n_6337),
.A2(n_5942),
.B(n_5982),
.C(n_6203),
.Y(n_7261)
);

NAND2xp33_ASAP7_75t_L g7262 ( 
.A(n_6069),
.B(n_5984),
.Y(n_7262)
);

NAND2xp5_ASAP7_75t_L g7263 ( 
.A(n_6803),
.B(n_5291),
.Y(n_7263)
);

INVxp67_ASAP7_75t_SL g7264 ( 
.A(n_6617),
.Y(n_7264)
);

INVx4_ASAP7_75t_L g7265 ( 
.A(n_6019),
.Y(n_7265)
);

AOI21xp5_ASAP7_75t_L g7266 ( 
.A1(n_6301),
.A2(n_5052),
.B(n_5046),
.Y(n_7266)
);

O2A1O1Ixp33_ASAP7_75t_L g7267 ( 
.A1(n_5982),
.A2(n_5759),
.B(n_5753),
.C(n_5663),
.Y(n_7267)
);

BUFx2_ASAP7_75t_L g7268 ( 
.A(n_6461),
.Y(n_7268)
);

AOI22xp33_ASAP7_75t_L g7269 ( 
.A1(n_6020),
.A2(n_4854),
.B1(n_4873),
.B2(n_4846),
.Y(n_7269)
);

NOR2xp33_ASAP7_75t_L g7270 ( 
.A(n_6191),
.B(n_5714),
.Y(n_7270)
);

OAI21xp33_ASAP7_75t_L g7271 ( 
.A1(n_6001),
.A2(n_5663),
.B(n_5662),
.Y(n_7271)
);

BUFx12f_ASAP7_75t_L g7272 ( 
.A(n_6861),
.Y(n_7272)
);

OAI221xp5_ASAP7_75t_L g7273 ( 
.A1(n_5988),
.A2(n_4763),
.B1(n_4732),
.B2(n_5664),
.C(n_5662),
.Y(n_7273)
);

AND2x2_ASAP7_75t_L g7274 ( 
.A(n_6096),
.B(n_4889),
.Y(n_7274)
);

NAND2xp33_ASAP7_75t_L g7275 ( 
.A(n_5984),
.B(n_6035),
.Y(n_7275)
);

NAND2xp5_ASAP7_75t_SL g7276 ( 
.A(n_6143),
.B(n_6079),
.Y(n_7276)
);

AND2x2_ASAP7_75t_L g7277 ( 
.A(n_6096),
.B(n_4889),
.Y(n_7277)
);

OR2x2_ASAP7_75t_L g7278 ( 
.A(n_6212),
.B(n_4889),
.Y(n_7278)
);

A2O1A1Ixp33_ASAP7_75t_L g7279 ( 
.A1(n_6143),
.A2(n_4804),
.B(n_4863),
.C(n_4795),
.Y(n_7279)
);

HB1xp67_ASAP7_75t_L g7280 ( 
.A(n_6332),
.Y(n_7280)
);

AOI21xp5_ASAP7_75t_L g7281 ( 
.A1(n_6293),
.A2(n_6154),
.B(n_6146),
.Y(n_7281)
);

OA22x2_ASAP7_75t_L g7282 ( 
.A1(n_6055),
.A2(n_4659),
.B1(n_4580),
.B2(n_4631),
.Y(n_7282)
);

BUFx2_ASAP7_75t_L g7283 ( 
.A(n_6461),
.Y(n_7283)
);

AOI21xp5_ASAP7_75t_L g7284 ( 
.A1(n_6293),
.A2(n_5052),
.B(n_5046),
.Y(n_7284)
);

NAND2xp5_ASAP7_75t_L g7285 ( 
.A(n_6803),
.B(n_5291),
.Y(n_7285)
);

AND2x2_ASAP7_75t_L g7286 ( 
.A(n_6106),
.B(n_4889),
.Y(n_7286)
);

OAI22xp5_ASAP7_75t_L g7287 ( 
.A1(n_6391),
.A2(n_5267),
.B1(n_5268),
.B2(n_5245),
.Y(n_7287)
);

AOI222xp33_ASAP7_75t_L g7288 ( 
.A1(n_6041),
.A2(n_5150),
.B1(n_5022),
.B2(n_5174),
.C1(n_5090),
.C2(n_5013),
.Y(n_7288)
);

BUFx2_ASAP7_75t_L g7289 ( 
.A(n_6461),
.Y(n_7289)
);

AOI21xp5_ASAP7_75t_L g7290 ( 
.A1(n_6295),
.A2(n_5075),
.B(n_5052),
.Y(n_7290)
);

AOI21xp5_ASAP7_75t_L g7291 ( 
.A1(n_6295),
.A2(n_6154),
.B(n_6146),
.Y(n_7291)
);

AOI21xp5_ASAP7_75t_L g7292 ( 
.A1(n_6163),
.A2(n_5075),
.B(n_5052),
.Y(n_7292)
);

INVx3_ASAP7_75t_SL g7293 ( 
.A(n_6082),
.Y(n_7293)
);

NAND2xp5_ASAP7_75t_SL g7294 ( 
.A(n_6079),
.B(n_5335),
.Y(n_7294)
);

BUFx12f_ASAP7_75t_L g7295 ( 
.A(n_6861),
.Y(n_7295)
);

OAI21x1_ASAP7_75t_SL g7296 ( 
.A1(n_6066),
.A2(n_5557),
.B(n_5547),
.Y(n_7296)
);

AOI21xp5_ASAP7_75t_L g7297 ( 
.A1(n_6309),
.A2(n_5075),
.B(n_5052),
.Y(n_7297)
);

AO21x1_ASAP7_75t_L g7298 ( 
.A1(n_6115),
.A2(n_6161),
.B(n_6010),
.Y(n_7298)
);

CKINVDCx8_ASAP7_75t_R g7299 ( 
.A(n_6111),
.Y(n_7299)
);

NAND2x1p5_ASAP7_75t_L g7300 ( 
.A(n_6028),
.B(n_4672),
.Y(n_7300)
);

BUFx2_ASAP7_75t_L g7301 ( 
.A(n_6469),
.Y(n_7301)
);

HB1xp67_ASAP7_75t_L g7302 ( 
.A(n_6332),
.Y(n_7302)
);

CKINVDCx8_ASAP7_75t_R g7303 ( 
.A(n_6124),
.Y(n_7303)
);

CKINVDCx5p33_ASAP7_75t_R g7304 ( 
.A(n_6162),
.Y(n_7304)
);

AOI21xp5_ASAP7_75t_L g7305 ( 
.A1(n_6363),
.A2(n_6163),
.B(n_6157),
.Y(n_7305)
);

NAND2x1p5_ASAP7_75t_L g7306 ( 
.A(n_6028),
.B(n_4672),
.Y(n_7306)
);

INVx1_ASAP7_75t_SL g7307 ( 
.A(n_6471),
.Y(n_7307)
);

AOI22xp5_ASAP7_75t_L g7308 ( 
.A1(n_6152),
.A2(n_4705),
.B1(n_4720),
.B2(n_4690),
.Y(n_7308)
);

BUFx12f_ASAP7_75t_L g7309 ( 
.A(n_6482),
.Y(n_7309)
);

NAND2xp5_ASAP7_75t_SL g7310 ( 
.A(n_6178),
.B(n_5335),
.Y(n_7310)
);

AOI22xp5_ASAP7_75t_L g7311 ( 
.A1(n_6152),
.A2(n_4705),
.B1(n_4720),
.B2(n_4690),
.Y(n_7311)
);

AOI21xp5_ASAP7_75t_L g7312 ( 
.A1(n_6197),
.A2(n_5075),
.B(n_5052),
.Y(n_7312)
);

AOI22xp33_ASAP7_75t_L g7313 ( 
.A1(n_5844),
.A2(n_4854),
.B1(n_4873),
.B2(n_4846),
.Y(n_7313)
);

CKINVDCx5p33_ASAP7_75t_R g7314 ( 
.A(n_6162),
.Y(n_7314)
);

AOI221xp5_ASAP7_75t_L g7315 ( 
.A1(n_6203),
.A2(n_5271),
.B1(n_5303),
.B2(n_5267),
.C(n_5245),
.Y(n_7315)
);

AO21x2_ASAP7_75t_L g7316 ( 
.A1(n_6130),
.A2(n_4574),
.B(n_4571),
.Y(n_7316)
);

INVxp67_ASAP7_75t_SL g7317 ( 
.A(n_6617),
.Y(n_7317)
);

BUFx12f_ASAP7_75t_L g7318 ( 
.A(n_6482),
.Y(n_7318)
);

NAND2xp5_ASAP7_75t_L g7319 ( 
.A(n_6714),
.B(n_5306),
.Y(n_7319)
);

NAND2xp5_ASAP7_75t_L g7320 ( 
.A(n_6714),
.B(n_5306),
.Y(n_7320)
);

O2A1O1Ixp5_ASAP7_75t_SL g7321 ( 
.A1(n_6099),
.A2(n_5695),
.B(n_5698),
.C(n_5696),
.Y(n_7321)
);

AND2x4_ASAP7_75t_L g7322 ( 
.A(n_6108),
.B(n_6134),
.Y(n_7322)
);

OR2x2_ASAP7_75t_L g7323 ( 
.A(n_6471),
.B(n_4935),
.Y(n_7323)
);

O2A1O1Ixp33_ASAP7_75t_SL g7324 ( 
.A1(n_5967),
.A2(n_6509),
.B(n_6501),
.C(n_6508),
.Y(n_7324)
);

O2A1O1Ixp33_ASAP7_75t_L g7325 ( 
.A1(n_6035),
.A2(n_5669),
.B(n_5670),
.C(n_5664),
.Y(n_7325)
);

NOR2xp33_ASAP7_75t_L g7326 ( 
.A(n_5844),
.B(n_5743),
.Y(n_7326)
);

BUFx2_ASAP7_75t_L g7327 ( 
.A(n_6469),
.Y(n_7327)
);

BUFx2_ASAP7_75t_L g7328 ( 
.A(n_6469),
.Y(n_7328)
);

BUFx2_ASAP7_75t_L g7329 ( 
.A(n_6469),
.Y(n_7329)
);

BUFx8_ASAP7_75t_SL g7330 ( 
.A(n_6211),
.Y(n_7330)
);

OR2x6_ASAP7_75t_L g7331 ( 
.A(n_5995),
.B(n_5682),
.Y(n_7331)
);

NAND2xp5_ASAP7_75t_L g7332 ( 
.A(n_6736),
.B(n_5306),
.Y(n_7332)
);

AOI21xp5_ASAP7_75t_L g7333 ( 
.A1(n_6363),
.A2(n_5075),
.B(n_5052),
.Y(n_7333)
);

NAND2xp33_ASAP7_75t_L g7334 ( 
.A(n_5801),
.B(n_5174),
.Y(n_7334)
);

AOI21xp5_ASAP7_75t_L g7335 ( 
.A1(n_6268),
.A2(n_6197),
.B(n_6157),
.Y(n_7335)
);

HB1xp67_ASAP7_75t_L g7336 ( 
.A(n_6342),
.Y(n_7336)
);

NOR2xp33_ASAP7_75t_SL g7337 ( 
.A(n_5859),
.B(n_5374),
.Y(n_7337)
);

BUFx2_ASAP7_75t_L g7338 ( 
.A(n_6469),
.Y(n_7338)
);

INVx1_ASAP7_75t_SL g7339 ( 
.A(n_6471),
.Y(n_7339)
);

OAI22xp5_ASAP7_75t_L g7340 ( 
.A1(n_6391),
.A2(n_5303),
.B1(n_5314),
.B2(n_5271),
.Y(n_7340)
);

NAND2xp5_ASAP7_75t_L g7341 ( 
.A(n_6736),
.B(n_5309),
.Y(n_7341)
);

AOI22xp5_ASAP7_75t_L g7342 ( 
.A1(n_6161),
.A2(n_4720),
.B1(n_4730),
.B2(n_4690),
.Y(n_7342)
);

NAND2xp5_ASAP7_75t_L g7343 ( 
.A(n_6270),
.B(n_5309),
.Y(n_7343)
);

AOI21xp5_ASAP7_75t_L g7344 ( 
.A1(n_6216),
.A2(n_5097),
.B(n_5075),
.Y(n_7344)
);

BUFx6f_ASAP7_75t_L g7345 ( 
.A(n_6036),
.Y(n_7345)
);

OAI21xp5_ASAP7_75t_L g7346 ( 
.A1(n_6297),
.A2(n_5501),
.B(n_5465),
.Y(n_7346)
);

CKINVDCx8_ASAP7_75t_R g7347 ( 
.A(n_6124),
.Y(n_7347)
);

INVxp67_ASAP7_75t_SL g7348 ( 
.A(n_6641),
.Y(n_7348)
);

NAND2xp5_ASAP7_75t_L g7349 ( 
.A(n_6270),
.B(n_5309),
.Y(n_7349)
);

OR2x2_ASAP7_75t_SL g7350 ( 
.A(n_5968),
.B(n_4846),
.Y(n_7350)
);

BUFx2_ASAP7_75t_L g7351 ( 
.A(n_6469),
.Y(n_7351)
);

BUFx2_ASAP7_75t_L g7352 ( 
.A(n_6535),
.Y(n_7352)
);

BUFx6f_ASAP7_75t_L g7353 ( 
.A(n_6036),
.Y(n_7353)
);

NAND2xp5_ASAP7_75t_SL g7354 ( 
.A(n_6178),
.B(n_5335),
.Y(n_7354)
);

BUFx6f_ASAP7_75t_L g7355 ( 
.A(n_6036),
.Y(n_7355)
);

INVx1_ASAP7_75t_SL g7356 ( 
.A(n_6515),
.Y(n_7356)
);

NAND2xp5_ASAP7_75t_L g7357 ( 
.A(n_6275),
.B(n_5309),
.Y(n_7357)
);

HB1xp67_ASAP7_75t_L g7358 ( 
.A(n_6342),
.Y(n_7358)
);

HB1xp67_ASAP7_75t_L g7359 ( 
.A(n_6366),
.Y(n_7359)
);

CKINVDCx5p33_ASAP7_75t_R g7360 ( 
.A(n_6449),
.Y(n_7360)
);

NAND2xp5_ASAP7_75t_SL g7361 ( 
.A(n_6115),
.B(n_5365),
.Y(n_7361)
);

NAND3xp33_ASAP7_75t_L g7362 ( 
.A(n_6066),
.B(n_5670),
.C(n_5669),
.Y(n_7362)
);

CKINVDCx5p33_ASAP7_75t_R g7363 ( 
.A(n_6449),
.Y(n_7363)
);

NAND2x1p5_ASAP7_75t_L g7364 ( 
.A(n_6036),
.B(n_4724),
.Y(n_7364)
);

NAND2xp5_ASAP7_75t_L g7365 ( 
.A(n_6275),
.B(n_5313),
.Y(n_7365)
);

BUFx6f_ASAP7_75t_L g7366 ( 
.A(n_6036),
.Y(n_7366)
);

BUFx6f_ASAP7_75t_L g7367 ( 
.A(n_6036),
.Y(n_7367)
);

AOI22xp33_ASAP7_75t_L g7368 ( 
.A1(n_6099),
.A2(n_4854),
.B1(n_4873),
.B2(n_4846),
.Y(n_7368)
);

NOR2x1_ASAP7_75t_L g7369 ( 
.A(n_6177),
.B(n_5715),
.Y(n_7369)
);

A2O1A1Ixp33_ASAP7_75t_L g7370 ( 
.A1(n_6078),
.A2(n_4804),
.B(n_4863),
.C(n_4795),
.Y(n_7370)
);

NOR2xp33_ASAP7_75t_L g7371 ( 
.A(n_6120),
.B(n_5743),
.Y(n_7371)
);

AOI22xp5_ASAP7_75t_L g7372 ( 
.A1(n_6156),
.A2(n_4755),
.B1(n_4777),
.B2(n_4730),
.Y(n_7372)
);

OR2x6_ASAP7_75t_L g7373 ( 
.A(n_5995),
.B(n_5682),
.Y(n_7373)
);

AOI22xp33_ASAP7_75t_L g7374 ( 
.A1(n_6138),
.A2(n_4873),
.B1(n_4854),
.B2(n_4755),
.Y(n_7374)
);

BUFx6f_ASAP7_75t_L g7375 ( 
.A(n_6043),
.Y(n_7375)
);

NAND2xp5_ASAP7_75t_L g7376 ( 
.A(n_6277),
.B(n_5318),
.Y(n_7376)
);

BUFx6f_ASAP7_75t_L g7377 ( 
.A(n_6043),
.Y(n_7377)
);

BUFx6f_ASAP7_75t_L g7378 ( 
.A(n_6043),
.Y(n_7378)
);

AOI22xp33_ASAP7_75t_L g7379 ( 
.A1(n_6138),
.A2(n_4873),
.B1(n_4854),
.B2(n_4755),
.Y(n_7379)
);

AOI21xp5_ASAP7_75t_L g7380 ( 
.A1(n_6279),
.A2(n_5097),
.B(n_5075),
.Y(n_7380)
);

BUFx8_ASAP7_75t_L g7381 ( 
.A(n_6585),
.Y(n_7381)
);

AOI21xp5_ASAP7_75t_L g7382 ( 
.A1(n_6279),
.A2(n_5097),
.B(n_5075),
.Y(n_7382)
);

OAI22xp5_ASAP7_75t_L g7383 ( 
.A1(n_6158),
.A2(n_5303),
.B1(n_5314),
.B2(n_5271),
.Y(n_7383)
);

OR2x6_ASAP7_75t_SL g7384 ( 
.A(n_6551),
.B(n_5300),
.Y(n_7384)
);

AND2x2_ASAP7_75t_SL g7385 ( 
.A(n_5766),
.B(n_5075),
.Y(n_7385)
);

A2O1A1Ixp33_ASAP7_75t_L g7386 ( 
.A1(n_6078),
.A2(n_6352),
.B(n_6297),
.C(n_6181),
.Y(n_7386)
);

CKINVDCx20_ASAP7_75t_R g7387 ( 
.A(n_6326),
.Y(n_7387)
);

NAND2xp5_ASAP7_75t_L g7388 ( 
.A(n_6277),
.B(n_5323),
.Y(n_7388)
);

AOI22xp33_ASAP7_75t_L g7389 ( 
.A1(n_6131),
.A2(n_4873),
.B1(n_4755),
.B2(n_4777),
.Y(n_7389)
);

INVxp67_ASAP7_75t_SL g7390 ( 
.A(n_6641),
.Y(n_7390)
);

AOI22xp33_ASAP7_75t_L g7391 ( 
.A1(n_6131),
.A2(n_4873),
.B1(n_4777),
.B2(n_4781),
.Y(n_7391)
);

OAI22xp5_ASAP7_75t_L g7392 ( 
.A1(n_6158),
.A2(n_6508),
.B1(n_6294),
.B2(n_6196),
.Y(n_7392)
);

NOR2xp33_ASAP7_75t_L g7393 ( 
.A(n_6120),
.B(n_5743),
.Y(n_7393)
);

AOI22xp33_ASAP7_75t_L g7394 ( 
.A1(n_6260),
.A2(n_4873),
.B1(n_4777),
.B2(n_4781),
.Y(n_7394)
);

CKINVDCx5p33_ASAP7_75t_R g7395 ( 
.A(n_6029),
.Y(n_7395)
);

AOI21xp5_ASAP7_75t_L g7396 ( 
.A1(n_6497),
.A2(n_5130),
.B(n_5097),
.Y(n_7396)
);

BUFx2_ASAP7_75t_L g7397 ( 
.A(n_6535),
.Y(n_7397)
);

CKINVDCx11_ASAP7_75t_R g7398 ( 
.A(n_5873),
.Y(n_7398)
);

AOI22xp5_ASAP7_75t_L g7399 ( 
.A1(n_6156),
.A2(n_4781),
.B1(n_4835),
.B2(n_4730),
.Y(n_7399)
);

AO21x1_ASAP7_75t_L g7400 ( 
.A1(n_6725),
.A2(n_4909),
.B(n_4903),
.Y(n_7400)
);

BUFx12f_ASAP7_75t_L g7401 ( 
.A(n_6640),
.Y(n_7401)
);

OR2x2_ASAP7_75t_L g7402 ( 
.A(n_6515),
.B(n_4935),
.Y(n_7402)
);

AOI22xp33_ASAP7_75t_L g7403 ( 
.A1(n_6260),
.A2(n_4873),
.B1(n_4781),
.B2(n_4835),
.Y(n_7403)
);

HB1xp67_ASAP7_75t_L g7404 ( 
.A(n_6366),
.Y(n_7404)
);

AOI21xp5_ASAP7_75t_L g7405 ( 
.A1(n_6268),
.A2(n_5130),
.B(n_5097),
.Y(n_7405)
);

OR2x6_ASAP7_75t_L g7406 ( 
.A(n_5995),
.B(n_4724),
.Y(n_7406)
);

NAND2xp5_ASAP7_75t_L g7407 ( 
.A(n_6328),
.B(n_5887),
.Y(n_7407)
);

BUFx6f_ASAP7_75t_SL g7408 ( 
.A(n_6324),
.Y(n_7408)
);

OR2x6_ASAP7_75t_L g7409 ( 
.A(n_6032),
.B(n_4724),
.Y(n_7409)
);

AOI22xp33_ASAP7_75t_L g7410 ( 
.A1(n_6353),
.A2(n_4835),
.B1(n_4852),
.B2(n_4730),
.Y(n_7410)
);

AOI21xp5_ASAP7_75t_L g7411 ( 
.A1(n_6257),
.A2(n_5130),
.B(n_5097),
.Y(n_7411)
);

OR2x6_ASAP7_75t_L g7412 ( 
.A(n_6032),
.B(n_4724),
.Y(n_7412)
);

AOI21xp5_ASAP7_75t_L g7413 ( 
.A1(n_6257),
.A2(n_5130),
.B(n_5097),
.Y(n_7413)
);

OAI22xp5_ASAP7_75t_L g7414 ( 
.A1(n_6294),
.A2(n_5345),
.B1(n_5336),
.B2(n_5312),
.Y(n_7414)
);

OAI21x1_ASAP7_75t_L g7415 ( 
.A1(n_6102),
.A2(n_6745),
.B(n_6216),
.Y(n_7415)
);

CKINVDCx16_ASAP7_75t_R g7416 ( 
.A(n_6585),
.Y(n_7416)
);

HB1xp67_ASAP7_75t_L g7417 ( 
.A(n_6368),
.Y(n_7417)
);

CKINVDCx20_ASAP7_75t_R g7418 ( 
.A(n_6831),
.Y(n_7418)
);

AOI22xp5_ASAP7_75t_L g7419 ( 
.A1(n_6055),
.A2(n_6411),
.B1(n_6077),
.B2(n_6582),
.Y(n_7419)
);

AOI22xp5_ASAP7_75t_L g7420 ( 
.A1(n_6411),
.A2(n_4835),
.B1(n_4852),
.B2(n_5748),
.Y(n_7420)
);

AOI21xp5_ASAP7_75t_L g7421 ( 
.A1(n_6385),
.A2(n_5133),
.B(n_5130),
.Y(n_7421)
);

NOR2xp33_ASAP7_75t_L g7422 ( 
.A(n_5967),
.B(n_5748),
.Y(n_7422)
);

AOI21x1_ASAP7_75t_L g7423 ( 
.A1(n_6255),
.A2(n_5700),
.B(n_5501),
.Y(n_7423)
);

INVx6_ASAP7_75t_L g7424 ( 
.A(n_6460),
.Y(n_7424)
);

AOI22xp5_ASAP7_75t_L g7425 ( 
.A1(n_6077),
.A2(n_4852),
.B1(n_5704),
.B2(n_5701),
.Y(n_7425)
);

BUFx2_ASAP7_75t_L g7426 ( 
.A(n_6535),
.Y(n_7426)
);

INVx8_ASAP7_75t_L g7427 ( 
.A(n_5908),
.Y(n_7427)
);

CKINVDCx5p33_ASAP7_75t_R g7428 ( 
.A(n_6029),
.Y(n_7428)
);

CKINVDCx5p33_ASAP7_75t_R g7429 ( 
.A(n_6029),
.Y(n_7429)
);

HB1xp67_ASAP7_75t_L g7430 ( 
.A(n_6368),
.Y(n_7430)
);

INVx5_ASAP7_75t_L g7431 ( 
.A(n_6050),
.Y(n_7431)
);

CKINVDCx8_ASAP7_75t_R g7432 ( 
.A(n_6336),
.Y(n_7432)
);

AND2x6_ASAP7_75t_L g7433 ( 
.A(n_5821),
.B(n_4852),
.Y(n_7433)
);

NOR2xp33_ASAP7_75t_L g7434 ( 
.A(n_6225),
.B(n_5104),
.Y(n_7434)
);

BUFx2_ASAP7_75t_L g7435 ( 
.A(n_6535),
.Y(n_7435)
);

BUFx3_ASAP7_75t_L g7436 ( 
.A(n_6370),
.Y(n_7436)
);

OR2x6_ASAP7_75t_L g7437 ( 
.A(n_6032),
.B(n_4724),
.Y(n_7437)
);

BUFx6f_ASAP7_75t_L g7438 ( 
.A(n_6050),
.Y(n_7438)
);

NAND2xp5_ASAP7_75t_SL g7439 ( 
.A(n_6556),
.B(n_5365),
.Y(n_7439)
);

BUFx3_ASAP7_75t_L g7440 ( 
.A(n_6370),
.Y(n_7440)
);

AOI22xp5_ASAP7_75t_L g7441 ( 
.A1(n_6582),
.A2(n_5701),
.B1(n_5705),
.B2(n_5704),
.Y(n_7441)
);

AOI22xp5_ASAP7_75t_L g7442 ( 
.A1(n_6287),
.A2(n_5705),
.B1(n_4763),
.B2(n_5345),
.Y(n_7442)
);

CKINVDCx5p33_ASAP7_75t_R g7443 ( 
.A(n_6039),
.Y(n_7443)
);

BUFx6f_ASAP7_75t_L g7444 ( 
.A(n_6050),
.Y(n_7444)
);

BUFx12f_ASAP7_75t_L g7445 ( 
.A(n_6640),
.Y(n_7445)
);

AOI21xp5_ASAP7_75t_L g7446 ( 
.A1(n_6309),
.A2(n_5133),
.B(n_5130),
.Y(n_7446)
);

AOI22xp33_ASAP7_75t_L g7447 ( 
.A1(n_6353),
.A2(n_5345),
.B1(n_5336),
.B2(n_5302),
.Y(n_7447)
);

AND2x2_ASAP7_75t_L g7448 ( 
.A(n_5868),
.B(n_5869),
.Y(n_7448)
);

A2O1A1Ixp33_ASAP7_75t_L g7449 ( 
.A1(n_6352),
.A2(n_4863),
.B(n_4933),
.C(n_4795),
.Y(n_7449)
);

BUFx2_ASAP7_75t_L g7450 ( 
.A(n_6535),
.Y(n_7450)
);

BUFx4f_ASAP7_75t_SL g7451 ( 
.A(n_5873),
.Y(n_7451)
);

BUFx2_ASAP7_75t_L g7452 ( 
.A(n_6535),
.Y(n_7452)
);

INVxp67_ASAP7_75t_L g7453 ( 
.A(n_6104),
.Y(n_7453)
);

AOI21xp5_ASAP7_75t_L g7454 ( 
.A1(n_6301),
.A2(n_5160),
.B(n_5133),
.Y(n_7454)
);

AOI22xp5_ASAP7_75t_L g7455 ( 
.A1(n_6287),
.A2(n_4763),
.B1(n_5336),
.B2(n_5520),
.Y(n_7455)
);

BUFx12f_ASAP7_75t_L g7456 ( 
.A(n_6644),
.Y(n_7456)
);

BUFx6f_ASAP7_75t_L g7457 ( 
.A(n_6050),
.Y(n_7457)
);

INVx3_ASAP7_75t_L g7458 ( 
.A(n_5868),
.Y(n_7458)
);

NOR2xp67_ASAP7_75t_L g7459 ( 
.A(n_6104),
.B(n_5721),
.Y(n_7459)
);

BUFx6f_ASAP7_75t_L g7460 ( 
.A(n_6050),
.Y(n_7460)
);

INVx3_ASAP7_75t_SL g7461 ( 
.A(n_6082),
.Y(n_7461)
);

NOR2xp33_ASAP7_75t_L g7462 ( 
.A(n_6225),
.B(n_5735),
.Y(n_7462)
);

INVx6_ASAP7_75t_L g7463 ( 
.A(n_6460),
.Y(n_7463)
);

INVx1_ASAP7_75t_SL g7464 ( 
.A(n_6531),
.Y(n_7464)
);

CKINVDCx5p33_ASAP7_75t_R g7465 ( 
.A(n_6039),
.Y(n_7465)
);

BUFx2_ASAP7_75t_L g7466 ( 
.A(n_6555),
.Y(n_7466)
);

O2A1O1Ixp33_ASAP7_75t_L g7467 ( 
.A1(n_6501),
.A2(n_5674),
.B(n_5312),
.C(n_5735),
.Y(n_7467)
);

BUFx2_ASAP7_75t_L g7468 ( 
.A(n_6555),
.Y(n_7468)
);

CKINVDCx8_ASAP7_75t_R g7469 ( 
.A(n_6336),
.Y(n_7469)
);

INVx3_ASAP7_75t_R g7470 ( 
.A(n_6813),
.Y(n_7470)
);

BUFx2_ASAP7_75t_R g7471 ( 
.A(n_6813),
.Y(n_7471)
);

INVx3_ASAP7_75t_L g7472 ( 
.A(n_5869),
.Y(n_7472)
);

NOR2xp33_ASAP7_75t_L g7473 ( 
.A(n_6564),
.B(n_5735),
.Y(n_7473)
);

INVxp67_ASAP7_75t_L g7474 ( 
.A(n_6104),
.Y(n_7474)
);

INVx1_ASAP7_75t_SL g7475 ( 
.A(n_6531),
.Y(n_7475)
);

CKINVDCx16_ASAP7_75t_R g7476 ( 
.A(n_6585),
.Y(n_7476)
);

A2O1A1Ixp33_ASAP7_75t_L g7477 ( 
.A1(n_6181),
.A2(n_4863),
.B(n_4933),
.C(n_4795),
.Y(n_7477)
);

AOI21xp5_ASAP7_75t_L g7478 ( 
.A1(n_6215),
.A2(n_5160),
.B(n_5133),
.Y(n_7478)
);

AOI21xp5_ASAP7_75t_L g7479 ( 
.A1(n_6215),
.A2(n_5160),
.B(n_5133),
.Y(n_7479)
);

AOI21xp5_ASAP7_75t_L g7480 ( 
.A1(n_6373),
.A2(n_5205),
.B(n_5160),
.Y(n_7480)
);

HB1xp67_ASAP7_75t_L g7481 ( 
.A(n_6491),
.Y(n_7481)
);

INVx2_ASAP7_75t_SL g7482 ( 
.A(n_6303),
.Y(n_7482)
);

AOI22xp33_ASAP7_75t_L g7483 ( 
.A1(n_5767),
.A2(n_5300),
.B1(n_4909),
.B2(n_4911),
.Y(n_7483)
);

CKINVDCx5p33_ASAP7_75t_R g7484 ( 
.A(n_6039),
.Y(n_7484)
);

NAND2xp33_ASAP7_75t_L g7485 ( 
.A(n_5801),
.B(n_5035),
.Y(n_7485)
);

BUFx2_ASAP7_75t_L g7486 ( 
.A(n_6555),
.Y(n_7486)
);

INVx6_ASAP7_75t_L g7487 ( 
.A(n_6873),
.Y(n_7487)
);

NAND2xp5_ASAP7_75t_SL g7488 ( 
.A(n_6566),
.B(n_5365),
.Y(n_7488)
);

AND2x2_ASAP7_75t_L g7489 ( 
.A(n_5869),
.B(n_5902),
.Y(n_7489)
);

NAND2xp5_ASAP7_75t_SL g7490 ( 
.A(n_6566),
.B(n_5365),
.Y(n_7490)
);

INVx2_ASAP7_75t_SL g7491 ( 
.A(n_6303),
.Y(n_7491)
);

BUFx2_ASAP7_75t_L g7492 ( 
.A(n_6555),
.Y(n_7492)
);

CKINVDCx5p33_ASAP7_75t_R g7493 ( 
.A(n_5973),
.Y(n_7493)
);

BUFx3_ASAP7_75t_L g7494 ( 
.A(n_6370),
.Y(n_7494)
);

CKINVDCx5p33_ASAP7_75t_R g7495 ( 
.A(n_5973),
.Y(n_7495)
);

NOR2xp33_ASAP7_75t_L g7496 ( 
.A(n_6564),
.B(n_5752),
.Y(n_7496)
);

INVx2_ASAP7_75t_SL g7497 ( 
.A(n_6303),
.Y(n_7497)
);

AOI22xp33_ASAP7_75t_L g7498 ( 
.A1(n_5767),
.A2(n_4909),
.B1(n_4911),
.B2(n_4903),
.Y(n_7498)
);

BUFx2_ASAP7_75t_L g7499 ( 
.A(n_6555),
.Y(n_7499)
);

A2O1A1Ixp33_ASAP7_75t_L g7500 ( 
.A1(n_5805),
.A2(n_4933),
.B(n_5103),
.C(n_4795),
.Y(n_7500)
);

HB1xp67_ASAP7_75t_L g7501 ( 
.A(n_6491),
.Y(n_7501)
);

BUFx2_ASAP7_75t_L g7502 ( 
.A(n_6555),
.Y(n_7502)
);

AOI21xp5_ASAP7_75t_L g7503 ( 
.A1(n_6520),
.A2(n_5205),
.B(n_5160),
.Y(n_7503)
);

INVx8_ASAP7_75t_L g7504 ( 
.A(n_5908),
.Y(n_7504)
);

AOI22xp33_ASAP7_75t_L g7505 ( 
.A1(n_5974),
.A2(n_4911),
.B1(n_4913),
.B2(n_4903),
.Y(n_7505)
);

NOR2x1_ASAP7_75t_SL g7506 ( 
.A(n_6801),
.B(n_5508),
.Y(n_7506)
);

CKINVDCx20_ASAP7_75t_R g7507 ( 
.A(n_6831),
.Y(n_7507)
);

OAI22xp33_ASAP7_75t_L g7508 ( 
.A1(n_6238),
.A2(n_5554),
.B1(n_5538),
.B2(n_4933),
.Y(n_7508)
);

INVx6_ASAP7_75t_SL g7509 ( 
.A(n_5811),
.Y(n_7509)
);

AOI221xp5_ASAP7_75t_L g7510 ( 
.A1(n_6247),
.A2(n_4923),
.B1(n_4934),
.B2(n_4918),
.C(n_4913),
.Y(n_7510)
);

AOI22xp5_ASAP7_75t_L g7511 ( 
.A1(n_5925),
.A2(n_5528),
.B1(n_5520),
.B2(n_5674),
.Y(n_7511)
);

AOI21xp33_ASAP7_75t_L g7512 ( 
.A1(n_6509),
.A2(n_5575),
.B(n_5712),
.Y(n_7512)
);

AOI22xp33_ASAP7_75t_L g7513 ( 
.A1(n_5974),
.A2(n_4918),
.B1(n_4923),
.B2(n_4913),
.Y(n_7513)
);

CKINVDCx16_ASAP7_75t_R g7514 ( 
.A(n_5826),
.Y(n_7514)
);

OA21x2_ASAP7_75t_L g7515 ( 
.A1(n_6102),
.A2(n_5723),
.B(n_5721),
.Y(n_7515)
);

NOR2xp33_ASAP7_75t_L g7516 ( 
.A(n_6592),
.B(n_5752),
.Y(n_7516)
);

CKINVDCx5p33_ASAP7_75t_R g7517 ( 
.A(n_5973),
.Y(n_7517)
);

AND2x4_ASAP7_75t_L g7518 ( 
.A(n_5811),
.B(n_5902),
.Y(n_7518)
);

BUFx6f_ASAP7_75t_L g7519 ( 
.A(n_6089),
.Y(n_7519)
);

AOI22xp5_ASAP7_75t_L g7520 ( 
.A1(n_5925),
.A2(n_5528),
.B1(n_5140),
.B2(n_5523),
.Y(n_7520)
);

BUFx2_ASAP7_75t_SL g7521 ( 
.A(n_6703),
.Y(n_7521)
);

INVx6_ASAP7_75t_L g7522 ( 
.A(n_6873),
.Y(n_7522)
);

AOI22xp33_ASAP7_75t_L g7523 ( 
.A1(n_6594),
.A2(n_4923),
.B1(n_4934),
.B2(n_4918),
.Y(n_7523)
);

AOI21xp5_ASAP7_75t_L g7524 ( 
.A1(n_6517),
.A2(n_6341),
.B(n_6296),
.Y(n_7524)
);

CKINVDCx5p33_ASAP7_75t_R g7525 ( 
.A(n_5779),
.Y(n_7525)
);

BUFx2_ASAP7_75t_SL g7526 ( 
.A(n_6703),
.Y(n_7526)
);

AOI21xp5_ASAP7_75t_L g7527 ( 
.A1(n_6500),
.A2(n_5205),
.B(n_5160),
.Y(n_7527)
);

BUFx3_ASAP7_75t_L g7528 ( 
.A(n_6703),
.Y(n_7528)
);

INVx5_ASAP7_75t_L g7529 ( 
.A(n_6089),
.Y(n_7529)
);

AOI21xp5_ASAP7_75t_L g7530 ( 
.A1(n_6385),
.A2(n_5258),
.B(n_5205),
.Y(n_7530)
);

BUFx6f_ASAP7_75t_L g7531 ( 
.A(n_6089),
.Y(n_7531)
);

CKINVDCx20_ASAP7_75t_R g7532 ( 
.A(n_6893),
.Y(n_7532)
);

AOI22xp5_ASAP7_75t_L g7533 ( 
.A1(n_6238),
.A2(n_5140),
.B1(n_5523),
.B2(n_5035),
.Y(n_7533)
);

OAI22xp5_ASAP7_75t_L g7534 ( 
.A1(n_6196),
.A2(n_5103),
.B1(n_5179),
.B2(n_4933),
.Y(n_7534)
);

BUFx6f_ASAP7_75t_SL g7535 ( 
.A(n_6324),
.Y(n_7535)
);

BUFx2_ASAP7_75t_L g7536 ( 
.A(n_6600),
.Y(n_7536)
);

AOI21xp5_ASAP7_75t_L g7537 ( 
.A1(n_6524),
.A2(n_5258),
.B(n_5205),
.Y(n_7537)
);

AOI21xp5_ASAP7_75t_L g7538 ( 
.A1(n_6341),
.A2(n_5258),
.B(n_5205),
.Y(n_7538)
);

BUFx12f_ASAP7_75t_L g7539 ( 
.A(n_6644),
.Y(n_7539)
);

AND2x2_ASAP7_75t_L g7540 ( 
.A(n_5940),
.B(n_5972),
.Y(n_7540)
);

CKINVDCx5p33_ASAP7_75t_R g7541 ( 
.A(n_6597),
.Y(n_7541)
);

BUFx3_ASAP7_75t_L g7542 ( 
.A(n_6819),
.Y(n_7542)
);

CKINVDCx5p33_ASAP7_75t_R g7543 ( 
.A(n_6731),
.Y(n_7543)
);

BUFx6f_ASAP7_75t_L g7544 ( 
.A(n_6155),
.Y(n_7544)
);

AOI22xp5_ASAP7_75t_L g7545 ( 
.A1(n_5877),
.A2(n_5140),
.B1(n_5523),
.B2(n_5035),
.Y(n_7545)
);

AOI22xp5_ASAP7_75t_L g7546 ( 
.A1(n_5877),
.A2(n_5140),
.B1(n_5523),
.B2(n_5035),
.Y(n_7546)
);

INVxp67_ASAP7_75t_SL g7547 ( 
.A(n_6492),
.Y(n_7547)
);

AOI21xp5_ASAP7_75t_L g7548 ( 
.A1(n_6477),
.A2(n_5258),
.B(n_5205),
.Y(n_7548)
);

INVx8_ASAP7_75t_L g7549 ( 
.A(n_5908),
.Y(n_7549)
);

CKINVDCx5p33_ASAP7_75t_R g7550 ( 
.A(n_6595),
.Y(n_7550)
);

BUFx2_ASAP7_75t_L g7551 ( 
.A(n_6600),
.Y(n_7551)
);

O2A1O1Ixp33_ASAP7_75t_L g7552 ( 
.A1(n_6024),
.A2(n_5755),
.B(n_5757),
.C(n_5752),
.Y(n_7552)
);

NOR2xp33_ASAP7_75t_L g7553 ( 
.A(n_6592),
.B(n_5755),
.Y(n_7553)
);

AOI21xp5_ASAP7_75t_L g7554 ( 
.A1(n_6296),
.A2(n_5283),
.B(n_5258),
.Y(n_7554)
);

O2A1O1Ixp33_ASAP7_75t_L g7555 ( 
.A1(n_6024),
.A2(n_5757),
.B(n_5758),
.C(n_5755),
.Y(n_7555)
);

BUFx2_ASAP7_75t_L g7556 ( 
.A(n_6600),
.Y(n_7556)
);

AOI21xp5_ASAP7_75t_L g7557 ( 
.A1(n_6373),
.A2(n_5283),
.B(n_5258),
.Y(n_7557)
);

AOI22xp33_ASAP7_75t_L g7558 ( 
.A1(n_6594),
.A2(n_4943),
.B1(n_4959),
.B2(n_4934),
.Y(n_7558)
);

INVx3_ASAP7_75t_L g7559 ( 
.A(n_5972),
.Y(n_7559)
);

AOI22xp33_ASAP7_75t_L g7560 ( 
.A1(n_6247),
.A2(n_4959),
.B1(n_4972),
.B2(n_4943),
.Y(n_7560)
);

AOI22xp5_ASAP7_75t_L g7561 ( 
.A1(n_5788),
.A2(n_5523),
.B1(n_5534),
.B2(n_5140),
.Y(n_7561)
);

INVx3_ASAP7_75t_SL g7562 ( 
.A(n_6082),
.Y(n_7562)
);

INVx3_ASAP7_75t_L g7563 ( 
.A(n_5972),
.Y(n_7563)
);

AOI22xp33_ASAP7_75t_L g7564 ( 
.A1(n_6330),
.A2(n_4959),
.B1(n_4972),
.B2(n_4943),
.Y(n_7564)
);

BUFx2_ASAP7_75t_L g7565 ( 
.A(n_6600),
.Y(n_7565)
);

INVx1_ASAP7_75t_SL g7566 ( 
.A(n_6557),
.Y(n_7566)
);

CKINVDCx5p33_ASAP7_75t_R g7567 ( 
.A(n_5825),
.Y(n_7567)
);

AOI21xp5_ASAP7_75t_L g7568 ( 
.A1(n_6403),
.A2(n_5283),
.B(n_5258),
.Y(n_7568)
);

O2A1O1Ixp5_ASAP7_75t_L g7569 ( 
.A1(n_6256),
.A2(n_4806),
.B(n_5179),
.C(n_5103),
.Y(n_7569)
);

A2O1A1Ixp33_ASAP7_75t_L g7570 ( 
.A1(n_5805),
.A2(n_5179),
.B(n_5279),
.C(n_5103),
.Y(n_7570)
);

AOI22xp33_ASAP7_75t_L g7571 ( 
.A1(n_6330),
.A2(n_4973),
.B1(n_4975),
.B2(n_4972),
.Y(n_7571)
);

BUFx8_ASAP7_75t_L g7572 ( 
.A(n_6906),
.Y(n_7572)
);

NOR2xp33_ASAP7_75t_L g7573 ( 
.A(n_6405),
.B(n_5757),
.Y(n_7573)
);

BUFx2_ASAP7_75t_SL g7574 ( 
.A(n_6819),
.Y(n_7574)
);

O2A1O1Ixp33_ASAP7_75t_L g7575 ( 
.A1(n_5793),
.A2(n_5760),
.B(n_5761),
.C(n_5758),
.Y(n_7575)
);

BUFx4f_ASAP7_75t_L g7576 ( 
.A(n_5978),
.Y(n_7576)
);

INVx5_ASAP7_75t_L g7577 ( 
.A(n_6249),
.Y(n_7577)
);

AOI22xp33_ASAP7_75t_L g7578 ( 
.A1(n_6395),
.A2(n_4975),
.B1(n_4976),
.B2(n_4973),
.Y(n_7578)
);

NAND3xp33_ASAP7_75t_L g7579 ( 
.A(n_6451),
.B(n_4975),
.C(n_4973),
.Y(n_7579)
);

AOI22xp33_ASAP7_75t_L g7580 ( 
.A1(n_6395),
.A2(n_4980),
.B1(n_4987),
.B2(n_4976),
.Y(n_7580)
);

BUFx2_ASAP7_75t_R g7581 ( 
.A(n_6003),
.Y(n_7581)
);

CKINVDCx8_ASAP7_75t_R g7582 ( 
.A(n_6376),
.Y(n_7582)
);

INVx1_ASAP7_75t_SL g7583 ( 
.A(n_6586),
.Y(n_7583)
);

INVx1_ASAP7_75t_SL g7584 ( 
.A(n_6586),
.Y(n_7584)
);

CKINVDCx12_ASAP7_75t_R g7585 ( 
.A(n_6685),
.Y(n_7585)
);

A2O1A1Ixp33_ASAP7_75t_L g7586 ( 
.A1(n_6256),
.A2(n_5179),
.B(n_5279),
.C(n_5103),
.Y(n_7586)
);

INVx5_ASAP7_75t_L g7587 ( 
.A(n_6249),
.Y(n_7587)
);

AOI22xp33_ASAP7_75t_L g7588 ( 
.A1(n_5774),
.A2(n_4980),
.B1(n_4987),
.B2(n_4976),
.Y(n_7588)
);

INVx3_ASAP7_75t_L g7589 ( 
.A(n_5980),
.Y(n_7589)
);

CKINVDCx5p33_ASAP7_75t_R g7590 ( 
.A(n_5843),
.Y(n_7590)
);

BUFx2_ASAP7_75t_L g7591 ( 
.A(n_6600),
.Y(n_7591)
);

NOR2xp33_ASAP7_75t_SL g7592 ( 
.A(n_5826),
.B(n_5538),
.Y(n_7592)
);

OAI22xp5_ASAP7_75t_L g7593 ( 
.A1(n_6554),
.A2(n_5279),
.B1(n_5297),
.B2(n_5179),
.Y(n_7593)
);

BUFx3_ASAP7_75t_L g7594 ( 
.A(n_6819),
.Y(n_7594)
);

INVx8_ASAP7_75t_L g7595 ( 
.A(n_5908),
.Y(n_7595)
);

BUFx4f_ASAP7_75t_L g7596 ( 
.A(n_5978),
.Y(n_7596)
);

INVx1_ASAP7_75t_SL g7597 ( 
.A(n_6586),
.Y(n_7597)
);

NOR2xp67_ASAP7_75t_SL g7598 ( 
.A(n_6003),
.B(n_5538),
.Y(n_7598)
);

BUFx6f_ASAP7_75t_L g7599 ( 
.A(n_6249),
.Y(n_7599)
);

BUFx8_ASAP7_75t_L g7600 ( 
.A(n_5780),
.Y(n_7600)
);

NAND2x1p5_ASAP7_75t_L g7601 ( 
.A(n_6249),
.B(n_4806),
.Y(n_7601)
);

INVx1_ASAP7_75t_SL g7602 ( 
.A(n_6709),
.Y(n_7602)
);

INVx3_ASAP7_75t_L g7603 ( 
.A(n_5980),
.Y(n_7603)
);

A2O1A1Ixp33_ASAP7_75t_L g7604 ( 
.A1(n_6676),
.A2(n_5297),
.B(n_5328),
.C(n_5279),
.Y(n_7604)
);

AOI22xp5_ASAP7_75t_L g7605 ( 
.A1(n_5788),
.A2(n_5523),
.B1(n_5534),
.B2(n_5140),
.Y(n_7605)
);

INVx3_ASAP7_75t_L g7606 ( 
.A(n_5980),
.Y(n_7606)
);

AOI22xp5_ASAP7_75t_L g7607 ( 
.A1(n_6378),
.A2(n_6588),
.B1(n_6574),
.B2(n_5770),
.Y(n_7607)
);

NOR2xp33_ASAP7_75t_L g7608 ( 
.A(n_6405),
.B(n_5758),
.Y(n_7608)
);

BUFx2_ASAP7_75t_L g7609 ( 
.A(n_6600),
.Y(n_7609)
);

BUFx4f_ASAP7_75t_L g7610 ( 
.A(n_5978),
.Y(n_7610)
);

BUFx2_ASAP7_75t_L g7611 ( 
.A(n_6604),
.Y(n_7611)
);

BUFx3_ASAP7_75t_L g7612 ( 
.A(n_6868),
.Y(n_7612)
);

AOI21xp5_ASAP7_75t_L g7613 ( 
.A1(n_6524),
.A2(n_5283),
.B(n_5297),
.Y(n_7613)
);

BUFx2_ASAP7_75t_L g7614 ( 
.A(n_6604),
.Y(n_7614)
);

INVx2_ASAP7_75t_SL g7615 ( 
.A(n_6701),
.Y(n_7615)
);

NOR2xp33_ASAP7_75t_L g7616 ( 
.A(n_6642),
.B(n_5760),
.Y(n_7616)
);

AOI21xp5_ASAP7_75t_L g7617 ( 
.A1(n_6403),
.A2(n_5328),
.B(n_5297),
.Y(n_7617)
);

OA21x2_ASAP7_75t_L g7618 ( 
.A1(n_6102),
.A2(n_5728),
.B(n_5723),
.Y(n_7618)
);

OAI22xp5_ASAP7_75t_L g7619 ( 
.A1(n_6554),
.A2(n_5328),
.B1(n_5443),
.B2(n_5297),
.Y(n_7619)
);

OAI21xp5_ASAP7_75t_L g7620 ( 
.A1(n_6451),
.A2(n_5465),
.B(n_5700),
.Y(n_7620)
);

OAI22xp5_ASAP7_75t_L g7621 ( 
.A1(n_6540),
.A2(n_5443),
.B1(n_5450),
.B2(n_5328),
.Y(n_7621)
);

NOR2x1_ASAP7_75t_R g7622 ( 
.A(n_6768),
.B(n_5538),
.Y(n_7622)
);

AOI21xp5_ASAP7_75t_L g7623 ( 
.A1(n_6500),
.A2(n_5450),
.B(n_5443),
.Y(n_7623)
);

AOI21xp5_ASAP7_75t_L g7624 ( 
.A1(n_6413),
.A2(n_5450),
.B(n_5443),
.Y(n_7624)
);

BUFx6f_ASAP7_75t_L g7625 ( 
.A(n_6249),
.Y(n_7625)
);

HB1xp67_ASAP7_75t_L g7626 ( 
.A(n_6236),
.Y(n_7626)
);

O2A1O1Ixp5_ASAP7_75t_L g7627 ( 
.A1(n_6100),
.A2(n_4806),
.B(n_5450),
.C(n_5443),
.Y(n_7627)
);

INVx8_ASAP7_75t_L g7628 ( 
.A(n_5908),
.Y(n_7628)
);

INVx2_ASAP7_75t_SL g7629 ( 
.A(n_6701),
.Y(n_7629)
);

OA21x2_ASAP7_75t_L g7630 ( 
.A1(n_6745),
.A2(n_5728),
.B(n_5723),
.Y(n_7630)
);

INVx2_ASAP7_75t_SL g7631 ( 
.A(n_6701),
.Y(n_7631)
);

HB1xp67_ASAP7_75t_L g7632 ( 
.A(n_6236),
.Y(n_7632)
);

AND2x4_ASAP7_75t_SL g7633 ( 
.A(n_6324),
.B(n_4568),
.Y(n_7633)
);

AOI22xp33_ASAP7_75t_L g7634 ( 
.A1(n_5774),
.A2(n_4987),
.B1(n_4991),
.B2(n_4980),
.Y(n_7634)
);

AOI21xp5_ASAP7_75t_L g7635 ( 
.A1(n_6413),
.A2(n_5703),
.B(n_5544),
.Y(n_7635)
);

NAND3xp33_ASAP7_75t_L g7636 ( 
.A(n_5787),
.B(n_4993),
.C(n_4991),
.Y(n_7636)
);

INVx1_ASAP7_75t_L g7637 ( 
.A(n_6160),
.Y(n_7637)
);

INVx1_ASAP7_75t_SL g7638 ( 
.A(n_6709),
.Y(n_7638)
);

A2O1A1Ixp33_ASAP7_75t_L g7639 ( 
.A1(n_6676),
.A2(n_5703),
.B(n_5544),
.C(n_4814),
.Y(n_7639)
);

OAI22xp5_ASAP7_75t_L g7640 ( 
.A1(n_6540),
.A2(n_6100),
.B1(n_6574),
.B2(n_6503),
.Y(n_7640)
);

A2O1A1Ixp33_ASAP7_75t_SL g7641 ( 
.A1(n_5807),
.A2(n_5589),
.B(n_5393),
.C(n_5725),
.Y(n_7641)
);

INVx1_ASAP7_75t_L g7642 ( 
.A(n_6160),
.Y(n_7642)
);

INVx1_ASAP7_75t_L g7643 ( 
.A(n_6166),
.Y(n_7643)
);

INVx1_ASAP7_75t_L g7644 ( 
.A(n_6166),
.Y(n_7644)
);

AOI21xp5_ASAP7_75t_L g7645 ( 
.A1(n_6497),
.A2(n_5703),
.B(n_5544),
.Y(n_7645)
);

OAI22xp33_ASAP7_75t_L g7646 ( 
.A1(n_5862),
.A2(n_5538),
.B1(n_5554),
.B2(n_5544),
.Y(n_7646)
);

INVx1_ASAP7_75t_L g7647 ( 
.A(n_6168),
.Y(n_7647)
);

AOI22xp33_ASAP7_75t_L g7648 ( 
.A1(n_6588),
.A2(n_6378),
.B1(n_6664),
.B2(n_6231),
.Y(n_7648)
);

INVx6_ASAP7_75t_L g7649 ( 
.A(n_6873),
.Y(n_7649)
);

CKINVDCx5p33_ASAP7_75t_R g7650 ( 
.A(n_6034),
.Y(n_7650)
);

BUFx2_ASAP7_75t_SL g7651 ( 
.A(n_6868),
.Y(n_7651)
);

NAND2xp5_ASAP7_75t_SL g7652 ( 
.A(n_6414),
.B(n_6457),
.Y(n_7652)
);

NAND2x1p5_ASAP7_75t_L g7653 ( 
.A(n_6333),
.B(n_5538),
.Y(n_7653)
);

OAI22xp5_ASAP7_75t_L g7654 ( 
.A1(n_6503),
.A2(n_5703),
.B1(n_4993),
.B2(n_5004),
.Y(n_7654)
);

INVx1_ASAP7_75t_L g7655 ( 
.A(n_6168),
.Y(n_7655)
);

AOI22xp33_ASAP7_75t_SL g7656 ( 
.A1(n_6233),
.A2(n_5534),
.B1(n_5523),
.B2(n_5508),
.Y(n_7656)
);

INVx1_ASAP7_75t_L g7657 ( 
.A(n_6173),
.Y(n_7657)
);

CKINVDCx5p33_ASAP7_75t_R g7658 ( 
.A(n_6037),
.Y(n_7658)
);

INVx5_ASAP7_75t_L g7659 ( 
.A(n_6333),
.Y(n_7659)
);

AOI21x1_ASAP7_75t_L g7660 ( 
.A1(n_6125),
.A2(n_5728),
.B(n_5763),
.Y(n_7660)
);

BUFx2_ASAP7_75t_L g7661 ( 
.A(n_6604),
.Y(n_7661)
);

OAI22xp5_ASAP7_75t_SL g7662 ( 
.A1(n_6003),
.A2(n_5365),
.B1(n_5414),
.B2(n_5382),
.Y(n_7662)
);

O2A1O1Ixp33_ASAP7_75t_L g7663 ( 
.A1(n_5793),
.A2(n_5761),
.B(n_5760),
.C(n_5426),
.Y(n_7663)
);

NOR2xp33_ASAP7_75t_SL g7664 ( 
.A(n_6868),
.B(n_5538),
.Y(n_7664)
);

INVx1_ASAP7_75t_L g7665 ( 
.A(n_6173),
.Y(n_7665)
);

INVx1_ASAP7_75t_L g7666 ( 
.A(n_6175),
.Y(n_7666)
);

NAND2xp5_ASAP7_75t_SL g7667 ( 
.A(n_6414),
.B(n_5365),
.Y(n_7667)
);

OR2x6_ASAP7_75t_L g7668 ( 
.A(n_6265),
.B(n_4894),
.Y(n_7668)
);

CKINVDCx5p33_ASAP7_75t_R g7669 ( 
.A(n_6085),
.Y(n_7669)
);

INVx1_ASAP7_75t_L g7670 ( 
.A(n_6175),
.Y(n_7670)
);

NAND2xp5_ASAP7_75t_L g7671 ( 
.A(n_6128),
.B(n_6213),
.Y(n_7671)
);

INVx1_ASAP7_75t_L g7672 ( 
.A(n_6179),
.Y(n_7672)
);

INVx1_ASAP7_75t_L g7673 ( 
.A(n_6179),
.Y(n_7673)
);

INVx1_ASAP7_75t_L g7674 ( 
.A(n_6187),
.Y(n_7674)
);

NOR2xp33_ASAP7_75t_L g7675 ( 
.A(n_6642),
.B(n_5761),
.Y(n_7675)
);

OR2x6_ASAP7_75t_L g7676 ( 
.A(n_6265),
.B(n_4894),
.Y(n_7676)
);

NAND2x1p5_ASAP7_75t_L g7677 ( 
.A(n_6333),
.B(n_5538),
.Y(n_7677)
);

AND2x2_ASAP7_75t_L g7678 ( 
.A(n_6603),
.B(n_6213),
.Y(n_7678)
);

INVx1_ASAP7_75t_L g7679 ( 
.A(n_6187),
.Y(n_7679)
);

A2O1A1Ixp33_ASAP7_75t_L g7680 ( 
.A1(n_5787),
.A2(n_4814),
.B(n_5652),
.C(n_5554),
.Y(n_7680)
);

INVx1_ASAP7_75t_L g7681 ( 
.A(n_6193),
.Y(n_7681)
);

AOI22xp33_ASAP7_75t_L g7682 ( 
.A1(n_6664),
.A2(n_4993),
.B1(n_5004),
.B2(n_4991),
.Y(n_7682)
);

AOI22xp5_ASAP7_75t_L g7683 ( 
.A1(n_5770),
.A2(n_5929),
.B1(n_5906),
.B2(n_5851),
.Y(n_7683)
);

OR2x6_ASAP7_75t_L g7684 ( 
.A(n_6658),
.B(n_4894),
.Y(n_7684)
);

AO21x2_ASAP7_75t_L g7685 ( 
.A1(n_6713),
.A2(n_6734),
.B(n_6717),
.Y(n_7685)
);

BUFx12f_ASAP7_75t_L g7686 ( 
.A(n_6768),
.Y(n_7686)
);

INVx1_ASAP7_75t_SL g7687 ( 
.A(n_6751),
.Y(n_7687)
);

INVx1_ASAP7_75t_L g7688 ( 
.A(n_6193),
.Y(n_7688)
);

INVx1_ASAP7_75t_L g7689 ( 
.A(n_6218),
.Y(n_7689)
);

INVx1_ASAP7_75t_L g7690 ( 
.A(n_6218),
.Y(n_7690)
);

INVx3_ASAP7_75t_SL g7691 ( 
.A(n_6082),
.Y(n_7691)
);

NAND2xp5_ASAP7_75t_SL g7692 ( 
.A(n_6457),
.B(n_5365),
.Y(n_7692)
);

INVx1_ASAP7_75t_SL g7693 ( 
.A(n_6751),
.Y(n_7693)
);

NOR2x1_ASAP7_75t_R g7694 ( 
.A(n_6080),
.B(n_5538),
.Y(n_7694)
);

BUFx2_ASAP7_75t_L g7695 ( 
.A(n_6604),
.Y(n_7695)
);

AOI21xp5_ASAP7_75t_L g7696 ( 
.A1(n_6444),
.A2(n_5554),
.B(n_5652),
.Y(n_7696)
);

AOI21xp5_ASAP7_75t_L g7697 ( 
.A1(n_6444),
.A2(n_5554),
.B(n_5652),
.Y(n_7697)
);

NOR2x1_ASAP7_75t_SL g7698 ( 
.A(n_6801),
.B(n_5554),
.Y(n_7698)
);

BUFx2_ASAP7_75t_L g7699 ( 
.A(n_6604),
.Y(n_7699)
);

INVx5_ASAP7_75t_L g7700 ( 
.A(n_6333),
.Y(n_7700)
);

AND2x4_ASAP7_75t_L g7701 ( 
.A(n_6887),
.B(n_6357),
.Y(n_7701)
);

NAND2xp5_ASAP7_75t_L g7702 ( 
.A(n_6214),
.B(n_6217),
.Y(n_7702)
);

HB1xp67_ASAP7_75t_L g7703 ( 
.A(n_6492),
.Y(n_7703)
);

OR2x6_ASAP7_75t_SL g7704 ( 
.A(n_6675),
.B(n_5547),
.Y(n_7704)
);

INVx6_ASAP7_75t_L g7705 ( 
.A(n_6873),
.Y(n_7705)
);

AND2x4_ASAP7_75t_L g7706 ( 
.A(n_6357),
.B(n_4568),
.Y(n_7706)
);

BUFx3_ASAP7_75t_L g7707 ( 
.A(n_6877),
.Y(n_7707)
);

HB1xp67_ASAP7_75t_L g7708 ( 
.A(n_6506),
.Y(n_7708)
);

INVx1_ASAP7_75t_L g7709 ( 
.A(n_6219),
.Y(n_7709)
);

OAI22xp5_ASAP7_75t_L g7710 ( 
.A1(n_6630),
.A2(n_5006),
.B1(n_5011),
.B2(n_5004),
.Y(n_7710)
);

BUFx6f_ASAP7_75t_L g7711 ( 
.A(n_6409),
.Y(n_7711)
);

HB1xp67_ASAP7_75t_L g7712 ( 
.A(n_6506),
.Y(n_7712)
);

OAI221xp5_ASAP7_75t_L g7713 ( 
.A1(n_5807),
.A2(n_5727),
.B1(n_5712),
.B2(n_5575),
.C(n_5037),
.Y(n_7713)
);

INVx1_ASAP7_75t_L g7714 ( 
.A(n_6219),
.Y(n_7714)
);

AOI22xp33_ASAP7_75t_L g7715 ( 
.A1(n_6229),
.A2(n_5011),
.B1(n_5037),
.B2(n_5006),
.Y(n_7715)
);

AOI21xp5_ASAP7_75t_L g7716 ( 
.A1(n_6477),
.A2(n_5554),
.B(n_5652),
.Y(n_7716)
);

AOI22xp5_ASAP7_75t_L g7717 ( 
.A1(n_5906),
.A2(n_5929),
.B1(n_5851),
.B2(n_6388),
.Y(n_7717)
);

BUFx2_ASAP7_75t_L g7718 ( 
.A(n_6604),
.Y(n_7718)
);

BUFx6f_ASAP7_75t_L g7719 ( 
.A(n_6409),
.Y(n_7719)
);

INVx4_ASAP7_75t_L g7720 ( 
.A(n_5978),
.Y(n_7720)
);

CKINVDCx5p33_ASAP7_75t_R g7721 ( 
.A(n_6186),
.Y(n_7721)
);

OR2x6_ASAP7_75t_L g7722 ( 
.A(n_6658),
.B(n_4814),
.Y(n_7722)
);

NAND2xp5_ASAP7_75t_L g7723 ( 
.A(n_6217),
.B(n_6243),
.Y(n_7723)
);

INVx1_ASAP7_75t_L g7724 ( 
.A(n_6220),
.Y(n_7724)
);

BUFx6f_ASAP7_75t_L g7725 ( 
.A(n_6409),
.Y(n_7725)
);

OAI22xp5_ASAP7_75t_L g7726 ( 
.A1(n_6630),
.A2(n_5011),
.B1(n_5037),
.B2(n_5006),
.Y(n_7726)
);

BUFx2_ASAP7_75t_L g7727 ( 
.A(n_6622),
.Y(n_7727)
);

CKINVDCx5p33_ASAP7_75t_R g7728 ( 
.A(n_6190),
.Y(n_7728)
);

NAND2xp5_ASAP7_75t_L g7729 ( 
.A(n_6243),
.B(n_6244),
.Y(n_7729)
);

INVx1_ASAP7_75t_L g7730 ( 
.A(n_6220),
.Y(n_7730)
);

AOI22xp5_ASAP7_75t_L g7731 ( 
.A1(n_6388),
.A2(n_5534),
.B1(n_5053),
.B2(n_5054),
.Y(n_7731)
);

AOI221xp5_ASAP7_75t_L g7732 ( 
.A1(n_6274),
.A2(n_5054),
.B1(n_5058),
.B2(n_5053),
.C(n_5047),
.Y(n_7732)
);

CKINVDCx5p33_ASAP7_75t_R g7733 ( 
.A(n_6550),
.Y(n_7733)
);

CKINVDCx6p67_ASAP7_75t_R g7734 ( 
.A(n_6063),
.Y(n_7734)
);

INVx1_ASAP7_75t_SL g7735 ( 
.A(n_6756),
.Y(n_7735)
);

BUFx6f_ASAP7_75t_L g7736 ( 
.A(n_6409),
.Y(n_7736)
);

O2A1O1Ixp33_ASAP7_75t_L g7737 ( 
.A1(n_6274),
.A2(n_5499),
.B(n_5699),
.C(n_5426),
.Y(n_7737)
);

AND2x4_ASAP7_75t_L g7738 ( 
.A(n_6357),
.B(n_4568),
.Y(n_7738)
);

CKINVDCx11_ASAP7_75t_R g7739 ( 
.A(n_6893),
.Y(n_7739)
);

INVx1_ASAP7_75t_L g7740 ( 
.A(n_6222),
.Y(n_7740)
);

AOI22xp33_ASAP7_75t_L g7741 ( 
.A1(n_6229),
.A2(n_5053),
.B1(n_5054),
.B2(n_5047),
.Y(n_7741)
);

BUFx3_ASAP7_75t_L g7742 ( 
.A(n_6877),
.Y(n_7742)
);

BUFx3_ASAP7_75t_L g7743 ( 
.A(n_6877),
.Y(n_7743)
);

INVx8_ASAP7_75t_L g7744 ( 
.A(n_5908),
.Y(n_7744)
);

AOI22xp5_ASAP7_75t_L g7745 ( 
.A1(n_6231),
.A2(n_5534),
.B1(n_5058),
.B2(n_5059),
.Y(n_7745)
);

INVx1_ASAP7_75t_L g7746 ( 
.A(n_6222),
.Y(n_7746)
);

INVx4_ASAP7_75t_L g7747 ( 
.A(n_5978),
.Y(n_7747)
);

NAND2x1p5_ASAP7_75t_L g7748 ( 
.A(n_6409),
.B(n_5554),
.Y(n_7748)
);

INVx1_ASAP7_75t_L g7749 ( 
.A(n_6223),
.Y(n_7749)
);

AOI22xp5_ASAP7_75t_L g7750 ( 
.A1(n_6240),
.A2(n_5534),
.B1(n_5058),
.B2(n_5059),
.Y(n_7750)
);

BUFx2_ASAP7_75t_L g7751 ( 
.A(n_6622),
.Y(n_7751)
);

HB1xp67_ASAP7_75t_L g7752 ( 
.A(n_5989),
.Y(n_7752)
);

AOI22xp33_ASAP7_75t_L g7753 ( 
.A1(n_6485),
.A2(n_5059),
.B1(n_5060),
.B2(n_5047),
.Y(n_7753)
);

INVx1_ASAP7_75t_L g7754 ( 
.A(n_6223),
.Y(n_7754)
);

A2O1A1Ixp33_ASAP7_75t_L g7755 ( 
.A1(n_5855),
.A2(n_5554),
.B(n_5742),
.C(n_5730),
.Y(n_7755)
);

NOR2xp33_ASAP7_75t_L g7756 ( 
.A(n_5790),
.B(n_5561),
.Y(n_7756)
);

BUFx3_ASAP7_75t_L g7757 ( 
.A(n_6462),
.Y(n_7757)
);

OAI21x1_ASAP7_75t_L g7758 ( 
.A1(n_6745),
.A2(n_4874),
.B(n_4865),
.Y(n_7758)
);

AOI22xp33_ASAP7_75t_L g7759 ( 
.A1(n_6485),
.A2(n_5063),
.B1(n_5064),
.B2(n_5060),
.Y(n_7759)
);

AOI22xp33_ASAP7_75t_L g7760 ( 
.A1(n_5820),
.A2(n_6562),
.B1(n_6233),
.B2(n_6422),
.Y(n_7760)
);

INVx1_ASAP7_75t_L g7761 ( 
.A(n_6235),
.Y(n_7761)
);

OAI22xp5_ASAP7_75t_L g7762 ( 
.A1(n_6177),
.A2(n_5063),
.B1(n_5064),
.B2(n_5060),
.Y(n_7762)
);

CKINVDCx6p67_ASAP7_75t_R g7763 ( 
.A(n_6063),
.Y(n_7763)
);

AOI22xp33_ASAP7_75t_L g7764 ( 
.A1(n_5820),
.A2(n_5064),
.B1(n_5068),
.B2(n_5063),
.Y(n_7764)
);

INVx1_ASAP7_75t_L g7765 ( 
.A(n_6235),
.Y(n_7765)
);

BUFx2_ASAP7_75t_L g7766 ( 
.A(n_6622),
.Y(n_7766)
);

BUFx2_ASAP7_75t_L g7767 ( 
.A(n_6622),
.Y(n_7767)
);

AOI22xp33_ASAP7_75t_L g7768 ( 
.A1(n_6562),
.A2(n_5083),
.B1(n_5086),
.B2(n_5068),
.Y(n_7768)
);

CKINVDCx20_ASAP7_75t_R g7769 ( 
.A(n_6453),
.Y(n_7769)
);

NAND2xp5_ASAP7_75t_SL g7770 ( 
.A(n_6470),
.B(n_5365),
.Y(n_7770)
);

INVx1_ASAP7_75t_L g7771 ( 
.A(n_6239),
.Y(n_7771)
);

NAND2xp5_ASAP7_75t_L g7772 ( 
.A(n_6252),
.B(n_6267),
.Y(n_7772)
);

AOI221xp5_ASAP7_75t_L g7773 ( 
.A1(n_6571),
.A2(n_5086),
.B1(n_5087),
.B2(n_5083),
.C(n_5068),
.Y(n_7773)
);

AND2x2_ASAP7_75t_SL g7774 ( 
.A(n_6502),
.B(n_5365),
.Y(n_7774)
);

OAI22xp5_ASAP7_75t_L g7775 ( 
.A1(n_6637),
.A2(n_5086),
.B1(n_5087),
.B2(n_5083),
.Y(n_7775)
);

INVx5_ASAP7_75t_L g7776 ( 
.A(n_6442),
.Y(n_7776)
);

AND2x4_ASAP7_75t_L g7777 ( 
.A(n_6357),
.B(n_4568),
.Y(n_7777)
);

AOI21xp5_ASAP7_75t_L g7778 ( 
.A1(n_6527),
.A2(n_5742),
.B(n_5730),
.Y(n_7778)
);

HB1xp67_ASAP7_75t_L g7779 ( 
.A(n_5989),
.Y(n_7779)
);

INVx5_ASAP7_75t_L g7780 ( 
.A(n_6442),
.Y(n_7780)
);

AND2x4_ASAP7_75t_L g7781 ( 
.A(n_6357),
.B(n_4568),
.Y(n_7781)
);

AND2x2_ASAP7_75t_L g7782 ( 
.A(n_6319),
.B(n_6507),
.Y(n_7782)
);

AOI22xp5_ASAP7_75t_L g7783 ( 
.A1(n_6240),
.A2(n_5534),
.B1(n_5091),
.B2(n_5102),
.Y(n_7783)
);

BUFx12f_ASAP7_75t_L g7784 ( 
.A(n_6900),
.Y(n_7784)
);

BUFx12f_ASAP7_75t_L g7785 ( 
.A(n_6878),
.Y(n_7785)
);

OAI22xp5_ASAP7_75t_L g7786 ( 
.A1(n_6637),
.A2(n_5091),
.B1(n_5102),
.B2(n_5087),
.Y(n_7786)
);

NOR2xp33_ASAP7_75t_L g7787 ( 
.A(n_5790),
.B(n_5563),
.Y(n_7787)
);

INVx1_ASAP7_75t_L g7788 ( 
.A(n_6239),
.Y(n_7788)
);

AOI21xp33_ASAP7_75t_L g7789 ( 
.A1(n_6679),
.A2(n_5727),
.B(n_5712),
.Y(n_7789)
);

BUFx3_ASAP7_75t_L g7790 ( 
.A(n_6462),
.Y(n_7790)
);

NOR2xp33_ASAP7_75t_L g7791 ( 
.A(n_6418),
.B(n_5563),
.Y(n_7791)
);

BUFx3_ASAP7_75t_L g7792 ( 
.A(n_6462),
.Y(n_7792)
);

BUFx2_ASAP7_75t_L g7793 ( 
.A(n_6622),
.Y(n_7793)
);

INVx1_ASAP7_75t_L g7794 ( 
.A(n_6251),
.Y(n_7794)
);

INVx5_ASAP7_75t_L g7795 ( 
.A(n_6442),
.Y(n_7795)
);

INVx1_ASAP7_75t_L g7796 ( 
.A(n_6251),
.Y(n_7796)
);

INVx3_ASAP7_75t_L g7797 ( 
.A(n_6895),
.Y(n_7797)
);

INVx4_ASAP7_75t_SL g7798 ( 
.A(n_6396),
.Y(n_7798)
);

OAI21xp5_ASAP7_75t_L g7799 ( 
.A1(n_6017),
.A2(n_5727),
.B(n_5709),
.Y(n_7799)
);

NAND3xp33_ASAP7_75t_SL g7800 ( 
.A(n_5838),
.B(n_5567),
.C(n_5565),
.Y(n_7800)
);

INVx8_ASAP7_75t_L g7801 ( 
.A(n_5917),
.Y(n_7801)
);

NAND2x1p5_ASAP7_75t_L g7802 ( 
.A(n_6442),
.B(n_4865),
.Y(n_7802)
);

BUFx6f_ASAP7_75t_L g7803 ( 
.A(n_6442),
.Y(n_7803)
);

BUFx4_ASAP7_75t_SL g7804 ( 
.A(n_6583),
.Y(n_7804)
);

AND2x2_ASAP7_75t_SL g7805 ( 
.A(n_6502),
.B(n_5382),
.Y(n_7805)
);

BUFx3_ASAP7_75t_L g7806 ( 
.A(n_6462),
.Y(n_7806)
);

AOI21xp5_ASAP7_75t_L g7807 ( 
.A1(n_6448),
.A2(n_5742),
.B(n_5730),
.Y(n_7807)
);

BUFx2_ASAP7_75t_L g7808 ( 
.A(n_6622),
.Y(n_7808)
);

CKINVDCx8_ASAP7_75t_R g7809 ( 
.A(n_6376),
.Y(n_7809)
);

INVx1_ASAP7_75t_SL g7810 ( 
.A(n_6756),
.Y(n_7810)
);

NOR2xp33_ASAP7_75t_L g7811 ( 
.A(n_6418),
.B(n_5565),
.Y(n_7811)
);

AOI22xp33_ASAP7_75t_L g7812 ( 
.A1(n_6422),
.A2(n_5102),
.B1(n_5124),
.B2(n_5091),
.Y(n_7812)
);

INVx3_ASAP7_75t_L g7813 ( 
.A(n_6895),
.Y(n_7813)
);

AOI21xp5_ASAP7_75t_L g7814 ( 
.A1(n_6448),
.A2(n_5742),
.B(n_5730),
.Y(n_7814)
);

INVx1_ASAP7_75t_L g7815 ( 
.A(n_6253),
.Y(n_7815)
);

NOR2xp33_ASAP7_75t_SL g7816 ( 
.A(n_6859),
.B(n_4674),
.Y(n_7816)
);

OAI21x1_ASAP7_75t_L g7817 ( 
.A1(n_6517),
.A2(n_4874),
.B(n_4865),
.Y(n_7817)
);

INVx1_ASAP7_75t_L g7818 ( 
.A(n_6253),
.Y(n_7818)
);

INVx3_ASAP7_75t_L g7819 ( 
.A(n_6895),
.Y(n_7819)
);

NOR2xp67_ASAP7_75t_L g7820 ( 
.A(n_6442),
.B(n_5731),
.Y(n_7820)
);

INVx3_ASAP7_75t_L g7821 ( 
.A(n_6895),
.Y(n_7821)
);

OAI22x1_ASAP7_75t_L g7822 ( 
.A1(n_6199),
.A2(n_5126),
.B1(n_5146),
.B2(n_5124),
.Y(n_7822)
);

CKINVDCx5p33_ASAP7_75t_R g7823 ( 
.A(n_6080),
.Y(n_7823)
);

INVx1_ASAP7_75t_SL g7824 ( 
.A(n_6904),
.Y(n_7824)
);

INVx1_ASAP7_75t_L g7825 ( 
.A(n_6269),
.Y(n_7825)
);

NAND2xp5_ASAP7_75t_L g7826 ( 
.A(n_6347),
.B(n_5568),
.Y(n_7826)
);

NOR2xp33_ASAP7_75t_L g7827 ( 
.A(n_6428),
.B(n_5568),
.Y(n_7827)
);

NAND2xp5_ASAP7_75t_L g7828 ( 
.A(n_6347),
.B(n_6350),
.Y(n_7828)
);

CKINVDCx5p33_ASAP7_75t_R g7829 ( 
.A(n_6080),
.Y(n_7829)
);

CKINVDCx20_ASAP7_75t_R g7830 ( 
.A(n_6583),
.Y(n_7830)
);

AOI22xp33_ASAP7_75t_L g7831 ( 
.A1(n_6428),
.A2(n_5126),
.B1(n_5146),
.B2(n_5124),
.Y(n_7831)
);

OAI22xp5_ASAP7_75t_L g7832 ( 
.A1(n_6510),
.A2(n_5146),
.B1(n_5152),
.B2(n_5126),
.Y(n_7832)
);

O2A1O1Ixp5_ASAP7_75t_SL g7833 ( 
.A1(n_6320),
.A2(n_5696),
.B(n_5698),
.C(n_5695),
.Y(n_7833)
);

AOI22xp33_ASAP7_75t_L g7834 ( 
.A1(n_5893),
.A2(n_5153),
.B1(n_5155),
.B2(n_5152),
.Y(n_7834)
);

INVx1_ASAP7_75t_L g7835 ( 
.A(n_6269),
.Y(n_7835)
);

NAND2xp5_ASAP7_75t_L g7836 ( 
.A(n_6350),
.B(n_5570),
.Y(n_7836)
);

BUFx3_ASAP7_75t_L g7837 ( 
.A(n_6462),
.Y(n_7837)
);

BUFx2_ASAP7_75t_L g7838 ( 
.A(n_6626),
.Y(n_7838)
);

AOI22xp5_ASAP7_75t_L g7839 ( 
.A1(n_6258),
.A2(n_5153),
.B1(n_5155),
.B2(n_5152),
.Y(n_7839)
);

AND2x4_ASAP7_75t_L g7840 ( 
.A(n_6153),
.B(n_6167),
.Y(n_7840)
);

INVx3_ASAP7_75t_L g7841 ( 
.A(n_6898),
.Y(n_7841)
);

INVx1_ASAP7_75t_L g7842 ( 
.A(n_6280),
.Y(n_7842)
);

NAND2xp5_ASAP7_75t_L g7843 ( 
.A(n_6381),
.B(n_5570),
.Y(n_7843)
);

INVx1_ASAP7_75t_L g7844 ( 
.A(n_6280),
.Y(n_7844)
);

INVx1_ASAP7_75t_L g7845 ( 
.A(n_6298),
.Y(n_7845)
);

OAI21x1_ASAP7_75t_L g7846 ( 
.A1(n_6520),
.A2(n_4874),
.B(n_4865),
.Y(n_7846)
);

NAND2xp5_ASAP7_75t_L g7847 ( 
.A(n_6381),
.B(n_5153),
.Y(n_7847)
);

CKINVDCx5p33_ASAP7_75t_R g7848 ( 
.A(n_6087),
.Y(n_7848)
);

INVx1_ASAP7_75t_L g7849 ( 
.A(n_6298),
.Y(n_7849)
);

INVx3_ASAP7_75t_L g7850 ( 
.A(n_6898),
.Y(n_7850)
);

BUFx3_ASAP7_75t_L g7851 ( 
.A(n_6686),
.Y(n_7851)
);

NAND2xp5_ASAP7_75t_L g7852 ( 
.A(n_6412),
.B(n_5155),
.Y(n_7852)
);

INVx1_ASAP7_75t_L g7853 ( 
.A(n_6305),
.Y(n_7853)
);

OAI22xp5_ASAP7_75t_L g7854 ( 
.A1(n_6510),
.A2(n_5175),
.B1(n_5177),
.B2(n_5156),
.Y(n_7854)
);

BUFx3_ASAP7_75t_L g7855 ( 
.A(n_6686),
.Y(n_7855)
);

OAI22xp5_ASAP7_75t_L g7856 ( 
.A1(n_6424),
.A2(n_5175),
.B1(n_5177),
.B2(n_5156),
.Y(n_7856)
);

INVx5_ASAP7_75t_L g7857 ( 
.A(n_6532),
.Y(n_7857)
);

INVx1_ASAP7_75t_L g7858 ( 
.A(n_6305),
.Y(n_7858)
);

INVx1_ASAP7_75t_SL g7859 ( 
.A(n_6904),
.Y(n_7859)
);

AOI22xp33_ASAP7_75t_L g7860 ( 
.A1(n_5893),
.A2(n_5175),
.B1(n_5177),
.B2(n_5156),
.Y(n_7860)
);

INVx1_ASAP7_75t_L g7861 ( 
.A(n_6313),
.Y(n_7861)
);

INVx3_ASAP7_75t_L g7862 ( 
.A(n_6898),
.Y(n_7862)
);

INVx1_ASAP7_75t_L g7863 ( 
.A(n_6313),
.Y(n_7863)
);

INVxp67_ASAP7_75t_SL g7864 ( 
.A(n_6519),
.Y(n_7864)
);

INVxp67_ASAP7_75t_L g7865 ( 
.A(n_6073),
.Y(n_7865)
);

OAI21xp33_ASAP7_75t_L g7866 ( 
.A1(n_6392),
.A2(n_5191),
.B(n_5181),
.Y(n_7866)
);

INVx5_ASAP7_75t_L g7867 ( 
.A(n_6532),
.Y(n_7867)
);

INVx4_ASAP7_75t_SL g7868 ( 
.A(n_6396),
.Y(n_7868)
);

OAI22xp5_ASAP7_75t_L g7869 ( 
.A1(n_6424),
.A2(n_5191),
.B1(n_5194),
.B2(n_5181),
.Y(n_7869)
);

NAND2xp5_ASAP7_75t_L g7870 ( 
.A(n_6412),
.B(n_5181),
.Y(n_7870)
);

O2A1O1Ixp33_ASAP7_75t_L g7871 ( 
.A1(n_5803),
.A2(n_5499),
.B(n_5699),
.C(n_5426),
.Y(n_7871)
);

AOI22xp5_ASAP7_75t_L g7872 ( 
.A1(n_6258),
.A2(n_6286),
.B1(n_6304),
.B2(n_6292),
.Y(n_7872)
);

NOR2xp33_ASAP7_75t_L g7873 ( 
.A(n_5961),
.B(n_5731),
.Y(n_7873)
);

BUFx2_ASAP7_75t_L g7874 ( 
.A(n_6626),
.Y(n_7874)
);

INVx1_ASAP7_75t_L g7875 ( 
.A(n_6322),
.Y(n_7875)
);

CKINVDCx5p33_ASAP7_75t_R g7876 ( 
.A(n_6087),
.Y(n_7876)
);

BUFx12f_ASAP7_75t_L g7877 ( 
.A(n_6087),
.Y(n_7877)
);

INVx1_ASAP7_75t_L g7878 ( 
.A(n_6322),
.Y(n_7878)
);

AOI21xp5_ASAP7_75t_L g7879 ( 
.A1(n_6527),
.A2(n_5742),
.B(n_5730),
.Y(n_7879)
);

INVx3_ASAP7_75t_L g7880 ( 
.A(n_6898),
.Y(n_7880)
);

BUFx2_ASAP7_75t_L g7881 ( 
.A(n_6626),
.Y(n_7881)
);

INVx1_ASAP7_75t_L g7882 ( 
.A(n_6325),
.Y(n_7882)
);

INVx1_ASAP7_75t_L g7883 ( 
.A(n_6325),
.Y(n_7883)
);

INVx3_ASAP7_75t_L g7884 ( 
.A(n_6898),
.Y(n_7884)
);

INVx1_ASAP7_75t_L g7885 ( 
.A(n_6327),
.Y(n_7885)
);

INVx1_ASAP7_75t_L g7886 ( 
.A(n_6327),
.Y(n_7886)
);

BUFx2_ASAP7_75t_L g7887 ( 
.A(n_6626),
.Y(n_7887)
);

BUFx2_ASAP7_75t_L g7888 ( 
.A(n_6626),
.Y(n_7888)
);

AOI21xp5_ASAP7_75t_L g7889 ( 
.A1(n_6529),
.A2(n_5775),
.B(n_6740),
.Y(n_7889)
);

AOI22xp5_ASAP7_75t_L g7890 ( 
.A1(n_6286),
.A2(n_5196),
.B1(n_5207),
.B2(n_5194),
.Y(n_7890)
);

OAI21xp5_ASAP7_75t_L g7891 ( 
.A1(n_6017),
.A2(n_6169),
.B(n_6057),
.Y(n_7891)
);

NAND3xp33_ASAP7_75t_SL g7892 ( 
.A(n_5838),
.B(n_5763),
.C(n_5741),
.Y(n_7892)
);

BUFx2_ASAP7_75t_L g7893 ( 
.A(n_6626),
.Y(n_7893)
);

BUFx3_ASAP7_75t_L g7894 ( 
.A(n_6686),
.Y(n_7894)
);

NOR2xp33_ASAP7_75t_R g7895 ( 
.A(n_6593),
.B(n_5276),
.Y(n_7895)
);

AOI21x1_ASAP7_75t_L g7896 ( 
.A1(n_6125),
.A2(n_5763),
.B(n_5741),
.Y(n_7896)
);

INVx3_ASAP7_75t_L g7897 ( 
.A(n_6905),
.Y(n_7897)
);

NAND2x1p5_ASAP7_75t_L g7898 ( 
.A(n_6532),
.B(n_4865),
.Y(n_7898)
);

BUFx2_ASAP7_75t_L g7899 ( 
.A(n_6628),
.Y(n_7899)
);

AOI22xp33_ASAP7_75t_L g7900 ( 
.A1(n_5926),
.A2(n_5207),
.B1(n_5216),
.B2(n_5196),
.Y(n_7900)
);

AOI22xp33_ASAP7_75t_L g7901 ( 
.A1(n_5926),
.A2(n_5216),
.B1(n_5230),
.B2(n_5207),
.Y(n_7901)
);

INVx1_ASAP7_75t_L g7902 ( 
.A(n_6331),
.Y(n_7902)
);

INVx5_ASAP7_75t_L g7903 ( 
.A(n_6532),
.Y(n_7903)
);

O2A1O1Ixp33_ASAP7_75t_SL g7904 ( 
.A1(n_6573),
.A2(n_4580),
.B(n_4631),
.C(n_4572),
.Y(n_7904)
);

BUFx3_ASAP7_75t_L g7905 ( 
.A(n_6686),
.Y(n_7905)
);

AOI22xp5_ASAP7_75t_L g7906 ( 
.A1(n_6292),
.A2(n_5232),
.B1(n_5238),
.B2(n_5230),
.Y(n_7906)
);

OAI21x1_ASAP7_75t_L g7907 ( 
.A1(n_7415),
.A2(n_6529),
.B(n_6805),
.Y(n_7907)
);

OAI21x1_ASAP7_75t_L g7908 ( 
.A1(n_7415),
.A2(n_7235),
.B(n_7233),
.Y(n_7908)
);

A2O1A1Ixp33_ASAP7_75t_L g7909 ( 
.A1(n_7275),
.A2(n_6897),
.B(n_6711),
.C(n_6717),
.Y(n_7909)
);

INVx1_ASAP7_75t_L g7910 ( 
.A(n_7637),
.Y(n_7910)
);

INVx1_ASAP7_75t_L g7911 ( 
.A(n_7637),
.Y(n_7911)
);

OA21x2_ASAP7_75t_L g7912 ( 
.A1(n_7233),
.A2(n_6711),
.B(n_6897),
.Y(n_7912)
);

OAI22xp33_ASAP7_75t_L g7913 ( 
.A1(n_7092),
.A2(n_5862),
.B1(n_6401),
.B2(n_5872),
.Y(n_7913)
);

AND2x4_ASAP7_75t_L g7914 ( 
.A(n_7518),
.B(n_6618),
.Y(n_7914)
);

NOR2xp33_ASAP7_75t_L g7915 ( 
.A(n_7022),
.B(n_6304),
.Y(n_7915)
);

INVx2_ASAP7_75t_SL g7916 ( 
.A(n_7431),
.Y(n_7916)
);

INVx2_ASAP7_75t_L g7917 ( 
.A(n_6931),
.Y(n_7917)
);

INVx1_ASAP7_75t_L g7918 ( 
.A(n_7637),
.Y(n_7918)
);

AOI22xp5_ASAP7_75t_L g7919 ( 
.A1(n_7275),
.A2(n_6655),
.B1(n_5803),
.B2(n_6308),
.Y(n_7919)
);

OAI21x1_ASAP7_75t_L g7920 ( 
.A1(n_7415),
.A2(n_6805),
.B(n_6825),
.Y(n_7920)
);

INVx2_ASAP7_75t_SL g7921 ( 
.A(n_7431),
.Y(n_7921)
);

OAI21xp5_ASAP7_75t_L g7922 ( 
.A1(n_7261),
.A2(n_6057),
.B(n_6017),
.Y(n_7922)
);

BUFx3_ASAP7_75t_L g7923 ( 
.A(n_7433),
.Y(n_7923)
);

INVx1_ASAP7_75t_L g7924 ( 
.A(n_7642),
.Y(n_7924)
);

OAI21xp5_ASAP7_75t_L g7925 ( 
.A1(n_7261),
.A2(n_6169),
.B(n_6057),
.Y(n_7925)
);

BUFx6f_ASAP7_75t_L g7926 ( 
.A(n_6940),
.Y(n_7926)
);

AOI22xp33_ASAP7_75t_L g7927 ( 
.A1(n_7092),
.A2(n_7071),
.B1(n_7217),
.B2(n_7022),
.Y(n_7927)
);

OA21x2_ASAP7_75t_L g7928 ( 
.A1(n_7235),
.A2(n_7257),
.B(n_7239),
.Y(n_7928)
);

NAND3xp33_ASAP7_75t_SL g7929 ( 
.A(n_7071),
.B(n_6655),
.C(n_6679),
.Y(n_7929)
);

INVx2_ASAP7_75t_L g7930 ( 
.A(n_6931),
.Y(n_7930)
);

AOI22xp5_ASAP7_75t_L g7931 ( 
.A1(n_7262),
.A2(n_6308),
.B1(n_5769),
.B2(n_5850),
.Y(n_7931)
);

OAI21x1_ASAP7_75t_L g7932 ( 
.A1(n_7415),
.A2(n_6805),
.B(n_6825),
.Y(n_7932)
);

CKINVDCx5p33_ASAP7_75t_R g7933 ( 
.A(n_7194),
.Y(n_7933)
);

BUFx3_ASAP7_75t_L g7934 ( 
.A(n_7433),
.Y(n_7934)
);

NAND2xp5_ASAP7_75t_L g7935 ( 
.A(n_6989),
.B(n_6507),
.Y(n_7935)
);

CKINVDCx5p33_ASAP7_75t_R g7936 ( 
.A(n_7194),
.Y(n_7936)
);

NAND2xp5_ASAP7_75t_L g7937 ( 
.A(n_6989),
.B(n_6992),
.Y(n_7937)
);

CKINVDCx16_ASAP7_75t_R g7938 ( 
.A(n_7219),
.Y(n_7938)
);

AOI22xp5_ASAP7_75t_L g7939 ( 
.A1(n_7262),
.A2(n_7092),
.B1(n_7217),
.B2(n_7137),
.Y(n_7939)
);

OA21x2_ASAP7_75t_L g7940 ( 
.A1(n_7239),
.A2(n_6615),
.B(n_6623),
.Y(n_7940)
);

AND2x2_ASAP7_75t_L g7941 ( 
.A(n_6907),
.B(n_6548),
.Y(n_7941)
);

NAND2x1p5_ASAP7_75t_L g7942 ( 
.A(n_7431),
.B(n_6532),
.Y(n_7942)
);

OA21x2_ASAP7_75t_L g7943 ( 
.A1(n_7257),
.A2(n_6615),
.B(n_6623),
.Y(n_7943)
);

INVxp67_ASAP7_75t_SL g7944 ( 
.A(n_7152),
.Y(n_7944)
);

AOI221xp5_ASAP7_75t_L g7945 ( 
.A1(n_7052),
.A2(n_6392),
.B1(n_6688),
.B2(n_6725),
.C(n_6537),
.Y(n_7945)
);

AND2x2_ASAP7_75t_L g7946 ( 
.A(n_6907),
.B(n_6548),
.Y(n_7946)
);

CKINVDCx5p33_ASAP7_75t_R g7947 ( 
.A(n_7330),
.Y(n_7947)
);

AND2x4_ASAP7_75t_L g7948 ( 
.A(n_7518),
.B(n_6618),
.Y(n_7948)
);

OA21x2_ASAP7_75t_L g7949 ( 
.A1(n_7266),
.A2(n_6638),
.B(n_6713),
.Y(n_7949)
);

AOI21xp5_ASAP7_75t_L g7950 ( 
.A1(n_7889),
.A2(n_5775),
.B(n_6740),
.Y(n_7950)
);

AOI21x1_ASAP7_75t_L g7951 ( 
.A1(n_6995),
.A2(n_6884),
.B(n_5890),
.Y(n_7951)
);

OAI21xp5_ASAP7_75t_L g7952 ( 
.A1(n_7276),
.A2(n_7052),
.B(n_7386),
.Y(n_7952)
);

INVx2_ASAP7_75t_L g7953 ( 
.A(n_6931),
.Y(n_7953)
);

OAI21x1_ASAP7_75t_L g7954 ( 
.A1(n_7266),
.A2(n_7290),
.B(n_7284),
.Y(n_7954)
);

OAI21x1_ASAP7_75t_L g7955 ( 
.A1(n_7284),
.A2(n_6825),
.B(n_6782),
.Y(n_7955)
);

OA21x2_ASAP7_75t_L g7956 ( 
.A1(n_7290),
.A2(n_6638),
.B(n_6734),
.Y(n_7956)
);

NAND2xp5_ASAP7_75t_SL g7957 ( 
.A(n_7219),
.B(n_6823),
.Y(n_7957)
);

INVx1_ASAP7_75t_L g7958 ( 
.A(n_7642),
.Y(n_7958)
);

OAI21x1_ASAP7_75t_L g7959 ( 
.A1(n_7292),
.A2(n_6782),
.B(n_6226),
.Y(n_7959)
);

AOI22xp33_ASAP7_75t_L g7960 ( 
.A1(n_7298),
.A2(n_6349),
.B1(n_6323),
.B2(n_6563),
.Y(n_7960)
);

INVx4_ASAP7_75t_L g7961 ( 
.A(n_7309),
.Y(n_7961)
);

OAI21x1_ASAP7_75t_L g7962 ( 
.A1(n_7292),
.A2(n_6782),
.B(n_6226),
.Y(n_7962)
);

NAND2xp5_ASAP7_75t_L g7963 ( 
.A(n_6989),
.B(n_6548),
.Y(n_7963)
);

OAI21x1_ASAP7_75t_L g7964 ( 
.A1(n_7297),
.A2(n_6226),
.B(n_6334),
.Y(n_7964)
);

INVx1_ASAP7_75t_L g7965 ( 
.A(n_7642),
.Y(n_7965)
);

AND2x2_ASAP7_75t_L g7966 ( 
.A(n_6907),
.B(n_6549),
.Y(n_7966)
);

INVx2_ASAP7_75t_L g7967 ( 
.A(n_6931),
.Y(n_7967)
);

O2A1O1Ixp33_ASAP7_75t_L g7968 ( 
.A1(n_7107),
.A2(n_6380),
.B(n_5915),
.C(n_6737),
.Y(n_7968)
);

NAND2xp33_ASAP7_75t_L g7969 ( 
.A(n_7386),
.B(n_6854),
.Y(n_7969)
);

OA21x2_ASAP7_75t_L g7970 ( 
.A1(n_7297),
.A2(n_6773),
.B(n_6737),
.Y(n_7970)
);

BUFx2_ASAP7_75t_SL g7971 ( 
.A(n_7431),
.Y(n_7971)
);

INVx1_ASAP7_75t_L g7972 ( 
.A(n_7643),
.Y(n_7972)
);

AO21x2_ASAP7_75t_L g7973 ( 
.A1(n_7891),
.A2(n_6227),
.B(n_6773),
.Y(n_7973)
);

OA21x2_ASAP7_75t_L g7974 ( 
.A1(n_7312),
.A2(n_6591),
.B(n_6227),
.Y(n_7974)
);

NOR2xp33_ASAP7_75t_L g7975 ( 
.A(n_7276),
.B(n_6318),
.Y(n_7975)
);

AOI22xp33_ASAP7_75t_L g7976 ( 
.A1(n_7298),
.A2(n_6349),
.B1(n_6323),
.B2(n_6563),
.Y(n_7976)
);

OAI22xp5_ASAP7_75t_L g7977 ( 
.A1(n_7419),
.A2(n_6401),
.B1(n_6844),
.B2(n_6575),
.Y(n_7977)
);

INVx2_ASAP7_75t_L g7978 ( 
.A(n_6941),
.Y(n_7978)
);

HB1xp67_ASAP7_75t_L g7979 ( 
.A(n_7152),
.Y(n_7979)
);

OA21x2_ASAP7_75t_L g7980 ( 
.A1(n_7312),
.A2(n_7344),
.B(n_7333),
.Y(n_7980)
);

AND2x2_ASAP7_75t_L g7981 ( 
.A(n_6907),
.B(n_6549),
.Y(n_7981)
);

OAI22xp5_ASAP7_75t_L g7982 ( 
.A1(n_7419),
.A2(n_6844),
.B1(n_6575),
.B2(n_6755),
.Y(n_7982)
);

OAI21x1_ASAP7_75t_L g7983 ( 
.A1(n_7333),
.A2(n_6334),
.B(n_6204),
.Y(n_7983)
);

NAND2x1p5_ASAP7_75t_L g7984 ( 
.A(n_7431),
.B(n_6532),
.Y(n_7984)
);

AND2x2_ASAP7_75t_L g7985 ( 
.A(n_7008),
.B(n_6603),
.Y(n_7985)
);

NOR2xp33_ASAP7_75t_L g7986 ( 
.A(n_6959),
.B(n_6318),
.Y(n_7986)
);

INVx1_ASAP7_75t_L g7987 ( 
.A(n_7643),
.Y(n_7987)
);

BUFx12f_ASAP7_75t_L g7988 ( 
.A(n_7398),
.Y(n_7988)
);

BUFx4f_ASAP7_75t_L g7989 ( 
.A(n_7309),
.Y(n_7989)
);

BUFx2_ASAP7_75t_L g7990 ( 
.A(n_7509),
.Y(n_7990)
);

AND2x4_ASAP7_75t_SL g7991 ( 
.A(n_7245),
.B(n_6324),
.Y(n_7991)
);

OA21x2_ASAP7_75t_L g7992 ( 
.A1(n_7344),
.A2(n_6591),
.B(n_6669),
.Y(n_7992)
);

OAI21x1_ASAP7_75t_L g7993 ( 
.A1(n_7380),
.A2(n_6334),
.B(n_6204),
.Y(n_7993)
);

OAI21x1_ASAP7_75t_L g7994 ( 
.A1(n_7380),
.A2(n_6200),
.B(n_6779),
.Y(n_7994)
);

AO21x2_ASAP7_75t_L g7995 ( 
.A1(n_7891),
.A2(n_6884),
.B(n_6205),
.Y(n_7995)
);

OAI21x1_ASAP7_75t_SL g7996 ( 
.A1(n_7296),
.A2(n_6343),
.B(n_6609),
.Y(n_7996)
);

INVx3_ASAP7_75t_SL g7997 ( 
.A(n_7000),
.Y(n_7997)
);

BUFx3_ASAP7_75t_L g7998 ( 
.A(n_7433),
.Y(n_7998)
);

INVx1_ASAP7_75t_L g7999 ( 
.A(n_7643),
.Y(n_7999)
);

OAI21x1_ASAP7_75t_L g8000 ( 
.A1(n_7195),
.A2(n_6707),
.B(n_6695),
.Y(n_8000)
);

INVx1_ASAP7_75t_L g8001 ( 
.A(n_7644),
.Y(n_8001)
);

NAND2x1p5_ASAP7_75t_L g8002 ( 
.A(n_7431),
.B(n_6532),
.Y(n_8002)
);

NAND2xp5_ASAP7_75t_L g8003 ( 
.A(n_6992),
.B(n_6627),
.Y(n_8003)
);

AOI22xp33_ASAP7_75t_L g8004 ( 
.A1(n_7298),
.A2(n_6073),
.B1(n_6675),
.B2(n_6406),
.Y(n_8004)
);

AOI22xp33_ASAP7_75t_SL g8005 ( 
.A1(n_7640),
.A2(n_5872),
.B1(n_5968),
.B2(n_6199),
.Y(n_8005)
);

AND2x2_ASAP7_75t_L g8006 ( 
.A(n_7008),
.B(n_7078),
.Y(n_8006)
);

NAND2x1p5_ASAP7_75t_L g8007 ( 
.A(n_7431),
.B(n_6546),
.Y(n_8007)
);

AOI21xp5_ASAP7_75t_L g8008 ( 
.A1(n_7889),
.A2(n_6058),
.B(n_6027),
.Y(n_8008)
);

INVx1_ASAP7_75t_L g8009 ( 
.A(n_7644),
.Y(n_8009)
);

INVx2_ASAP7_75t_L g8010 ( 
.A(n_6941),
.Y(n_8010)
);

AND2x2_ASAP7_75t_L g8011 ( 
.A(n_7008),
.B(n_6631),
.Y(n_8011)
);

OAI21xp5_ASAP7_75t_L g8012 ( 
.A1(n_7052),
.A2(n_6169),
.B(n_6688),
.Y(n_8012)
);

AO31x2_ASAP7_75t_L g8013 ( 
.A1(n_7400),
.A2(n_5861),
.A3(n_6300),
.B(n_6530),
.Y(n_8013)
);

AO21x2_ASAP7_75t_L g8014 ( 
.A1(n_7891),
.A2(n_6205),
.B(n_6148),
.Y(n_8014)
);

OAI22xp5_ASAP7_75t_L g8015 ( 
.A1(n_7419),
.A2(n_6755),
.B1(n_5857),
.B2(n_6649),
.Y(n_8015)
);

HB1xp67_ASAP7_75t_L g8016 ( 
.A(n_7177),
.Y(n_8016)
);

NAND2xp33_ASAP7_75t_L g8017 ( 
.A(n_7895),
.B(n_6854),
.Y(n_8017)
);

NOR2xp33_ASAP7_75t_SL g8018 ( 
.A(n_7581),
.B(n_6023),
.Y(n_8018)
);

AND2x6_ASAP7_75t_L g8019 ( 
.A(n_7706),
.B(n_5234),
.Y(n_8019)
);

AOI21xp33_ASAP7_75t_L g8020 ( 
.A1(n_7640),
.A2(n_6823),
.B(n_6795),
.Y(n_8020)
);

AOI21xp5_ASAP7_75t_L g8021 ( 
.A1(n_7034),
.A2(n_7324),
.B(n_6928),
.Y(n_8021)
);

NAND2xp5_ASAP7_75t_L g8022 ( 
.A(n_6992),
.B(n_6631),
.Y(n_8022)
);

INVx2_ASAP7_75t_L g8023 ( 
.A(n_6941),
.Y(n_8023)
);

AOI22x1_ASAP7_75t_L g8024 ( 
.A1(n_7219),
.A2(n_7107),
.B1(n_7296),
.B2(n_7173),
.Y(n_8024)
);

AOI22x1_ASAP7_75t_L g8025 ( 
.A1(n_7107),
.A2(n_5966),
.B1(n_5861),
.B2(n_5879),
.Y(n_8025)
);

BUFx6f_ASAP7_75t_L g8026 ( 
.A(n_6940),
.Y(n_8026)
);

BUFx2_ASAP7_75t_L g8027 ( 
.A(n_7509),
.Y(n_8027)
);

NAND2xp5_ASAP7_75t_L g8028 ( 
.A(n_6959),
.B(n_6631),
.Y(n_8028)
);

INVx1_ASAP7_75t_L g8029 ( 
.A(n_7644),
.Y(n_8029)
);

OR2x2_ASAP7_75t_L g8030 ( 
.A(n_7350),
.B(n_6228),
.Y(n_8030)
);

INVx1_ASAP7_75t_L g8031 ( 
.A(n_7647),
.Y(n_8031)
);

INVx2_ASAP7_75t_L g8032 ( 
.A(n_6941),
.Y(n_8032)
);

INVx2_ASAP7_75t_L g8033 ( 
.A(n_6953),
.Y(n_8033)
);

INVxp67_ASAP7_75t_L g8034 ( 
.A(n_7462),
.Y(n_8034)
);

INVx2_ASAP7_75t_SL g8035 ( 
.A(n_7431),
.Y(n_8035)
);

AO21x2_ASAP7_75t_L g8036 ( 
.A1(n_7175),
.A2(n_6516),
.B(n_6148),
.Y(n_8036)
);

O2A1O1Ixp33_ASAP7_75t_SL g8037 ( 
.A1(n_7652),
.A2(n_7830),
.B(n_7035),
.C(n_7279),
.Y(n_8037)
);

INVxp67_ASAP7_75t_L g8038 ( 
.A(n_7462),
.Y(n_8038)
);

AOI22xp33_ASAP7_75t_SL g8039 ( 
.A1(n_7640),
.A2(n_5968),
.B1(n_6502),
.B2(n_6569),
.Y(n_8039)
);

INVx1_ASAP7_75t_L g8040 ( 
.A(n_7647),
.Y(n_8040)
);

AND2x4_ASAP7_75t_L g8041 ( 
.A(n_7518),
.B(n_6421),
.Y(n_8041)
);

BUFx3_ASAP7_75t_L g8042 ( 
.A(n_7433),
.Y(n_8042)
);

AND2x4_ASAP7_75t_L g8043 ( 
.A(n_7518),
.B(n_6421),
.Y(n_8043)
);

OA21x2_ASAP7_75t_L g8044 ( 
.A1(n_7382),
.A2(n_6669),
.B(n_6530),
.Y(n_8044)
);

OAI21x1_ASAP7_75t_L g8045 ( 
.A1(n_6918),
.A2(n_7660),
.B(n_7396),
.Y(n_8045)
);

BUFx3_ASAP7_75t_L g8046 ( 
.A(n_7433),
.Y(n_8046)
);

AND2x2_ASAP7_75t_L g8047 ( 
.A(n_7008),
.B(n_6648),
.Y(n_8047)
);

AO21x2_ASAP7_75t_L g8048 ( 
.A1(n_7175),
.A2(n_6516),
.B(n_6744),
.Y(n_8048)
);

AO21x2_ASAP7_75t_L g8049 ( 
.A1(n_7191),
.A2(n_7225),
.B(n_7197),
.Y(n_8049)
);

INVxp67_ASAP7_75t_SL g8050 ( 
.A(n_7177),
.Y(n_8050)
);

NAND2xp5_ASAP7_75t_L g8051 ( 
.A(n_6959),
.B(n_6648),
.Y(n_8051)
);

OAI21x1_ASAP7_75t_L g8052 ( 
.A1(n_6918),
.A2(n_6767),
.B(n_6511),
.Y(n_8052)
);

INVx2_ASAP7_75t_SL g8053 ( 
.A(n_7431),
.Y(n_8053)
);

AOI22xp33_ASAP7_75t_L g8054 ( 
.A1(n_7298),
.A2(n_6406),
.B1(n_6426),
.B2(n_6339),
.Y(n_8054)
);

NAND2xp5_ASAP7_75t_L g8055 ( 
.A(n_6956),
.B(n_6657),
.Y(n_8055)
);

NOR2xp67_ASAP7_75t_L g8056 ( 
.A(n_7579),
.B(n_5861),
.Y(n_8056)
);

AOI21x1_ASAP7_75t_L g8057 ( 
.A1(n_6995),
.A2(n_5890),
.B(n_6398),
.Y(n_8057)
);

BUFx2_ASAP7_75t_L g8058 ( 
.A(n_7509),
.Y(n_8058)
);

AOI21x1_ASAP7_75t_L g8059 ( 
.A1(n_6995),
.A2(n_6481),
.B(n_6398),
.Y(n_8059)
);

AND2x4_ASAP7_75t_L g8060 ( 
.A(n_7518),
.B(n_6264),
.Y(n_8060)
);

AND2x4_ASAP7_75t_L g8061 ( 
.A(n_7518),
.B(n_6264),
.Y(n_8061)
);

INVx2_ASAP7_75t_L g8062 ( 
.A(n_6953),
.Y(n_8062)
);

INVx1_ASAP7_75t_L g8063 ( 
.A(n_7647),
.Y(n_8063)
);

HB1xp67_ASAP7_75t_L g8064 ( 
.A(n_7188),
.Y(n_8064)
);

NAND2xp5_ASAP7_75t_L g8065 ( 
.A(n_6956),
.B(n_6657),
.Y(n_8065)
);

OAI21x1_ASAP7_75t_L g8066 ( 
.A1(n_6918),
.A2(n_7660),
.B(n_7396),
.Y(n_8066)
);

OAI21x1_ASAP7_75t_L g8067 ( 
.A1(n_6918),
.A2(n_6767),
.B(n_6511),
.Y(n_8067)
);

OAI21x1_ASAP7_75t_L g8068 ( 
.A1(n_7660),
.A2(n_6511),
.B(n_6779),
.Y(n_8068)
);

INVx2_ASAP7_75t_L g8069 ( 
.A(n_6953),
.Y(n_8069)
);

AOI22xp33_ASAP7_75t_L g8070 ( 
.A1(n_7137),
.A2(n_6426),
.B1(n_6493),
.B2(n_6339),
.Y(n_8070)
);

OAI21x1_ASAP7_75t_L g8071 ( 
.A1(n_7382),
.A2(n_6787),
.B(n_6780),
.Y(n_8071)
);

INVx4_ASAP7_75t_L g8072 ( 
.A(n_7309),
.Y(n_8072)
);

INVx1_ASAP7_75t_SL g8073 ( 
.A(n_7181),
.Y(n_8073)
);

CKINVDCx11_ASAP7_75t_R g8074 ( 
.A(n_7309),
.Y(n_8074)
);

CKINVDCx8_ASAP7_75t_R g8075 ( 
.A(n_7000),
.Y(n_8075)
);

AOI22xp5_ASAP7_75t_L g8076 ( 
.A1(n_7607),
.A2(n_5769),
.B1(n_5850),
.B2(n_6573),
.Y(n_8076)
);

OA21x2_ASAP7_75t_L g8077 ( 
.A1(n_7405),
.A2(n_6781),
.B(n_6744),
.Y(n_8077)
);

INVx2_ASAP7_75t_L g8078 ( 
.A(n_6953),
.Y(n_8078)
);

AND2x4_ASAP7_75t_L g8079 ( 
.A(n_6913),
.B(n_6264),
.Y(n_8079)
);

AO221x2_ASAP7_75t_L g8080 ( 
.A1(n_7392),
.A2(n_6778),
.B1(n_6571),
.B2(n_6845),
.C(n_6828),
.Y(n_8080)
);

OAI21x1_ASAP7_75t_L g8081 ( 
.A1(n_7405),
.A2(n_7413),
.B(n_7411),
.Y(n_8081)
);

AND2x4_ASAP7_75t_L g8082 ( 
.A(n_6913),
.B(n_6264),
.Y(n_8082)
);

INVx2_ASAP7_75t_L g8083 ( 
.A(n_6962),
.Y(n_8083)
);

AO21x2_ASAP7_75t_L g8084 ( 
.A1(n_7191),
.A2(n_6772),
.B(n_6135),
.Y(n_8084)
);

OAI21xp5_ASAP7_75t_L g8085 ( 
.A1(n_7652),
.A2(n_7324),
.B(n_7607),
.Y(n_8085)
);

AOI21xp5_ASAP7_75t_L g8086 ( 
.A1(n_7034),
.A2(n_6058),
.B(n_6027),
.Y(n_8086)
);

INVx6_ASAP7_75t_L g8087 ( 
.A(n_7572),
.Y(n_8087)
);

CKINVDCx5p33_ASAP7_75t_R g8088 ( 
.A(n_7330),
.Y(n_8088)
);

INVx1_ASAP7_75t_L g8089 ( 
.A(n_7655),
.Y(n_8089)
);

OAI21x1_ASAP7_75t_L g8090 ( 
.A1(n_7411),
.A2(n_6787),
.B(n_6780),
.Y(n_8090)
);

AOI221xp5_ASAP7_75t_SL g8091 ( 
.A1(n_7648),
.A2(n_6828),
.B1(n_6778),
.B2(n_6245),
.C(n_6234),
.Y(n_8091)
);

INVxp67_ASAP7_75t_SL g8092 ( 
.A(n_7188),
.Y(n_8092)
);

INVx2_ASAP7_75t_L g8093 ( 
.A(n_6962),
.Y(n_8093)
);

OAI22xp5_ASAP7_75t_L g8094 ( 
.A1(n_7760),
.A2(n_5857),
.B1(n_6649),
.B2(n_5832),
.Y(n_8094)
);

BUFx6f_ASAP7_75t_L g8095 ( 
.A(n_6940),
.Y(n_8095)
);

AO21x2_ASAP7_75t_L g8096 ( 
.A1(n_7197),
.A2(n_6772),
.B(n_6135),
.Y(n_8096)
);

CKINVDCx6p67_ASAP7_75t_R g8097 ( 
.A(n_7009),
.Y(n_8097)
);

OAI21x1_ASAP7_75t_L g8098 ( 
.A1(n_7413),
.A2(n_6793),
.B(n_6789),
.Y(n_8098)
);

OAI21x1_ASAP7_75t_L g8099 ( 
.A1(n_7421),
.A2(n_6793),
.B(n_6789),
.Y(n_8099)
);

AND2x2_ASAP7_75t_L g8100 ( 
.A(n_7078),
.B(n_6657),
.Y(n_8100)
);

OAI21x1_ASAP7_75t_L g8101 ( 
.A1(n_7421),
.A2(n_6871),
.B(n_6856),
.Y(n_8101)
);

BUFx8_ASAP7_75t_L g8102 ( 
.A(n_7318),
.Y(n_8102)
);

OA21x2_ASAP7_75t_L g8103 ( 
.A1(n_7446),
.A2(n_7478),
.B(n_7454),
.Y(n_8103)
);

AND2x2_ASAP7_75t_L g8104 ( 
.A(n_7078),
.B(n_6689),
.Y(n_8104)
);

INVx1_ASAP7_75t_L g8105 ( 
.A(n_7655),
.Y(n_8105)
);

HB1xp67_ASAP7_75t_L g8106 ( 
.A(n_7201),
.Y(n_8106)
);

INVx1_ASAP7_75t_SL g8107 ( 
.A(n_7181),
.Y(n_8107)
);

INVx1_ASAP7_75t_L g8108 ( 
.A(n_7655),
.Y(n_8108)
);

OAI21x1_ASAP7_75t_L g8109 ( 
.A1(n_7446),
.A2(n_6871),
.B(n_6856),
.Y(n_8109)
);

INVx2_ASAP7_75t_L g8110 ( 
.A(n_6962),
.Y(n_8110)
);

INVx2_ASAP7_75t_L g8111 ( 
.A(n_6962),
.Y(n_8111)
);

INVx1_ASAP7_75t_SL g8112 ( 
.A(n_7181),
.Y(n_8112)
);

INVx1_ASAP7_75t_L g8113 ( 
.A(n_7657),
.Y(n_8113)
);

NAND2x1p5_ASAP7_75t_L g8114 ( 
.A(n_7431),
.B(n_6546),
.Y(n_8114)
);

OA21x2_ASAP7_75t_L g8115 ( 
.A1(n_7454),
.A2(n_6781),
.B(n_6552),
.Y(n_8115)
);

CKINVDCx16_ASAP7_75t_R g8116 ( 
.A(n_6921),
.Y(n_8116)
);

OAI21x1_ASAP7_75t_L g8117 ( 
.A1(n_7478),
.A2(n_6881),
.B(n_6875),
.Y(n_8117)
);

OAI21x1_ASAP7_75t_L g8118 ( 
.A1(n_7479),
.A2(n_6881),
.B(n_6875),
.Y(n_8118)
);

INVx3_ASAP7_75t_L g8119 ( 
.A(n_7509),
.Y(n_8119)
);

BUFx3_ASAP7_75t_L g8120 ( 
.A(n_7433),
.Y(n_8120)
);

AOI22xp33_ASAP7_75t_L g8121 ( 
.A1(n_7648),
.A2(n_6495),
.B1(n_6498),
.B2(n_6493),
.Y(n_8121)
);

INVx1_ASAP7_75t_L g8122 ( 
.A(n_7657),
.Y(n_8122)
);

INVx1_ASAP7_75t_L g8123 ( 
.A(n_7657),
.Y(n_8123)
);

INVx2_ASAP7_75t_L g8124 ( 
.A(n_6975),
.Y(n_8124)
);

OA21x2_ASAP7_75t_L g8125 ( 
.A1(n_7479),
.A2(n_7503),
.B(n_7480),
.Y(n_8125)
);

INVx2_ASAP7_75t_L g8126 ( 
.A(n_6975),
.Y(n_8126)
);

OAI21x1_ASAP7_75t_L g8127 ( 
.A1(n_7480),
.A2(n_6888),
.B(n_6886),
.Y(n_8127)
);

NAND2xp5_ASAP7_75t_L g8128 ( 
.A(n_7791),
.B(n_6689),
.Y(n_8128)
);

INVx2_ASAP7_75t_L g8129 ( 
.A(n_6975),
.Y(n_8129)
);

OAI22xp5_ASAP7_75t_L g8130 ( 
.A1(n_7760),
.A2(n_5832),
.B1(n_5968),
.B2(n_6846),
.Y(n_8130)
);

AO31x2_ASAP7_75t_L g8131 ( 
.A1(n_7400),
.A2(n_6300),
.A3(n_6552),
.B(n_6245),
.Y(n_8131)
);

OAI22xp5_ASAP7_75t_L g8132 ( 
.A1(n_7607),
.A2(n_5968),
.B1(n_6846),
.B2(n_6429),
.Y(n_8132)
);

INVx1_ASAP7_75t_L g8133 ( 
.A(n_7665),
.Y(n_8133)
);

OAI21x1_ASAP7_75t_L g8134 ( 
.A1(n_7503),
.A2(n_6888),
.B(n_6886),
.Y(n_8134)
);

AOI22xp33_ASAP7_75t_L g8135 ( 
.A1(n_7107),
.A2(n_6495),
.B1(n_6498),
.B2(n_6408),
.Y(n_8135)
);

AOI21xp5_ASAP7_75t_L g8136 ( 
.A1(n_6917),
.A2(n_6577),
.B(n_6025),
.Y(n_8136)
);

AOI21xp5_ASAP7_75t_L g8137 ( 
.A1(n_6917),
.A2(n_6928),
.B(n_7755),
.Y(n_8137)
);

INVx2_ASAP7_75t_SL g8138 ( 
.A(n_7529),
.Y(n_8138)
);

NAND2xp5_ASAP7_75t_SL g8139 ( 
.A(n_7514),
.B(n_6795),
.Y(n_8139)
);

OAI21x1_ASAP7_75t_L g8140 ( 
.A1(n_7527),
.A2(n_7537),
.B(n_7530),
.Y(n_8140)
);

AND2x2_ASAP7_75t_L g8141 ( 
.A(n_7078),
.B(n_6722),
.Y(n_8141)
);

BUFx6f_ASAP7_75t_L g8142 ( 
.A(n_6940),
.Y(n_8142)
);

OAI21xp5_ASAP7_75t_L g8143 ( 
.A1(n_7392),
.A2(n_6344),
.B(n_6316),
.Y(n_8143)
);

NAND2xp5_ASAP7_75t_L g8144 ( 
.A(n_7791),
.B(n_6722),
.Y(n_8144)
);

INVx1_ASAP7_75t_L g8145 ( 
.A(n_7665),
.Y(n_8145)
);

BUFx2_ASAP7_75t_L g8146 ( 
.A(n_7509),
.Y(n_8146)
);

INVx1_ASAP7_75t_L g8147 ( 
.A(n_7665),
.Y(n_8147)
);

INVx1_ASAP7_75t_L g8148 ( 
.A(n_7666),
.Y(n_8148)
);

INVx2_ASAP7_75t_L g8149 ( 
.A(n_6975),
.Y(n_8149)
);

AO21x2_ASAP7_75t_L g8150 ( 
.A1(n_7225),
.A2(n_6132),
.B(n_5949),
.Y(n_8150)
);

OA21x2_ASAP7_75t_L g8151 ( 
.A1(n_7527),
.A2(n_6892),
.B(n_6537),
.Y(n_8151)
);

BUFx3_ASAP7_75t_L g8152 ( 
.A(n_7433),
.Y(n_8152)
);

INVx1_ASAP7_75t_L g8153 ( 
.A(n_7666),
.Y(n_8153)
);

NOR2xp33_ASAP7_75t_L g8154 ( 
.A(n_7037),
.B(n_5813),
.Y(n_8154)
);

NAND2xp5_ASAP7_75t_SL g8155 ( 
.A(n_7514),
.B(n_6502),
.Y(n_8155)
);

AOI22xp33_ASAP7_75t_L g8156 ( 
.A1(n_7107),
.A2(n_6408),
.B1(n_5776),
.B2(n_5896),
.Y(n_8156)
);

AND2x2_ASAP7_75t_L g8157 ( 
.A(n_7678),
.B(n_6722),
.Y(n_8157)
);

NAND2xp5_ASAP7_75t_L g8158 ( 
.A(n_7811),
.B(n_6724),
.Y(n_8158)
);

OAI21xp5_ASAP7_75t_L g8159 ( 
.A1(n_7392),
.A2(n_7168),
.B(n_7683),
.Y(n_8159)
);

AO21x2_ASAP7_75t_L g8160 ( 
.A1(n_7227),
.A2(n_7232),
.B(n_7530),
.Y(n_8160)
);

AOI22xp5_ASAP7_75t_L g8161 ( 
.A1(n_7683),
.A2(n_5782),
.B1(n_5765),
.B2(n_5898),
.Y(n_8161)
);

CKINVDCx20_ASAP7_75t_R g8162 ( 
.A(n_7418),
.Y(n_8162)
);

OAI21x1_ASAP7_75t_L g8163 ( 
.A1(n_7537),
.A2(n_6892),
.B(n_6577),
.Y(n_8163)
);

INVx2_ASAP7_75t_SL g8164 ( 
.A(n_7529),
.Y(n_8164)
);

NAND2xp5_ASAP7_75t_L g8165 ( 
.A(n_7811),
.B(n_6724),
.Y(n_8165)
);

INVx1_ASAP7_75t_SL g8166 ( 
.A(n_7196),
.Y(n_8166)
);

INVx1_ASAP7_75t_L g8167 ( 
.A(n_7666),
.Y(n_8167)
);

AND2x2_ASAP7_75t_L g8168 ( 
.A(n_7678),
.B(n_6724),
.Y(n_8168)
);

BUFx12f_ASAP7_75t_L g8169 ( 
.A(n_7398),
.Y(n_8169)
);

OAI21x1_ASAP7_75t_L g8170 ( 
.A1(n_7538),
.A2(n_5949),
.B(n_6021),
.Y(n_8170)
);

OAI21x1_ASAP7_75t_L g8171 ( 
.A1(n_7538),
.A2(n_6025),
.B(n_6021),
.Y(n_8171)
);

INVx2_ASAP7_75t_SL g8172 ( 
.A(n_7529),
.Y(n_8172)
);

INVx1_ASAP7_75t_L g8173 ( 
.A(n_7670),
.Y(n_8173)
);

INVx1_ASAP7_75t_L g8174 ( 
.A(n_7670),
.Y(n_8174)
);

AOI21xp5_ASAP7_75t_L g8175 ( 
.A1(n_7755),
.A2(n_6344),
.B(n_6316),
.Y(n_8175)
);

HB1xp67_ASAP7_75t_L g8176 ( 
.A(n_7201),
.Y(n_8176)
);

INVx1_ASAP7_75t_L g8177 ( 
.A(n_7670),
.Y(n_8177)
);

INVx2_ASAP7_75t_L g8178 ( 
.A(n_6980),
.Y(n_8178)
);

BUFx3_ASAP7_75t_L g8179 ( 
.A(n_7433),
.Y(n_8179)
);

AO32x2_ASAP7_75t_L g8180 ( 
.A1(n_7241),
.A2(n_6842),
.A3(n_6840),
.B1(n_6835),
.B2(n_5791),
.Y(n_8180)
);

INVx1_ASAP7_75t_L g8181 ( 
.A(n_7672),
.Y(n_8181)
);

OR2x2_ASAP7_75t_L g8182 ( 
.A(n_7350),
.B(n_6228),
.Y(n_8182)
);

AND2x4_ASAP7_75t_L g8183 ( 
.A(n_6913),
.B(n_6924),
.Y(n_8183)
);

INVxp67_ASAP7_75t_L g8184 ( 
.A(n_7434),
.Y(n_8184)
);

AO21x2_ASAP7_75t_L g8185 ( 
.A1(n_7227),
.A2(n_6132),
.B(n_6320),
.Y(n_8185)
);

INVx1_ASAP7_75t_L g8186 ( 
.A(n_7672),
.Y(n_8186)
);

AND2x2_ASAP7_75t_L g8187 ( 
.A(n_7678),
.B(n_6754),
.Y(n_8187)
);

AO21x2_ASAP7_75t_L g8188 ( 
.A1(n_7232),
.A2(n_5842),
.B(n_6896),
.Y(n_8188)
);

OAI22xp5_ASAP7_75t_L g8189 ( 
.A1(n_7012),
.A2(n_6429),
.B1(n_6593),
.B2(n_5839),
.Y(n_8189)
);

INVx1_ASAP7_75t_L g8190 ( 
.A(n_7672),
.Y(n_8190)
);

NOR2xp33_ASAP7_75t_L g8191 ( 
.A(n_7037),
.B(n_5813),
.Y(n_8191)
);

NAND2xp5_ASAP7_75t_L g8192 ( 
.A(n_7827),
.B(n_6754),
.Y(n_8192)
);

INVx1_ASAP7_75t_L g8193 ( 
.A(n_7673),
.Y(n_8193)
);

CKINVDCx20_ASAP7_75t_R g8194 ( 
.A(n_7418),
.Y(n_8194)
);

A2O1A1Ixp33_ASAP7_75t_L g8195 ( 
.A1(n_7146),
.A2(n_6234),
.B(n_5855),
.C(n_5810),
.Y(n_8195)
);

INVx2_ASAP7_75t_L g8196 ( 
.A(n_6980),
.Y(n_8196)
);

NAND2xp5_ASAP7_75t_SL g8197 ( 
.A(n_7514),
.B(n_6850),
.Y(n_8197)
);

INVx1_ASAP7_75t_L g8198 ( 
.A(n_7673),
.Y(n_8198)
);

INVx1_ASAP7_75t_L g8199 ( 
.A(n_7673),
.Y(n_8199)
);

INVx1_ASAP7_75t_L g8200 ( 
.A(n_7674),
.Y(n_8200)
);

BUFx12f_ASAP7_75t_L g8201 ( 
.A(n_7009),
.Y(n_8201)
);

INVx1_ASAP7_75t_L g8202 ( 
.A(n_7674),
.Y(n_8202)
);

OAI21x1_ASAP7_75t_L g8203 ( 
.A1(n_7548),
.A2(n_6200),
.B(n_6723),
.Y(n_8203)
);

OAI21x1_ASAP7_75t_L g8204 ( 
.A1(n_7548),
.A2(n_6200),
.B(n_6723),
.Y(n_8204)
);

OAI21x1_ASAP7_75t_L g8205 ( 
.A1(n_7554),
.A2(n_6723),
.B(n_5848),
.Y(n_8205)
);

INVx1_ASAP7_75t_L g8206 ( 
.A(n_7674),
.Y(n_8206)
);

NAND2xp5_ASAP7_75t_L g8207 ( 
.A(n_7827),
.B(n_6754),
.Y(n_8207)
);

NAND2x1p5_ASAP7_75t_L g8208 ( 
.A(n_7529),
.B(n_6546),
.Y(n_8208)
);

OAI21x1_ASAP7_75t_L g8209 ( 
.A1(n_7554),
.A2(n_6723),
.B(n_5848),
.Y(n_8209)
);

BUFx10_ASAP7_75t_L g8210 ( 
.A(n_7408),
.Y(n_8210)
);

BUFx2_ASAP7_75t_L g8211 ( 
.A(n_7509),
.Y(n_8211)
);

OR2x2_ASAP7_75t_L g8212 ( 
.A(n_7350),
.B(n_6266),
.Y(n_8212)
);

NAND2xp5_ASAP7_75t_L g8213 ( 
.A(n_7073),
.B(n_6266),
.Y(n_8213)
);

OAI21x1_ASAP7_75t_L g8214 ( 
.A1(n_7557),
.A2(n_6723),
.B(n_6698),
.Y(n_8214)
);

OAI21x1_ASAP7_75t_L g8215 ( 
.A1(n_7557),
.A2(n_6698),
.B(n_6496),
.Y(n_8215)
);

AOI22xp33_ASAP7_75t_SL g8216 ( 
.A1(n_6921),
.A2(n_6569),
.B1(n_6763),
.B2(n_6685),
.Y(n_8216)
);

CKINVDCx6p67_ASAP7_75t_R g8217 ( 
.A(n_7009),
.Y(n_8217)
);

BUFx2_ASAP7_75t_L g8218 ( 
.A(n_7509),
.Y(n_8218)
);

INVx3_ASAP7_75t_L g8219 ( 
.A(n_6940),
.Y(n_8219)
);

AOI222xp33_ASAP7_75t_L g8220 ( 
.A1(n_7012),
.A2(n_6764),
.B1(n_6589),
.B2(n_6122),
.C1(n_5879),
.C2(n_5898),
.Y(n_8220)
);

INVx1_ASAP7_75t_SL g8221 ( 
.A(n_7196),
.Y(n_8221)
);

AOI22xp33_ASAP7_75t_L g8222 ( 
.A1(n_7146),
.A2(n_5896),
.B1(n_5782),
.B2(n_5765),
.Y(n_8222)
);

AOI31xp67_ASAP7_75t_L g8223 ( 
.A1(n_7713),
.A2(n_7282),
.A3(n_7354),
.B(n_7310),
.Y(n_8223)
);

AOI22xp33_ASAP7_75t_L g8224 ( 
.A1(n_7146),
.A2(n_5961),
.B1(n_6230),
.B2(n_6764),
.Y(n_8224)
);

AOI21xp33_ASAP7_75t_L g8225 ( 
.A1(n_7467),
.A2(n_6665),
.B(n_6489),
.Y(n_8225)
);

AOI22xp5_ASAP7_75t_L g8226 ( 
.A1(n_7683),
.A2(n_7012),
.B1(n_6947),
.B2(n_7717),
.Y(n_8226)
);

BUFx3_ASAP7_75t_L g8227 ( 
.A(n_7433),
.Y(n_8227)
);

AOI21x1_ASAP7_75t_L g8228 ( 
.A1(n_7896),
.A2(n_6496),
.B(n_6481),
.Y(n_8228)
);

AND2x2_ASAP7_75t_L g8229 ( 
.A(n_7678),
.B(n_6259),
.Y(n_8229)
);

OAI21x1_ASAP7_75t_L g8230 ( 
.A1(n_7568),
.A2(n_6645),
.B(n_6539),
.Y(n_8230)
);

OAI21x1_ASAP7_75t_SL g8231 ( 
.A1(n_7296),
.A2(n_6343),
.B(n_7698),
.Y(n_8231)
);

INVx2_ASAP7_75t_L g8232 ( 
.A(n_6980),
.Y(n_8232)
);

OAI21x1_ASAP7_75t_L g8233 ( 
.A1(n_7568),
.A2(n_6645),
.B(n_6539),
.Y(n_8233)
);

OAI21xp5_ASAP7_75t_L g8234 ( 
.A1(n_7168),
.A2(n_5939),
.B(n_5810),
.Y(n_8234)
);

OAI21x1_ASAP7_75t_L g8235 ( 
.A1(n_7896),
.A2(n_6810),
.B(n_6766),
.Y(n_8235)
);

INVx1_ASAP7_75t_L g8236 ( 
.A(n_7679),
.Y(n_8236)
);

INVx2_ASAP7_75t_L g8237 ( 
.A(n_6980),
.Y(n_8237)
);

AO31x2_ASAP7_75t_L g8238 ( 
.A1(n_7400),
.A2(n_7832),
.A3(n_7854),
.B(n_7822),
.Y(n_8238)
);

INVx1_ASAP7_75t_L g8239 ( 
.A(n_7679),
.Y(n_8239)
);

INVx2_ASAP7_75t_L g8240 ( 
.A(n_6983),
.Y(n_8240)
);

NOR2xp33_ASAP7_75t_L g8241 ( 
.A(n_7037),
.B(n_5815),
.Y(n_8241)
);

INVx2_ASAP7_75t_L g8242 ( 
.A(n_6983),
.Y(n_8242)
);

AOI22xp33_ASAP7_75t_L g8243 ( 
.A1(n_7394),
.A2(n_6230),
.B1(n_6526),
.B2(n_6589),
.Y(n_8243)
);

AND2x4_ASAP7_75t_L g8244 ( 
.A(n_6913),
.B(n_6421),
.Y(n_8244)
);

OAI21x1_ASAP7_75t_L g8245 ( 
.A1(n_7896),
.A2(n_6810),
.B(n_6766),
.Y(n_8245)
);

AOI21x1_ASAP7_75t_L g8246 ( 
.A1(n_7423),
.A2(n_7692),
.B(n_7667),
.Y(n_8246)
);

CKINVDCx5p33_ASAP7_75t_R g8247 ( 
.A(n_7251),
.Y(n_8247)
);

INVx1_ASAP7_75t_L g8248 ( 
.A(n_7679),
.Y(n_8248)
);

INVx1_ASAP7_75t_L g8249 ( 
.A(n_7681),
.Y(n_8249)
);

AO21x2_ASAP7_75t_L g8250 ( 
.A1(n_7174),
.A2(n_5842),
.B(n_6896),
.Y(n_8250)
);

OAI21x1_ASAP7_75t_L g8251 ( 
.A1(n_7100),
.A2(n_6834),
.B(n_6811),
.Y(n_8251)
);

OAI21x1_ASAP7_75t_L g8252 ( 
.A1(n_7100),
.A2(n_6834),
.B(n_6811),
.Y(n_8252)
);

OR2x6_ASAP7_75t_L g8253 ( 
.A(n_7427),
.B(n_6601),
.Y(n_8253)
);

INVx2_ASAP7_75t_L g8254 ( 
.A(n_6983),
.Y(n_8254)
);

INVx2_ASAP7_75t_SL g8255 ( 
.A(n_7529),
.Y(n_8255)
);

OAI21x1_ASAP7_75t_L g8256 ( 
.A1(n_7281),
.A2(n_6614),
.B(n_6526),
.Y(n_8256)
);

INVx1_ASAP7_75t_L g8257 ( 
.A(n_7681),
.Y(n_8257)
);

NAND2xp5_ASAP7_75t_L g8258 ( 
.A(n_7073),
.B(n_6281),
.Y(n_8258)
);

OAI21x1_ASAP7_75t_L g8259 ( 
.A1(n_7281),
.A2(n_6614),
.B(n_6874),
.Y(n_8259)
);

OAI21x1_ASAP7_75t_SL g8260 ( 
.A1(n_7698),
.A2(n_6609),
.B(n_6879),
.Y(n_8260)
);

INVx1_ASAP7_75t_L g8261 ( 
.A(n_7681),
.Y(n_8261)
);

AND4x1_ASAP7_75t_L g8262 ( 
.A(n_6921),
.B(n_6023),
.C(n_6729),
.D(n_6699),
.Y(n_8262)
);

CKINVDCx5p33_ASAP7_75t_R g8263 ( 
.A(n_7251),
.Y(n_8263)
);

INVx2_ASAP7_75t_L g8264 ( 
.A(n_6983),
.Y(n_8264)
);

NAND2xp5_ASAP7_75t_SL g8265 ( 
.A(n_7044),
.B(n_6850),
.Y(n_8265)
);

OR2x2_ASAP7_75t_L g8266 ( 
.A(n_7350),
.B(n_6964),
.Y(n_8266)
);

OAI21x1_ASAP7_75t_L g8267 ( 
.A1(n_7291),
.A2(n_6889),
.B(n_6874),
.Y(n_8267)
);

HB1xp67_ASAP7_75t_L g8268 ( 
.A(n_7214),
.Y(n_8268)
);

INVx3_ASAP7_75t_L g8269 ( 
.A(n_6940),
.Y(n_8269)
);

INVx2_ASAP7_75t_L g8270 ( 
.A(n_6988),
.Y(n_8270)
);

AOI21x1_ASAP7_75t_L g8271 ( 
.A1(n_7423),
.A2(n_6869),
.B(n_5914),
.Y(n_8271)
);

OAI21x1_ASAP7_75t_L g8272 ( 
.A1(n_7291),
.A2(n_6889),
.B(n_6650),
.Y(n_8272)
);

INVx2_ASAP7_75t_L g8273 ( 
.A(n_6988),
.Y(n_8273)
);

INVx4_ASAP7_75t_L g8274 ( 
.A(n_7318),
.Y(n_8274)
);

OAI221xp5_ASAP7_75t_L g8275 ( 
.A1(n_7717),
.A2(n_6732),
.B1(n_6836),
.B2(n_6699),
.C(n_6796),
.Y(n_8275)
);

INVx2_ASAP7_75t_L g8276 ( 
.A(n_6988),
.Y(n_8276)
);

BUFx3_ASAP7_75t_L g8277 ( 
.A(n_7433),
.Y(n_8277)
);

A2O1A1Ixp33_ASAP7_75t_L g8278 ( 
.A1(n_6925),
.A2(n_5952),
.B(n_6665),
.C(n_5966),
.Y(n_8278)
);

INVx1_ASAP7_75t_L g8279 ( 
.A(n_7688),
.Y(n_8279)
);

INVx2_ASAP7_75t_L g8280 ( 
.A(n_6988),
.Y(n_8280)
);

NAND3xp33_ASAP7_75t_L g8281 ( 
.A(n_7168),
.B(n_6489),
.C(n_6470),
.Y(n_8281)
);

NAND2xp5_ASAP7_75t_L g8282 ( 
.A(n_7073),
.B(n_7084),
.Y(n_8282)
);

OAI21x1_ASAP7_75t_L g8283 ( 
.A1(n_7305),
.A2(n_6650),
.B(n_5895),
.Y(n_8283)
);

OAI21xp5_ASAP7_75t_L g8284 ( 
.A1(n_6982),
.A2(n_5939),
.B(n_5915),
.Y(n_8284)
);

OAI21x1_ASAP7_75t_L g8285 ( 
.A1(n_7305),
.A2(n_5895),
.B(n_6869),
.Y(n_8285)
);

OAI21x1_ASAP7_75t_L g8286 ( 
.A1(n_7335),
.A2(n_6747),
.B(n_6733),
.Y(n_8286)
);

OAI21x1_ASAP7_75t_L g8287 ( 
.A1(n_7335),
.A2(n_6747),
.B(n_6733),
.Y(n_8287)
);

OA21x2_ASAP7_75t_L g8288 ( 
.A1(n_7524),
.A2(n_7161),
.B(n_7090),
.Y(n_8288)
);

INVx2_ASAP7_75t_L g8289 ( 
.A(n_7001),
.Y(n_8289)
);

OAI21x1_ASAP7_75t_L g8290 ( 
.A1(n_7524),
.A2(n_6747),
.B(n_6733),
.Y(n_8290)
);

OAI21x1_ASAP7_75t_L g8291 ( 
.A1(n_7090),
.A2(n_6747),
.B(n_6733),
.Y(n_8291)
);

INVx1_ASAP7_75t_L g8292 ( 
.A(n_7688),
.Y(n_8292)
);

CKINVDCx16_ASAP7_75t_R g8293 ( 
.A(n_7384),
.Y(n_8293)
);

INVx1_ASAP7_75t_L g8294 ( 
.A(n_7688),
.Y(n_8294)
);

BUFx6f_ASAP7_75t_L g8295 ( 
.A(n_6940),
.Y(n_8295)
);

INVx6_ASAP7_75t_L g8296 ( 
.A(n_7572),
.Y(n_8296)
);

OAI21xp5_ASAP7_75t_L g8297 ( 
.A1(n_6982),
.A2(n_5939),
.B(n_5778),
.Y(n_8297)
);

CKINVDCx5p33_ASAP7_75t_R g8298 ( 
.A(n_7739),
.Y(n_8298)
);

AO31x2_ASAP7_75t_L g8299 ( 
.A1(n_7400),
.A2(n_6567),
.A3(n_6879),
.B(n_6882),
.Y(n_8299)
);

OAI21x1_ASAP7_75t_SL g8300 ( 
.A1(n_7698),
.A2(n_5952),
.B(n_6443),
.Y(n_8300)
);

OAI21x1_ASAP7_75t_L g8301 ( 
.A1(n_7161),
.A2(n_5883),
.B(n_6098),
.Y(n_8301)
);

NAND2xp5_ASAP7_75t_L g8302 ( 
.A(n_7084),
.B(n_6281),
.Y(n_8302)
);

OAI21x1_ASAP7_75t_L g8303 ( 
.A1(n_7696),
.A2(n_5883),
.B(n_6098),
.Y(n_8303)
);

INVx2_ASAP7_75t_SL g8304 ( 
.A(n_7529),
.Y(n_8304)
);

INVx1_ASAP7_75t_L g8305 ( 
.A(n_7689),
.Y(n_8305)
);

INVx1_ASAP7_75t_L g8306 ( 
.A(n_7689),
.Y(n_8306)
);

A2O1A1Ixp33_ASAP7_75t_L g8307 ( 
.A1(n_6925),
.A2(n_5778),
.B(n_6567),
.C(n_6859),
.Y(n_8307)
);

OAI22xp5_ASAP7_75t_L g8308 ( 
.A1(n_7717),
.A2(n_5839),
.B1(n_5954),
.B2(n_6732),
.Y(n_8308)
);

OAI221xp5_ASAP7_75t_L g8309 ( 
.A1(n_7483),
.A2(n_6836),
.B1(n_6796),
.B2(n_6729),
.C(n_6785),
.Y(n_8309)
);

INVx1_ASAP7_75t_L g8310 ( 
.A(n_7689),
.Y(n_8310)
);

OAI21x1_ASAP7_75t_L g8311 ( 
.A1(n_7696),
.A2(n_6113),
.B(n_5829),
.Y(n_8311)
);

INVx1_ASAP7_75t_L g8312 ( 
.A(n_7690),
.Y(n_8312)
);

OAI21x1_ASAP7_75t_L g8313 ( 
.A1(n_7697),
.A2(n_6113),
.B(n_5829),
.Y(n_8313)
);

INVx2_ASAP7_75t_L g8314 ( 
.A(n_7001),
.Y(n_8314)
);

OAI21x1_ASAP7_75t_L g8315 ( 
.A1(n_7697),
.A2(n_5963),
.B(n_5823),
.Y(n_8315)
);

NAND2xp5_ASAP7_75t_L g8316 ( 
.A(n_7084),
.B(n_6372),
.Y(n_8316)
);

INVx2_ASAP7_75t_L g8317 ( 
.A(n_7001),
.Y(n_8317)
);

CKINVDCx20_ASAP7_75t_R g8318 ( 
.A(n_7507),
.Y(n_8318)
);

INVx2_ASAP7_75t_L g8319 ( 
.A(n_7001),
.Y(n_8319)
);

AO21x2_ASAP7_75t_L g8320 ( 
.A1(n_7174),
.A2(n_6818),
.B(n_5919),
.Y(n_8320)
);

INVx1_ASAP7_75t_L g8321 ( 
.A(n_7690),
.Y(n_8321)
);

OAI21x1_ASAP7_75t_L g8322 ( 
.A1(n_7716),
.A2(n_5963),
.B(n_5823),
.Y(n_8322)
);

CKINVDCx6p67_ASAP7_75t_R g8323 ( 
.A(n_7009),
.Y(n_8323)
);

OAI21x1_ASAP7_75t_L g8324 ( 
.A1(n_7716),
.A2(n_5963),
.B(n_6230),
.Y(n_8324)
);

INVx6_ASAP7_75t_L g8325 ( 
.A(n_7572),
.Y(n_8325)
);

INVx1_ASAP7_75t_L g8326 ( 
.A(n_7690),
.Y(n_8326)
);

OAI21x1_ASAP7_75t_SL g8327 ( 
.A1(n_7871),
.A2(n_6443),
.B(n_6749),
.Y(n_8327)
);

AO21x1_ASAP7_75t_L g8328 ( 
.A1(n_7667),
.A2(n_6870),
.B(n_5957),
.Y(n_8328)
);

NAND2x1p5_ASAP7_75t_L g8329 ( 
.A(n_7529),
.B(n_6546),
.Y(n_8329)
);

OAI21x1_ASAP7_75t_L g8330 ( 
.A1(n_7162),
.A2(n_5870),
.B(n_5912),
.Y(n_8330)
);

AOI222xp33_ASAP7_75t_L g8331 ( 
.A1(n_7271),
.A2(n_6528),
.B1(n_6533),
.B2(n_5888),
.C1(n_5881),
.C2(n_5991),
.Y(n_8331)
);

AOI21x1_ASAP7_75t_L g8332 ( 
.A1(n_7423),
.A2(n_5914),
.B(n_6848),
.Y(n_8332)
);

OAI21x1_ASAP7_75t_SL g8333 ( 
.A1(n_7871),
.A2(n_6749),
.B(n_5786),
.Y(n_8333)
);

INVx2_ASAP7_75t_L g8334 ( 
.A(n_7006),
.Y(n_8334)
);

INVx1_ASAP7_75t_L g8335 ( 
.A(n_7902),
.Y(n_8335)
);

HB1xp67_ASAP7_75t_L g8336 ( 
.A(n_7214),
.Y(n_8336)
);

NOR2xp67_ASAP7_75t_SL g8337 ( 
.A(n_7318),
.B(n_6809),
.Y(n_8337)
);

BUFx10_ASAP7_75t_L g8338 ( 
.A(n_7408),
.Y(n_8338)
);

OAI21x1_ASAP7_75t_L g8339 ( 
.A1(n_7162),
.A2(n_7082),
.B(n_7080),
.Y(n_8339)
);

INVx2_ASAP7_75t_L g8340 ( 
.A(n_7006),
.Y(n_8340)
);

INVx1_ASAP7_75t_L g8341 ( 
.A(n_7902),
.Y(n_8341)
);

AOI22xp33_ASAP7_75t_L g8342 ( 
.A1(n_7394),
.A2(n_6230),
.B1(n_5888),
.B2(n_5881),
.Y(n_8342)
);

OAI22xp5_ASAP7_75t_L g8343 ( 
.A1(n_7704),
.A2(n_5954),
.B1(n_6864),
.B2(n_5953),
.Y(n_8343)
);

AOI21xp5_ASAP7_75t_L g8344 ( 
.A1(n_7080),
.A2(n_5870),
.B(n_6184),
.Y(n_8344)
);

AOI22xp33_ASAP7_75t_L g8345 ( 
.A1(n_7403),
.A2(n_6230),
.B1(n_6607),
.B2(n_5943),
.Y(n_8345)
);

INVx1_ASAP7_75t_L g8346 ( 
.A(n_7902),
.Y(n_8346)
);

NOR2xp33_ASAP7_75t_L g8347 ( 
.A(n_7872),
.B(n_5815),
.Y(n_8347)
);

INVx1_ASAP7_75t_L g8348 ( 
.A(n_7709),
.Y(n_8348)
);

AND2x4_ASAP7_75t_L g8349 ( 
.A(n_6913),
.B(n_6264),
.Y(n_8349)
);

OAI221xp5_ASAP7_75t_L g8350 ( 
.A1(n_7483),
.A2(n_6785),
.B1(n_6830),
.B2(n_6821),
.C(n_6513),
.Y(n_8350)
);

OAI21xp5_ASAP7_75t_L g8351 ( 
.A1(n_7636),
.A2(n_5849),
.B(n_5794),
.Y(n_8351)
);

OAI21x1_ASAP7_75t_SL g8352 ( 
.A1(n_7346),
.A2(n_5786),
.B(n_6870),
.Y(n_8352)
);

INVx2_ASAP7_75t_SL g8353 ( 
.A(n_7529),
.Y(n_8353)
);

CKINVDCx12_ASAP7_75t_R g8354 ( 
.A(n_7804),
.Y(n_8354)
);

INVx2_ASAP7_75t_L g8355 ( 
.A(n_7006),
.Y(n_8355)
);

INVx1_ASAP7_75t_L g8356 ( 
.A(n_7709),
.Y(n_8356)
);

OAI21x1_ASAP7_75t_L g8357 ( 
.A1(n_7082),
.A2(n_5918),
.B(n_5912),
.Y(n_8357)
);

OA21x2_ASAP7_75t_L g8358 ( 
.A1(n_7086),
.A2(n_6818),
.B(n_5919),
.Y(n_8358)
);

AOI21x1_ASAP7_75t_L g8359 ( 
.A1(n_7692),
.A2(n_6848),
.B(n_6681),
.Y(n_8359)
);

OAI21x1_ASAP7_75t_L g8360 ( 
.A1(n_7086),
.A2(n_5928),
.B(n_5918),
.Y(n_8360)
);

OAI21x1_ASAP7_75t_L g8361 ( 
.A1(n_7817),
.A2(n_5928),
.B(n_5957),
.Y(n_8361)
);

AND2x2_ASAP7_75t_L g8362 ( 
.A(n_7782),
.B(n_6259),
.Y(n_8362)
);

OAI22xp33_ASAP7_75t_L g8363 ( 
.A1(n_6943),
.A2(n_5837),
.B1(n_6315),
.B2(n_6183),
.Y(n_8363)
);

AO32x2_ASAP7_75t_L g8364 ( 
.A1(n_7241),
.A2(n_5791),
.A3(n_5933),
.B1(n_5876),
.B2(n_5852),
.Y(n_8364)
);

OAI21x1_ASAP7_75t_L g8365 ( 
.A1(n_7817),
.A2(n_5941),
.B(n_6365),
.Y(n_8365)
);

INVxp33_ASAP7_75t_L g8366 ( 
.A(n_7739),
.Y(n_8366)
);

CKINVDCx20_ASAP7_75t_R g8367 ( 
.A(n_7507),
.Y(n_8367)
);

NAND2xp5_ASAP7_75t_L g8368 ( 
.A(n_7093),
.B(n_6372),
.Y(n_8368)
);

INVx1_ASAP7_75t_L g8369 ( 
.A(n_7709),
.Y(n_8369)
);

OAI21x1_ASAP7_75t_L g8370 ( 
.A1(n_7817),
.A2(n_5941),
.B(n_6365),
.Y(n_8370)
);

OAI22xp33_ASAP7_75t_L g8371 ( 
.A1(n_6943),
.A2(n_5837),
.B1(n_6315),
.B2(n_6183),
.Y(n_8371)
);

AO21x2_ASAP7_75t_L g8372 ( 
.A1(n_7134),
.A2(n_6084),
.B(n_5856),
.Y(n_8372)
);

AND2x2_ASAP7_75t_L g8373 ( 
.A(n_7782),
.B(n_6262),
.Y(n_8373)
);

OA21x2_ASAP7_75t_L g8374 ( 
.A1(n_7164),
.A2(n_6084),
.B(n_5856),
.Y(n_8374)
);

OAI22xp5_ASAP7_75t_L g8375 ( 
.A1(n_7704),
.A2(n_6864),
.B1(n_5953),
.B2(n_6763),
.Y(n_8375)
);

INVx1_ASAP7_75t_L g8376 ( 
.A(n_7714),
.Y(n_8376)
);

OA21x2_ASAP7_75t_L g8377 ( 
.A1(n_7164),
.A2(n_6389),
.B(n_6137),
.Y(n_8377)
);

AOI221xp5_ASAP7_75t_L g8378 ( 
.A1(n_7361),
.A2(n_6542),
.B1(n_6514),
.B2(n_6513),
.C(n_6576),
.Y(n_8378)
);

OR2x6_ASAP7_75t_L g8379 ( 
.A(n_7427),
.B(n_6601),
.Y(n_8379)
);

CKINVDCx20_ASAP7_75t_R g8380 ( 
.A(n_6951),
.Y(n_8380)
);

NAND2x1p5_ASAP7_75t_L g8381 ( 
.A(n_7529),
.B(n_6546),
.Y(n_8381)
);

INVx1_ASAP7_75t_L g8382 ( 
.A(n_7714),
.Y(n_8382)
);

OAI21x1_ASAP7_75t_L g8383 ( 
.A1(n_7817),
.A2(n_5944),
.B(n_5794),
.Y(n_8383)
);

INVx1_ASAP7_75t_L g8384 ( 
.A(n_7714),
.Y(n_8384)
);

AOI22xp5_ASAP7_75t_L g8385 ( 
.A1(n_6947),
.A2(n_5828),
.B1(n_5885),
.B2(n_5867),
.Y(n_8385)
);

OA21x2_ASAP7_75t_L g8386 ( 
.A1(n_7789),
.A2(n_6389),
.B(n_6137),
.Y(n_8386)
);

OAI21x1_ASAP7_75t_L g8387 ( 
.A1(n_7846),
.A2(n_7758),
.B(n_7613),
.Y(n_8387)
);

INVx2_ASAP7_75t_L g8388 ( 
.A(n_7006),
.Y(n_8388)
);

INVx1_ASAP7_75t_L g8389 ( 
.A(n_7724),
.Y(n_8389)
);

CKINVDCx20_ASAP7_75t_R g8390 ( 
.A(n_6951),
.Y(n_8390)
);

INVx1_ASAP7_75t_L g8391 ( 
.A(n_7724),
.Y(n_8391)
);

BUFx2_ASAP7_75t_SL g8392 ( 
.A(n_7529),
.Y(n_8392)
);

INVx1_ASAP7_75t_L g8393 ( 
.A(n_7724),
.Y(n_8393)
);

INVx1_ASAP7_75t_L g8394 ( 
.A(n_7730),
.Y(n_8394)
);

BUFx3_ASAP7_75t_L g8395 ( 
.A(n_7433),
.Y(n_8395)
);

INVx2_ASAP7_75t_L g8396 ( 
.A(n_7015),
.Y(n_8396)
);

NOR2xp33_ASAP7_75t_L g8397 ( 
.A(n_7872),
.B(n_5969),
.Y(n_8397)
);

AOI22x1_ASAP7_75t_L g8398 ( 
.A1(n_7173),
.A2(n_6809),
.B1(n_6683),
.B2(n_6396),
.Y(n_8398)
);

OAI21x1_ASAP7_75t_L g8399 ( 
.A1(n_7846),
.A2(n_5944),
.B(n_5792),
.Y(n_8399)
);

NOR2xp33_ASAP7_75t_L g8400 ( 
.A(n_7872),
.B(n_5969),
.Y(n_8400)
);

NAND2xp5_ASAP7_75t_L g8401 ( 
.A(n_7093),
.B(n_6394),
.Y(n_8401)
);

BUFx3_ASAP7_75t_L g8402 ( 
.A(n_7433),
.Y(n_8402)
);

OAI21x1_ASAP7_75t_L g8403 ( 
.A1(n_7846),
.A2(n_5944),
.B(n_5792),
.Y(n_8403)
);

AOI22xp5_ASAP7_75t_L g8404 ( 
.A1(n_7585),
.A2(n_5828),
.B1(n_5885),
.B2(n_5867),
.Y(n_8404)
);

OAI21x1_ASAP7_75t_L g8405 ( 
.A1(n_7846),
.A2(n_7758),
.B(n_7613),
.Y(n_8405)
);

O2A1O1Ixp33_ASAP7_75t_L g8406 ( 
.A1(n_7361),
.A2(n_6380),
.B(n_6569),
.C(n_5849),
.Y(n_8406)
);

OAI21x1_ASAP7_75t_SL g8407 ( 
.A1(n_7346),
.A2(n_6830),
.B(n_5913),
.Y(n_8407)
);

OA21x2_ASAP7_75t_L g8408 ( 
.A1(n_7789),
.A2(n_6839),
.B(n_6807),
.Y(n_8408)
);

AOI22xp5_ASAP7_75t_L g8409 ( 
.A1(n_7585),
.A2(n_6845),
.B1(n_6759),
.B2(n_6821),
.Y(n_8409)
);

INVx3_ASAP7_75t_L g8410 ( 
.A(n_6940),
.Y(n_8410)
);

AND2x2_ASAP7_75t_L g8411 ( 
.A(n_7782),
.B(n_6262),
.Y(n_8411)
);

AND2x4_ASAP7_75t_L g8412 ( 
.A(n_6913),
.B(n_6311),
.Y(n_8412)
);

INVx2_ASAP7_75t_L g8413 ( 
.A(n_7015),
.Y(n_8413)
);

BUFx3_ASAP7_75t_L g8414 ( 
.A(n_7318),
.Y(n_8414)
);

AOI21x1_ASAP7_75t_L g8415 ( 
.A1(n_7770),
.A2(n_7820),
.B(n_7354),
.Y(n_8415)
);

NAND3xp33_ASAP7_75t_L g8416 ( 
.A(n_7467),
.B(n_6542),
.C(n_6514),
.Y(n_8416)
);

AOI22x1_ASAP7_75t_L g8417 ( 
.A1(n_7173),
.A2(n_7288),
.B1(n_7033),
.B2(n_7822),
.Y(n_8417)
);

OR2x2_ASAP7_75t_L g8418 ( 
.A(n_6964),
.B(n_7196),
.Y(n_8418)
);

INVxp33_ASAP7_75t_L g8419 ( 
.A(n_7895),
.Y(n_8419)
);

BUFx3_ASAP7_75t_L g8420 ( 
.A(n_7401),
.Y(n_8420)
);

INVx2_ASAP7_75t_L g8421 ( 
.A(n_7015),
.Y(n_8421)
);

NOR2xp67_ASAP7_75t_L g8422 ( 
.A(n_7579),
.B(n_6271),
.Y(n_8422)
);

NAND2xp5_ASAP7_75t_L g8423 ( 
.A(n_7093),
.B(n_6394),
.Y(n_8423)
);

AND2x4_ASAP7_75t_L g8424 ( 
.A(n_6913),
.B(n_6311),
.Y(n_8424)
);

BUFx3_ASAP7_75t_L g8425 ( 
.A(n_7401),
.Y(n_8425)
);

INVx2_ASAP7_75t_SL g8426 ( 
.A(n_7577),
.Y(n_8426)
);

NAND2x1p5_ASAP7_75t_L g8427 ( 
.A(n_7577),
.B(n_6546),
.Y(n_8427)
);

BUFx3_ASAP7_75t_L g8428 ( 
.A(n_7401),
.Y(n_8428)
);

AOI22xp33_ASAP7_75t_L g8429 ( 
.A1(n_7403),
.A2(n_6607),
.B1(n_5943),
.B2(n_5983),
.Y(n_8429)
);

BUFx6f_ASAP7_75t_L g8430 ( 
.A(n_6940),
.Y(n_8430)
);

AO21x2_ASAP7_75t_L g8431 ( 
.A1(n_7134),
.A2(n_6899),
.B(n_6681),
.Y(n_8431)
);

BUFx2_ASAP7_75t_SL g8432 ( 
.A(n_7577),
.Y(n_8432)
);

OAI21x1_ASAP7_75t_L g8433 ( 
.A1(n_7758),
.A2(n_7677),
.B(n_7653),
.Y(n_8433)
);

AOI22xp33_ASAP7_75t_L g8434 ( 
.A1(n_7004),
.A2(n_7200),
.B1(n_6929),
.B2(n_7032),
.Y(n_8434)
);

NAND2x1p5_ASAP7_75t_L g8435 ( 
.A(n_7577),
.B(n_6546),
.Y(n_8435)
);

AOI22xp33_ASAP7_75t_L g8436 ( 
.A1(n_7004),
.A2(n_5983),
.B1(n_5991),
.B2(n_5927),
.Y(n_8436)
);

INVx8_ASAP7_75t_L g8437 ( 
.A(n_7401),
.Y(n_8437)
);

NOR4xp25_ASAP7_75t_L g8438 ( 
.A(n_7800),
.B(n_5875),
.C(n_5913),
.D(n_5871),
.Y(n_8438)
);

OR2x2_ASAP7_75t_L g8439 ( 
.A(n_6964),
.B(n_6458),
.Y(n_8439)
);

AO21x2_ASAP7_75t_L g8440 ( 
.A1(n_7134),
.A2(n_6899),
.B(n_6643),
.Y(n_8440)
);

OAI21x1_ASAP7_75t_L g8441 ( 
.A1(n_7653),
.A2(n_6849),
.B(n_6826),
.Y(n_8441)
);

INVx1_ASAP7_75t_L g8442 ( 
.A(n_7730),
.Y(n_8442)
);

BUFx2_ASAP7_75t_L g8443 ( 
.A(n_7237),
.Y(n_8443)
);

AOI22xp33_ASAP7_75t_L g8444 ( 
.A1(n_7004),
.A2(n_5992),
.B1(n_6007),
.B2(n_5927),
.Y(n_8444)
);

NAND3xp33_ASAP7_75t_L g8445 ( 
.A(n_6929),
.B(n_5871),
.C(n_6576),
.Y(n_8445)
);

A2O1A1Ixp33_ASAP7_75t_L g8446 ( 
.A1(n_7044),
.A2(n_6759),
.B(n_6901),
.C(n_6876),
.Y(n_8446)
);

BUFx2_ASAP7_75t_L g8447 ( 
.A(n_7237),
.Y(n_8447)
);

OAI21x1_ASAP7_75t_L g8448 ( 
.A1(n_7653),
.A2(n_6849),
.B(n_6826),
.Y(n_8448)
);

AOI21x1_ASAP7_75t_L g8449 ( 
.A1(n_7770),
.A2(n_6643),
.B(n_6653),
.Y(n_8449)
);

A2O1A1Ixp33_ASAP7_75t_L g8450 ( 
.A1(n_7044),
.A2(n_6876),
.B(n_6901),
.C(n_6757),
.Y(n_8450)
);

OAI21x1_ASAP7_75t_L g8451 ( 
.A1(n_7653),
.A2(n_6849),
.B(n_6826),
.Y(n_8451)
);

OAI21x1_ASAP7_75t_L g8452 ( 
.A1(n_7653),
.A2(n_6849),
.B(n_6826),
.Y(n_8452)
);

AOI21xp33_ASAP7_75t_L g8453 ( 
.A1(n_7575),
.A2(n_5875),
.B(n_6611),
.Y(n_8453)
);

NOR2xp33_ASAP7_75t_SL g8454 ( 
.A(n_7581),
.B(n_6063),
.Y(n_8454)
);

AOI22xp33_ASAP7_75t_L g8455 ( 
.A1(n_7200),
.A2(n_6007),
.B1(n_6015),
.B2(n_5992),
.Y(n_8455)
);

OR2x2_ASAP7_75t_L g8456 ( 
.A(n_6964),
.B(n_6458),
.Y(n_8456)
);

O2A1O1Ixp33_ASAP7_75t_L g8457 ( 
.A1(n_6934),
.A2(n_6380),
.B(n_6569),
.C(n_5836),
.Y(n_8457)
);

OAI21x1_ASAP7_75t_SL g8458 ( 
.A1(n_7346),
.A2(n_6882),
.B(n_6611),
.Y(n_8458)
);

OAI21x1_ASAP7_75t_L g8459 ( 
.A1(n_7677),
.A2(n_6826),
.B(n_6904),
.Y(n_8459)
);

CKINVDCx16_ASAP7_75t_R g8460 ( 
.A(n_7384),
.Y(n_8460)
);

OAI21x1_ASAP7_75t_L g8461 ( 
.A1(n_7677),
.A2(n_6354),
.B(n_6903),
.Y(n_8461)
);

OAI21x1_ASAP7_75t_L g8462 ( 
.A1(n_7677),
.A2(n_7748),
.B(n_7802),
.Y(n_8462)
);

INVx4_ASAP7_75t_L g8463 ( 
.A(n_7445),
.Y(n_8463)
);

HB1xp67_ASAP7_75t_L g8464 ( 
.A(n_7260),
.Y(n_8464)
);

INVx2_ASAP7_75t_SL g8465 ( 
.A(n_7577),
.Y(n_8465)
);

OAI21x1_ASAP7_75t_L g8466 ( 
.A1(n_7677),
.A2(n_6354),
.B(n_6903),
.Y(n_8466)
);

OAI21x1_ASAP7_75t_L g8467 ( 
.A1(n_7748),
.A2(n_6763),
.B(n_6866),
.Y(n_8467)
);

BUFx6f_ASAP7_75t_L g8468 ( 
.A(n_6940),
.Y(n_8468)
);

INVx6_ASAP7_75t_L g8469 ( 
.A(n_7572),
.Y(n_8469)
);

OAI21xp5_ASAP7_75t_L g8470 ( 
.A1(n_7636),
.A2(n_5956),
.B(n_5836),
.Y(n_8470)
);

AOI222xp33_ASAP7_75t_L g8471 ( 
.A1(n_7271),
.A2(n_6934),
.B1(n_7764),
.B2(n_7773),
.C1(n_7005),
.C2(n_7362),
.Y(n_8471)
);

BUFx8_ASAP7_75t_L g8472 ( 
.A(n_7445),
.Y(n_8472)
);

XNOR2xp5_ASAP7_75t_L g8473 ( 
.A(n_7255),
.B(n_7830),
.Y(n_8473)
);

AO31x2_ASAP7_75t_L g8474 ( 
.A1(n_7832),
.A2(n_6866),
.A3(n_6757),
.B(n_6761),
.Y(n_8474)
);

INVx2_ASAP7_75t_L g8475 ( 
.A(n_7015),
.Y(n_8475)
);

OAI21x1_ASAP7_75t_L g8476 ( 
.A1(n_7748),
.A2(n_6763),
.B(n_6237),
.Y(n_8476)
);

OAI21x1_ASAP7_75t_L g8477 ( 
.A1(n_7748),
.A2(n_6237),
.B(n_6857),
.Y(n_8477)
);

OAI21xp5_ASAP7_75t_L g8478 ( 
.A1(n_7636),
.A2(n_7311),
.B(n_7308),
.Y(n_8478)
);

AOI22xp33_ASAP7_75t_L g8479 ( 
.A1(n_7032),
.A2(n_7189),
.B1(n_7764),
.B2(n_7773),
.Y(n_8479)
);

AND2x2_ASAP7_75t_L g8480 ( 
.A(n_7782),
.B(n_6291),
.Y(n_8480)
);

BUFx6f_ASAP7_75t_L g8481 ( 
.A(n_6949),
.Y(n_8481)
);

INVx1_ASAP7_75t_L g8482 ( 
.A(n_7730),
.Y(n_8482)
);

INVx1_ASAP7_75t_SL g8483 ( 
.A(n_7687),
.Y(n_8483)
);

NAND2xp5_ASAP7_75t_L g8484 ( 
.A(n_7099),
.B(n_6369),
.Y(n_8484)
);

INVx2_ASAP7_75t_L g8485 ( 
.A(n_7042),
.Y(n_8485)
);

INVx2_ASAP7_75t_L g8486 ( 
.A(n_7042),
.Y(n_8486)
);

INVx1_ASAP7_75t_L g8487 ( 
.A(n_7740),
.Y(n_8487)
);

AO21x2_ASAP7_75t_L g8488 ( 
.A1(n_7134),
.A2(n_6899),
.B(n_6807),
.Y(n_8488)
);

AO21x2_ASAP7_75t_L g8489 ( 
.A1(n_7134),
.A2(n_6899),
.B(n_6812),
.Y(n_8489)
);

AND2x2_ASAP7_75t_L g8490 ( 
.A(n_7824),
.B(n_6291),
.Y(n_8490)
);

NAND2xp5_ASAP7_75t_L g8491 ( 
.A(n_7099),
.B(n_6369),
.Y(n_8491)
);

BUFx6f_ASAP7_75t_L g8492 ( 
.A(n_6949),
.Y(n_8492)
);

OR2x2_ASAP7_75t_L g8493 ( 
.A(n_7055),
.B(n_6832),
.Y(n_8493)
);

OAI21x1_ASAP7_75t_L g8494 ( 
.A1(n_7748),
.A2(n_6857),
.B(n_6815),
.Y(n_8494)
);

OAI22xp5_ASAP7_75t_L g8495 ( 
.A1(n_7704),
.A2(n_6656),
.B1(n_6646),
.B2(n_6806),
.Y(n_8495)
);

CKINVDCx6p67_ASAP7_75t_R g8496 ( 
.A(n_7135),
.Y(n_8496)
);

AO21x2_ASAP7_75t_L g8497 ( 
.A1(n_7134),
.A2(n_6899),
.B(n_6812),
.Y(n_8497)
);

INVx1_ASAP7_75t_L g8498 ( 
.A(n_7740),
.Y(n_8498)
);

INVx3_ASAP7_75t_L g8499 ( 
.A(n_6949),
.Y(n_8499)
);

AND2x4_ASAP7_75t_L g8500 ( 
.A(n_6913),
.B(n_6364),
.Y(n_8500)
);

INVx1_ASAP7_75t_L g8501 ( 
.A(n_7740),
.Y(n_8501)
);

NOR2xp33_ASAP7_75t_L g8502 ( 
.A(n_7011),
.B(n_5971),
.Y(n_8502)
);

NAND2xp5_ASAP7_75t_L g8503 ( 
.A(n_7099),
.B(n_6463),
.Y(n_8503)
);

INVx1_ASAP7_75t_L g8504 ( 
.A(n_7746),
.Y(n_8504)
);

AOI22xp5_ASAP7_75t_L g8505 ( 
.A1(n_7308),
.A2(n_6761),
.B1(n_6315),
.B2(n_6183),
.Y(n_8505)
);

INVx4_ASAP7_75t_L g8506 ( 
.A(n_7445),
.Y(n_8506)
);

INVx2_ASAP7_75t_L g8507 ( 
.A(n_7042),
.Y(n_8507)
);

AND2x4_ASAP7_75t_L g8508 ( 
.A(n_6913),
.B(n_6435),
.Y(n_8508)
);

INVx2_ASAP7_75t_SL g8509 ( 
.A(n_7577),
.Y(n_8509)
);

OAI21x1_ASAP7_75t_L g8510 ( 
.A1(n_7140),
.A2(n_6774),
.B(n_6770),
.Y(n_8510)
);

INVx2_ASAP7_75t_L g8511 ( 
.A(n_7042),
.Y(n_8511)
);

INVx2_ASAP7_75t_SL g8512 ( 
.A(n_7577),
.Y(n_8512)
);

OAI21x1_ASAP7_75t_L g8513 ( 
.A1(n_7140),
.A2(n_7833),
.B(n_7321),
.Y(n_8513)
);

AO21x2_ASAP7_75t_L g8514 ( 
.A1(n_7789),
.A2(n_6797),
.B(n_6544),
.Y(n_8514)
);

O2A1O1Ixp33_ASAP7_75t_SL g8515 ( 
.A1(n_7035),
.A2(n_6804),
.B(n_6610),
.C(n_6005),
.Y(n_8515)
);

OAI21x1_ASAP7_75t_L g8516 ( 
.A1(n_7140),
.A2(n_7833),
.B(n_7321),
.Y(n_8516)
);

AOI21xp5_ASAP7_75t_L g8517 ( 
.A1(n_6976),
.A2(n_7007),
.B(n_6987),
.Y(n_8517)
);

AO21x2_ASAP7_75t_L g8518 ( 
.A1(n_7641),
.A2(n_7892),
.B(n_7799),
.Y(n_8518)
);

OAI22xp5_ASAP7_75t_L g8519 ( 
.A1(n_7704),
.A2(n_6656),
.B1(n_6646),
.B2(n_6806),
.Y(n_8519)
);

AND2x2_ASAP7_75t_L g8520 ( 
.A(n_7824),
.B(n_6317),
.Y(n_8520)
);

INVx1_ASAP7_75t_L g8521 ( 
.A(n_7746),
.Y(n_8521)
);

INVx1_ASAP7_75t_L g8522 ( 
.A(n_7746),
.Y(n_8522)
);

INVx1_ASAP7_75t_L g8523 ( 
.A(n_7749),
.Y(n_8523)
);

AOI221xp5_ASAP7_75t_L g8524 ( 
.A1(n_7710),
.A2(n_6797),
.B1(n_6533),
.B2(n_6528),
.C(n_6605),
.Y(n_8524)
);

NAND2x1p5_ASAP7_75t_L g8525 ( 
.A(n_7577),
.B(n_6546),
.Y(n_8525)
);

AOI22xp33_ASAP7_75t_L g8526 ( 
.A1(n_7032),
.A2(n_7189),
.B1(n_7271),
.B2(n_7488),
.Y(n_8526)
);

INVx1_ASAP7_75t_L g8527 ( 
.A(n_7749),
.Y(n_8527)
);

BUFx2_ASAP7_75t_L g8528 ( 
.A(n_7237),
.Y(n_8528)
);

A2O1A1Ixp33_ASAP7_75t_L g8529 ( 
.A1(n_7044),
.A2(n_6380),
.B(n_5910),
.C(n_5935),
.Y(n_8529)
);

OAI221xp5_ASAP7_75t_L g8530 ( 
.A1(n_7308),
.A2(n_5772),
.B1(n_6015),
.B2(n_6051),
.C(n_6022),
.Y(n_8530)
);

OAI21x1_ASAP7_75t_L g8531 ( 
.A1(n_7833),
.A2(n_6777),
.B(n_6770),
.Y(n_8531)
);

OAI21x1_ASAP7_75t_L g8532 ( 
.A1(n_7321),
.A2(n_6798),
.B(n_6777),
.Y(n_8532)
);

AO31x2_ASAP7_75t_L g8533 ( 
.A1(n_7832),
.A2(n_5824),
.A3(n_5845),
.B(n_5796),
.Y(n_8533)
);

AOI21xp5_ASAP7_75t_L g8534 ( 
.A1(n_6976),
.A2(n_6184),
.B(n_5956),
.Y(n_8534)
);

OAI22xp33_ASAP7_75t_L g8535 ( 
.A1(n_6943),
.A2(n_6683),
.B1(n_6396),
.B2(n_6691),
.Y(n_8535)
);

AOI21xp5_ASAP7_75t_L g8536 ( 
.A1(n_6987),
.A2(n_7024),
.B(n_7007),
.Y(n_8536)
);

AOI22xp5_ASAP7_75t_L g8537 ( 
.A1(n_7311),
.A2(n_7420),
.B1(n_7442),
.B2(n_7342),
.Y(n_8537)
);

A2O1A1Ixp33_ASAP7_75t_L g8538 ( 
.A1(n_7044),
.A2(n_5910),
.B(n_5935),
.C(n_5921),
.Y(n_8538)
);

CKINVDCx6p67_ASAP7_75t_R g8539 ( 
.A(n_7135),
.Y(n_8539)
);

OAI21xp5_ASAP7_75t_L g8540 ( 
.A1(n_7311),
.A2(n_5923),
.B(n_5924),
.Y(n_8540)
);

O2A1O1Ixp33_ASAP7_75t_SL g8541 ( 
.A1(n_7279),
.A2(n_6610),
.B(n_6005),
.C(n_6013),
.Y(n_8541)
);

INVx1_ASAP7_75t_L g8542 ( 
.A(n_7749),
.Y(n_8542)
);

OAI22xp33_ASAP7_75t_L g8543 ( 
.A1(n_7442),
.A2(n_7420),
.B1(n_7441),
.B2(n_7342),
.Y(n_8543)
);

AOI22xp33_ASAP7_75t_L g8544 ( 
.A1(n_7488),
.A2(n_6051),
.B1(n_6064),
.B2(n_6022),
.Y(n_8544)
);

AO31x2_ASAP7_75t_L g8545 ( 
.A1(n_7854),
.A2(n_5824),
.A3(n_5845),
.B(n_5796),
.Y(n_8545)
);

AO21x2_ASAP7_75t_L g8546 ( 
.A1(n_7641),
.A2(n_6544),
.B(n_6519),
.Y(n_8546)
);

OAI21x1_ASAP7_75t_L g8547 ( 
.A1(n_7898),
.A2(n_6288),
.B(n_6283),
.Y(n_8547)
);

CKINVDCx11_ASAP7_75t_R g8548 ( 
.A(n_7445),
.Y(n_8548)
);

OAI21x1_ASAP7_75t_L g8549 ( 
.A1(n_7898),
.A2(n_7024),
.B(n_7125),
.Y(n_8549)
);

NOR2xp67_ASAP7_75t_L g8550 ( 
.A(n_7579),
.B(n_7892),
.Y(n_8550)
);

INVx3_ASAP7_75t_L g8551 ( 
.A(n_6949),
.Y(n_8551)
);

AOI21x1_ASAP7_75t_L g8552 ( 
.A1(n_7820),
.A2(n_6853),
.B(n_6653),
.Y(n_8552)
);

OAI21x1_ASAP7_75t_L g8553 ( 
.A1(n_7898),
.A2(n_6288),
.B(n_6283),
.Y(n_8553)
);

AO21x2_ASAP7_75t_L g8554 ( 
.A1(n_7799),
.A2(n_6565),
.B(n_6758),
.Y(n_8554)
);

AOI21xp5_ASAP7_75t_L g8555 ( 
.A1(n_6978),
.A2(n_6184),
.B(n_6853),
.Y(n_8555)
);

BUFx2_ASAP7_75t_L g8556 ( 
.A(n_7237),
.Y(n_8556)
);

NAND2xp5_ASAP7_75t_L g8557 ( 
.A(n_7038),
.B(n_6463),
.Y(n_8557)
);

OAI21xp5_ASAP7_75t_L g8558 ( 
.A1(n_7663),
.A2(n_5923),
.B(n_5924),
.Y(n_8558)
);

AO21x1_ASAP7_75t_L g8559 ( 
.A1(n_7439),
.A2(n_6817),
.B(n_5921),
.Y(n_8559)
);

OAI21xp5_ASAP7_75t_L g8560 ( 
.A1(n_7663),
.A2(n_5772),
.B(n_6505),
.Y(n_8560)
);

OAI21x1_ASAP7_75t_L g8561 ( 
.A1(n_7898),
.A2(n_6288),
.B(n_6283),
.Y(n_8561)
);

CKINVDCx5p33_ASAP7_75t_R g8562 ( 
.A(n_7105),
.Y(n_8562)
);

INVx3_ASAP7_75t_L g8563 ( 
.A(n_6949),
.Y(n_8563)
);

AND2x2_ASAP7_75t_L g8564 ( 
.A(n_7824),
.B(n_7859),
.Y(n_8564)
);

OAI21x1_ASAP7_75t_L g8565 ( 
.A1(n_7125),
.A2(n_6288),
.B(n_6283),
.Y(n_8565)
);

NOR2x1_ASAP7_75t_SL g8566 ( 
.A(n_7521),
.B(n_6792),
.Y(n_8566)
);

AND2x2_ASAP7_75t_L g8567 ( 
.A(n_7859),
.B(n_6317),
.Y(n_8567)
);

INVx1_ASAP7_75t_L g8568 ( 
.A(n_7754),
.Y(n_8568)
);

INVx2_ASAP7_75t_L g8569 ( 
.A(n_7054),
.Y(n_8569)
);

OAI21xp5_ASAP7_75t_L g8570 ( 
.A1(n_7342),
.A2(n_6522),
.B(n_6505),
.Y(n_8570)
);

OAI22xp5_ASAP7_75t_L g8571 ( 
.A1(n_7588),
.A2(n_6822),
.B1(n_6824),
.B2(n_6814),
.Y(n_8571)
);

OA21x2_ASAP7_75t_L g8572 ( 
.A1(n_7680),
.A2(n_6335),
.B(n_6331),
.Y(n_8572)
);

INVx2_ASAP7_75t_L g8573 ( 
.A(n_7054),
.Y(n_8573)
);

AO21x2_ASAP7_75t_L g8574 ( 
.A1(n_7799),
.A2(n_6565),
.B(n_6758),
.Y(n_8574)
);

NAND2xp5_ASAP7_75t_L g8575 ( 
.A(n_7038),
.B(n_5840),
.Y(n_8575)
);

INVx2_ASAP7_75t_L g8576 ( 
.A(n_7054),
.Y(n_8576)
);

INVx2_ASAP7_75t_L g8577 ( 
.A(n_7054),
.Y(n_8577)
);

INVx2_ASAP7_75t_L g8578 ( 
.A(n_7061),
.Y(n_8578)
);

AND2x4_ASAP7_75t_L g8579 ( 
.A(n_6913),
.B(n_6374),
.Y(n_8579)
);

INVx2_ASAP7_75t_L g8580 ( 
.A(n_7061),
.Y(n_8580)
);

AND2x2_ASAP7_75t_L g8581 ( 
.A(n_7859),
.B(n_6402),
.Y(n_8581)
);

OAI21x1_ASAP7_75t_L g8582 ( 
.A1(n_7125),
.A2(n_6314),
.B(n_6283),
.Y(n_8582)
);

AO21x2_ASAP7_75t_L g8583 ( 
.A1(n_7685),
.A2(n_7203),
.B(n_7182),
.Y(n_8583)
);

INVx1_ASAP7_75t_L g8584 ( 
.A(n_7754),
.Y(n_8584)
);

OAI21x1_ASAP7_75t_L g8585 ( 
.A1(n_7125),
.A2(n_6383),
.B(n_6314),
.Y(n_8585)
);

OAI21x1_ASAP7_75t_L g8586 ( 
.A1(n_7125),
.A2(n_6383),
.B(n_6314),
.Y(n_8586)
);

AOI22xp5_ASAP7_75t_L g8587 ( 
.A1(n_7420),
.A2(n_6064),
.B1(n_6072),
.B2(n_6067),
.Y(n_8587)
);

OA21x2_ASAP7_75t_L g8588 ( 
.A1(n_7680),
.A2(n_6345),
.B(n_6335),
.Y(n_8588)
);

NAND2xp33_ASAP7_75t_L g8589 ( 
.A(n_7033),
.B(n_6683),
.Y(n_8589)
);

AND2x2_ASAP7_75t_L g8590 ( 
.A(n_7448),
.B(n_6402),
.Y(n_8590)
);

AOI21x1_ASAP7_75t_L g8591 ( 
.A1(n_7820),
.A2(n_7310),
.B(n_7459),
.Y(n_8591)
);

AOI21xp5_ASAP7_75t_L g8592 ( 
.A1(n_6978),
.A2(n_6184),
.B(n_6891),
.Y(n_8592)
);

OAI21x1_ASAP7_75t_L g8593 ( 
.A1(n_7199),
.A2(n_6383),
.B(n_6314),
.Y(n_8593)
);

OAI22xp33_ASAP7_75t_L g8594 ( 
.A1(n_7442),
.A2(n_6683),
.B1(n_6784),
.B2(n_6691),
.Y(n_8594)
);

OAI22xp33_ASAP7_75t_L g8595 ( 
.A1(n_7441),
.A2(n_6784),
.B1(n_6189),
.B2(n_6207),
.Y(n_8595)
);

O2A1O1Ixp33_ASAP7_75t_SL g8596 ( 
.A1(n_7172),
.A2(n_5971),
.B(n_6014),
.C(n_6013),
.Y(n_8596)
);

AOI21x1_ASAP7_75t_L g8597 ( 
.A1(n_7459),
.A2(n_6891),
.B(n_6865),
.Y(n_8597)
);

AO21x2_ASAP7_75t_L g8598 ( 
.A1(n_7685),
.A2(n_7203),
.B(n_7182),
.Y(n_8598)
);

AOI21xp33_ASAP7_75t_SL g8599 ( 
.A1(n_7395),
.A2(n_5931),
.B(n_6432),
.Y(n_8599)
);

OAI21x1_ASAP7_75t_SL g8600 ( 
.A1(n_7506),
.A2(n_5771),
.B(n_5768),
.Y(n_8600)
);

OAI21x1_ASAP7_75t_L g8601 ( 
.A1(n_7199),
.A2(n_6383),
.B(n_6314),
.Y(n_8601)
);

CKINVDCx14_ASAP7_75t_R g8602 ( 
.A(n_7105),
.Y(n_8602)
);

OAI21x1_ASAP7_75t_L g8603 ( 
.A1(n_7199),
.A2(n_6393),
.B(n_6383),
.Y(n_8603)
);

BUFx3_ASAP7_75t_L g8604 ( 
.A(n_7456),
.Y(n_8604)
);

NAND2xp33_ASAP7_75t_L g8605 ( 
.A(n_7370),
.B(n_5780),
.Y(n_8605)
);

CKINVDCx6p67_ASAP7_75t_R g8606 ( 
.A(n_7135),
.Y(n_8606)
);

OAI21x1_ASAP7_75t_L g8607 ( 
.A1(n_7199),
.A2(n_6410),
.B(n_6393),
.Y(n_8607)
);

BUFx6f_ASAP7_75t_L g8608 ( 
.A(n_6949),
.Y(n_8608)
);

NAND2x1p5_ASAP7_75t_L g8609 ( 
.A(n_7577),
.B(n_6708),
.Y(n_8609)
);

A2O1A1Ixp33_ASAP7_75t_L g8610 ( 
.A1(n_7044),
.A2(n_6865),
.B(n_6659),
.C(n_6750),
.Y(n_8610)
);

OAI22xp5_ASAP7_75t_L g8611 ( 
.A1(n_7588),
.A2(n_6822),
.B1(n_6824),
.B2(n_6814),
.Y(n_8611)
);

NOR2x1_ASAP7_75t_SL g8612 ( 
.A(n_7521),
.B(n_6792),
.Y(n_8612)
);

INVx1_ASAP7_75t_SL g8613 ( 
.A(n_7687),
.Y(n_8613)
);

INVx1_ASAP7_75t_L g8614 ( 
.A(n_7754),
.Y(n_8614)
);

AND2x4_ASAP7_75t_L g8615 ( 
.A(n_6924),
.B(n_6311),
.Y(n_8615)
);

AOI222xp33_ASAP7_75t_L g8616 ( 
.A1(n_7005),
.A2(n_6095),
.B1(n_6067),
.B2(n_6127),
.C1(n_6116),
.C2(n_6072),
.Y(n_8616)
);

BUFx3_ASAP7_75t_L g8617 ( 
.A(n_7456),
.Y(n_8617)
);

AOI22xp33_ASAP7_75t_L g8618 ( 
.A1(n_7490),
.A2(n_6093),
.B1(n_6116),
.B2(n_6095),
.Y(n_8618)
);

INVx1_ASAP7_75t_L g8619 ( 
.A(n_7761),
.Y(n_8619)
);

INVx2_ASAP7_75t_L g8620 ( 
.A(n_7061),
.Y(n_8620)
);

A2O1A1Ixp33_ASAP7_75t_L g8621 ( 
.A1(n_7051),
.A2(n_6659),
.B(n_6750),
.C(n_6670),
.Y(n_8621)
);

OAI21x1_ASAP7_75t_L g8622 ( 
.A1(n_7199),
.A2(n_6410),
.B(n_6393),
.Y(n_8622)
);

AOI21xp5_ASAP7_75t_L g8623 ( 
.A1(n_6978),
.A2(n_6184),
.B(n_6794),
.Y(n_8623)
);

AND2x4_ASAP7_75t_L g8624 ( 
.A(n_6924),
.B(n_6311),
.Y(n_8624)
);

INVx1_ASAP7_75t_L g8625 ( 
.A(n_7761),
.Y(n_8625)
);

AO21x2_ASAP7_75t_L g8626 ( 
.A1(n_7685),
.A2(n_6620),
.B(n_6619),
.Y(n_8626)
);

OAI21x1_ASAP7_75t_L g8627 ( 
.A1(n_7223),
.A2(n_6410),
.B(n_6393),
.Y(n_8627)
);

AOI22xp33_ASAP7_75t_L g8628 ( 
.A1(n_7490),
.A2(n_6093),
.B1(n_6136),
.B2(n_6127),
.Y(n_8628)
);

AO31x2_ASAP7_75t_L g8629 ( 
.A1(n_7854),
.A2(n_5979),
.A3(n_6026),
.B(n_5858),
.Y(n_8629)
);

OAI21x1_ASAP7_75t_L g8630 ( 
.A1(n_7223),
.A2(n_6410),
.B(n_6393),
.Y(n_8630)
);

OAI21x1_ASAP7_75t_L g8631 ( 
.A1(n_7223),
.A2(n_6431),
.B(n_6410),
.Y(n_8631)
);

NAND2xp5_ASAP7_75t_SL g8632 ( 
.A(n_7051),
.B(n_6311),
.Y(n_8632)
);

BUFx3_ASAP7_75t_L g8633 ( 
.A(n_7456),
.Y(n_8633)
);

INVx1_ASAP7_75t_L g8634 ( 
.A(n_7761),
.Y(n_8634)
);

OAI22xp33_ASAP7_75t_L g8635 ( 
.A1(n_7441),
.A2(n_6273),
.B1(n_6289),
.B2(n_6192),
.Y(n_8635)
);

OAI21xp5_ASAP7_75t_L g8636 ( 
.A1(n_7800),
.A2(n_6522),
.B(n_6139),
.Y(n_8636)
);

OAI21x1_ASAP7_75t_L g8637 ( 
.A1(n_7223),
.A2(n_6441),
.B(n_6431),
.Y(n_8637)
);

OAI21x1_ASAP7_75t_L g8638 ( 
.A1(n_7223),
.A2(n_6441),
.B(n_6431),
.Y(n_8638)
);

BUFx6f_ASAP7_75t_L g8639 ( 
.A(n_6949),
.Y(n_8639)
);

INVx2_ASAP7_75t_L g8640 ( 
.A(n_7061),
.Y(n_8640)
);

AO21x2_ASAP7_75t_L g8641 ( 
.A1(n_7685),
.A2(n_6620),
.B(n_6619),
.Y(n_8641)
);

INVx1_ASAP7_75t_L g8642 ( 
.A(n_7765),
.Y(n_8642)
);

INVx2_ASAP7_75t_SL g8643 ( 
.A(n_7577),
.Y(n_8643)
);

OAI22xp5_ASAP7_75t_L g8644 ( 
.A1(n_7634),
.A2(n_7091),
.B1(n_6952),
.B2(n_7581),
.Y(n_8644)
);

AND2x2_ASAP7_75t_L g8645 ( 
.A(n_7448),
.B(n_6407),
.Y(n_8645)
);

OA21x2_ASAP7_75t_L g8646 ( 
.A1(n_7453),
.A2(n_6346),
.B(n_6345),
.Y(n_8646)
);

HB1xp67_ASAP7_75t_L g8647 ( 
.A(n_7260),
.Y(n_8647)
);

INVx1_ASAP7_75t_L g8648 ( 
.A(n_7765),
.Y(n_8648)
);

INVx1_ASAP7_75t_L g8649 ( 
.A(n_7765),
.Y(n_8649)
);

AND2x2_ASAP7_75t_L g8650 ( 
.A(n_7448),
.B(n_6407),
.Y(n_8650)
);

INVx6_ASAP7_75t_L g8651 ( 
.A(n_7572),
.Y(n_8651)
);

AND2x2_ASAP7_75t_L g8652 ( 
.A(n_7448),
.B(n_7489),
.Y(n_8652)
);

BUFx2_ASAP7_75t_L g8653 ( 
.A(n_7237),
.Y(n_8653)
);

HB1xp67_ASAP7_75t_L g8654 ( 
.A(n_7280),
.Y(n_8654)
);

AO21x2_ASAP7_75t_L g8655 ( 
.A1(n_7685),
.A2(n_6625),
.B(n_6624),
.Y(n_8655)
);

OAI21x1_ASAP7_75t_L g8656 ( 
.A1(n_7259),
.A2(n_7306),
.B(n_7300),
.Y(n_8656)
);

AO21x2_ASAP7_75t_L g8657 ( 
.A1(n_7685),
.A2(n_6625),
.B(n_6624),
.Y(n_8657)
);

INVx2_ASAP7_75t_L g8658 ( 
.A(n_7068),
.Y(n_8658)
);

O2A1O1Ixp33_ASAP7_75t_L g8659 ( 
.A1(n_7016),
.A2(n_6817),
.B(n_5970),
.C(n_6059),
.Y(n_8659)
);

INVx2_ASAP7_75t_L g8660 ( 
.A(n_7068),
.Y(n_8660)
);

AO22x2_ASAP7_75t_L g8661 ( 
.A1(n_7241),
.A2(n_6170),
.B1(n_6167),
.B2(n_6361),
.Y(n_8661)
);

AOI22xp33_ASAP7_75t_SL g8662 ( 
.A1(n_6972),
.A2(n_6760),
.B1(n_6686),
.B2(n_6109),
.Y(n_8662)
);

INVx2_ASAP7_75t_L g8663 ( 
.A(n_7068),
.Y(n_8663)
);

INVx1_ASAP7_75t_L g8664 ( 
.A(n_7771),
.Y(n_8664)
);

AO21x2_ASAP7_75t_L g8665 ( 
.A1(n_7182),
.A2(n_6651),
.B(n_6636),
.Y(n_8665)
);

AND2x2_ASAP7_75t_L g8666 ( 
.A(n_7489),
.B(n_6440),
.Y(n_8666)
);

INVx1_ASAP7_75t_SL g8667 ( 
.A(n_7687),
.Y(n_8667)
);

INVx3_ASAP7_75t_L g8668 ( 
.A(n_6949),
.Y(n_8668)
);

AO21x1_ASAP7_75t_L g8669 ( 
.A1(n_7439),
.A2(n_5970),
.B(n_6184),
.Y(n_8669)
);

INVx2_ASAP7_75t_L g8670 ( 
.A(n_7068),
.Y(n_8670)
);

INVx2_ASAP7_75t_SL g8671 ( 
.A(n_7587),
.Y(n_8671)
);

INVx3_ASAP7_75t_L g8672 ( 
.A(n_6949),
.Y(n_8672)
);

INVx2_ASAP7_75t_L g8673 ( 
.A(n_7072),
.Y(n_8673)
);

CKINVDCx20_ASAP7_75t_R g8674 ( 
.A(n_7255),
.Y(n_8674)
);

AOI21xp5_ASAP7_75t_L g8675 ( 
.A1(n_7592),
.A2(n_6184),
.B(n_6794),
.Y(n_8675)
);

AOI21xp5_ASAP7_75t_L g8676 ( 
.A1(n_7592),
.A2(n_6799),
.B(n_6794),
.Y(n_8676)
);

CKINVDCx5p33_ASAP7_75t_R g8677 ( 
.A(n_7129),
.Y(n_8677)
);

INVx2_ASAP7_75t_L g8678 ( 
.A(n_7072),
.Y(n_8678)
);

INVx2_ASAP7_75t_L g8679 ( 
.A(n_7072),
.Y(n_8679)
);

AOI21xp5_ASAP7_75t_L g8680 ( 
.A1(n_7592),
.A2(n_6799),
.B(n_6794),
.Y(n_8680)
);

BUFx2_ASAP7_75t_L g8681 ( 
.A(n_7237),
.Y(n_8681)
);

NAND2xp5_ASAP7_75t_L g8682 ( 
.A(n_7038),
.B(n_5840),
.Y(n_8682)
);

INVx3_ASAP7_75t_L g8683 ( 
.A(n_6949),
.Y(n_8683)
);

BUFx3_ASAP7_75t_L g8684 ( 
.A(n_7456),
.Y(n_8684)
);

INVx4_ASAP7_75t_L g8685 ( 
.A(n_7539),
.Y(n_8685)
);

AND2x4_ASAP7_75t_L g8686 ( 
.A(n_6924),
.B(n_6364),
.Y(n_8686)
);

INVx1_ASAP7_75t_L g8687 ( 
.A(n_7771),
.Y(n_8687)
);

INVx3_ASAP7_75t_L g8688 ( 
.A(n_6973),
.Y(n_8688)
);

NAND2xp5_ASAP7_75t_L g8689 ( 
.A(n_7055),
.B(n_6694),
.Y(n_8689)
);

INVx1_ASAP7_75t_L g8690 ( 
.A(n_7771),
.Y(n_8690)
);

NAND2xp5_ASAP7_75t_L g8691 ( 
.A(n_7055),
.B(n_6694),
.Y(n_8691)
);

A2O1A1Ixp33_ASAP7_75t_L g8692 ( 
.A1(n_7051),
.A2(n_6670),
.B(n_6690),
.C(n_6663),
.Y(n_8692)
);

INVx5_ASAP7_75t_SL g8693 ( 
.A(n_7013),
.Y(n_8693)
);

OR2x2_ASAP7_75t_L g8694 ( 
.A(n_6911),
.B(n_6832),
.Y(n_8694)
);

CKINVDCx16_ASAP7_75t_R g8695 ( 
.A(n_7384),
.Y(n_8695)
);

INVx8_ASAP7_75t_L g8696 ( 
.A(n_7539),
.Y(n_8696)
);

INVx1_ASAP7_75t_L g8697 ( 
.A(n_7788),
.Y(n_8697)
);

AOI21xp5_ASAP7_75t_L g8698 ( 
.A1(n_7136),
.A2(n_6799),
.B(n_6794),
.Y(n_8698)
);

AO21x2_ASAP7_75t_L g8699 ( 
.A1(n_7203),
.A2(n_6651),
.B(n_6636),
.Y(n_8699)
);

AOI22xp33_ASAP7_75t_SL g8700 ( 
.A1(n_6972),
.A2(n_6760),
.B1(n_6109),
.B2(n_6241),
.Y(n_8700)
);

INVx2_ASAP7_75t_L g8701 ( 
.A(n_7072),
.Y(n_8701)
);

OAI22xp5_ASAP7_75t_L g8702 ( 
.A1(n_7634),
.A2(n_7091),
.B1(n_6952),
.B2(n_7315),
.Y(n_8702)
);

INVx1_ASAP7_75t_L g8703 ( 
.A(n_7788),
.Y(n_8703)
);

AO31x2_ASAP7_75t_L g8704 ( 
.A1(n_7822),
.A2(n_5979),
.A3(n_6026),
.B(n_5858),
.Y(n_8704)
);

OAI21x1_ASAP7_75t_SL g8705 ( 
.A1(n_7506),
.A2(n_5771),
.B(n_5768),
.Y(n_8705)
);

OA21x2_ASAP7_75t_L g8706 ( 
.A1(n_7453),
.A2(n_6356),
.B(n_6346),
.Y(n_8706)
);

INVx2_ASAP7_75t_L g8707 ( 
.A(n_7076),
.Y(n_8707)
);

INVx1_ASAP7_75t_SL g8708 ( 
.A(n_7693),
.Y(n_8708)
);

AO21x2_ASAP7_75t_L g8709 ( 
.A1(n_7169),
.A2(n_6660),
.B(n_6652),
.Y(n_8709)
);

OAI22xp5_ASAP7_75t_L g8710 ( 
.A1(n_7315),
.A2(n_6880),
.B1(n_6894),
.B2(n_6852),
.Y(n_8710)
);

HB1xp67_ASAP7_75t_L g8711 ( 
.A(n_7280),
.Y(n_8711)
);

AOI22xp33_ASAP7_75t_L g8712 ( 
.A1(n_7231),
.A2(n_6139),
.B1(n_6145),
.B2(n_6136),
.Y(n_8712)
);

AOI21xp5_ASAP7_75t_L g8713 ( 
.A1(n_7136),
.A2(n_7337),
.B(n_7586),
.Y(n_8713)
);

INVx2_ASAP7_75t_SL g8714 ( 
.A(n_7587),
.Y(n_8714)
);

OR2x2_ASAP7_75t_L g8715 ( 
.A(n_6911),
.B(n_6986),
.Y(n_8715)
);

AO31x2_ASAP7_75t_L g8716 ( 
.A1(n_7822),
.A2(n_6053),
.A3(n_6065),
.B(n_6038),
.Y(n_8716)
);

BUFx3_ASAP7_75t_L g8717 ( 
.A(n_7539),
.Y(n_8717)
);

OR2x2_ASAP7_75t_L g8718 ( 
.A(n_6911),
.B(n_6841),
.Y(n_8718)
);

OAI21xp5_ASAP7_75t_L g8719 ( 
.A1(n_7575),
.A2(n_6151),
.B(n_6145),
.Y(n_8719)
);

NAND2xp5_ASAP7_75t_L g8720 ( 
.A(n_7070),
.B(n_6735),
.Y(n_8720)
);

AND2x2_ASAP7_75t_L g8721 ( 
.A(n_7489),
.B(n_7540),
.Y(n_8721)
);

CKINVDCx16_ASAP7_75t_R g8722 ( 
.A(n_7384),
.Y(n_8722)
);

OAI21x1_ASAP7_75t_L g8723 ( 
.A1(n_7300),
.A2(n_7364),
.B(n_7306),
.Y(n_8723)
);

NAND2xp5_ASAP7_75t_L g8724 ( 
.A(n_7070),
.B(n_7027),
.Y(n_8724)
);

INVx1_ASAP7_75t_SL g8725 ( 
.A(n_7693),
.Y(n_8725)
);

INVx2_ASAP7_75t_L g8726 ( 
.A(n_7076),
.Y(n_8726)
);

INVx2_ASAP7_75t_L g8727 ( 
.A(n_7076),
.Y(n_8727)
);

INVxp67_ASAP7_75t_SL g8728 ( 
.A(n_7302),
.Y(n_8728)
);

AOI22xp33_ASAP7_75t_L g8729 ( 
.A1(n_7231),
.A2(n_6151),
.B1(n_6189),
.B2(n_6172),
.Y(n_8729)
);

AOI22xp33_ASAP7_75t_SL g8730 ( 
.A1(n_6972),
.A2(n_6760),
.B1(n_6109),
.B2(n_6241),
.Y(n_8730)
);

AND2x2_ASAP7_75t_L g8731 ( 
.A(n_7489),
.B(n_6440),
.Y(n_8731)
);

AO21x2_ASAP7_75t_L g8732 ( 
.A1(n_7169),
.A2(n_6660),
.B(n_6652),
.Y(n_8732)
);

INVx1_ASAP7_75t_L g8733 ( 
.A(n_7788),
.Y(n_8733)
);

OA21x2_ASAP7_75t_L g8734 ( 
.A1(n_7474),
.A2(n_6968),
.B(n_7627),
.Y(n_8734)
);

AOI21xp5_ASAP7_75t_L g8735 ( 
.A1(n_7136),
.A2(n_6799),
.B(n_6794),
.Y(n_8735)
);

AND2x2_ASAP7_75t_L g8736 ( 
.A(n_7540),
.B(n_6446),
.Y(n_8736)
);

OR2x2_ASAP7_75t_L g8737 ( 
.A(n_6986),
.B(n_6841),
.Y(n_8737)
);

NAND2xp5_ASAP7_75t_L g8738 ( 
.A(n_7070),
.B(n_6735),
.Y(n_8738)
);

OAI21x1_ASAP7_75t_SL g8739 ( 
.A1(n_7506),
.A2(n_5771),
.B(n_5768),
.Y(n_8739)
);

CKINVDCx5p33_ASAP7_75t_R g8740 ( 
.A(n_7129),
.Y(n_8740)
);

INVx2_ASAP7_75t_L g8741 ( 
.A(n_7076),
.Y(n_8741)
);

INVx1_ASAP7_75t_L g8742 ( 
.A(n_7794),
.Y(n_8742)
);

AND2x2_ASAP7_75t_L g8743 ( 
.A(n_7540),
.B(n_6446),
.Y(n_8743)
);

BUFx3_ASAP7_75t_L g8744 ( 
.A(n_7539),
.Y(n_8744)
);

AND2x4_ASAP7_75t_L g8745 ( 
.A(n_6924),
.B(n_6416),
.Y(n_8745)
);

INVx2_ASAP7_75t_L g8746 ( 
.A(n_7083),
.Y(n_8746)
);

NAND2x1p5_ASAP7_75t_L g8747 ( 
.A(n_7587),
.B(n_6708),
.Y(n_8747)
);

AO21x2_ASAP7_75t_L g8748 ( 
.A1(n_7169),
.A2(n_6667),
.B(n_6662),
.Y(n_8748)
);

INVxp67_ASAP7_75t_SL g8749 ( 
.A(n_7302),
.Y(n_8749)
);

OAI22xp33_ASAP7_75t_L g8750 ( 
.A1(n_7455),
.A2(n_6338),
.B1(n_6261),
.B2(n_6172),
.Y(n_8750)
);

AO31x2_ASAP7_75t_L g8751 ( 
.A1(n_7762),
.A2(n_6053),
.A3(n_6065),
.B(n_6038),
.Y(n_8751)
);

BUFx10_ASAP7_75t_L g8752 ( 
.A(n_7408),
.Y(n_8752)
);

BUFx3_ASAP7_75t_L g8753 ( 
.A(n_7686),
.Y(n_8753)
);

INVx3_ASAP7_75t_L g8754 ( 
.A(n_6973),
.Y(n_8754)
);

OAI21xp5_ASAP7_75t_L g8755 ( 
.A1(n_7066),
.A2(n_6194),
.B(n_6192),
.Y(n_8755)
);

BUFx3_ASAP7_75t_L g8756 ( 
.A(n_7686),
.Y(n_8756)
);

AO21x2_ASAP7_75t_L g8757 ( 
.A1(n_7459),
.A2(n_6667),
.B(n_6662),
.Y(n_8757)
);

INVx5_ASAP7_75t_L g8758 ( 
.A(n_6973),
.Y(n_8758)
);

NOR3xp33_ASAP7_75t_SL g8759 ( 
.A(n_7139),
.B(n_5958),
.C(n_5950),
.Y(n_8759)
);

AO21x2_ASAP7_75t_L g8760 ( 
.A1(n_7512),
.A2(n_6671),
.B(n_6668),
.Y(n_8760)
);

INVx1_ASAP7_75t_L g8761 ( 
.A(n_7794),
.Y(n_8761)
);

AO21x2_ASAP7_75t_L g8762 ( 
.A1(n_7512),
.A2(n_6671),
.B(n_6668),
.Y(n_8762)
);

BUFx2_ASAP7_75t_L g8763 ( 
.A(n_7237),
.Y(n_8763)
);

INVx5_ASAP7_75t_L g8764 ( 
.A(n_6973),
.Y(n_8764)
);

AND2x4_ASAP7_75t_L g8765 ( 
.A(n_6924),
.B(n_6374),
.Y(n_8765)
);

AOI21xp5_ASAP7_75t_SL g8766 ( 
.A1(n_7370),
.A2(n_6799),
.B(n_5917),
.Y(n_8766)
);

AND2x4_ASAP7_75t_L g8767 ( 
.A(n_6924),
.B(n_6374),
.Y(n_8767)
);

NAND2x1p5_ASAP7_75t_L g8768 ( 
.A(n_7587),
.B(n_6708),
.Y(n_8768)
);

INVxp67_ASAP7_75t_L g8769 ( 
.A(n_7434),
.Y(n_8769)
);

HB1xp67_ASAP7_75t_L g8770 ( 
.A(n_7336),
.Y(n_8770)
);

A2O1A1Ixp33_ASAP7_75t_L g8771 ( 
.A1(n_7051),
.A2(n_6690),
.B(n_6663),
.C(n_6605),
.Y(n_8771)
);

AO21x1_ASAP7_75t_L g8772 ( 
.A1(n_7066),
.A2(n_5789),
.B(n_5932),
.Y(n_8772)
);

INVx2_ASAP7_75t_L g8773 ( 
.A(n_7083),
.Y(n_8773)
);

INVx3_ASAP7_75t_L g8774 ( 
.A(n_6973),
.Y(n_8774)
);

INVx2_ASAP7_75t_L g8775 ( 
.A(n_7083),
.Y(n_8775)
);

INVx1_ASAP7_75t_SL g8776 ( 
.A(n_7693),
.Y(n_8776)
);

INVx1_ASAP7_75t_L g8777 ( 
.A(n_7794),
.Y(n_8777)
);

NOR2x1_ASAP7_75t_SL g8778 ( 
.A(n_7521),
.B(n_6792),
.Y(n_8778)
);

INVx1_ASAP7_75t_L g8779 ( 
.A(n_7796),
.Y(n_8779)
);

BUFx3_ASAP7_75t_L g8780 ( 
.A(n_7686),
.Y(n_8780)
);

NAND2x1p5_ASAP7_75t_L g8781 ( 
.A(n_7587),
.B(n_6708),
.Y(n_8781)
);

AOI21x1_ASAP7_75t_L g8782 ( 
.A1(n_7116),
.A2(n_6719),
.B(n_6697),
.Y(n_8782)
);

NOR2xp33_ASAP7_75t_L g8783 ( 
.A(n_7011),
.B(n_6014),
.Y(n_8783)
);

AOI21xp5_ASAP7_75t_L g8784 ( 
.A1(n_7337),
.A2(n_6799),
.B(n_6792),
.Y(n_8784)
);

AO21x2_ASAP7_75t_L g8785 ( 
.A1(n_7512),
.A2(n_6693),
.B(n_6680),
.Y(n_8785)
);

INVx1_ASAP7_75t_L g8786 ( 
.A(n_7796),
.Y(n_8786)
);

O2A1O1Ixp33_ASAP7_75t_L g8787 ( 
.A1(n_7016),
.A2(n_6059),
.B(n_6202),
.C(n_6194),
.Y(n_8787)
);

INVx5_ASAP7_75t_L g8788 ( 
.A(n_6973),
.Y(n_8788)
);

OA21x2_ASAP7_75t_L g8789 ( 
.A1(n_7474),
.A2(n_6358),
.B(n_6356),
.Y(n_8789)
);

AO21x2_ASAP7_75t_L g8790 ( 
.A1(n_7249),
.A2(n_6693),
.B(n_6680),
.Y(n_8790)
);

A2O1A1Ixp33_ASAP7_75t_L g8791 ( 
.A1(n_7051),
.A2(n_6599),
.B(n_6207),
.C(n_6224),
.Y(n_8791)
);

BUFx2_ASAP7_75t_L g8792 ( 
.A(n_7237),
.Y(n_8792)
);

AND2x2_ASAP7_75t_L g8793 ( 
.A(n_7540),
.B(n_6455),
.Y(n_8793)
);

AO21x2_ASAP7_75t_L g8794 ( 
.A1(n_7249),
.A2(n_6705),
.B(n_6700),
.Y(n_8794)
);

INVx1_ASAP7_75t_L g8795 ( 
.A(n_7796),
.Y(n_8795)
);

INVx2_ASAP7_75t_SL g8796 ( 
.A(n_7587),
.Y(n_8796)
);

BUFx4f_ASAP7_75t_L g8797 ( 
.A(n_7686),
.Y(n_8797)
);

INVx1_ASAP7_75t_L g8798 ( 
.A(n_7815),
.Y(n_8798)
);

OAI21xp5_ASAP7_75t_L g8799 ( 
.A1(n_7500),
.A2(n_6224),
.B(n_6202),
.Y(n_8799)
);

NAND2x1p5_ASAP7_75t_L g8800 ( 
.A(n_7587),
.B(n_6708),
.Y(n_8800)
);

AO21x2_ASAP7_75t_L g8801 ( 
.A1(n_7249),
.A2(n_6968),
.B(n_7243),
.Y(n_8801)
);

OA21x2_ASAP7_75t_L g8802 ( 
.A1(n_6968),
.A2(n_6360),
.B(n_6358),
.Y(n_8802)
);

INVx1_ASAP7_75t_L g8803 ( 
.A(n_7815),
.Y(n_8803)
);

AND2x4_ASAP7_75t_L g8804 ( 
.A(n_6924),
.B(n_6399),
.Y(n_8804)
);

AO31x2_ASAP7_75t_L g8805 ( 
.A1(n_7762),
.A2(n_6133),
.A3(n_6141),
.B(n_6086),
.Y(n_8805)
);

OR2x2_ASAP7_75t_L g8806 ( 
.A(n_6986),
.B(n_7030),
.Y(n_8806)
);

INVx2_ASAP7_75t_L g8807 ( 
.A(n_7083),
.Y(n_8807)
);

OAI22xp33_ASAP7_75t_SL g8808 ( 
.A1(n_7156),
.A2(n_6250),
.B1(n_6261),
.B2(n_6242),
.Y(n_8808)
);

NAND2xp5_ASAP7_75t_L g8809 ( 
.A(n_7027),
.B(n_6820),
.Y(n_8809)
);

NAND3xp33_ASAP7_75t_L g8810 ( 
.A(n_7016),
.B(n_6250),
.C(n_6242),
.Y(n_8810)
);

AOI22xp33_ASAP7_75t_L g8811 ( 
.A1(n_7250),
.A2(n_6263),
.B1(n_6284),
.B2(n_6273),
.Y(n_8811)
);

NOR2xp33_ASAP7_75t_L g8812 ( 
.A(n_7190),
.B(n_6263),
.Y(n_8812)
);

INVx4_ASAP7_75t_L g8813 ( 
.A(n_7734),
.Y(n_8813)
);

CKINVDCx5p33_ASAP7_75t_R g8814 ( 
.A(n_7804),
.Y(n_8814)
);

NOR2xp33_ASAP7_75t_L g8815 ( 
.A(n_7190),
.B(n_6284),
.Y(n_8815)
);

INVx2_ASAP7_75t_L g8816 ( 
.A(n_7094),
.Y(n_8816)
);

BUFx4_ASAP7_75t_SL g8817 ( 
.A(n_7139),
.Y(n_8817)
);

NAND2xp5_ASAP7_75t_L g8818 ( 
.A(n_7027),
.B(n_6820),
.Y(n_8818)
);

AOI21xp5_ASAP7_75t_L g8819 ( 
.A1(n_7337),
.A2(n_6792),
.B(n_6771),
.Y(n_8819)
);

INVx1_ASAP7_75t_L g8820 ( 
.A(n_7815),
.Y(n_8820)
);

OAI21x1_ASAP7_75t_L g8821 ( 
.A1(n_7601),
.A2(n_7623),
.B(n_7617),
.Y(n_8821)
);

NOR2xp33_ASAP7_75t_L g8822 ( 
.A(n_7206),
.B(n_6289),
.Y(n_8822)
);

INVx1_ASAP7_75t_L g8823 ( 
.A(n_7818),
.Y(n_8823)
);

AND2x4_ASAP7_75t_L g8824 ( 
.A(n_6924),
.B(n_6364),
.Y(n_8824)
);

OAI21xp5_ASAP7_75t_L g8825 ( 
.A1(n_7500),
.A2(n_6306),
.B(n_6302),
.Y(n_8825)
);

NAND2xp5_ASAP7_75t_L g8826 ( 
.A(n_7573),
.B(n_6827),
.Y(n_8826)
);

INVx1_ASAP7_75t_L g8827 ( 
.A(n_7818),
.Y(n_8827)
);

INVx2_ASAP7_75t_L g8828 ( 
.A(n_7094),
.Y(n_8828)
);

INVx3_ASAP7_75t_L g8829 ( 
.A(n_6973),
.Y(n_8829)
);

INVx1_ASAP7_75t_L g8830 ( 
.A(n_7818),
.Y(n_8830)
);

OAI22xp5_ASAP7_75t_SL g8831 ( 
.A1(n_7470),
.A2(n_6480),
.B1(n_6487),
.B2(n_6159),
.Y(n_8831)
);

OA21x2_ASAP7_75t_L g8832 ( 
.A1(n_7627),
.A2(n_6362),
.B(n_6360),
.Y(n_8832)
);

INVx2_ASAP7_75t_SL g8833 ( 
.A(n_7587),
.Y(n_8833)
);

NAND2x1p5_ASAP7_75t_L g8834 ( 
.A(n_7587),
.B(n_6708),
.Y(n_8834)
);

AOI21xp33_ASAP7_75t_L g8835 ( 
.A1(n_7209),
.A2(n_6827),
.B(n_6306),
.Y(n_8835)
);

NOR2x1_ASAP7_75t_R g8836 ( 
.A(n_7135),
.B(n_6159),
.Y(n_8836)
);

AO22x1_ASAP7_75t_L g8837 ( 
.A1(n_7369),
.A2(n_6760),
.B1(n_6109),
.B2(n_6241),
.Y(n_8837)
);

BUFx6f_ASAP7_75t_L g8838 ( 
.A(n_6973),
.Y(n_8838)
);

INVx2_ASAP7_75t_L g8839 ( 
.A(n_7094),
.Y(n_8839)
);

INVx2_ASAP7_75t_L g8840 ( 
.A(n_7094),
.Y(n_8840)
);

INVxp67_ASAP7_75t_SL g8841 ( 
.A(n_7336),
.Y(n_8841)
);

BUFx3_ASAP7_75t_L g8842 ( 
.A(n_7141),
.Y(n_8842)
);

INVx1_ASAP7_75t_L g8843 ( 
.A(n_7825),
.Y(n_8843)
);

AND2x4_ASAP7_75t_L g8844 ( 
.A(n_6924),
.B(n_6416),
.Y(n_8844)
);

OAI21x1_ASAP7_75t_L g8845 ( 
.A1(n_7624),
.A2(n_7645),
.B(n_7635),
.Y(n_8845)
);

OR2x6_ASAP7_75t_L g8846 ( 
.A(n_7427),
.B(n_6792),
.Y(n_8846)
);

AO21x2_ASAP7_75t_L g8847 ( 
.A1(n_7243),
.A2(n_6705),
.B(n_6700),
.Y(n_8847)
);

AOI21xp33_ASAP7_75t_L g8848 ( 
.A1(n_7209),
.A2(n_6321),
.B(n_6302),
.Y(n_8848)
);

NAND2x1_ASAP7_75t_L g8849 ( 
.A(n_7598),
.B(n_5917),
.Y(n_8849)
);

AOI221xp5_ASAP7_75t_L g8850 ( 
.A1(n_7710),
.A2(n_6599),
.B1(n_6329),
.B2(n_6340),
.C(n_6338),
.Y(n_8850)
);

CKINVDCx8_ASAP7_75t_R g8851 ( 
.A(n_7526),
.Y(n_8851)
);

AOI21x1_ASAP7_75t_L g8852 ( 
.A1(n_7116),
.A2(n_6719),
.B(n_6697),
.Y(n_8852)
);

OAI21x1_ASAP7_75t_L g8853 ( 
.A1(n_7515),
.A2(n_6351),
.B(n_6348),
.Y(n_8853)
);

NAND2xp5_ASAP7_75t_L g8854 ( 
.A(n_7573),
.B(n_6867),
.Y(n_8854)
);

AOI21x1_ASAP7_75t_L g8855 ( 
.A1(n_7156),
.A2(n_6741),
.B(n_6420),
.Y(n_8855)
);

OAI21x1_ASAP7_75t_L g8856 ( 
.A1(n_7515),
.A2(n_6367),
.B(n_6351),
.Y(n_8856)
);

OA21x2_ASAP7_75t_L g8857 ( 
.A1(n_7778),
.A2(n_6371),
.B(n_6362),
.Y(n_8857)
);

CKINVDCx20_ASAP7_75t_R g8858 ( 
.A(n_7532),
.Y(n_8858)
);

OAI21x1_ASAP7_75t_L g8859 ( 
.A1(n_7515),
.A2(n_6382),
.B(n_6367),
.Y(n_8859)
);

BUFx2_ASAP7_75t_R g8860 ( 
.A(n_7171),
.Y(n_8860)
);

OAI22xp5_ASAP7_75t_L g8861 ( 
.A1(n_7455),
.A2(n_6880),
.B1(n_6894),
.B2(n_6852),
.Y(n_8861)
);

AND2x4_ASAP7_75t_L g8862 ( 
.A(n_6977),
.B(n_6994),
.Y(n_8862)
);

OAI21x1_ASAP7_75t_L g8863 ( 
.A1(n_7569),
.A2(n_6441),
.B(n_6431),
.Y(n_8863)
);

INVx2_ASAP7_75t_L g8864 ( 
.A(n_7097),
.Y(n_8864)
);

A2O1A1Ixp33_ASAP7_75t_L g8865 ( 
.A1(n_7051),
.A2(n_6321),
.B(n_6359),
.C(n_6340),
.Y(n_8865)
);

OAI21x1_ASAP7_75t_L g8866 ( 
.A1(n_7569),
.A2(n_6441),
.B(n_6431),
.Y(n_8866)
);

HB1xp67_ASAP7_75t_L g8867 ( 
.A(n_7358),
.Y(n_8867)
);

NAND2x1p5_ASAP7_75t_L g8868 ( 
.A(n_7587),
.B(n_6708),
.Y(n_8868)
);

O2A1O1Ixp33_ASAP7_75t_SL g8869 ( 
.A1(n_7172),
.A2(n_6359),
.B(n_6390),
.C(n_6329),
.Y(n_8869)
);

AOI21xp5_ASAP7_75t_L g8870 ( 
.A1(n_7586),
.A2(n_6771),
.B(n_6708),
.Y(n_8870)
);

OAI22xp5_ASAP7_75t_L g8871 ( 
.A1(n_7455),
.A2(n_6390),
.B1(n_6404),
.B2(n_6397),
.Y(n_8871)
);

INVx2_ASAP7_75t_L g8872 ( 
.A(n_7097),
.Y(n_8872)
);

AO31x2_ASAP7_75t_L g8873 ( 
.A1(n_7762),
.A2(n_6133),
.A3(n_6141),
.B(n_6086),
.Y(n_8873)
);

AOI21xp5_ASAP7_75t_L g8874 ( 
.A1(n_7604),
.A2(n_6776),
.B(n_6771),
.Y(n_8874)
);

AOI21x1_ASAP7_75t_L g8875 ( 
.A1(n_7185),
.A2(n_6741),
.B(n_6420),
.Y(n_8875)
);

AOI22xp33_ASAP7_75t_SL g8876 ( 
.A1(n_6910),
.A2(n_6760),
.B1(n_6109),
.B2(n_6241),
.Y(n_8876)
);

INVx1_ASAP7_75t_L g8877 ( 
.A(n_7825),
.Y(n_8877)
);

AO32x2_ASAP7_75t_L g8878 ( 
.A1(n_7662),
.A2(n_5791),
.A3(n_5933),
.B1(n_5876),
.B2(n_5852),
.Y(n_8878)
);

NOR2x1_ASAP7_75t_SL g8879 ( 
.A(n_7526),
.B(n_5917),
.Y(n_8879)
);

AOI221xp5_ASAP7_75t_L g8880 ( 
.A1(n_7710),
.A2(n_6404),
.B1(n_6433),
.B2(n_6425),
.C(n_6397),
.Y(n_8880)
);

INVx5_ASAP7_75t_L g8881 ( 
.A(n_6973),
.Y(n_8881)
);

INVx2_ASAP7_75t_L g8882 ( 
.A(n_7097),
.Y(n_8882)
);

BUFx6f_ASAP7_75t_L g8883 ( 
.A(n_6973),
.Y(n_8883)
);

OAI21xp5_ASAP7_75t_L g8884 ( 
.A1(n_7570),
.A2(n_6433),
.B(n_6425),
.Y(n_8884)
);

INVx1_ASAP7_75t_L g8885 ( 
.A(n_7825),
.Y(n_8885)
);

OAI22xp5_ASAP7_75t_L g8886 ( 
.A1(n_7511),
.A2(n_6450),
.B1(n_6454),
.B2(n_6452),
.Y(n_8886)
);

OAI21x1_ASAP7_75t_L g8887 ( 
.A1(n_7515),
.A2(n_6472),
.B(n_6447),
.Y(n_8887)
);

CKINVDCx6p67_ASAP7_75t_R g8888 ( 
.A(n_7141),
.Y(n_8888)
);

CKINVDCx11_ASAP7_75t_R g8889 ( 
.A(n_7769),
.Y(n_8889)
);

BUFx2_ASAP7_75t_L g8890 ( 
.A(n_7237),
.Y(n_8890)
);

BUFx8_ASAP7_75t_L g8891 ( 
.A(n_7141),
.Y(n_8891)
);

INVx2_ASAP7_75t_SL g8892 ( 
.A(n_7659),
.Y(n_8892)
);

AO21x2_ASAP7_75t_L g8893 ( 
.A1(n_7243),
.A2(n_6712),
.B(n_6710),
.Y(n_8893)
);

AND2x4_ASAP7_75t_L g8894 ( 
.A(n_6977),
.B(n_6435),
.Y(n_8894)
);

AO21x2_ASAP7_75t_L g8895 ( 
.A1(n_7185),
.A2(n_6712),
.B(n_6710),
.Y(n_8895)
);

INVx2_ASAP7_75t_L g8896 ( 
.A(n_7097),
.Y(n_8896)
);

OAI21x1_ASAP7_75t_L g8897 ( 
.A1(n_7515),
.A2(n_6472),
.B(n_6447),
.Y(n_8897)
);

AND2x2_ASAP7_75t_L g8898 ( 
.A(n_7589),
.B(n_6455),
.Y(n_8898)
);

OAI22xp33_ASAP7_75t_L g8899 ( 
.A1(n_7511),
.A2(n_6450),
.B1(n_6454),
.B2(n_6452),
.Y(n_8899)
);

OAI21x1_ASAP7_75t_L g8900 ( 
.A1(n_7515),
.A2(n_7618),
.B(n_7369),
.Y(n_8900)
);

OAI21x1_ASAP7_75t_L g8901 ( 
.A1(n_7515),
.A2(n_6472),
.B(n_6447),
.Y(n_8901)
);

OAI22xp5_ASAP7_75t_L g8902 ( 
.A1(n_7511),
.A2(n_6465),
.B1(n_6488),
.B2(n_6475),
.Y(n_8902)
);

OR2x2_ASAP7_75t_L g8903 ( 
.A(n_7030),
.B(n_6578),
.Y(n_8903)
);

INVx2_ASAP7_75t_SL g8904 ( 
.A(n_7659),
.Y(n_8904)
);

INVx1_ASAP7_75t_L g8905 ( 
.A(n_7835),
.Y(n_8905)
);

NAND2xp33_ASAP7_75t_L g8906 ( 
.A(n_6909),
.B(n_5780),
.Y(n_8906)
);

BUFx3_ASAP7_75t_L g8907 ( 
.A(n_7141),
.Y(n_8907)
);

OAI21x1_ASAP7_75t_L g8908 ( 
.A1(n_7618),
.A2(n_6525),
.B(n_6472),
.Y(n_8908)
);

AO31x2_ASAP7_75t_L g8909 ( 
.A1(n_7103),
.A2(n_6150),
.A3(n_6206),
.B(n_6149),
.Y(n_8909)
);

AND2x4_ASAP7_75t_L g8910 ( 
.A(n_6977),
.B(n_6435),
.Y(n_8910)
);

OAI22xp33_ASAP7_75t_L g8911 ( 
.A1(n_7273),
.A2(n_6488),
.B1(n_6475),
.B2(n_6465),
.Y(n_8911)
);

INVx1_ASAP7_75t_L g8912 ( 
.A(n_7835),
.Y(n_8912)
);

INVx2_ASAP7_75t_SL g8913 ( 
.A(n_7659),
.Y(n_8913)
);

NOR2xp67_ASAP7_75t_L g8914 ( 
.A(n_7659),
.B(n_6271),
.Y(n_8914)
);

OA21x2_ASAP7_75t_L g8915 ( 
.A1(n_7778),
.A2(n_6375),
.B(n_6371),
.Y(n_8915)
);

INVxp67_ASAP7_75t_SL g8916 ( 
.A(n_7358),
.Y(n_8916)
);

BUFx3_ASAP7_75t_L g8917 ( 
.A(n_7244),
.Y(n_8917)
);

INVx1_ASAP7_75t_L g8918 ( 
.A(n_7835),
.Y(n_8918)
);

OA21x2_ASAP7_75t_L g8919 ( 
.A1(n_7807),
.A2(n_6377),
.B(n_6375),
.Y(n_8919)
);

INVx1_ASAP7_75t_L g8920 ( 
.A(n_7842),
.Y(n_8920)
);

INVxp67_ASAP7_75t_L g8921 ( 
.A(n_7608),
.Y(n_8921)
);

AOI22xp33_ASAP7_75t_L g8922 ( 
.A1(n_7250),
.A2(n_6147),
.B1(n_5946),
.B2(n_5947),
.Y(n_8922)
);

NAND2xp5_ASAP7_75t_L g8923 ( 
.A(n_7608),
.B(n_6867),
.Y(n_8923)
);

OAI21x1_ASAP7_75t_L g8924 ( 
.A1(n_7618),
.A2(n_7814),
.B(n_7807),
.Y(n_8924)
);

INVx2_ASAP7_75t_L g8925 ( 
.A(n_7106),
.Y(n_8925)
);

OAI21xp5_ASAP7_75t_L g8926 ( 
.A1(n_7570),
.A2(n_5789),
.B(n_6558),
.Y(n_8926)
);

OAI21x1_ASAP7_75t_L g8927 ( 
.A1(n_7618),
.A2(n_6545),
.B(n_6525),
.Y(n_8927)
);

NOR2xp33_ASAP7_75t_L g8928 ( 
.A(n_7206),
.B(n_6716),
.Y(n_8928)
);

O2A1O1Ixp33_ASAP7_75t_L g8929 ( 
.A1(n_7273),
.A2(n_7064),
.B(n_7713),
.C(n_7555),
.Y(n_8929)
);

NOR2xp33_ASAP7_75t_SL g8930 ( 
.A(n_7694),
.B(n_6147),
.Y(n_8930)
);

AND2x2_ASAP7_75t_L g8931 ( 
.A(n_7589),
.B(n_6521),
.Y(n_8931)
);

INVx2_ASAP7_75t_SL g8932 ( 
.A(n_7659),
.Y(n_8932)
);

AO32x2_ASAP7_75t_L g8933 ( 
.A1(n_7662),
.A2(n_5933),
.A3(n_5996),
.B1(n_5876),
.B2(n_5852),
.Y(n_8933)
);

BUFx6f_ASAP7_75t_L g8934 ( 
.A(n_6981),
.Y(n_8934)
);

AND2x2_ASAP7_75t_L g8935 ( 
.A(n_7589),
.B(n_6521),
.Y(n_8935)
);

INVx1_ASAP7_75t_L g8936 ( 
.A(n_7842),
.Y(n_8936)
);

AOI22xp33_ASAP7_75t_L g8937 ( 
.A1(n_7288),
.A2(n_6147),
.B1(n_5946),
.B2(n_5947),
.Y(n_8937)
);

OAI21xp5_ASAP7_75t_L g8938 ( 
.A1(n_7552),
.A2(n_6559),
.B(n_6558),
.Y(n_8938)
);

BUFx6f_ASAP7_75t_L g8939 ( 
.A(n_6981),
.Y(n_8939)
);

AOI21x1_ASAP7_75t_L g8940 ( 
.A1(n_7369),
.A2(n_6420),
.B(n_6379),
.Y(n_8940)
);

NOR2xp33_ASAP7_75t_L g8941 ( 
.A(n_7865),
.B(n_6716),
.Y(n_8941)
);

OAI222xp33_ASAP7_75t_L g8942 ( 
.A1(n_6970),
.A2(n_5917),
.B1(n_6718),
.B2(n_6728),
.C1(n_6726),
.C2(n_6721),
.Y(n_8942)
);

A2O1A1Ixp33_ASAP7_75t_L g8943 ( 
.A1(n_7449),
.A2(n_6909),
.B(n_7023),
.C(n_7064),
.Y(n_8943)
);

NAND2x1p5_ASAP7_75t_L g8944 ( 
.A(n_7659),
.B(n_6771),
.Y(n_8944)
);

INVx1_ASAP7_75t_L g8945 ( 
.A(n_7842),
.Y(n_8945)
);

OAI21x1_ASAP7_75t_L g8946 ( 
.A1(n_7618),
.A2(n_6382),
.B(n_6367),
.Y(n_8946)
);

O2A1O1Ixp33_ASAP7_75t_L g8947 ( 
.A1(n_7273),
.A2(n_5958),
.B(n_5950),
.C(n_5899),
.Y(n_8947)
);

A2O1A1Ixp33_ASAP7_75t_L g8948 ( 
.A1(n_7449),
.A2(n_6312),
.B(n_6726),
.C(n_6718),
.Y(n_8948)
);

INVx2_ASAP7_75t_L g8949 ( 
.A(n_7106),
.Y(n_8949)
);

O2A1O1Ixp33_ASAP7_75t_L g8950 ( 
.A1(n_7713),
.A2(n_5899),
.B(n_5878),
.C(n_6721),
.Y(n_8950)
);

INVx2_ASAP7_75t_SL g8951 ( 
.A(n_7659),
.Y(n_8951)
);

AOI21x1_ASAP7_75t_L g8952 ( 
.A1(n_7598),
.A2(n_6474),
.B(n_6379),
.Y(n_8952)
);

NOR2xp33_ASAP7_75t_L g8953 ( 
.A(n_7865),
.B(n_7026),
.Y(n_8953)
);

INVx1_ASAP7_75t_L g8954 ( 
.A(n_7844),
.Y(n_8954)
);

INVx2_ASAP7_75t_L g8955 ( 
.A(n_7106),
.Y(n_8955)
);

BUFx3_ASAP7_75t_L g8956 ( 
.A(n_7244),
.Y(n_8956)
);

AO31x2_ASAP7_75t_L g8957 ( 
.A1(n_7103),
.A2(n_6150),
.A3(n_6206),
.B(n_6149),
.Y(n_8957)
);

OAI21x1_ASAP7_75t_L g8958 ( 
.A1(n_7618),
.A2(n_6419),
.B(n_6382),
.Y(n_8958)
);

INVx2_ASAP7_75t_L g8959 ( 
.A(n_7106),
.Y(n_8959)
);

AND2x2_ASAP7_75t_L g8960 ( 
.A(n_7589),
.B(n_6538),
.Y(n_8960)
);

OAI21xp33_ASAP7_75t_SL g8961 ( 
.A1(n_7774),
.A2(n_6276),
.B(n_6271),
.Y(n_8961)
);

O2A1O1Ixp33_ASAP7_75t_SL g8962 ( 
.A1(n_7242),
.A2(n_6584),
.B(n_6587),
.C(n_6578),
.Y(n_8962)
);

OAI21x1_ASAP7_75t_L g8963 ( 
.A1(n_7618),
.A2(n_6430),
.B(n_6419),
.Y(n_8963)
);

OA21x2_ASAP7_75t_L g8964 ( 
.A1(n_7814),
.A2(n_6387),
.B(n_6377),
.Y(n_8964)
);

INVx4_ASAP7_75t_L g8965 ( 
.A(n_7734),
.Y(n_8965)
);

O2A1O1Ixp33_ASAP7_75t_SL g8966 ( 
.A1(n_7242),
.A2(n_6587),
.B(n_6584),
.C(n_6728),
.Y(n_8966)
);

BUFx8_ASAP7_75t_SL g8967 ( 
.A(n_7171),
.Y(n_8967)
);

A2O1A1Ixp33_ASAP7_75t_L g8968 ( 
.A1(n_6909),
.A2(n_6312),
.B(n_6739),
.C(n_6738),
.Y(n_8968)
);

OAI21x1_ASAP7_75t_L g8969 ( 
.A1(n_7620),
.A2(n_6430),
.B(n_6419),
.Y(n_8969)
);

A2O1A1Ixp33_ASAP7_75t_L g8970 ( 
.A1(n_7023),
.A2(n_6312),
.B(n_6746),
.C(n_6739),
.Y(n_8970)
);

NOR2xp67_ASAP7_75t_L g8971 ( 
.A(n_7659),
.B(n_6276),
.Y(n_8971)
);

OAI21x1_ASAP7_75t_L g8972 ( 
.A1(n_7620),
.A2(n_6439),
.B(n_6430),
.Y(n_8972)
);

NAND2xp5_ASAP7_75t_L g8973 ( 
.A(n_7407),
.B(n_5891),
.Y(n_8973)
);

OAI21xp5_ASAP7_75t_L g8974 ( 
.A1(n_7552),
.A2(n_6559),
.B(n_5878),
.Y(n_8974)
);

OAI21x1_ASAP7_75t_L g8975 ( 
.A1(n_7620),
.A2(n_6445),
.B(n_6439),
.Y(n_8975)
);

OAI21x1_ASAP7_75t_L g8976 ( 
.A1(n_7180),
.A2(n_6445),
.B(n_6439),
.Y(n_8976)
);

INVx2_ASAP7_75t_L g8977 ( 
.A(n_7110),
.Y(n_8977)
);

INVx1_ASAP7_75t_SL g8978 ( 
.A(n_7735),
.Y(n_8978)
);

AO21x2_ASAP7_75t_L g8979 ( 
.A1(n_7096),
.A2(n_6743),
.B(n_6727),
.Y(n_8979)
);

INVx3_ASAP7_75t_L g8980 ( 
.A(n_6981),
.Y(n_8980)
);

INVx1_ASAP7_75t_L g8981 ( 
.A(n_7844),
.Y(n_8981)
);

OA21x2_ASAP7_75t_L g8982 ( 
.A1(n_7879),
.A2(n_6400),
.B(n_6387),
.Y(n_8982)
);

OAI21x1_ASAP7_75t_L g8983 ( 
.A1(n_7180),
.A2(n_6456),
.B(n_6445),
.Y(n_8983)
);

NOR2x1_ASAP7_75t_R g8984 ( 
.A(n_7244),
.B(n_6159),
.Y(n_8984)
);

AO21x2_ASAP7_75t_L g8985 ( 
.A1(n_7096),
.A2(n_6743),
.B(n_6727),
.Y(n_8985)
);

NOR2xp33_ASAP7_75t_L g8986 ( 
.A(n_7026),
.B(n_6738),
.Y(n_8986)
);

NAND2xp5_ASAP7_75t_SL g8987 ( 
.A(n_7774),
.B(n_6361),
.Y(n_8987)
);

OAI221xp5_ASAP7_75t_SL g8988 ( 
.A1(n_7682),
.A2(n_6746),
.B1(n_5853),
.B2(n_5808),
.C(n_5830),
.Y(n_8988)
);

NAND2xp5_ASAP7_75t_L g8989 ( 
.A(n_7407),
.B(n_5891),
.Y(n_8989)
);

AOI22xp33_ASAP7_75t_L g8990 ( 
.A1(n_7288),
.A2(n_5946),
.B1(n_5947),
.B2(n_5945),
.Y(n_8990)
);

HB1xp67_ASAP7_75t_L g8991 ( 
.A(n_7359),
.Y(n_8991)
);

INVx2_ASAP7_75t_L g8992 ( 
.A(n_7110),
.Y(n_8992)
);

AOI21xp5_ASAP7_75t_L g8993 ( 
.A1(n_7604),
.A2(n_6776),
.B(n_6771),
.Y(n_8993)
);

NOR2xp67_ASAP7_75t_L g8994 ( 
.A(n_7659),
.B(n_6276),
.Y(n_8994)
);

INVx1_ASAP7_75t_L g8995 ( 
.A(n_7844),
.Y(n_8995)
);

INVx1_ASAP7_75t_L g8996 ( 
.A(n_7845),
.Y(n_8996)
);

A2O1A1Ixp33_ASAP7_75t_L g8997 ( 
.A1(n_7555),
.A2(n_6285),
.B(n_6282),
.C(n_6883),
.Y(n_8997)
);

OAI22xp5_ASAP7_75t_L g8998 ( 
.A1(n_7498),
.A2(n_7103),
.B1(n_7731),
.B2(n_6971),
.Y(n_8998)
);

NAND2xp5_ASAP7_75t_L g8999 ( 
.A(n_7407),
.B(n_5907),
.Y(n_8999)
);

O2A1O1Ixp33_ASAP7_75t_SL g9000 ( 
.A1(n_7477),
.A2(n_5907),
.B(n_6232),
.C(n_6165),
.Y(n_9000)
);

OA21x2_ASAP7_75t_L g9001 ( 
.A1(n_7879),
.A2(n_6415),
.B(n_6400),
.Y(n_9001)
);

CKINVDCx5p33_ASAP7_75t_R g9002 ( 
.A(n_7205),
.Y(n_9002)
);

INVx1_ASAP7_75t_L g9003 ( 
.A(n_7845),
.Y(n_9003)
);

OAI21xp5_ASAP7_75t_L g9004 ( 
.A1(n_7362),
.A2(n_5932),
.B(n_6634),
.Y(n_9004)
);

BUFx3_ASAP7_75t_L g9005 ( 
.A(n_7244),
.Y(n_9005)
);

OAI21x1_ASAP7_75t_L g9006 ( 
.A1(n_7180),
.A2(n_6464),
.B(n_6456),
.Y(n_9006)
);

AO21x2_ASAP7_75t_L g9007 ( 
.A1(n_7096),
.A2(n_6762),
.B(n_6752),
.Y(n_9007)
);

OAI22xp33_ASAP7_75t_L g9008 ( 
.A1(n_6970),
.A2(n_5917),
.B1(n_6715),
.B2(n_6628),
.Y(n_9008)
);

OAI21x1_ASAP7_75t_L g9009 ( 
.A1(n_7180),
.A2(n_6464),
.B(n_6456),
.Y(n_9009)
);

NAND2xp5_ASAP7_75t_L g9010 ( 
.A(n_7756),
.B(n_6165),
.Y(n_9010)
);

OAI21x1_ASAP7_75t_L g9011 ( 
.A1(n_7180),
.A2(n_6473),
.B(n_6464),
.Y(n_9011)
);

AND2x2_ASAP7_75t_L g9012 ( 
.A(n_7589),
.B(n_6538),
.Y(n_9012)
);

OAI22xp33_ASAP7_75t_L g9013 ( 
.A1(n_6970),
.A2(n_6628),
.B1(n_6765),
.B2(n_6715),
.Y(n_9013)
);

AND2x4_ASAP7_75t_L g9014 ( 
.A(n_6977),
.B(n_6994),
.Y(n_9014)
);

AND2x2_ASAP7_75t_L g9015 ( 
.A(n_7589),
.B(n_6560),
.Y(n_9015)
);

OAI21x1_ASAP7_75t_L g9016 ( 
.A1(n_7180),
.A2(n_7630),
.B(n_7282),
.Y(n_9016)
);

CKINVDCx20_ASAP7_75t_R g9017 ( 
.A(n_7532),
.Y(n_9017)
);

OAI21x1_ASAP7_75t_L g9018 ( 
.A1(n_7180),
.A2(n_6499),
.B(n_6473),
.Y(n_9018)
);

HB1xp67_ASAP7_75t_L g9019 ( 
.A(n_7359),
.Y(n_9019)
);

AO21x2_ASAP7_75t_L g9020 ( 
.A1(n_7096),
.A2(n_6762),
.B(n_6752),
.Y(n_9020)
);

OAI21x1_ASAP7_75t_L g9021 ( 
.A1(n_7630),
.A2(n_6499),
.B(n_6473),
.Y(n_9021)
);

INVx3_ASAP7_75t_L g9022 ( 
.A(n_6981),
.Y(n_9022)
);

AOI21xp33_ASAP7_75t_L g9023 ( 
.A1(n_7267),
.A2(n_5853),
.B(n_5802),
.Y(n_9023)
);

NAND2x1p5_ASAP7_75t_L g9024 ( 
.A(n_7659),
.B(n_6771),
.Y(n_9024)
);

AOI21x1_ASAP7_75t_L g9025 ( 
.A1(n_7598),
.A2(n_6474),
.B(n_6379),
.Y(n_9025)
);

AND2x4_ASAP7_75t_L g9026 ( 
.A(n_6977),
.B(n_6384),
.Y(n_9026)
);

OAI21x1_ASAP7_75t_L g9027 ( 
.A1(n_7630),
.A2(n_6512),
.B(n_6499),
.Y(n_9027)
);

INVx1_ASAP7_75t_L g9028 ( 
.A(n_7845),
.Y(n_9028)
);

OAI22xp5_ASAP7_75t_L g9029 ( 
.A1(n_7498),
.A2(n_6753),
.B1(n_6696),
.B2(n_6704),
.Y(n_9029)
);

INVx2_ASAP7_75t_L g9030 ( 
.A(n_7110),
.Y(n_9030)
);

OAI21x1_ASAP7_75t_L g9031 ( 
.A1(n_7630),
.A2(n_6518),
.B(n_6512),
.Y(n_9031)
);

OAI22x1_ASAP7_75t_L g9032 ( 
.A1(n_7745),
.A2(n_6012),
.B1(n_6119),
.B2(n_5996),
.Y(n_9032)
);

OAI21x1_ASAP7_75t_L g9033 ( 
.A1(n_7630),
.A2(n_6518),
.B(n_6512),
.Y(n_9033)
);

OAI21x1_ASAP7_75t_L g9034 ( 
.A1(n_7630),
.A2(n_6523),
.B(n_6518),
.Y(n_9034)
);

HB1xp67_ASAP7_75t_L g9035 ( 
.A(n_7404),
.Y(n_9035)
);

INVx1_ASAP7_75t_L g9036 ( 
.A(n_7849),
.Y(n_9036)
);

OAI21x1_ASAP7_75t_L g9037 ( 
.A1(n_7630),
.A2(n_6541),
.B(n_6523),
.Y(n_9037)
);

AOI21xp5_ASAP7_75t_L g9038 ( 
.A1(n_6966),
.A2(n_6776),
.B(n_6771),
.Y(n_9038)
);

AOI22xp33_ASAP7_75t_L g9039 ( 
.A1(n_7383),
.A2(n_5959),
.B1(n_5945),
.B2(n_5894),
.Y(n_9039)
);

AO21x1_ASAP7_75t_L g9040 ( 
.A1(n_7294),
.A2(n_6639),
.B(n_6634),
.Y(n_9040)
);

OAI21x1_ASAP7_75t_L g9041 ( 
.A1(n_7282),
.A2(n_7294),
.B(n_7654),
.Y(n_9041)
);

NOR2xp33_ASAP7_75t_L g9042 ( 
.A(n_7473),
.B(n_6560),
.Y(n_9042)
);

INVx2_ASAP7_75t_L g9043 ( 
.A(n_7110),
.Y(n_9043)
);

BUFx8_ASAP7_75t_L g9044 ( 
.A(n_7272),
.Y(n_9044)
);

INVx1_ASAP7_75t_L g9045 ( 
.A(n_7849),
.Y(n_9045)
);

INVx1_ASAP7_75t_L g9046 ( 
.A(n_7849),
.Y(n_9046)
);

INVx2_ASAP7_75t_SL g9047 ( 
.A(n_7700),
.Y(n_9047)
);

BUFx10_ASAP7_75t_L g9048 ( 
.A(n_7408),
.Y(n_9048)
);

INVx2_ASAP7_75t_L g9049 ( 
.A(n_7119),
.Y(n_9049)
);

AND2x2_ASAP7_75t_L g9050 ( 
.A(n_7603),
.B(n_6596),
.Y(n_9050)
);

OA21x2_ASAP7_75t_L g9051 ( 
.A1(n_7866),
.A2(n_6417),
.B(n_6415),
.Y(n_9051)
);

NAND2xp5_ASAP7_75t_L g9052 ( 
.A(n_7756),
.B(n_6232),
.Y(n_9052)
);

BUFx10_ASAP7_75t_L g9053 ( 
.A(n_7408),
.Y(n_9053)
);

HB1xp67_ASAP7_75t_L g9054 ( 
.A(n_7404),
.Y(n_9054)
);

NAND2x1_ASAP7_75t_L g9055 ( 
.A(n_7237),
.B(n_6628),
.Y(n_9055)
);

BUFx3_ASAP7_75t_L g9056 ( 
.A(n_7272),
.Y(n_9056)
);

OAI21x1_ASAP7_75t_L g9057 ( 
.A1(n_7282),
.A2(n_7654),
.B(n_7472),
.Y(n_9057)
);

OA21x2_ASAP7_75t_L g9058 ( 
.A1(n_7866),
.A2(n_6423),
.B(n_6417),
.Y(n_9058)
);

OA21x2_ASAP7_75t_L g9059 ( 
.A1(n_7866),
.A2(n_6434),
.B(n_6423),
.Y(n_9059)
);

OA21x2_ASAP7_75t_L g9060 ( 
.A1(n_7639),
.A2(n_6437),
.B(n_6434),
.Y(n_9060)
);

AND2x2_ASAP7_75t_L g9061 ( 
.A(n_7603),
.B(n_6596),
.Y(n_9061)
);

INVx2_ASAP7_75t_L g9062 ( 
.A(n_7119),
.Y(n_9062)
);

AOI21xp5_ASAP7_75t_L g9063 ( 
.A1(n_6966),
.A2(n_6776),
.B(n_6771),
.Y(n_9063)
);

OAI21x1_ASAP7_75t_SL g9064 ( 
.A1(n_7737),
.A2(n_5771),
.B(n_5768),
.Y(n_9064)
);

INVx3_ASAP7_75t_L g9065 ( 
.A(n_6981),
.Y(n_9065)
);

INVx1_ASAP7_75t_L g9066 ( 
.A(n_7853),
.Y(n_9066)
);

AO31x2_ASAP7_75t_L g9067 ( 
.A1(n_7775),
.A2(n_6541),
.A3(n_6547),
.B(n_6523),
.Y(n_9067)
);

INVx2_ASAP7_75t_L g9068 ( 
.A(n_7119),
.Y(n_9068)
);

AOI21x1_ASAP7_75t_L g9069 ( 
.A1(n_7722),
.A2(n_6478),
.B(n_6474),
.Y(n_9069)
);

INVx1_ASAP7_75t_L g9070 ( 
.A(n_7853),
.Y(n_9070)
);

INVx1_ASAP7_75t_SL g9071 ( 
.A(n_7735),
.Y(n_9071)
);

NAND2x1p5_ASAP7_75t_L g9072 ( 
.A(n_7700),
.B(n_6776),
.Y(n_9072)
);

INVx1_ASAP7_75t_L g9073 ( 
.A(n_7853),
.Y(n_9073)
);

INVx4_ASAP7_75t_L g9074 ( 
.A(n_7734),
.Y(n_9074)
);

AND2x4_ASAP7_75t_L g9075 ( 
.A(n_6977),
.B(n_6361),
.Y(n_9075)
);

OAI21x1_ASAP7_75t_L g9076 ( 
.A1(n_7282),
.A2(n_6547),
.B(n_6541),
.Y(n_9076)
);

AO21x2_ASAP7_75t_L g9077 ( 
.A1(n_7096),
.A2(n_6786),
.B(n_6769),
.Y(n_9077)
);

AND2x4_ASAP7_75t_L g9078 ( 
.A(n_6977),
.B(n_6361),
.Y(n_9078)
);

INVx1_ASAP7_75t_L g9079 ( 
.A(n_7858),
.Y(n_9079)
);

AO21x2_ASAP7_75t_L g9080 ( 
.A1(n_7096),
.A2(n_6786),
.B(n_6769),
.Y(n_9080)
);

BUFx6f_ASAP7_75t_L g9081 ( 
.A(n_6981),
.Y(n_9081)
);

INVx6_ASAP7_75t_SL g9082 ( 
.A(n_7109),
.Y(n_9082)
);

INVxp67_ASAP7_75t_L g9083 ( 
.A(n_7616),
.Y(n_9083)
);

INVx2_ASAP7_75t_SL g9084 ( 
.A(n_7700),
.Y(n_9084)
);

INVx1_ASAP7_75t_L g9085 ( 
.A(n_7858),
.Y(n_9085)
);

OA21x2_ASAP7_75t_L g9086 ( 
.A1(n_7639),
.A2(n_6438),
.B(n_6437),
.Y(n_9086)
);

AOI21x1_ASAP7_75t_L g9087 ( 
.A1(n_7722),
.A2(n_6486),
.B(n_6478),
.Y(n_9087)
);

NAND2xp5_ASAP7_75t_L g9088 ( 
.A(n_7787),
.B(n_5846),
.Y(n_9088)
);

AOI22xp33_ASAP7_75t_SL g9089 ( 
.A1(n_6910),
.A2(n_6241),
.B1(n_5886),
.B2(n_6788),
.Y(n_9089)
);

INVx1_ASAP7_75t_L g9090 ( 
.A(n_7858),
.Y(n_9090)
);

INVx1_ASAP7_75t_L g9091 ( 
.A(n_7861),
.Y(n_9091)
);

OA21x2_ASAP7_75t_L g9092 ( 
.A1(n_7750),
.A2(n_6459),
.B(n_6438),
.Y(n_9092)
);

CKINVDCx5p33_ASAP7_75t_R g9093 ( 
.A(n_7205),
.Y(n_9093)
);

NAND2xp5_ASAP7_75t_L g9094 ( 
.A(n_7787),
.B(n_5846),
.Y(n_9094)
);

AND2x2_ASAP7_75t_L g9095 ( 
.A(n_7603),
.B(n_6616),
.Y(n_9095)
);

CKINVDCx20_ASAP7_75t_R g9096 ( 
.A(n_7769),
.Y(n_9096)
);

OAI21x1_ASAP7_75t_L g9097 ( 
.A1(n_7458),
.A2(n_6545),
.B(n_6525),
.Y(n_9097)
);

INVx2_ASAP7_75t_L g9098 ( 
.A(n_7119),
.Y(n_9098)
);

INVx1_ASAP7_75t_SL g9099 ( 
.A(n_7735),
.Y(n_9099)
);

AND2x2_ASAP7_75t_L g9100 ( 
.A(n_7603),
.B(n_6616),
.Y(n_9100)
);

OAI21xp5_ASAP7_75t_L g9101 ( 
.A1(n_7362),
.A2(n_6639),
.B(n_5802),
.Y(n_9101)
);

INVx2_ASAP7_75t_L g9102 ( 
.A(n_7122),
.Y(n_9102)
);

INVx2_ASAP7_75t_L g9103 ( 
.A(n_7122),
.Y(n_9103)
);

INVx1_ASAP7_75t_L g9104 ( 
.A(n_7861),
.Y(n_9104)
);

OAI21xp5_ASAP7_75t_L g9105 ( 
.A1(n_7002),
.A2(n_7737),
.B(n_7151),
.Y(n_9105)
);

INVx1_ASAP7_75t_L g9106 ( 
.A(n_7861),
.Y(n_9106)
);

INVx1_ASAP7_75t_L g9107 ( 
.A(n_7863),
.Y(n_9107)
);

INVx1_ASAP7_75t_L g9108 ( 
.A(n_7863),
.Y(n_9108)
);

HB1xp67_ASAP7_75t_L g9109 ( 
.A(n_7417),
.Y(n_9109)
);

AOI221xp5_ASAP7_75t_L g9110 ( 
.A1(n_7726),
.A2(n_5835),
.B1(n_5847),
.B2(n_5818),
.C(n_5799),
.Y(n_9110)
);

AOI22xp33_ASAP7_75t_L g9111 ( 
.A1(n_7383),
.A2(n_5959),
.B1(n_5945),
.B2(n_5894),
.Y(n_9111)
);

INVx2_ASAP7_75t_L g9112 ( 
.A(n_7122),
.Y(n_9112)
);

NAND2xp5_ASAP7_75t_L g9113 ( 
.A(n_7826),
.B(n_5846),
.Y(n_9113)
);

OA21x2_ASAP7_75t_L g9114 ( 
.A1(n_7750),
.A2(n_6466),
.B(n_6459),
.Y(n_9114)
);

HB1xp67_ASAP7_75t_L g9115 ( 
.A(n_7417),
.Y(n_9115)
);

AOI22xp33_ASAP7_75t_L g9116 ( 
.A1(n_7383),
.A2(n_5959),
.B1(n_5894),
.B2(n_5916),
.Y(n_9116)
);

A2O1A1Ixp33_ASAP7_75t_L g9117 ( 
.A1(n_7325),
.A2(n_6285),
.B(n_6282),
.C(n_6776),
.Y(n_9117)
);

AND2x2_ASAP7_75t_SL g9118 ( 
.A(n_7774),
.B(n_6632),
.Y(n_9118)
);

NOR2xp33_ASAP7_75t_L g9119 ( 
.A(n_7473),
.B(n_6632),
.Y(n_9119)
);

INVx1_ASAP7_75t_L g9120 ( 
.A(n_7863),
.Y(n_9120)
);

OAI22xp33_ASAP7_75t_L g9121 ( 
.A1(n_7057),
.A2(n_6628),
.B1(n_6765),
.B2(n_6715),
.Y(n_9121)
);

NAND3xp33_ASAP7_75t_L g9122 ( 
.A(n_7021),
.B(n_5818),
.C(n_5799),
.Y(n_9122)
);

BUFx2_ASAP7_75t_L g9123 ( 
.A(n_7237),
.Y(n_9123)
);

INVx1_ASAP7_75t_L g9124 ( 
.A(n_7875),
.Y(n_9124)
);

INVx2_ASAP7_75t_L g9125 ( 
.A(n_7122),
.Y(n_9125)
);

CKINVDCx20_ASAP7_75t_R g9126 ( 
.A(n_7387),
.Y(n_9126)
);

INVx2_ASAP7_75t_L g9127 ( 
.A(n_7131),
.Y(n_9127)
);

INVx1_ASAP7_75t_L g9128 ( 
.A(n_7875),
.Y(n_9128)
);

AOI21x1_ASAP7_75t_L g9129 ( 
.A1(n_7722),
.A2(n_6486),
.B(n_6478),
.Y(n_9129)
);

OR2x2_ASAP7_75t_L g9130 ( 
.A(n_7030),
.B(n_5901),
.Y(n_9130)
);

INVx2_ASAP7_75t_SL g9131 ( 
.A(n_7700),
.Y(n_9131)
);

HB1xp67_ASAP7_75t_L g9132 ( 
.A(n_7430),
.Y(n_9132)
);

AND3x2_ASAP7_75t_L g9133 ( 
.A(n_7664),
.B(n_6210),
.C(n_6209),
.Y(n_9133)
);

NAND2x1p5_ASAP7_75t_L g9134 ( 
.A(n_7700),
.B(n_6776),
.Y(n_9134)
);

NAND2xp5_ASAP7_75t_L g9135 ( 
.A(n_7826),
.B(n_6009),
.Y(n_9135)
);

INVx1_ASAP7_75t_L g9136 ( 
.A(n_7875),
.Y(n_9136)
);

INVx1_ASAP7_75t_L g9137 ( 
.A(n_7878),
.Y(n_9137)
);

BUFx2_ASAP7_75t_L g9138 ( 
.A(n_7237),
.Y(n_9138)
);

INVx2_ASAP7_75t_L g9139 ( 
.A(n_7131),
.Y(n_9139)
);

AND2x2_ASAP7_75t_L g9140 ( 
.A(n_7603),
.B(n_7606),
.Y(n_9140)
);

INVx1_ASAP7_75t_L g9141 ( 
.A(n_7878),
.Y(n_9141)
);

OAI21xp5_ASAP7_75t_L g9142 ( 
.A1(n_7002),
.A2(n_5847),
.B(n_5835),
.Y(n_9142)
);

INVx1_ASAP7_75t_L g9143 ( 
.A(n_7878),
.Y(n_9143)
);

AOI211xp5_ASAP7_75t_L g9144 ( 
.A1(n_7228),
.A2(n_5853),
.B(n_5830),
.C(n_5808),
.Y(n_9144)
);

OAI21xp5_ASAP7_75t_L g9145 ( 
.A1(n_7151),
.A2(n_6753),
.B(n_6696),
.Y(n_9145)
);

OAI21x1_ASAP7_75t_SL g9146 ( 
.A1(n_7534),
.A2(n_5771),
.B(n_5768),
.Y(n_9146)
);

INVx1_ASAP7_75t_L g9147 ( 
.A(n_7882),
.Y(n_9147)
);

OAI22xp5_ASAP7_75t_L g9148 ( 
.A1(n_7731),
.A2(n_6702),
.B1(n_6704),
.B2(n_5978),
.Y(n_9148)
);

BUFx3_ASAP7_75t_L g9149 ( 
.A(n_7272),
.Y(n_9149)
);

INVx1_ASAP7_75t_L g9150 ( 
.A(n_7882),
.Y(n_9150)
);

AO31x2_ASAP7_75t_L g9151 ( 
.A1(n_7775),
.A2(n_6661),
.A3(n_6672),
.B(n_6635),
.Y(n_9151)
);

NAND2xp5_ASAP7_75t_L g9152 ( 
.A(n_7826),
.B(n_6009),
.Y(n_9152)
);

INVx2_ASAP7_75t_L g9153 ( 
.A(n_7131),
.Y(n_9153)
);

INVx2_ASAP7_75t_L g9154 ( 
.A(n_7131),
.Y(n_9154)
);

AOI21xp5_ASAP7_75t_L g9155 ( 
.A1(n_6966),
.A2(n_7664),
.B(n_7477),
.Y(n_9155)
);

AO21x1_ASAP7_75t_L g9156 ( 
.A1(n_7786),
.A2(n_6570),
.B(n_6568),
.Y(n_9156)
);

NAND2xp5_ASAP7_75t_L g9157 ( 
.A(n_7836),
.B(n_6018),
.Y(n_9157)
);

BUFx2_ASAP7_75t_L g9158 ( 
.A(n_7240),
.Y(n_9158)
);

INVx2_ASAP7_75t_L g9159 ( 
.A(n_7145),
.Y(n_9159)
);

AOI21x1_ASAP7_75t_L g9160 ( 
.A1(n_7722),
.A2(n_6553),
.B(n_6486),
.Y(n_9160)
);

AND2x2_ASAP7_75t_L g9161 ( 
.A(n_7603),
.B(n_6666),
.Y(n_9161)
);

AND2x2_ASAP7_75t_L g9162 ( 
.A(n_7606),
.B(n_6666),
.Y(n_9162)
);

NAND2xp33_ASAP7_75t_SL g9163 ( 
.A(n_7470),
.B(n_6282),
.Y(n_9163)
);

AOI21xp5_ASAP7_75t_L g9164 ( 
.A1(n_6966),
.A2(n_6802),
.B(n_6776),
.Y(n_9164)
);

AO21x2_ASAP7_75t_L g9165 ( 
.A1(n_7316),
.A2(n_6800),
.B(n_6790),
.Y(n_9165)
);

AND2x2_ASAP7_75t_L g9166 ( 
.A(n_7606),
.B(n_6692),
.Y(n_9166)
);

NAND2xp5_ASAP7_75t_L g9167 ( 
.A(n_7836),
.B(n_6018),
.Y(n_9167)
);

OAI21xp5_ASAP7_75t_SL g9168 ( 
.A1(n_7142),
.A2(n_6833),
.B(n_6720),
.Y(n_9168)
);

CKINVDCx5p33_ASAP7_75t_R g9169 ( 
.A(n_7211),
.Y(n_9169)
);

AOI22xp5_ASAP7_75t_L g9170 ( 
.A1(n_7619),
.A2(n_7593),
.B1(n_7534),
.B2(n_7422),
.Y(n_9170)
);

OA21x2_ASAP7_75t_L g9171 ( 
.A1(n_7750),
.A2(n_7783),
.B(n_7049),
.Y(n_9171)
);

AND2x4_ASAP7_75t_L g9172 ( 
.A(n_6977),
.B(n_6994),
.Y(n_9172)
);

OAI221xp5_ASAP7_75t_L g9173 ( 
.A1(n_7142),
.A2(n_5830),
.B1(n_6628),
.B2(n_6765),
.C(n_6715),
.Y(n_9173)
);

BUFx2_ASAP7_75t_L g9174 ( 
.A(n_7240),
.Y(n_9174)
);

INVx1_ASAP7_75t_L g9175 ( 
.A(n_7882),
.Y(n_9175)
);

INVx1_ASAP7_75t_L g9176 ( 
.A(n_7883),
.Y(n_9176)
);

HB1xp67_ASAP7_75t_L g9177 ( 
.A(n_7430),
.Y(n_9177)
);

AND2x4_ASAP7_75t_L g9178 ( 
.A(n_6977),
.B(n_6621),
.Y(n_9178)
);

OA21x2_ASAP7_75t_L g9179 ( 
.A1(n_7783),
.A2(n_6467),
.B(n_6466),
.Y(n_9179)
);

AND2x4_ASAP7_75t_L g9180 ( 
.A(n_6977),
.B(n_6361),
.Y(n_9180)
);

OAI22xp5_ASAP7_75t_L g9181 ( 
.A1(n_7731),
.A2(n_6702),
.B1(n_6783),
.B2(n_6706),
.Y(n_9181)
);

INVx2_ASAP7_75t_L g9182 ( 
.A(n_7145),
.Y(n_9182)
);

OA21x2_ASAP7_75t_L g9183 ( 
.A1(n_7783),
.A2(n_7049),
.B(n_6984),
.Y(n_9183)
);

INVx2_ASAP7_75t_L g9184 ( 
.A(n_7145),
.Y(n_9184)
);

OAI21xp5_ASAP7_75t_L g9185 ( 
.A1(n_7151),
.A2(n_6164),
.B(n_6045),
.Y(n_9185)
);

BUFx2_ASAP7_75t_L g9186 ( 
.A(n_7240),
.Y(n_9186)
);

OA21x2_ASAP7_75t_L g9187 ( 
.A1(n_6984),
.A2(n_6468),
.B(n_6467),
.Y(n_9187)
);

INVx2_ASAP7_75t_L g9188 ( 
.A(n_7145),
.Y(n_9188)
);

OAI22xp5_ASAP7_75t_L g9189 ( 
.A1(n_6971),
.A2(n_6783),
.B1(n_6706),
.B2(n_6858),
.Y(n_9189)
);

OAI222xp33_ASAP7_75t_L g9190 ( 
.A1(n_6910),
.A2(n_6765),
.B1(n_6775),
.B2(n_6715),
.C1(n_6692),
.C2(n_6788),
.Y(n_9190)
);

OA21x2_ASAP7_75t_L g9191 ( 
.A1(n_6984),
.A2(n_6476),
.B(n_6468),
.Y(n_9191)
);

A2O1A1Ixp33_ASAP7_75t_L g9192 ( 
.A1(n_7325),
.A2(n_6285),
.B(n_6883),
.C(n_6843),
.Y(n_9192)
);

INVx2_ASAP7_75t_L g9193 ( 
.A(n_7147),
.Y(n_9193)
);

INVx2_ASAP7_75t_L g9194 ( 
.A(n_7147),
.Y(n_9194)
);

AOI22x1_ASAP7_75t_L g9195 ( 
.A1(n_7272),
.A2(n_6487),
.B1(n_6633),
.B2(n_6480),
.Y(n_9195)
);

BUFx2_ASAP7_75t_L g9196 ( 
.A(n_7240),
.Y(n_9196)
);

OA21x2_ASAP7_75t_L g9197 ( 
.A1(n_7049),
.A2(n_6479),
.B(n_6476),
.Y(n_9197)
);

AOI21xp5_ASAP7_75t_L g9198 ( 
.A1(n_6966),
.A2(n_6843),
.B(n_6802),
.Y(n_9198)
);

INVx2_ASAP7_75t_SL g9199 ( 
.A(n_7700),
.Y(n_9199)
);

NOR2xp33_ASAP7_75t_L g9200 ( 
.A(n_7496),
.B(n_6905),
.Y(n_9200)
);

INVx1_ASAP7_75t_L g9201 ( 
.A(n_7883),
.Y(n_9201)
);

OA21x2_ASAP7_75t_L g9202 ( 
.A1(n_7069),
.A2(n_6483),
.B(n_6479),
.Y(n_9202)
);

CKINVDCx20_ASAP7_75t_R g9203 ( 
.A(n_7387),
.Y(n_9203)
);

AOI221x1_ASAP7_75t_L g9204 ( 
.A1(n_7025),
.A2(n_5756),
.B1(n_5741),
.B2(n_5731),
.C(n_5238),
.Y(n_9204)
);

INVx3_ASAP7_75t_L g9205 ( 
.A(n_6981),
.Y(n_9205)
);

AND2x2_ASAP7_75t_L g9206 ( 
.A(n_7606),
.B(n_6715),
.Y(n_9206)
);

INVx2_ASAP7_75t_L g9207 ( 
.A(n_7147),
.Y(n_9207)
);

OAI22xp5_ASAP7_75t_L g9208 ( 
.A1(n_7682),
.A2(n_6783),
.B1(n_6858),
.B2(n_6706),
.Y(n_9208)
);

NAND2x1p5_ASAP7_75t_L g9209 ( 
.A(n_7700),
.B(n_7776),
.Y(n_9209)
);

AND2x4_ASAP7_75t_L g9210 ( 
.A(n_6994),
.B(n_6374),
.Y(n_9210)
);

INVx1_ASAP7_75t_L g9211 ( 
.A(n_7883),
.Y(n_9211)
);

NAND2x1p5_ASAP7_75t_L g9212 ( 
.A(n_7700),
.B(n_6802),
.Y(n_9212)
);

OAI21x1_ASAP7_75t_L g9213 ( 
.A1(n_7559),
.A2(n_7563),
.B(n_7856),
.Y(n_9213)
);

AOI22x1_ASAP7_75t_L g9214 ( 
.A1(n_7295),
.A2(n_7211),
.B1(n_7252),
.B2(n_7221),
.Y(n_9214)
);

AND2x4_ASAP7_75t_L g9215 ( 
.A(n_6994),
.B(n_6374),
.Y(n_9215)
);

INVx2_ASAP7_75t_SL g9216 ( 
.A(n_7700),
.Y(n_9216)
);

INVx1_ASAP7_75t_L g9217 ( 
.A(n_7885),
.Y(n_9217)
);

NAND2xp5_ASAP7_75t_L g9218 ( 
.A(n_7836),
.B(n_6045),
.Y(n_9218)
);

INVx1_ASAP7_75t_L g9219 ( 
.A(n_7885),
.Y(n_9219)
);

BUFx2_ASAP7_75t_L g9220 ( 
.A(n_7240),
.Y(n_9220)
);

BUFx8_ASAP7_75t_L g9221 ( 
.A(n_7295),
.Y(n_9221)
);

HB1xp67_ASAP7_75t_L g9222 ( 
.A(n_7481),
.Y(n_9222)
);

NOR2xp67_ASAP7_75t_L g9223 ( 
.A(n_7700),
.B(n_6905),
.Y(n_9223)
);

INVxp67_ASAP7_75t_L g9224 ( 
.A(n_7616),
.Y(n_9224)
);

AND2x4_ASAP7_75t_L g9225 ( 
.A(n_6994),
.B(n_6384),
.Y(n_9225)
);

BUFx6f_ASAP7_75t_L g9226 ( 
.A(n_6981),
.Y(n_9226)
);

INVx1_ASAP7_75t_L g9227 ( 
.A(n_7885),
.Y(n_9227)
);

INVx1_ASAP7_75t_L g9228 ( 
.A(n_7886),
.Y(n_9228)
);

NAND2xp5_ASAP7_75t_L g9229 ( 
.A(n_7843),
.B(n_6164),
.Y(n_9229)
);

OAI21x1_ASAP7_75t_L g9230 ( 
.A1(n_7559),
.A2(n_7563),
.B(n_7797),
.Y(n_9230)
);

CKINVDCx20_ASAP7_75t_R g9231 ( 
.A(n_7470),
.Y(n_9231)
);

HB1xp67_ASAP7_75t_L g9232 ( 
.A(n_7481),
.Y(n_9232)
);

OA21x2_ASAP7_75t_L g9233 ( 
.A1(n_7069),
.A2(n_6484),
.B(n_6483),
.Y(n_9233)
);

INVx6_ASAP7_75t_L g9234 ( 
.A(n_7572),
.Y(n_9234)
);

O2A1O1Ixp5_ASAP7_75t_L g9235 ( 
.A1(n_7534),
.A2(n_6278),
.B(n_6290),
.C(n_6171),
.Y(n_9235)
);

AOI22xp5_ASAP7_75t_L g9236 ( 
.A1(n_7593),
.A2(n_5936),
.B1(n_6788),
.B2(n_6783),
.Y(n_9236)
);

INVx2_ASAP7_75t_L g9237 ( 
.A(n_7147),
.Y(n_9237)
);

OA21x2_ASAP7_75t_L g9238 ( 
.A1(n_7069),
.A2(n_6490),
.B(n_6484),
.Y(n_9238)
);

OAI21x1_ASAP7_75t_L g9239 ( 
.A1(n_7559),
.A2(n_6545),
.B(n_6525),
.Y(n_9239)
);

NOR2xp33_ASAP7_75t_L g9240 ( 
.A(n_7496),
.B(n_6905),
.Y(n_9240)
);

OR2x6_ASAP7_75t_L g9241 ( 
.A(n_7427),
.B(n_5806),
.Y(n_9241)
);

INVx1_ASAP7_75t_L g9242 ( 
.A(n_7886),
.Y(n_9242)
);

A2O1A1Ixp33_ASAP7_75t_L g9243 ( 
.A1(n_7745),
.A2(n_6883),
.B(n_6843),
.C(n_6862),
.Y(n_9243)
);

NOR2xp33_ASAP7_75t_L g9244 ( 
.A(n_7516),
.B(n_6905),
.Y(n_9244)
);

BUFx6f_ASAP7_75t_L g9245 ( 
.A(n_6981),
.Y(n_9245)
);

OAI21x1_ASAP7_75t_L g9246 ( 
.A1(n_7563),
.A2(n_6545),
.B(n_6525),
.Y(n_9246)
);

INVx1_ASAP7_75t_SL g9247 ( 
.A(n_7810),
.Y(n_9247)
);

AOI22xp33_ASAP7_75t_L g9248 ( 
.A1(n_7021),
.A2(n_5916),
.B1(n_5936),
.B2(n_5897),
.Y(n_9248)
);

HB1xp67_ASAP7_75t_L g9249 ( 
.A(n_7501),
.Y(n_9249)
);

NAND2xp5_ASAP7_75t_L g9250 ( 
.A(n_7843),
.B(n_5916),
.Y(n_9250)
);

NOR2xp33_ASAP7_75t_L g9251 ( 
.A(n_7516),
.B(n_6364),
.Y(n_9251)
);

INVx1_ASAP7_75t_L g9252 ( 
.A(n_7886),
.Y(n_9252)
);

OAI21xp5_ASAP7_75t_L g9253 ( 
.A1(n_7138),
.A2(n_7860),
.B(n_7834),
.Y(n_9253)
);

AOI21x1_ASAP7_75t_L g9254 ( 
.A1(n_7722),
.A2(n_6581),
.B(n_6553),
.Y(n_9254)
);

AOI221xp5_ASAP7_75t_L g9255 ( 
.A1(n_7726),
.A2(n_5238),
.B1(n_5253),
.B2(n_5232),
.C(n_5230),
.Y(n_9255)
);

OAI22xp33_ASAP7_75t_L g9256 ( 
.A1(n_7057),
.A2(n_6765),
.B1(n_6775),
.B2(n_6706),
.Y(n_9256)
);

INVx1_ASAP7_75t_L g9257 ( 
.A(n_6908),
.Y(n_9257)
);

INVx1_ASAP7_75t_L g9258 ( 
.A(n_6908),
.Y(n_9258)
);

INVx1_ASAP7_75t_L g9259 ( 
.A(n_6908),
.Y(n_9259)
);

NOR2xp33_ASAP7_75t_L g9260 ( 
.A(n_7553),
.B(n_6364),
.Y(n_9260)
);

BUFx6f_ASAP7_75t_L g9261 ( 
.A(n_6981),
.Y(n_9261)
);

NAND2xp5_ASAP7_75t_L g9262 ( 
.A(n_7843),
.B(n_6847),
.Y(n_9262)
);

NOR2xp33_ASAP7_75t_L g9263 ( 
.A(n_7553),
.B(n_6384),
.Y(n_9263)
);

O2A1O1Ixp33_ASAP7_75t_L g9264 ( 
.A1(n_7726),
.A2(n_5122),
.B(n_5166),
.C(n_5106),
.Y(n_9264)
);

INVx1_ASAP7_75t_L g9265 ( 
.A(n_6923),
.Y(n_9265)
);

CKINVDCx5p33_ASAP7_75t_R g9266 ( 
.A(n_7525),
.Y(n_9266)
);

INVx2_ASAP7_75t_L g9267 ( 
.A(n_7148),
.Y(n_9267)
);

HB1xp67_ASAP7_75t_L g9268 ( 
.A(n_7501),
.Y(n_9268)
);

HB1xp67_ASAP7_75t_L g9269 ( 
.A(n_7703),
.Y(n_9269)
);

BUFx3_ASAP7_75t_L g9270 ( 
.A(n_7295),
.Y(n_9270)
);

INVx1_ASAP7_75t_L g9271 ( 
.A(n_6923),
.Y(n_9271)
);

OR2x6_ASAP7_75t_L g9272 ( 
.A(n_7504),
.B(n_5806),
.Y(n_9272)
);

HB1xp67_ASAP7_75t_L g9273 ( 
.A(n_7703),
.Y(n_9273)
);

OA21x2_ASAP7_75t_L g9274 ( 
.A1(n_7074),
.A2(n_6494),
.B(n_6490),
.Y(n_9274)
);

AOI22x1_ASAP7_75t_L g9275 ( 
.A1(n_7295),
.A2(n_6487),
.B1(n_6633),
.B2(n_6480),
.Y(n_9275)
);

AND2x4_ASAP7_75t_L g9276 ( 
.A(n_6994),
.B(n_6416),
.Y(n_9276)
);

NAND2xp5_ASAP7_75t_SL g9277 ( 
.A(n_7774),
.B(n_6384),
.Y(n_9277)
);

INVx8_ASAP7_75t_L g9278 ( 
.A(n_7877),
.Y(n_9278)
);

NAND2xp5_ASAP7_75t_L g9279 ( 
.A(n_7675),
.B(n_6847),
.Y(n_9279)
);

INVx1_ASAP7_75t_L g9280 ( 
.A(n_6923),
.Y(n_9280)
);

AOI22xp33_ASAP7_75t_L g9281 ( 
.A1(n_6985),
.A2(n_5936),
.B1(n_5960),
.B2(n_5897),
.Y(n_9281)
);

NAND2x1p5_ASAP7_75t_L g9282 ( 
.A(n_7776),
.B(n_6802),
.Y(n_9282)
);

AOI22xp33_ASAP7_75t_L g9283 ( 
.A1(n_6985),
.A2(n_5960),
.B1(n_5897),
.B2(n_6633),
.Y(n_9283)
);

INVx1_ASAP7_75t_L g9284 ( 
.A(n_6942),
.Y(n_9284)
);

OAI22xp33_ASAP7_75t_L g9285 ( 
.A1(n_7057),
.A2(n_6765),
.B1(n_6775),
.B2(n_6706),
.Y(n_9285)
);

AOI22xp33_ASAP7_75t_SL g9286 ( 
.A1(n_7774),
.A2(n_5886),
.B1(n_5784),
.B2(n_5814),
.Y(n_9286)
);

NAND2x1p5_ASAP7_75t_L g9287 ( 
.A(n_7776),
.B(n_6802),
.Y(n_9287)
);

INVx1_ASAP7_75t_SL g9288 ( 
.A(n_7810),
.Y(n_9288)
);

INVx1_ASAP7_75t_SL g9289 ( 
.A(n_7810),
.Y(n_9289)
);

AND2x4_ASAP7_75t_L g9290 ( 
.A(n_6994),
.B(n_6421),
.Y(n_9290)
);

INVx1_ASAP7_75t_L g9291 ( 
.A(n_6942),
.Y(n_9291)
);

AND2x4_ASAP7_75t_L g9292 ( 
.A(n_6994),
.B(n_6421),
.Y(n_9292)
);

INVx1_ASAP7_75t_L g9293 ( 
.A(n_6942),
.Y(n_9293)
);

AOI22xp33_ASAP7_75t_L g9294 ( 
.A1(n_6993),
.A2(n_5960),
.B1(n_5897),
.B2(n_6677),
.Y(n_9294)
);

INVx1_ASAP7_75t_L g9295 ( 
.A(n_6944),
.Y(n_9295)
);

OR2x2_ASAP7_75t_L g9296 ( 
.A(n_7036),
.B(n_5901),
.Y(n_9296)
);

AOI21x1_ASAP7_75t_L g9297 ( 
.A1(n_7722),
.A2(n_6581),
.B(n_6553),
.Y(n_9297)
);

CKINVDCx20_ASAP7_75t_R g9298 ( 
.A(n_7525),
.Y(n_9298)
);

INVx2_ASAP7_75t_L g9299 ( 
.A(n_7148),
.Y(n_9299)
);

AOI21xp5_ASAP7_75t_L g9300 ( 
.A1(n_6966),
.A2(n_6843),
.B(n_6802),
.Y(n_9300)
);

INVx2_ASAP7_75t_L g9301 ( 
.A(n_7148),
.Y(n_9301)
);

BUFx4_ASAP7_75t_SL g9302 ( 
.A(n_7395),
.Y(n_9302)
);

INVx1_ASAP7_75t_L g9303 ( 
.A(n_6944),
.Y(n_9303)
);

INVx2_ASAP7_75t_SL g9304 ( 
.A(n_7776),
.Y(n_9304)
);

INVx1_ASAP7_75t_L g9305 ( 
.A(n_6944),
.Y(n_9305)
);

INVx1_ASAP7_75t_L g9306 ( 
.A(n_6954),
.Y(n_9306)
);

INVx1_ASAP7_75t_L g9307 ( 
.A(n_6954),
.Y(n_9307)
);

AOI21xp5_ASAP7_75t_L g9308 ( 
.A1(n_6966),
.A2(n_6843),
.B(n_6802),
.Y(n_9308)
);

NOR2xp33_ASAP7_75t_L g9309 ( 
.A(n_6932),
.B(n_6967),
.Y(n_9309)
);

NOR2xp33_ASAP7_75t_L g9310 ( 
.A(n_6932),
.B(n_6384),
.Y(n_9310)
);

CKINVDCx6p67_ASAP7_75t_R g9311 ( 
.A(n_7877),
.Y(n_9311)
);

CKINVDCx20_ASAP7_75t_R g9312 ( 
.A(n_7048),
.Y(n_9312)
);

INVx1_ASAP7_75t_L g9313 ( 
.A(n_9257),
.Y(n_9313)
);

AOI22xp33_ASAP7_75t_L g9314 ( 
.A1(n_8080),
.A2(n_7969),
.B1(n_8159),
.B2(n_8143),
.Y(n_9314)
);

AOI22xp33_ASAP7_75t_L g9315 ( 
.A1(n_8080),
.A2(n_6990),
.B1(n_7385),
.B2(n_7805),
.Y(n_9315)
);

OAI21xp5_ASAP7_75t_SL g9316 ( 
.A1(n_7939),
.A2(n_7236),
.B(n_7138),
.Y(n_9316)
);

BUFx6f_ASAP7_75t_L g9317 ( 
.A(n_8074),
.Y(n_9317)
);

OAI22xp5_ASAP7_75t_L g9318 ( 
.A1(n_7939),
.A2(n_7520),
.B1(n_7605),
.B2(n_7561),
.Y(n_9318)
);

INVx1_ASAP7_75t_L g9319 ( 
.A(n_9257),
.Y(n_9319)
);

BUFx6f_ASAP7_75t_L g9320 ( 
.A(n_8074),
.Y(n_9320)
);

CKINVDCx5p33_ASAP7_75t_R g9321 ( 
.A(n_8889),
.Y(n_9321)
);

INVx1_ASAP7_75t_L g9322 ( 
.A(n_9257),
.Y(n_9322)
);

INVx2_ASAP7_75t_L g9323 ( 
.A(n_9187),
.Y(n_9323)
);

OR2x6_ASAP7_75t_L g9324 ( 
.A(n_8021),
.B(n_7526),
.Y(n_9324)
);

BUFx2_ASAP7_75t_L g9325 ( 
.A(n_9082),
.Y(n_9325)
);

INVx2_ASAP7_75t_L g9326 ( 
.A(n_9187),
.Y(n_9326)
);

INVx1_ASAP7_75t_SL g9327 ( 
.A(n_8889),
.Y(n_9327)
);

INVx2_ASAP7_75t_SL g9328 ( 
.A(n_8437),
.Y(n_9328)
);

INVx1_ASAP7_75t_L g9329 ( 
.A(n_9258),
.Y(n_9329)
);

OAI22xp33_ASAP7_75t_L g9330 ( 
.A1(n_8226),
.A2(n_7520),
.B1(n_7816),
.B2(n_7605),
.Y(n_9330)
);

BUFx6f_ASAP7_75t_L g9331 ( 
.A(n_8548),
.Y(n_9331)
);

INVx2_ASAP7_75t_L g9332 ( 
.A(n_9187),
.Y(n_9332)
);

OAI22xp5_ASAP7_75t_L g9333 ( 
.A1(n_7927),
.A2(n_7520),
.B1(n_7605),
.B2(n_7561),
.Y(n_9333)
);

NAND2xp5_ASAP7_75t_L g9334 ( 
.A(n_7986),
.B(n_7326),
.Y(n_9334)
);

AOI22xp33_ASAP7_75t_L g9335 ( 
.A1(n_8080),
.A2(n_7969),
.B1(n_8159),
.B2(n_8143),
.Y(n_9335)
);

OR2x6_ASAP7_75t_L g9336 ( 
.A(n_8021),
.B(n_7574),
.Y(n_9336)
);

INVx1_ASAP7_75t_L g9337 ( 
.A(n_9258),
.Y(n_9337)
);

INVx2_ASAP7_75t_L g9338 ( 
.A(n_9187),
.Y(n_9338)
);

BUFx3_ASAP7_75t_L g9339 ( 
.A(n_8102),
.Y(n_9339)
);

AOI22xp33_ASAP7_75t_L g9340 ( 
.A1(n_8080),
.A2(n_7929),
.B1(n_8085),
.B2(n_7952),
.Y(n_9340)
);

INVx5_ASAP7_75t_L g9341 ( 
.A(n_7988),
.Y(n_9341)
);

INVx1_ASAP7_75t_L g9342 ( 
.A(n_9258),
.Y(n_9342)
);

INVx4_ASAP7_75t_L g9343 ( 
.A(n_7988),
.Y(n_9343)
);

INVx1_ASAP7_75t_L g9344 ( 
.A(n_9259),
.Y(n_9344)
);

AND2x2_ASAP7_75t_L g9345 ( 
.A(n_8006),
.B(n_7840),
.Y(n_9345)
);

AOI22xp33_ASAP7_75t_SL g9346 ( 
.A1(n_8085),
.A2(n_7385),
.B1(n_6990),
.B2(n_7805),
.Y(n_9346)
);

AND2x2_ASAP7_75t_L g9347 ( 
.A(n_8006),
.B(n_7840),
.Y(n_9347)
);

INVx2_ASAP7_75t_L g9348 ( 
.A(n_9187),
.Y(n_9348)
);

INVx1_ASAP7_75t_SL g9349 ( 
.A(n_8860),
.Y(n_9349)
);

INVx3_ASAP7_75t_L g9350 ( 
.A(n_7923),
.Y(n_9350)
);

AO21x2_ASAP7_75t_L g9351 ( 
.A1(n_9156),
.A2(n_7285),
.B(n_7263),
.Y(n_9351)
);

INVx2_ASAP7_75t_L g9352 ( 
.A(n_9187),
.Y(n_9352)
);

BUFx2_ASAP7_75t_L g9353 ( 
.A(n_9082),
.Y(n_9353)
);

INVx3_ASAP7_75t_L g9354 ( 
.A(n_7923),
.Y(n_9354)
);

CKINVDCx6p67_ASAP7_75t_R g9355 ( 
.A(n_8354),
.Y(n_9355)
);

INVx1_ASAP7_75t_SL g9356 ( 
.A(n_8860),
.Y(n_9356)
);

BUFx6f_ASAP7_75t_L g9357 ( 
.A(n_8548),
.Y(n_9357)
);

AOI22xp5_ASAP7_75t_L g9358 ( 
.A1(n_7927),
.A2(n_8226),
.B1(n_7919),
.B2(n_8220),
.Y(n_9358)
);

INVx1_ASAP7_75t_L g9359 ( 
.A(n_9259),
.Y(n_9359)
);

BUFx2_ASAP7_75t_L g9360 ( 
.A(n_9082),
.Y(n_9360)
);

OR2x2_ASAP7_75t_L g9361 ( 
.A(n_8418),
.B(n_7671),
.Y(n_9361)
);

INVx1_ASAP7_75t_L g9362 ( 
.A(n_9259),
.Y(n_9362)
);

INVx2_ASAP7_75t_L g9363 ( 
.A(n_9191),
.Y(n_9363)
);

INVx3_ASAP7_75t_L g9364 ( 
.A(n_7923),
.Y(n_9364)
);

INVx1_ASAP7_75t_L g9365 ( 
.A(n_9265),
.Y(n_9365)
);

INVx1_ASAP7_75t_L g9366 ( 
.A(n_9265),
.Y(n_9366)
);

INVx1_ASAP7_75t_L g9367 ( 
.A(n_9265),
.Y(n_9367)
);

NAND2xp5_ASAP7_75t_L g9368 ( 
.A(n_7986),
.B(n_7326),
.Y(n_9368)
);

OA21x2_ASAP7_75t_L g9369 ( 
.A1(n_8900),
.A2(n_7081),
.B(n_7074),
.Y(n_9369)
);

OAI21x1_ASAP7_75t_L g9370 ( 
.A1(n_9038),
.A2(n_7819),
.B(n_7813),
.Y(n_9370)
);

AOI22xp33_ASAP7_75t_SL g9371 ( 
.A1(n_8080),
.A2(n_7385),
.B1(n_6990),
.B2(n_7805),
.Y(n_9371)
);

INVx1_ASAP7_75t_L g9372 ( 
.A(n_9271),
.Y(n_9372)
);

CKINVDCx20_ASAP7_75t_R g9373 ( 
.A(n_9126),
.Y(n_9373)
);

AND2x2_ASAP7_75t_L g9374 ( 
.A(n_8006),
.B(n_7840),
.Y(n_9374)
);

OAI22xp33_ASAP7_75t_SL g9375 ( 
.A1(n_7957),
.A2(n_6993),
.B1(n_7429),
.B2(n_7428),
.Y(n_9375)
);

INVx2_ASAP7_75t_L g9376 ( 
.A(n_9191),
.Y(n_9376)
);

NOR2x1_ASAP7_75t_SL g9377 ( 
.A(n_8987),
.B(n_7574),
.Y(n_9377)
);

OAI21x1_ASAP7_75t_L g9378 ( 
.A1(n_9038),
.A2(n_9164),
.B(n_9063),
.Y(n_9378)
);

AND2x2_ASAP7_75t_L g9379 ( 
.A(n_7938),
.B(n_7840),
.Y(n_9379)
);

INVx1_ASAP7_75t_L g9380 ( 
.A(n_9271),
.Y(n_9380)
);

INVx2_ASAP7_75t_L g9381 ( 
.A(n_9191),
.Y(n_9381)
);

NOR2xp33_ASAP7_75t_L g9382 ( 
.A(n_8366),
.B(n_7428),
.Y(n_9382)
);

NAND2xp5_ASAP7_75t_L g9383 ( 
.A(n_7975),
.B(n_8034),
.Y(n_9383)
);

BUFx3_ASAP7_75t_L g9384 ( 
.A(n_8102),
.Y(n_9384)
);

INVx1_ASAP7_75t_L g9385 ( 
.A(n_9271),
.Y(n_9385)
);

INVx3_ASAP7_75t_L g9386 ( 
.A(n_7923),
.Y(n_9386)
);

AND2x2_ASAP7_75t_L g9387 ( 
.A(n_7938),
.B(n_7840),
.Y(n_9387)
);

INVx1_ASAP7_75t_L g9388 ( 
.A(n_9280),
.Y(n_9388)
);

INVx1_ASAP7_75t_L g9389 ( 
.A(n_9280),
.Y(n_9389)
);

INVx6_ASAP7_75t_L g9390 ( 
.A(n_8102),
.Y(n_9390)
);

INVx1_ASAP7_75t_L g9391 ( 
.A(n_9280),
.Y(n_9391)
);

AO21x2_ASAP7_75t_L g9392 ( 
.A1(n_9156),
.A2(n_7285),
.B(n_7263),
.Y(n_9392)
);

INVx2_ASAP7_75t_L g9393 ( 
.A(n_9191),
.Y(n_9393)
);

INVx2_ASAP7_75t_L g9394 ( 
.A(n_9191),
.Y(n_9394)
);

BUFx6f_ASAP7_75t_L g9395 ( 
.A(n_7988),
.Y(n_9395)
);

INVx2_ASAP7_75t_L g9396 ( 
.A(n_9191),
.Y(n_9396)
);

AO21x1_ASAP7_75t_L g9397 ( 
.A1(n_7952),
.A2(n_7155),
.B(n_7025),
.Y(n_9397)
);

INVx1_ASAP7_75t_L g9398 ( 
.A(n_9284),
.Y(n_9398)
);

NAND2xp5_ASAP7_75t_L g9399 ( 
.A(n_7975),
.B(n_7371),
.Y(n_9399)
);

AND2x2_ASAP7_75t_L g9400 ( 
.A(n_7938),
.B(n_7840),
.Y(n_9400)
);

INVx2_ASAP7_75t_L g9401 ( 
.A(n_9197),
.Y(n_9401)
);

BUFx4f_ASAP7_75t_SL g9402 ( 
.A(n_9298),
.Y(n_9402)
);

INVx1_ASAP7_75t_L g9403 ( 
.A(n_9284),
.Y(n_9403)
);

CKINVDCx16_ASAP7_75t_R g9404 ( 
.A(n_7988),
.Y(n_9404)
);

INVx1_ASAP7_75t_L g9405 ( 
.A(n_9284),
.Y(n_9405)
);

AND2x2_ASAP7_75t_L g9406 ( 
.A(n_8041),
.B(n_7133),
.Y(n_9406)
);

INVx1_ASAP7_75t_L g9407 ( 
.A(n_9291),
.Y(n_9407)
);

INVx1_ASAP7_75t_L g9408 ( 
.A(n_9291),
.Y(n_9408)
);

INVx2_ASAP7_75t_L g9409 ( 
.A(n_9197),
.Y(n_9409)
);

INVx2_ASAP7_75t_L g9410 ( 
.A(n_9197),
.Y(n_9410)
);

OR2x6_ASAP7_75t_L g9411 ( 
.A(n_8175),
.B(n_7574),
.Y(n_9411)
);

NAND2xp5_ASAP7_75t_L g9412 ( 
.A(n_8034),
.B(n_7371),
.Y(n_9412)
);

INVx1_ASAP7_75t_L g9413 ( 
.A(n_9291),
.Y(n_9413)
);

AND2x4_ASAP7_75t_L g9414 ( 
.A(n_7934),
.B(n_7998),
.Y(n_9414)
);

INVx2_ASAP7_75t_L g9415 ( 
.A(n_9197),
.Y(n_9415)
);

BUFx6f_ASAP7_75t_L g9416 ( 
.A(n_8169),
.Y(n_9416)
);

BUFx4f_ASAP7_75t_SL g9417 ( 
.A(n_9298),
.Y(n_9417)
);

INVx2_ASAP7_75t_SL g9418 ( 
.A(n_8437),
.Y(n_9418)
);

BUFx12f_ASAP7_75t_L g9419 ( 
.A(n_8169),
.Y(n_9419)
);

CKINVDCx5p33_ASAP7_75t_R g9420 ( 
.A(n_8967),
.Y(n_9420)
);

OAI21xp5_ASAP7_75t_L g9421 ( 
.A1(n_8054),
.A2(n_7236),
.B(n_7138),
.Y(n_9421)
);

INVx1_ASAP7_75t_SL g9422 ( 
.A(n_7997),
.Y(n_9422)
);

INVx1_ASAP7_75t_L g9423 ( 
.A(n_9293),
.Y(n_9423)
);

AOI22xp33_ASAP7_75t_L g9424 ( 
.A1(n_8080),
.A2(n_6990),
.B1(n_7385),
.B2(n_7805),
.Y(n_9424)
);

INVx2_ASAP7_75t_L g9425 ( 
.A(n_9197),
.Y(n_9425)
);

INVx2_ASAP7_75t_SL g9426 ( 
.A(n_8437),
.Y(n_9426)
);

AOI22xp33_ASAP7_75t_L g9427 ( 
.A1(n_7929),
.A2(n_6990),
.B1(n_7385),
.B2(n_7805),
.Y(n_9427)
);

AOI21x1_ASAP7_75t_L g9428 ( 
.A1(n_8337),
.A2(n_7154),
.B(n_7148),
.Y(n_9428)
);

BUFx3_ASAP7_75t_L g9429 ( 
.A(n_8102),
.Y(n_9429)
);

INVx1_ASAP7_75t_L g9430 ( 
.A(n_9293),
.Y(n_9430)
);

INVx1_ASAP7_75t_L g9431 ( 
.A(n_9293),
.Y(n_9431)
);

CKINVDCx11_ASAP7_75t_R g9432 ( 
.A(n_8075),
.Y(n_9432)
);

INVx1_ASAP7_75t_L g9433 ( 
.A(n_9295),
.Y(n_9433)
);

BUFx6f_ASAP7_75t_L g9434 ( 
.A(n_8169),
.Y(n_9434)
);

BUFx2_ASAP7_75t_L g9435 ( 
.A(n_9082),
.Y(n_9435)
);

AND2x4_ASAP7_75t_L g9436 ( 
.A(n_7934),
.B(n_6926),
.Y(n_9436)
);

CKINVDCx20_ASAP7_75t_R g9437 ( 
.A(n_9126),
.Y(n_9437)
);

INVx1_ASAP7_75t_L g9438 ( 
.A(n_9295),
.Y(n_9438)
);

NAND2x1p5_ASAP7_75t_L g9439 ( 
.A(n_7974),
.B(n_7776),
.Y(n_9439)
);

INVx1_ASAP7_75t_L g9440 ( 
.A(n_9295),
.Y(n_9440)
);

INVx1_ASAP7_75t_L g9441 ( 
.A(n_9303),
.Y(n_9441)
);

INVx5_ASAP7_75t_SL g9442 ( 
.A(n_8097),
.Y(n_9442)
);

INVx2_ASAP7_75t_L g9443 ( 
.A(n_9197),
.Y(n_9443)
);

INVx1_ASAP7_75t_L g9444 ( 
.A(n_9303),
.Y(n_9444)
);

INVx2_ASAP7_75t_L g9445 ( 
.A(n_9202),
.Y(n_9445)
);

INVx1_ASAP7_75t_L g9446 ( 
.A(n_9303),
.Y(n_9446)
);

AND2x4_ASAP7_75t_L g9447 ( 
.A(n_7934),
.B(n_7998),
.Y(n_9447)
);

INVx1_ASAP7_75t_L g9448 ( 
.A(n_9305),
.Y(n_9448)
);

INVx1_ASAP7_75t_L g9449 ( 
.A(n_9305),
.Y(n_9449)
);

AND2x2_ASAP7_75t_L g9450 ( 
.A(n_8041),
.B(n_7133),
.Y(n_9450)
);

HB1xp67_ASAP7_75t_L g9451 ( 
.A(n_8418),
.Y(n_9451)
);

INVx1_ASAP7_75t_L g9452 ( 
.A(n_9305),
.Y(n_9452)
);

INVx1_ASAP7_75t_L g9453 ( 
.A(n_9306),
.Y(n_9453)
);

INVx1_ASAP7_75t_L g9454 ( 
.A(n_9306),
.Y(n_9454)
);

AOI22xp33_ASAP7_75t_L g9455 ( 
.A1(n_8417),
.A2(n_7593),
.B1(n_7619),
.B2(n_7621),
.Y(n_9455)
);

INVx1_ASAP7_75t_L g9456 ( 
.A(n_9306),
.Y(n_9456)
);

BUFx2_ASAP7_75t_L g9457 ( 
.A(n_9082),
.Y(n_9457)
);

AOI22xp33_ASAP7_75t_L g9458 ( 
.A1(n_8417),
.A2(n_7619),
.B1(n_7621),
.B2(n_7422),
.Y(n_9458)
);

INVx1_ASAP7_75t_L g9459 ( 
.A(n_9307),
.Y(n_9459)
);

INVx2_ASAP7_75t_L g9460 ( 
.A(n_9202),
.Y(n_9460)
);

OAI21x1_ASAP7_75t_L g9461 ( 
.A1(n_9063),
.A2(n_7819),
.B(n_7813),
.Y(n_9461)
);

HB1xp67_ASAP7_75t_L g9462 ( 
.A(n_8418),
.Y(n_9462)
);

OAI22xp5_ASAP7_75t_L g9463 ( 
.A1(n_8054),
.A2(n_7561),
.B1(n_7533),
.B2(n_7391),
.Y(n_9463)
);

BUFx2_ASAP7_75t_R g9464 ( 
.A(n_8967),
.Y(n_9464)
);

OAI22xp5_ASAP7_75t_L g9465 ( 
.A1(n_7919),
.A2(n_7533),
.B1(n_7391),
.B2(n_7389),
.Y(n_9465)
);

INVx1_ASAP7_75t_L g9466 ( 
.A(n_9307),
.Y(n_9466)
);

INVx2_ASAP7_75t_L g9467 ( 
.A(n_9202),
.Y(n_9467)
);

OAI21xp5_ASAP7_75t_SL g9468 ( 
.A1(n_9170),
.A2(n_7075),
.B(n_7745),
.Y(n_9468)
);

NAND2xp5_ASAP7_75t_L g9469 ( 
.A(n_8038),
.B(n_7393),
.Y(n_9469)
);

INVx2_ASAP7_75t_L g9470 ( 
.A(n_9202),
.Y(n_9470)
);

OAI22xp5_ASAP7_75t_L g9471 ( 
.A1(n_7931),
.A2(n_7533),
.B1(n_7389),
.B2(n_7545),
.Y(n_9471)
);

BUFx6f_ASAP7_75t_L g9472 ( 
.A(n_8169),
.Y(n_9472)
);

OA21x2_ASAP7_75t_L g9473 ( 
.A1(n_8900),
.A2(n_7081),
.B(n_7074),
.Y(n_9473)
);

INVx1_ASAP7_75t_L g9474 ( 
.A(n_9307),
.Y(n_9474)
);

INVx1_ASAP7_75t_L g9475 ( 
.A(n_7910),
.Y(n_9475)
);

INVx1_ASAP7_75t_L g9476 ( 
.A(n_7910),
.Y(n_9476)
);

AOI22xp33_ASAP7_75t_L g9477 ( 
.A1(n_8417),
.A2(n_7621),
.B1(n_7113),
.B2(n_6969),
.Y(n_9477)
);

INVx2_ASAP7_75t_L g9478 ( 
.A(n_9202),
.Y(n_9478)
);

INVx1_ASAP7_75t_L g9479 ( 
.A(n_7910),
.Y(n_9479)
);

HB1xp67_ASAP7_75t_L g9480 ( 
.A(n_8073),
.Y(n_9480)
);

INVx1_ASAP7_75t_L g9481 ( 
.A(n_7911),
.Y(n_9481)
);

INVx2_ASAP7_75t_L g9482 ( 
.A(n_9202),
.Y(n_9482)
);

INVx6_ASAP7_75t_L g9483 ( 
.A(n_8102),
.Y(n_9483)
);

INVx3_ASAP7_75t_L g9484 ( 
.A(n_7934),
.Y(n_9484)
);

INVx2_ASAP7_75t_L g9485 ( 
.A(n_9233),
.Y(n_9485)
);

INVx1_ASAP7_75t_L g9486 ( 
.A(n_7911),
.Y(n_9486)
);

INVx1_ASAP7_75t_SL g9487 ( 
.A(n_7997),
.Y(n_9487)
);

INVx2_ASAP7_75t_L g9488 ( 
.A(n_9233),
.Y(n_9488)
);

INVx1_ASAP7_75t_L g9489 ( 
.A(n_7911),
.Y(n_9489)
);

NAND2x1p5_ASAP7_75t_L g9490 ( 
.A(n_7974),
.B(n_7776),
.Y(n_9490)
);

OAI22xp33_ASAP7_75t_L g9491 ( 
.A1(n_8076),
.A2(n_7931),
.B1(n_8409),
.B2(n_8404),
.Y(n_9491)
);

INVx2_ASAP7_75t_L g9492 ( 
.A(n_9233),
.Y(n_9492)
);

INVx2_ASAP7_75t_L g9493 ( 
.A(n_9233),
.Y(n_9493)
);

HB1xp67_ASAP7_75t_L g9494 ( 
.A(n_8073),
.Y(n_9494)
);

INVx1_ASAP7_75t_L g9495 ( 
.A(n_7918),
.Y(n_9495)
);

BUFx2_ASAP7_75t_SL g9496 ( 
.A(n_9231),
.Y(n_9496)
);

INVx1_ASAP7_75t_L g9497 ( 
.A(n_7918),
.Y(n_9497)
);

INVx1_ASAP7_75t_L g9498 ( 
.A(n_7918),
.Y(n_9498)
);

INVx4_ASAP7_75t_L g9499 ( 
.A(n_8201),
.Y(n_9499)
);

OAI22xp5_ASAP7_75t_L g9500 ( 
.A1(n_8076),
.A2(n_7546),
.B1(n_7545),
.B2(n_7204),
.Y(n_9500)
);

BUFx6f_ASAP7_75t_L g9501 ( 
.A(n_7989),
.Y(n_9501)
);

AOI22xp33_ASAP7_75t_L g9502 ( 
.A1(n_8015),
.A2(n_7113),
.B1(n_6969),
.B2(n_7427),
.Y(n_9502)
);

AOI21x1_ASAP7_75t_L g9503 ( 
.A1(n_8337),
.A2(n_8059),
.B(n_7957),
.Y(n_9503)
);

INVx2_ASAP7_75t_L g9504 ( 
.A(n_9233),
.Y(n_9504)
);

OAI22xp5_ASAP7_75t_L g9505 ( 
.A1(n_8436),
.A2(n_7546),
.B1(n_7545),
.B2(n_7204),
.Y(n_9505)
);

OR2x6_ASAP7_75t_L g9506 ( 
.A(n_8175),
.B(n_7651),
.Y(n_9506)
);

INVx2_ASAP7_75t_L g9507 ( 
.A(n_9233),
.Y(n_9507)
);

OR2x2_ASAP7_75t_L g9508 ( 
.A(n_7937),
.B(n_7671),
.Y(n_9508)
);

INVx1_ASAP7_75t_L g9509 ( 
.A(n_7924),
.Y(n_9509)
);

INVx2_ASAP7_75t_SL g9510 ( 
.A(n_8437),
.Y(n_9510)
);

INVx2_ASAP7_75t_L g9511 ( 
.A(n_9238),
.Y(n_9511)
);

NAND2x1p5_ASAP7_75t_L g9512 ( 
.A(n_7974),
.B(n_7776),
.Y(n_9512)
);

CKINVDCx5p33_ASAP7_75t_R g9513 ( 
.A(n_8817),
.Y(n_9513)
);

AOI22xp33_ASAP7_75t_L g9514 ( 
.A1(n_8015),
.A2(n_7427),
.B1(n_7549),
.B2(n_7504),
.Y(n_9514)
);

OAI22xp5_ASAP7_75t_L g9515 ( 
.A1(n_8436),
.A2(n_7546),
.B1(n_7204),
.B2(n_7410),
.Y(n_9515)
);

INVx2_ASAP7_75t_L g9516 ( 
.A(n_9238),
.Y(n_9516)
);

INVx1_ASAP7_75t_L g9517 ( 
.A(n_7924),
.Y(n_9517)
);

HB1xp67_ASAP7_75t_L g9518 ( 
.A(n_8107),
.Y(n_9518)
);

INVx1_ASAP7_75t_L g9519 ( 
.A(n_7924),
.Y(n_9519)
);

INVx2_ASAP7_75t_L g9520 ( 
.A(n_9238),
.Y(n_9520)
);

AND2x2_ASAP7_75t_L g9521 ( 
.A(n_8041),
.B(n_7133),
.Y(n_9521)
);

INVx1_ASAP7_75t_L g9522 ( 
.A(n_7958),
.Y(n_9522)
);

INVx2_ASAP7_75t_L g9523 ( 
.A(n_9238),
.Y(n_9523)
);

AOI22xp33_ASAP7_75t_L g9524 ( 
.A1(n_8024),
.A2(n_8094),
.B1(n_8189),
.B2(n_8899),
.Y(n_9524)
);

AND2x2_ASAP7_75t_L g9525 ( 
.A(n_8041),
.B(n_7133),
.Y(n_9525)
);

INVx1_ASAP7_75t_L g9526 ( 
.A(n_7958),
.Y(n_9526)
);

AOI22xp33_ASAP7_75t_SL g9527 ( 
.A1(n_8024),
.A2(n_7662),
.B1(n_7816),
.B2(n_7025),
.Y(n_9527)
);

INVx2_ASAP7_75t_L g9528 ( 
.A(n_9238),
.Y(n_9528)
);

CKINVDCx5p33_ASAP7_75t_R g9529 ( 
.A(n_8817),
.Y(n_9529)
);

NOR2x1_ASAP7_75t_R g9530 ( 
.A(n_7961),
.B(n_7877),
.Y(n_9530)
);

INVx2_ASAP7_75t_L g9531 ( 
.A(n_9238),
.Y(n_9531)
);

INVx1_ASAP7_75t_L g9532 ( 
.A(n_7958),
.Y(n_9532)
);

BUFx3_ASAP7_75t_L g9533 ( 
.A(n_8102),
.Y(n_9533)
);

NAND2x1p5_ASAP7_75t_L g9534 ( 
.A(n_7974),
.B(n_7776),
.Y(n_9534)
);

AND2x4_ASAP7_75t_L g9535 ( 
.A(n_7998),
.B(n_6926),
.Y(n_9535)
);

INVx1_ASAP7_75t_L g9536 ( 
.A(n_7965),
.Y(n_9536)
);

INVx1_ASAP7_75t_L g9537 ( 
.A(n_7965),
.Y(n_9537)
);

AO21x2_ASAP7_75t_L g9538 ( 
.A1(n_9156),
.A2(n_7285),
.B(n_7263),
.Y(n_9538)
);

AOI22xp33_ASAP7_75t_SL g9539 ( 
.A1(n_8024),
.A2(n_7816),
.B1(n_7127),
.B2(n_7155),
.Y(n_9539)
);

AND2x2_ASAP7_75t_L g9540 ( 
.A(n_8041),
.B(n_7133),
.Y(n_9540)
);

AOI22xp5_ASAP7_75t_L g9541 ( 
.A1(n_8220),
.A2(n_7127),
.B1(n_7228),
.B2(n_7374),
.Y(n_9541)
);

AOI222xp33_ASAP7_75t_L g9542 ( 
.A1(n_8886),
.A2(n_8902),
.B1(n_8445),
.B2(n_9253),
.C1(n_8899),
.C2(n_8702),
.Y(n_9542)
);

BUFx2_ASAP7_75t_R g9543 ( 
.A(n_8814),
.Y(n_9543)
);

AND2x2_ASAP7_75t_L g9544 ( 
.A(n_8041),
.B(n_7133),
.Y(n_9544)
);

INVx2_ASAP7_75t_L g9545 ( 
.A(n_9274),
.Y(n_9545)
);

OAI21xp5_ASAP7_75t_L g9546 ( 
.A1(n_8281),
.A2(n_7425),
.B(n_6955),
.Y(n_9546)
);

INVx1_ASAP7_75t_L g9547 ( 
.A(n_7965),
.Y(n_9547)
);

INVx1_ASAP7_75t_SL g9548 ( 
.A(n_7997),
.Y(n_9548)
);

INVx1_ASAP7_75t_L g9549 ( 
.A(n_7972),
.Y(n_9549)
);

NAND2x1p5_ASAP7_75t_L g9550 ( 
.A(n_7974),
.B(n_7776),
.Y(n_9550)
);

AOI22xp33_ASAP7_75t_SL g9551 ( 
.A1(n_8886),
.A2(n_7127),
.B1(n_7155),
.B2(n_7416),
.Y(n_9551)
);

AND2x2_ASAP7_75t_L g9552 ( 
.A(n_8043),
.B(n_7207),
.Y(n_9552)
);

INVx2_ASAP7_75t_L g9553 ( 
.A(n_9274),
.Y(n_9553)
);

CKINVDCx20_ASAP7_75t_R g9554 ( 
.A(n_9203),
.Y(n_9554)
);

INVx3_ASAP7_75t_L g9555 ( 
.A(n_7998),
.Y(n_9555)
);

BUFx2_ASAP7_75t_L g9556 ( 
.A(n_9082),
.Y(n_9556)
);

BUFx6f_ASAP7_75t_L g9557 ( 
.A(n_7989),
.Y(n_9557)
);

CKINVDCx6p67_ASAP7_75t_R g9558 ( 
.A(n_7997),
.Y(n_9558)
);

AOI22xp5_ASAP7_75t_L g9559 ( 
.A1(n_7982),
.A2(n_8094),
.B1(n_8902),
.B2(n_8091),
.Y(n_9559)
);

BUFx3_ASAP7_75t_L g9560 ( 
.A(n_8472),
.Y(n_9560)
);

INVx1_ASAP7_75t_SL g9561 ( 
.A(n_8247),
.Y(n_9561)
);

AND2x2_ASAP7_75t_L g9562 ( 
.A(n_8043),
.B(n_7207),
.Y(n_9562)
);

AOI22xp33_ASAP7_75t_SL g9563 ( 
.A1(n_8025),
.A2(n_7476),
.B1(n_7416),
.B2(n_7121),
.Y(n_9563)
);

INVx3_ASAP7_75t_L g9564 ( 
.A(n_8042),
.Y(n_9564)
);

AOI22xp33_ASAP7_75t_L g9565 ( 
.A1(n_8189),
.A2(n_7427),
.B1(n_7549),
.B2(n_7504),
.Y(n_9565)
);

INVx2_ASAP7_75t_L g9566 ( 
.A(n_9274),
.Y(n_9566)
);

AOI22xp33_ASAP7_75t_L g9567 ( 
.A1(n_7982),
.A2(n_7427),
.B1(n_7549),
.B2(n_7504),
.Y(n_9567)
);

INVx2_ASAP7_75t_L g9568 ( 
.A(n_9274),
.Y(n_9568)
);

INVx2_ASAP7_75t_L g9569 ( 
.A(n_9274),
.Y(n_9569)
);

AOI22xp5_ASAP7_75t_L g9570 ( 
.A1(n_8091),
.A2(n_7379),
.B1(n_7374),
.B2(n_7334),
.Y(n_9570)
);

AOI22xp33_ASAP7_75t_L g9571 ( 
.A1(n_8216),
.A2(n_7504),
.B1(n_7595),
.B2(n_7549),
.Y(n_9571)
);

OAI22xp5_ASAP7_75t_L g9572 ( 
.A1(n_8444),
.A2(n_7410),
.B1(n_7372),
.B2(n_7399),
.Y(n_9572)
);

INVx1_ASAP7_75t_L g9573 ( 
.A(n_7972),
.Y(n_9573)
);

INVx1_ASAP7_75t_L g9574 ( 
.A(n_7972),
.Y(n_9574)
);

INVx1_ASAP7_75t_L g9575 ( 
.A(n_7987),
.Y(n_9575)
);

INVx2_ASAP7_75t_SL g9576 ( 
.A(n_8437),
.Y(n_9576)
);

AOI22xp33_ASAP7_75t_L g9577 ( 
.A1(n_8216),
.A2(n_7504),
.B1(n_7595),
.B2(n_7549),
.Y(n_9577)
);

INVx1_ASAP7_75t_L g9578 ( 
.A(n_7987),
.Y(n_9578)
);

INVx1_ASAP7_75t_L g9579 ( 
.A(n_7987),
.Y(n_9579)
);

INVx3_ASAP7_75t_L g9580 ( 
.A(n_8042),
.Y(n_9580)
);

INVx1_ASAP7_75t_L g9581 ( 
.A(n_7999),
.Y(n_9581)
);

INVx1_ASAP7_75t_L g9582 ( 
.A(n_7999),
.Y(n_9582)
);

BUFx8_ASAP7_75t_L g9583 ( 
.A(n_8201),
.Y(n_9583)
);

BUFx6f_ASAP7_75t_L g9584 ( 
.A(n_7989),
.Y(n_9584)
);

INVx2_ASAP7_75t_L g9585 ( 
.A(n_9274),
.Y(n_9585)
);

INVx2_ASAP7_75t_L g9586 ( 
.A(n_9021),
.Y(n_9586)
);

OAI22xp5_ASAP7_75t_L g9587 ( 
.A1(n_8444),
.A2(n_7372),
.B1(n_7399),
.B2(n_7187),
.Y(n_9587)
);

INVx2_ASAP7_75t_L g9588 ( 
.A(n_9021),
.Y(n_9588)
);

INVx2_ASAP7_75t_L g9589 ( 
.A(n_9021),
.Y(n_9589)
);

NAND2xp5_ASAP7_75t_L g9590 ( 
.A(n_8038),
.B(n_7393),
.Y(n_9590)
);

OAI22xp5_ASAP7_75t_L g9591 ( 
.A1(n_8224),
.A2(n_7372),
.B1(n_7399),
.B2(n_7187),
.Y(n_9591)
);

OAI21x1_ASAP7_75t_L g9592 ( 
.A1(n_9164),
.A2(n_7819),
.B(n_7813),
.Y(n_9592)
);

BUFx2_ASAP7_75t_L g9593 ( 
.A(n_9163),
.Y(n_9593)
);

INVx2_ASAP7_75t_L g9594 ( 
.A(n_9027),
.Y(n_9594)
);

NAND2xp5_ASAP7_75t_L g9595 ( 
.A(n_8941),
.B(n_7675),
.Y(n_9595)
);

INVxp67_ASAP7_75t_L g9596 ( 
.A(n_8953),
.Y(n_9596)
);

INVx1_ASAP7_75t_L g9597 ( 
.A(n_7999),
.Y(n_9597)
);

AND2x2_ASAP7_75t_L g9598 ( 
.A(n_8043),
.B(n_7207),
.Y(n_9598)
);

OAI22xp5_ASAP7_75t_L g9599 ( 
.A1(n_8224),
.A2(n_7187),
.B1(n_7075),
.B2(n_7269),
.Y(n_9599)
);

OAI22xp5_ASAP7_75t_L g9600 ( 
.A1(n_8004),
.A2(n_7075),
.B1(n_7269),
.B2(n_7379),
.Y(n_9600)
);

INVx11_ASAP7_75t_L g9601 ( 
.A(n_8472),
.Y(n_9601)
);

AOI21xp5_ASAP7_75t_L g9602 ( 
.A1(n_8195),
.A2(n_7968),
.B(n_8307),
.Y(n_9602)
);

INVx2_ASAP7_75t_L g9603 ( 
.A(n_9027),
.Y(n_9603)
);

BUFx2_ASAP7_75t_R g9604 ( 
.A(n_8814),
.Y(n_9604)
);

INVxp67_ASAP7_75t_SL g9605 ( 
.A(n_8422),
.Y(n_9605)
);

BUFx3_ASAP7_75t_L g9606 ( 
.A(n_8472),
.Y(n_9606)
);

BUFx3_ASAP7_75t_L g9607 ( 
.A(n_8472),
.Y(n_9607)
);

CKINVDCx20_ASAP7_75t_R g9608 ( 
.A(n_9203),
.Y(n_9608)
);

INVx1_ASAP7_75t_L g9609 ( 
.A(n_8001),
.Y(n_9609)
);

CKINVDCx11_ASAP7_75t_R g9610 ( 
.A(n_8075),
.Y(n_9610)
);

INVx2_ASAP7_75t_L g9611 ( 
.A(n_9027),
.Y(n_9611)
);

OAI21xp5_ASAP7_75t_L g9612 ( 
.A1(n_8281),
.A2(n_7425),
.B(n_6955),
.Y(n_9612)
);

AO21x1_ASAP7_75t_L g9613 ( 
.A1(n_8495),
.A2(n_7340),
.B(n_7287),
.Y(n_9613)
);

OA21x2_ASAP7_75t_L g9614 ( 
.A1(n_8900),
.A2(n_7108),
.B(n_7081),
.Y(n_9614)
);

INVx2_ASAP7_75t_SL g9615 ( 
.A(n_8437),
.Y(n_9615)
);

AOI22xp33_ASAP7_75t_L g9616 ( 
.A1(n_8998),
.A2(n_7504),
.B1(n_7595),
.B2(n_7549),
.Y(n_9616)
);

AND2x2_ASAP7_75t_L g9617 ( 
.A(n_8043),
.B(n_7207),
.Y(n_9617)
);

INVx1_ASAP7_75t_L g9618 ( 
.A(n_8001),
.Y(n_9618)
);

OR2x6_ASAP7_75t_L g9619 ( 
.A(n_8766),
.B(n_7651),
.Y(n_9619)
);

INVx3_ASAP7_75t_L g9620 ( 
.A(n_8042),
.Y(n_9620)
);

NAND2x1p5_ASAP7_75t_L g9621 ( 
.A(n_7974),
.B(n_7776),
.Y(n_9621)
);

INVx2_ASAP7_75t_L g9622 ( 
.A(n_9031),
.Y(n_9622)
);

BUFx2_ASAP7_75t_L g9623 ( 
.A(n_9163),
.Y(n_9623)
);

INVx1_ASAP7_75t_L g9624 ( 
.A(n_8001),
.Y(n_9624)
);

INVx2_ASAP7_75t_L g9625 ( 
.A(n_9031),
.Y(n_9625)
);

NOR2xp33_ASAP7_75t_L g9626 ( 
.A(n_8366),
.B(n_7429),
.Y(n_9626)
);

INVx1_ASAP7_75t_L g9627 ( 
.A(n_8009),
.Y(n_9627)
);

AOI22xp5_ASAP7_75t_L g9628 ( 
.A1(n_8308),
.A2(n_7334),
.B1(n_7062),
.B2(n_7425),
.Y(n_9628)
);

INVx3_ASAP7_75t_L g9629 ( 
.A(n_8042),
.Y(n_9629)
);

HB1xp67_ASAP7_75t_L g9630 ( 
.A(n_8107),
.Y(n_9630)
);

INVx1_ASAP7_75t_L g9631 ( 
.A(n_8009),
.Y(n_9631)
);

CKINVDCx6p67_ASAP7_75t_R g9632 ( 
.A(n_8201),
.Y(n_9632)
);

AOI22xp33_ASAP7_75t_L g9633 ( 
.A1(n_8998),
.A2(n_7504),
.B1(n_7595),
.B2(n_7549),
.Y(n_9633)
);

BUFx8_ASAP7_75t_SL g9634 ( 
.A(n_7933),
.Y(n_9634)
);

INVx1_ASAP7_75t_L g9635 ( 
.A(n_8009),
.Y(n_9635)
);

INVx1_ASAP7_75t_L g9636 ( 
.A(n_8029),
.Y(n_9636)
);

AOI22xp33_ASAP7_75t_L g9637 ( 
.A1(n_8434),
.A2(n_7549),
.B1(n_7628),
.B2(n_7595),
.Y(n_9637)
);

INVx2_ASAP7_75t_L g9638 ( 
.A(n_9031),
.Y(n_9638)
);

INVx1_ASAP7_75t_L g9639 ( 
.A(n_8029),
.Y(n_9639)
);

HB1xp67_ASAP7_75t_L g9640 ( 
.A(n_8112),
.Y(n_9640)
);

INVx2_ASAP7_75t_SL g9641 ( 
.A(n_8437),
.Y(n_9641)
);

OAI21x1_ASAP7_75t_L g9642 ( 
.A1(n_9198),
.A2(n_9308),
.B(n_9300),
.Y(n_9642)
);

INVx1_ASAP7_75t_L g9643 ( 
.A(n_8029),
.Y(n_9643)
);

OR2x6_ASAP7_75t_L g9644 ( 
.A(n_8837),
.B(n_7651),
.Y(n_9644)
);

INVx2_ASAP7_75t_SL g9645 ( 
.A(n_8696),
.Y(n_9645)
);

OAI22xp5_ASAP7_75t_L g9646 ( 
.A1(n_8004),
.A2(n_7098),
.B1(n_7299),
.B2(n_7047),
.Y(n_9646)
);

INVx2_ASAP7_75t_L g9647 ( 
.A(n_9033),
.Y(n_9647)
);

AOI22xp33_ASAP7_75t_SL g9648 ( 
.A1(n_8025),
.A2(n_7476),
.B1(n_7416),
.B2(n_7121),
.Y(n_9648)
);

HB1xp67_ASAP7_75t_L g9649 ( 
.A(n_8112),
.Y(n_9649)
);

INVx2_ASAP7_75t_SL g9650 ( 
.A(n_8696),
.Y(n_9650)
);

INVx1_ASAP7_75t_L g9651 ( 
.A(n_8031),
.Y(n_9651)
);

AO21x1_ASAP7_75t_L g9652 ( 
.A1(n_8495),
.A2(n_7340),
.B(n_7287),
.Y(n_9652)
);

INVx2_ASAP7_75t_L g9653 ( 
.A(n_9033),
.Y(n_9653)
);

BUFx2_ASAP7_75t_L g9654 ( 
.A(n_8472),
.Y(n_9654)
);

OAI21x1_ASAP7_75t_L g9655 ( 
.A1(n_9198),
.A2(n_7819),
.B(n_7813),
.Y(n_9655)
);

INVx1_ASAP7_75t_L g9656 ( 
.A(n_8031),
.Y(n_9656)
);

INVx1_ASAP7_75t_L g9657 ( 
.A(n_8031),
.Y(n_9657)
);

AND2x2_ASAP7_75t_L g9658 ( 
.A(n_8043),
.B(n_7207),
.Y(n_9658)
);

INVx1_ASAP7_75t_L g9659 ( 
.A(n_8040),
.Y(n_9659)
);

INVx1_ASAP7_75t_L g9660 ( 
.A(n_8040),
.Y(n_9660)
);

AOI22xp33_ASAP7_75t_SL g9661 ( 
.A1(n_8025),
.A2(n_7476),
.B1(n_7121),
.B2(n_7128),
.Y(n_9661)
);

AOI22xp33_ASAP7_75t_L g9662 ( 
.A1(n_8434),
.A2(n_7595),
.B1(n_7744),
.B2(n_7628),
.Y(n_9662)
);

CKINVDCx11_ASAP7_75t_R g9663 ( 
.A(n_8075),
.Y(n_9663)
);

INVx4_ASAP7_75t_L g9664 ( 
.A(n_8201),
.Y(n_9664)
);

INVx3_ASAP7_75t_L g9665 ( 
.A(n_8046),
.Y(n_9665)
);

INVx1_ASAP7_75t_L g9666 ( 
.A(n_8040),
.Y(n_9666)
);

INVx1_ASAP7_75t_L g9667 ( 
.A(n_8063),
.Y(n_9667)
);

BUFx12f_ASAP7_75t_L g9668 ( 
.A(n_7933),
.Y(n_9668)
);

NAND2x1p5_ASAP7_75t_L g9669 ( 
.A(n_7992),
.B(n_7780),
.Y(n_9669)
);

NAND2xp5_ASAP7_75t_L g9670 ( 
.A(n_8941),
.B(n_7256),
.Y(n_9670)
);

INVx1_ASAP7_75t_L g9671 ( 
.A(n_8063),
.Y(n_9671)
);

AND2x2_ASAP7_75t_L g9672 ( 
.A(n_8043),
.B(n_7207),
.Y(n_9672)
);

INVx2_ASAP7_75t_L g9673 ( 
.A(n_9033),
.Y(n_9673)
);

INVx2_ASAP7_75t_SL g9674 ( 
.A(n_8696),
.Y(n_9674)
);

OAI22xp33_ASAP7_75t_L g9675 ( 
.A1(n_8409),
.A2(n_7088),
.B1(n_7098),
.B2(n_7118),
.Y(n_9675)
);

INVx1_ASAP7_75t_L g9676 ( 
.A(n_8063),
.Y(n_9676)
);

HB1xp67_ASAP7_75t_L g9677 ( 
.A(n_8166),
.Y(n_9677)
);

AOI21x1_ASAP7_75t_L g9678 ( 
.A1(n_8337),
.A2(n_7158),
.B(n_7154),
.Y(n_9678)
);

AOI22xp33_ASAP7_75t_L g9679 ( 
.A1(n_8039),
.A2(n_7595),
.B1(n_7744),
.B2(n_7628),
.Y(n_9679)
);

OAI21xp5_ASAP7_75t_L g9680 ( 
.A1(n_8445),
.A2(n_6955),
.B(n_7088),
.Y(n_9680)
);

AND2x2_ASAP7_75t_L g9681 ( 
.A(n_8060),
.B(n_8061),
.Y(n_9681)
);

INVx2_ASAP7_75t_L g9682 ( 
.A(n_9034),
.Y(n_9682)
);

AND2x2_ASAP7_75t_L g9683 ( 
.A(n_8060),
.B(n_7322),
.Y(n_9683)
);

BUFx2_ASAP7_75t_L g9684 ( 
.A(n_8472),
.Y(n_9684)
);

INVx2_ASAP7_75t_L g9685 ( 
.A(n_9034),
.Y(n_9685)
);

BUFx3_ASAP7_75t_L g9686 ( 
.A(n_8891),
.Y(n_9686)
);

INVx2_ASAP7_75t_L g9687 ( 
.A(n_9034),
.Y(n_9687)
);

INVx1_ASAP7_75t_L g9688 ( 
.A(n_8089),
.Y(n_9688)
);

INVx2_ASAP7_75t_L g9689 ( 
.A(n_9037),
.Y(n_9689)
);

NAND2xp5_ASAP7_75t_L g9690 ( 
.A(n_8347),
.B(n_7256),
.Y(n_9690)
);

INVx1_ASAP7_75t_L g9691 ( 
.A(n_8089),
.Y(n_9691)
);

INVx1_ASAP7_75t_L g9692 ( 
.A(n_8089),
.Y(n_9692)
);

INVx1_ASAP7_75t_L g9693 ( 
.A(n_8105),
.Y(n_9693)
);

AOI22xp33_ASAP7_75t_L g9694 ( 
.A1(n_8039),
.A2(n_7595),
.B1(n_7744),
.B2(n_7628),
.Y(n_9694)
);

INVx1_ASAP7_75t_L g9695 ( 
.A(n_8105),
.Y(n_9695)
);

INVx1_ASAP7_75t_L g9696 ( 
.A(n_8105),
.Y(n_9696)
);

INVx1_ASAP7_75t_L g9697 ( 
.A(n_8108),
.Y(n_9697)
);

OAI22xp5_ASAP7_75t_L g9698 ( 
.A1(n_8070),
.A2(n_7098),
.B1(n_7299),
.B2(n_7047),
.Y(n_9698)
);

BUFx2_ASAP7_75t_R g9699 ( 
.A(n_7936),
.Y(n_9699)
);

AOI22xp33_ASAP7_75t_L g9700 ( 
.A1(n_8471),
.A2(n_7628),
.B1(n_7801),
.B2(n_7744),
.Y(n_9700)
);

AOI22xp33_ASAP7_75t_L g9701 ( 
.A1(n_8471),
.A2(n_7628),
.B1(n_7801),
.B2(n_7744),
.Y(n_9701)
);

AND2x2_ASAP7_75t_L g9702 ( 
.A(n_8060),
.B(n_8061),
.Y(n_9702)
);

AOI22xp33_ASAP7_75t_L g9703 ( 
.A1(n_8543),
.A2(n_7628),
.B1(n_7801),
.B2(n_7744),
.Y(n_9703)
);

INVx2_ASAP7_75t_SL g9704 ( 
.A(n_8696),
.Y(n_9704)
);

INVx2_ASAP7_75t_L g9705 ( 
.A(n_9037),
.Y(n_9705)
);

BUFx2_ASAP7_75t_L g9706 ( 
.A(n_8878),
.Y(n_9706)
);

AOI22xp33_ASAP7_75t_L g9707 ( 
.A1(n_8543),
.A2(n_7628),
.B1(n_7801),
.B2(n_7744),
.Y(n_9707)
);

NAND2x1p5_ASAP7_75t_L g9708 ( 
.A(n_7992),
.B(n_7780),
.Y(n_9708)
);

NOR2xp33_ASAP7_75t_L g9709 ( 
.A(n_7961),
.B(n_7443),
.Y(n_9709)
);

OAI22xp5_ASAP7_75t_SL g9710 ( 
.A1(n_8293),
.A2(n_7465),
.B1(n_7484),
.B2(n_7443),
.Y(n_9710)
);

INVx1_ASAP7_75t_L g9711 ( 
.A(n_8108),
.Y(n_9711)
);

AND2x4_ASAP7_75t_L g9712 ( 
.A(n_8046),
.B(n_8120),
.Y(n_9712)
);

INVx1_ASAP7_75t_L g9713 ( 
.A(n_8108),
.Y(n_9713)
);

INVx4_ASAP7_75t_L g9714 ( 
.A(n_8696),
.Y(n_9714)
);

INVx2_ASAP7_75t_L g9715 ( 
.A(n_9037),
.Y(n_9715)
);

INVx2_ASAP7_75t_L g9716 ( 
.A(n_8853),
.Y(n_9716)
);

INVx1_ASAP7_75t_L g9717 ( 
.A(n_8113),
.Y(n_9717)
);

BUFx4f_ASAP7_75t_SL g9718 ( 
.A(n_9096),
.Y(n_9718)
);

INVx5_ASAP7_75t_L g9719 ( 
.A(n_7926),
.Y(n_9719)
);

AOI22xp5_ASAP7_75t_L g9720 ( 
.A1(n_8308),
.A2(n_7062),
.B1(n_7118),
.B2(n_6958),
.Y(n_9720)
);

INVx2_ASAP7_75t_SL g9721 ( 
.A(n_8696),
.Y(n_9721)
);

INVx3_ASAP7_75t_L g9722 ( 
.A(n_8046),
.Y(n_9722)
);

BUFx4f_ASAP7_75t_L g9723 ( 
.A(n_8097),
.Y(n_9723)
);

INVx1_ASAP7_75t_SL g9724 ( 
.A(n_8247),
.Y(n_9724)
);

INVx2_ASAP7_75t_L g9725 ( 
.A(n_8853),
.Y(n_9725)
);

INVx1_ASAP7_75t_L g9726 ( 
.A(n_8113),
.Y(n_9726)
);

AOI22xp33_ASAP7_75t_L g9727 ( 
.A1(n_8020),
.A2(n_7801),
.B1(n_7744),
.B2(n_7176),
.Y(n_9727)
);

INVx1_ASAP7_75t_L g9728 ( 
.A(n_8113),
.Y(n_9728)
);

INVx2_ASAP7_75t_L g9729 ( 
.A(n_8853),
.Y(n_9729)
);

NAND2xp5_ASAP7_75t_L g9730 ( 
.A(n_8347),
.B(n_7270),
.Y(n_9730)
);

AO21x1_ASAP7_75t_SL g9731 ( 
.A1(n_8470),
.A2(n_7860),
.B(n_7834),
.Y(n_9731)
);

INVx1_ASAP7_75t_L g9732 ( 
.A(n_8122),
.Y(n_9732)
);

INVxp33_ASAP7_75t_L g9733 ( 
.A(n_8473),
.Y(n_9733)
);

INVx3_ASAP7_75t_L g9734 ( 
.A(n_8046),
.Y(n_9734)
);

AOI22xp33_ASAP7_75t_L g9735 ( 
.A1(n_8020),
.A2(n_7801),
.B1(n_7176),
.B2(n_7088),
.Y(n_9735)
);

INVx1_ASAP7_75t_L g9736 ( 
.A(n_8122),
.Y(n_9736)
);

INVx1_ASAP7_75t_L g9737 ( 
.A(n_8122),
.Y(n_9737)
);

AOI21x1_ASAP7_75t_L g9738 ( 
.A1(n_8059),
.A2(n_7158),
.B(n_7154),
.Y(n_9738)
);

BUFx2_ASAP7_75t_R g9739 ( 
.A(n_7936),
.Y(n_9739)
);

INVx1_ASAP7_75t_L g9740 ( 
.A(n_8123),
.Y(n_9740)
);

BUFx2_ASAP7_75t_L g9741 ( 
.A(n_8878),
.Y(n_9741)
);

AOI22xp33_ASAP7_75t_SL g9742 ( 
.A1(n_8519),
.A2(n_7121),
.B1(n_7128),
.B2(n_7079),
.Y(n_9742)
);

INVx2_ASAP7_75t_L g9743 ( 
.A(n_8856),
.Y(n_9743)
);

AOI22xp33_ASAP7_75t_SL g9744 ( 
.A1(n_8519),
.A2(n_7121),
.B1(n_7128),
.B2(n_7079),
.Y(n_9744)
);

BUFx2_ASAP7_75t_R g9745 ( 
.A(n_7947),
.Y(n_9745)
);

INVx2_ASAP7_75t_SL g9746 ( 
.A(n_8696),
.Y(n_9746)
);

OA21x2_ASAP7_75t_L g9747 ( 
.A1(n_7954),
.A2(n_7112),
.B(n_7108),
.Y(n_9747)
);

INVx2_ASAP7_75t_L g9748 ( 
.A(n_8856),
.Y(n_9748)
);

AOI22xp33_ASAP7_75t_L g9749 ( 
.A1(n_8265),
.A2(n_7801),
.B1(n_7176),
.B2(n_7238),
.Y(n_9749)
);

INVx2_ASAP7_75t_L g9750 ( 
.A(n_8856),
.Y(n_9750)
);

BUFx12f_ASAP7_75t_L g9751 ( 
.A(n_9002),
.Y(n_9751)
);

INVx1_ASAP7_75t_L g9752 ( 
.A(n_8123),
.Y(n_9752)
);

INVx1_ASAP7_75t_L g9753 ( 
.A(n_8123),
.Y(n_9753)
);

INVx3_ASAP7_75t_L g9754 ( 
.A(n_8120),
.Y(n_9754)
);

CKINVDCx11_ASAP7_75t_R g9755 ( 
.A(n_9096),
.Y(n_9755)
);

INVx1_ASAP7_75t_L g9756 ( 
.A(n_8133),
.Y(n_9756)
);

INVx1_ASAP7_75t_L g9757 ( 
.A(n_8133),
.Y(n_9757)
);

HB1xp67_ASAP7_75t_L g9758 ( 
.A(n_8166),
.Y(n_9758)
);

INVx2_ASAP7_75t_L g9759 ( 
.A(n_8859),
.Y(n_9759)
);

NAND2xp5_ASAP7_75t_SL g9760 ( 
.A(n_7989),
.B(n_7465),
.Y(n_9760)
);

BUFx6f_ASAP7_75t_L g9761 ( 
.A(n_7989),
.Y(n_9761)
);

BUFx3_ASAP7_75t_L g9762 ( 
.A(n_8891),
.Y(n_9762)
);

INVx2_ASAP7_75t_L g9763 ( 
.A(n_8859),
.Y(n_9763)
);

INVx2_ASAP7_75t_SL g9764 ( 
.A(n_8414),
.Y(n_9764)
);

OAI22xp5_ASAP7_75t_L g9765 ( 
.A1(n_8070),
.A2(n_7299),
.B1(n_7303),
.B2(n_7047),
.Y(n_9765)
);

BUFx3_ASAP7_75t_L g9766 ( 
.A(n_8891),
.Y(n_9766)
);

INVx3_ASAP7_75t_L g9767 ( 
.A(n_8120),
.Y(n_9767)
);

BUFx2_ASAP7_75t_SL g9768 ( 
.A(n_9231),
.Y(n_9768)
);

OAI22xp5_ASAP7_75t_L g9769 ( 
.A1(n_8404),
.A2(n_7299),
.B1(n_7303),
.B2(n_7047),
.Y(n_9769)
);

INVx2_ASAP7_75t_L g9770 ( 
.A(n_8859),
.Y(n_9770)
);

INVx1_ASAP7_75t_L g9771 ( 
.A(n_8133),
.Y(n_9771)
);

INVx1_ASAP7_75t_L g9772 ( 
.A(n_8145),
.Y(n_9772)
);

AND2x2_ASAP7_75t_L g9773 ( 
.A(n_8060),
.B(n_7322),
.Y(n_9773)
);

INVx2_ASAP7_75t_L g9774 ( 
.A(n_8946),
.Y(n_9774)
);

INVx1_ASAP7_75t_L g9775 ( 
.A(n_8145),
.Y(n_9775)
);

AND2x4_ASAP7_75t_L g9776 ( 
.A(n_8120),
.B(n_6926),
.Y(n_9776)
);

INVx1_ASAP7_75t_L g9777 ( 
.A(n_8145),
.Y(n_9777)
);

NAND2xp5_ASAP7_75t_L g9778 ( 
.A(n_8397),
.B(n_7270),
.Y(n_9778)
);

OAI21x1_ASAP7_75t_L g9779 ( 
.A1(n_9300),
.A2(n_7821),
.B(n_7819),
.Y(n_9779)
);

AOI22xp33_ASAP7_75t_L g9780 ( 
.A1(n_8265),
.A2(n_7801),
.B1(n_7176),
.B2(n_7238),
.Y(n_9780)
);

AOI22xp33_ASAP7_75t_SL g9781 ( 
.A1(n_8116),
.A2(n_7121),
.B1(n_7128),
.B2(n_7079),
.Y(n_9781)
);

INVx2_ASAP7_75t_L g9782 ( 
.A(n_8946),
.Y(n_9782)
);

OAI22xp33_ASAP7_75t_L g9783 ( 
.A1(n_8385),
.A2(n_7118),
.B1(n_7013),
.B2(n_7664),
.Y(n_9783)
);

BUFx2_ASAP7_75t_SL g9784 ( 
.A(n_8422),
.Y(n_9784)
);

INVx3_ASAP7_75t_L g9785 ( 
.A(n_8152),
.Y(n_9785)
);

INVx2_ASAP7_75t_SL g9786 ( 
.A(n_8414),
.Y(n_9786)
);

HB1xp67_ASAP7_75t_L g9787 ( 
.A(n_8221),
.Y(n_9787)
);

INVx1_ASAP7_75t_L g9788 ( 
.A(n_8147),
.Y(n_9788)
);

AOI22xp33_ASAP7_75t_SL g9789 ( 
.A1(n_8116),
.A2(n_7128),
.B1(n_7246),
.B2(n_7079),
.Y(n_9789)
);

INVx1_ASAP7_75t_L g9790 ( 
.A(n_8147),
.Y(n_9790)
);

AOI222xp33_ASAP7_75t_L g9791 ( 
.A1(n_9253),
.A2(n_7017),
.B1(n_7340),
.B2(n_7287),
.C1(n_7414),
.C2(n_6967),
.Y(n_9791)
);

INVx1_ASAP7_75t_L g9792 ( 
.A(n_8147),
.Y(n_9792)
);

BUFx2_ASAP7_75t_L g9793 ( 
.A(n_8878),
.Y(n_9793)
);

AOI22xp33_ASAP7_75t_L g9794 ( 
.A1(n_8275),
.A2(n_7176),
.B1(n_7238),
.B2(n_7213),
.Y(n_9794)
);

INVx2_ASAP7_75t_L g9795 ( 
.A(n_8946),
.Y(n_9795)
);

AO21x1_ASAP7_75t_SL g9796 ( 
.A1(n_8470),
.A2(n_7513),
.B(n_7505),
.Y(n_9796)
);

BUFx2_ASAP7_75t_L g9797 ( 
.A(n_8878),
.Y(n_9797)
);

INVx1_ASAP7_75t_L g9798 ( 
.A(n_8148),
.Y(n_9798)
);

BUFx4f_ASAP7_75t_L g9799 ( 
.A(n_8097),
.Y(n_9799)
);

INVx2_ASAP7_75t_L g9800 ( 
.A(n_8958),
.Y(n_9800)
);

BUFx3_ASAP7_75t_L g9801 ( 
.A(n_8891),
.Y(n_9801)
);

AND2x4_ASAP7_75t_L g9802 ( 
.A(n_8152),
.B(n_6926),
.Y(n_9802)
);

INVx1_ASAP7_75t_L g9803 ( 
.A(n_8148),
.Y(n_9803)
);

AOI21x1_ASAP7_75t_L g9804 ( 
.A1(n_8059),
.A2(n_7158),
.B(n_7154),
.Y(n_9804)
);

BUFx2_ASAP7_75t_L g9805 ( 
.A(n_8878),
.Y(n_9805)
);

BUFx3_ASAP7_75t_L g9806 ( 
.A(n_8891),
.Y(n_9806)
);

OAI22xp33_ASAP7_75t_SL g9807 ( 
.A1(n_8139),
.A2(n_7484),
.B1(n_7461),
.B2(n_7293),
.Y(n_9807)
);

INVx5_ASAP7_75t_L g9808 ( 
.A(n_7926),
.Y(n_9808)
);

INVx2_ASAP7_75t_L g9809 ( 
.A(n_8958),
.Y(n_9809)
);

BUFx3_ASAP7_75t_L g9810 ( 
.A(n_8891),
.Y(n_9810)
);

INVx1_ASAP7_75t_L g9811 ( 
.A(n_8148),
.Y(n_9811)
);

AOI22xp33_ASAP7_75t_L g9812 ( 
.A1(n_8275),
.A2(n_7176),
.B1(n_7253),
.B2(n_7213),
.Y(n_9812)
);

INVx1_ASAP7_75t_L g9813 ( 
.A(n_8153),
.Y(n_9813)
);

INVx2_ASAP7_75t_L g9814 ( 
.A(n_8958),
.Y(n_9814)
);

INVx1_ASAP7_75t_L g9815 ( 
.A(n_8153),
.Y(n_9815)
);

AOI22xp33_ASAP7_75t_L g9816 ( 
.A1(n_8398),
.A2(n_7176),
.B1(n_7253),
.B2(n_7213),
.Y(n_9816)
);

AOI22xp33_ASAP7_75t_L g9817 ( 
.A1(n_8398),
.A2(n_7176),
.B1(n_7268),
.B2(n_7253),
.Y(n_9817)
);

BUFx6f_ASAP7_75t_L g9818 ( 
.A(n_8797),
.Y(n_9818)
);

AOI22xp33_ASAP7_75t_L g9819 ( 
.A1(n_8398),
.A2(n_7283),
.B1(n_7289),
.B2(n_7268),
.Y(n_9819)
);

INVx8_ASAP7_75t_L g9820 ( 
.A(n_9278),
.Y(n_9820)
);

HB1xp67_ASAP7_75t_L g9821 ( 
.A(n_8221),
.Y(n_9821)
);

INVx1_ASAP7_75t_L g9822 ( 
.A(n_8153),
.Y(n_9822)
);

INVx2_ASAP7_75t_L g9823 ( 
.A(n_8963),
.Y(n_9823)
);

BUFx6f_ASAP7_75t_L g9824 ( 
.A(n_8797),
.Y(n_9824)
);

INVx1_ASAP7_75t_L g9825 ( 
.A(n_8167),
.Y(n_9825)
);

OAI21x1_ASAP7_75t_L g9826 ( 
.A1(n_9308),
.A2(n_7821),
.B(n_7819),
.Y(n_9826)
);

AND2x2_ASAP7_75t_L g9827 ( 
.A(n_8060),
.B(n_7322),
.Y(n_9827)
);

BUFx8_ASAP7_75t_SL g9828 ( 
.A(n_9002),
.Y(n_9828)
);

AOI22xp33_ASAP7_75t_L g9829 ( 
.A1(n_8526),
.A2(n_7283),
.B1(n_7289),
.B2(n_7268),
.Y(n_9829)
);

INVx1_ASAP7_75t_L g9830 ( 
.A(n_8167),
.Y(n_9830)
);

AND2x4_ASAP7_75t_L g9831 ( 
.A(n_8152),
.B(n_6930),
.Y(n_9831)
);

AOI21x1_ASAP7_75t_L g9832 ( 
.A1(n_8228),
.A2(n_7159),
.B(n_7158),
.Y(n_9832)
);

AND2x2_ASAP7_75t_L g9833 ( 
.A(n_8060),
.B(n_7322),
.Y(n_9833)
);

AND2x2_ASAP7_75t_L g9834 ( 
.A(n_8061),
.B(n_7322),
.Y(n_9834)
);

NAND2xp5_ASAP7_75t_L g9835 ( 
.A(n_8397),
.B(n_7873),
.Y(n_9835)
);

INVx2_ASAP7_75t_SL g9836 ( 
.A(n_8414),
.Y(n_9836)
);

INVx2_ASAP7_75t_L g9837 ( 
.A(n_8963),
.Y(n_9837)
);

INVx1_ASAP7_75t_L g9838 ( 
.A(n_8167),
.Y(n_9838)
);

OAI22xp5_ASAP7_75t_SL g9839 ( 
.A1(n_8293),
.A2(n_7252),
.B1(n_7304),
.B2(n_7221),
.Y(n_9839)
);

INVx1_ASAP7_75t_L g9840 ( 
.A(n_8173),
.Y(n_9840)
);

INVx2_ASAP7_75t_L g9841 ( 
.A(n_8963),
.Y(n_9841)
);

AOI22xp33_ASAP7_75t_L g9842 ( 
.A1(n_8526),
.A2(n_7289),
.B1(n_7301),
.B2(n_7283),
.Y(n_9842)
);

HB1xp67_ASAP7_75t_L g9843 ( 
.A(n_9269),
.Y(n_9843)
);

INVxp67_ASAP7_75t_L g9844 ( 
.A(n_8953),
.Y(n_9844)
);

INVx2_ASAP7_75t_L g9845 ( 
.A(n_9076),
.Y(n_9845)
);

INVx1_ASAP7_75t_L g9846 ( 
.A(n_8173),
.Y(n_9846)
);

OAI21x1_ASAP7_75t_L g9847 ( 
.A1(n_8940),
.A2(n_7841),
.B(n_7821),
.Y(n_9847)
);

AO21x2_ASAP7_75t_L g9848 ( 
.A1(n_8550),
.A2(n_7646),
.B(n_7508),
.Y(n_9848)
);

HB1xp67_ASAP7_75t_L g9849 ( 
.A(n_9269),
.Y(n_9849)
);

AOI22xp33_ASAP7_75t_SL g9850 ( 
.A1(n_8116),
.A2(n_7079),
.B1(n_7246),
.B2(n_7128),
.Y(n_9850)
);

INVx1_ASAP7_75t_L g9851 ( 
.A(n_8173),
.Y(n_9851)
);

AND2x2_ASAP7_75t_L g9852 ( 
.A(n_8061),
.B(n_7322),
.Y(n_9852)
);

BUFx12f_ASAP7_75t_L g9853 ( 
.A(n_9093),
.Y(n_9853)
);

HB1xp67_ASAP7_75t_L g9854 ( 
.A(n_9273),
.Y(n_9854)
);

AO21x2_ASAP7_75t_L g9855 ( 
.A1(n_8550),
.A2(n_7646),
.B(n_7508),
.Y(n_9855)
);

OAI21x1_ASAP7_75t_SL g9856 ( 
.A1(n_8559),
.A2(n_6919),
.B(n_6915),
.Y(n_9856)
);

INVx1_ASAP7_75t_L g9857 ( 
.A(n_8174),
.Y(n_9857)
);

BUFx10_ASAP7_75t_L g9858 ( 
.A(n_8263),
.Y(n_9858)
);

INVx1_ASAP7_75t_L g9859 ( 
.A(n_8174),
.Y(n_9859)
);

OAI21x1_ASAP7_75t_L g9860 ( 
.A1(n_8940),
.A2(n_7841),
.B(n_7821),
.Y(n_9860)
);

BUFx3_ASAP7_75t_L g9861 ( 
.A(n_9044),
.Y(n_9861)
);

BUFx3_ASAP7_75t_L g9862 ( 
.A(n_9044),
.Y(n_9862)
);

BUFx2_ASAP7_75t_L g9863 ( 
.A(n_8878),
.Y(n_9863)
);

AOI22xp33_ASAP7_75t_SL g9864 ( 
.A1(n_8375),
.A2(n_7977),
.B1(n_8460),
.B2(n_8293),
.Y(n_9864)
);

INVx2_ASAP7_75t_L g9865 ( 
.A(n_9076),
.Y(n_9865)
);

BUFx12f_ASAP7_75t_L g9866 ( 
.A(n_9093),
.Y(n_9866)
);

OAI22xp33_ASAP7_75t_L g9867 ( 
.A1(n_8385),
.A2(n_8537),
.B1(n_9170),
.B2(n_8161),
.Y(n_9867)
);

NAND2xp5_ASAP7_75t_L g9868 ( 
.A(n_8400),
.B(n_7873),
.Y(n_9868)
);

BUFx2_ASAP7_75t_R g9869 ( 
.A(n_7947),
.Y(n_9869)
);

INVx1_ASAP7_75t_L g9870 ( 
.A(n_8174),
.Y(n_9870)
);

INVx1_ASAP7_75t_L g9871 ( 
.A(n_8177),
.Y(n_9871)
);

AOI22xp33_ASAP7_75t_SL g9872 ( 
.A1(n_8375),
.A2(n_7977),
.B1(n_8695),
.B2(n_8460),
.Y(n_9872)
);

AOI22xp33_ASAP7_75t_SL g9873 ( 
.A1(n_8460),
.A2(n_8722),
.B1(n_8695),
.B2(n_8808),
.Y(n_9873)
);

OAI21x1_ASAP7_75t_L g9874 ( 
.A1(n_8940),
.A2(n_7841),
.B(n_7821),
.Y(n_9874)
);

INVx2_ASAP7_75t_L g9875 ( 
.A(n_9076),
.Y(n_9875)
);

AO21x1_ASAP7_75t_L g9876 ( 
.A1(n_8139),
.A2(n_8808),
.B(n_7925),
.Y(n_9876)
);

OR2x6_ASAP7_75t_L g9877 ( 
.A(n_8837),
.B(n_7109),
.Y(n_9877)
);

CKINVDCx5p33_ASAP7_75t_R g9878 ( 
.A(n_8263),
.Y(n_9878)
);

INVx1_ASAP7_75t_L g9879 ( 
.A(n_8177),
.Y(n_9879)
);

CKINVDCx20_ASAP7_75t_R g9880 ( 
.A(n_8162),
.Y(n_9880)
);

INVx1_ASAP7_75t_L g9881 ( 
.A(n_8177),
.Y(n_9881)
);

INVx1_ASAP7_75t_L g9882 ( 
.A(n_8181),
.Y(n_9882)
);

INVx1_ASAP7_75t_L g9883 ( 
.A(n_8181),
.Y(n_9883)
);

INVx2_ASAP7_75t_SL g9884 ( 
.A(n_8414),
.Y(n_9884)
);

BUFx2_ASAP7_75t_L g9885 ( 
.A(n_8878),
.Y(n_9885)
);

INVx1_ASAP7_75t_L g9886 ( 
.A(n_8181),
.Y(n_9886)
);

INVx2_ASAP7_75t_L g9887 ( 
.A(n_8646),
.Y(n_9887)
);

BUFx2_ASAP7_75t_L g9888 ( 
.A(n_8878),
.Y(n_9888)
);

INVx6_ASAP7_75t_L g9889 ( 
.A(n_9044),
.Y(n_9889)
);

BUFx6f_ASAP7_75t_L g9890 ( 
.A(n_8797),
.Y(n_9890)
);

BUFx3_ASAP7_75t_L g9891 ( 
.A(n_9044),
.Y(n_9891)
);

BUFx2_ASAP7_75t_R g9892 ( 
.A(n_8088),
.Y(n_9892)
);

INVx2_ASAP7_75t_L g9893 ( 
.A(n_8646),
.Y(n_9893)
);

INVx2_ASAP7_75t_L g9894 ( 
.A(n_8646),
.Y(n_9894)
);

INVx2_ASAP7_75t_L g9895 ( 
.A(n_8646),
.Y(n_9895)
);

BUFx4f_ASAP7_75t_SL g9896 ( 
.A(n_9312),
.Y(n_9896)
);

INVx2_ASAP7_75t_L g9897 ( 
.A(n_8646),
.Y(n_9897)
);

BUFx10_ASAP7_75t_L g9898 ( 
.A(n_8562),
.Y(n_9898)
);

AOI22xp33_ASAP7_75t_L g9899 ( 
.A1(n_8702),
.A2(n_7327),
.B1(n_7328),
.B2(n_7301),
.Y(n_9899)
);

AOI22xp5_ASAP7_75t_L g9900 ( 
.A1(n_8644),
.A2(n_6958),
.B1(n_7414),
.B2(n_7368),
.Y(n_9900)
);

INVx2_ASAP7_75t_L g9901 ( 
.A(n_8646),
.Y(n_9901)
);

INVx1_ASAP7_75t_SL g9902 ( 
.A(n_9302),
.Y(n_9902)
);

AOI22xp33_ASAP7_75t_L g9903 ( 
.A1(n_8644),
.A2(n_7327),
.B1(n_7328),
.B2(n_7301),
.Y(n_9903)
);

INVx1_ASAP7_75t_L g9904 ( 
.A(n_8186),
.Y(n_9904)
);

INVx2_ASAP7_75t_L g9905 ( 
.A(n_8706),
.Y(n_9905)
);

OAI21x1_ASAP7_75t_L g9906 ( 
.A1(n_7954),
.A2(n_7841),
.B(n_7821),
.Y(n_9906)
);

AOI22xp33_ASAP7_75t_L g9907 ( 
.A1(n_8559),
.A2(n_7328),
.B1(n_7329),
.B2(n_7327),
.Y(n_9907)
);

INVx2_ASAP7_75t_L g9908 ( 
.A(n_8706),
.Y(n_9908)
);

INVx1_ASAP7_75t_L g9909 ( 
.A(n_8186),
.Y(n_9909)
);

INVx2_ASAP7_75t_SL g9910 ( 
.A(n_8420),
.Y(n_9910)
);

INVx2_ASAP7_75t_L g9911 ( 
.A(n_8706),
.Y(n_9911)
);

NOR2x1_ASAP7_75t_SL g9912 ( 
.A(n_8987),
.B(n_6915),
.Y(n_9912)
);

INVx6_ASAP7_75t_L g9913 ( 
.A(n_9044),
.Y(n_9913)
);

INVx1_ASAP7_75t_L g9914 ( 
.A(n_8186),
.Y(n_9914)
);

INVx2_ASAP7_75t_L g9915 ( 
.A(n_8706),
.Y(n_9915)
);

BUFx12f_ASAP7_75t_L g9916 ( 
.A(n_8562),
.Y(n_9916)
);

INVx1_ASAP7_75t_L g9917 ( 
.A(n_8190),
.Y(n_9917)
);

INVx2_ASAP7_75t_L g9918 ( 
.A(n_8706),
.Y(n_9918)
);

BUFx8_ASAP7_75t_L g9919 ( 
.A(n_8420),
.Y(n_9919)
);

BUFx3_ASAP7_75t_L g9920 ( 
.A(n_9044),
.Y(n_9920)
);

AOI22xp33_ASAP7_75t_L g9921 ( 
.A1(n_8559),
.A2(n_7338),
.B1(n_7351),
.B2(n_7329),
.Y(n_9921)
);

BUFx6f_ASAP7_75t_L g9922 ( 
.A(n_8797),
.Y(n_9922)
);

INVx2_ASAP7_75t_L g9923 ( 
.A(n_8706),
.Y(n_9923)
);

INVx1_ASAP7_75t_L g9924 ( 
.A(n_8190),
.Y(n_9924)
);

OAI22xp5_ASAP7_75t_L g9925 ( 
.A1(n_8121),
.A2(n_7347),
.B1(n_7432),
.B2(n_7303),
.Y(n_9925)
);

BUFx2_ASAP7_75t_L g9926 ( 
.A(n_8878),
.Y(n_9926)
);

AO21x2_ASAP7_75t_L g9927 ( 
.A1(n_8012),
.A2(n_7166),
.B(n_6965),
.Y(n_9927)
);

OR2x2_ASAP7_75t_L g9928 ( 
.A(n_7937),
.B(n_7671),
.Y(n_9928)
);

AND2x2_ASAP7_75t_L g9929 ( 
.A(n_8061),
.B(n_7941),
.Y(n_9929)
);

INVx2_ASAP7_75t_L g9930 ( 
.A(n_8789),
.Y(n_9930)
);

AOI22xp33_ASAP7_75t_L g9931 ( 
.A1(n_8478),
.A2(n_7338),
.B1(n_7351),
.B2(n_7329),
.Y(n_9931)
);

NAND2xp5_ASAP7_75t_L g9932 ( 
.A(n_8400),
.B(n_7212),
.Y(n_9932)
);

INVx1_ASAP7_75t_L g9933 ( 
.A(n_8190),
.Y(n_9933)
);

AOI22xp33_ASAP7_75t_L g9934 ( 
.A1(n_8478),
.A2(n_7351),
.B1(n_7352),
.B2(n_7338),
.Y(n_9934)
);

INVx1_ASAP7_75t_SL g9935 ( 
.A(n_9302),
.Y(n_9935)
);

INVx1_ASAP7_75t_L g9936 ( 
.A(n_8193),
.Y(n_9936)
);

INVx1_ASAP7_75t_SL g9937 ( 
.A(n_9169),
.Y(n_9937)
);

AOI22xp33_ASAP7_75t_SL g9938 ( 
.A1(n_8695),
.A2(n_8722),
.B1(n_9118),
.B2(n_8132),
.Y(n_9938)
);

OAI21x1_ASAP7_75t_L g9939 ( 
.A1(n_7954),
.A2(n_7850),
.B(n_7841),
.Y(n_9939)
);

NAND2x1p5_ASAP7_75t_L g9940 ( 
.A(n_7992),
.B(n_7780),
.Y(n_9940)
);

BUFx2_ASAP7_75t_L g9941 ( 
.A(n_8933),
.Y(n_9941)
);

BUFx2_ASAP7_75t_L g9942 ( 
.A(n_8933),
.Y(n_9942)
);

AOI22xp5_ASAP7_75t_SL g9943 ( 
.A1(n_8473),
.A2(n_7829),
.B1(n_7848),
.B2(n_7823),
.Y(n_9943)
);

OAI22xp33_ASAP7_75t_L g9944 ( 
.A1(n_8537),
.A2(n_7013),
.B1(n_7347),
.B2(n_7303),
.Y(n_9944)
);

AOI22xp33_ASAP7_75t_SL g9945 ( 
.A1(n_8722),
.A2(n_9118),
.B1(n_8132),
.B2(n_8416),
.Y(n_9945)
);

INVx1_ASAP7_75t_L g9946 ( 
.A(n_8193),
.Y(n_9946)
);

NAND2xp5_ASAP7_75t_L g9947 ( 
.A(n_8184),
.B(n_7212),
.Y(n_9947)
);

INVx1_ASAP7_75t_L g9948 ( 
.A(n_8193),
.Y(n_9948)
);

AND2x4_ASAP7_75t_L g9949 ( 
.A(n_8152),
.B(n_6930),
.Y(n_9949)
);

INVx1_ASAP7_75t_L g9950 ( 
.A(n_8198),
.Y(n_9950)
);

INVx2_ASAP7_75t_L g9951 ( 
.A(n_8789),
.Y(n_9951)
);

INVx1_ASAP7_75t_L g9952 ( 
.A(n_8198),
.Y(n_9952)
);

OAI22xp5_ASAP7_75t_L g9953 ( 
.A1(n_8121),
.A2(n_7432),
.B1(n_7469),
.B2(n_7347),
.Y(n_9953)
);

INVx2_ASAP7_75t_L g9954 ( 
.A(n_8789),
.Y(n_9954)
);

INVx1_ASAP7_75t_L g9955 ( 
.A(n_8198),
.Y(n_9955)
);

OAI21x1_ASAP7_75t_L g9956 ( 
.A1(n_7954),
.A2(n_7850),
.B(n_7841),
.Y(n_9956)
);

BUFx3_ASAP7_75t_L g9957 ( 
.A(n_9221),
.Y(n_9957)
);

INVx2_ASAP7_75t_L g9958 ( 
.A(n_8789),
.Y(n_9958)
);

NAND2xp5_ASAP7_75t_L g9959 ( 
.A(n_8184),
.B(n_7059),
.Y(n_9959)
);

AND2x2_ASAP7_75t_L g9960 ( 
.A(n_8061),
.B(n_6915),
.Y(n_9960)
);

BUFx10_ASAP7_75t_L g9961 ( 
.A(n_8677),
.Y(n_9961)
);

AND2x2_ASAP7_75t_L g9962 ( 
.A(n_7941),
.B(n_6915),
.Y(n_9962)
);

AO21x1_ASAP7_75t_L g9963 ( 
.A1(n_7922),
.A2(n_7925),
.B(n_7968),
.Y(n_9963)
);

INVx1_ASAP7_75t_L g9964 ( 
.A(n_8199),
.Y(n_9964)
);

AOI22xp33_ASAP7_75t_L g9965 ( 
.A1(n_8343),
.A2(n_7397),
.B1(n_7426),
.B2(n_7352),
.Y(n_9965)
);

AOI22xp33_ASAP7_75t_L g9966 ( 
.A1(n_8343),
.A2(n_8309),
.B1(n_8371),
.B2(n_8363),
.Y(n_9966)
);

INVx1_ASAP7_75t_L g9967 ( 
.A(n_8199),
.Y(n_9967)
);

AND2x2_ASAP7_75t_L g9968 ( 
.A(n_7941),
.B(n_6919),
.Y(n_9968)
);

INVx1_ASAP7_75t_L g9969 ( 
.A(n_8199),
.Y(n_9969)
);

INVx2_ASAP7_75t_L g9970 ( 
.A(n_8789),
.Y(n_9970)
);

INVx3_ASAP7_75t_L g9971 ( 
.A(n_8179),
.Y(n_9971)
);

NAND2xp5_ASAP7_75t_L g9972 ( 
.A(n_8769),
.B(n_7059),
.Y(n_9972)
);

AND2x4_ASAP7_75t_L g9973 ( 
.A(n_8179),
.B(n_6930),
.Y(n_9973)
);

OAI21x1_ASAP7_75t_L g9974 ( 
.A1(n_8081),
.A2(n_8140),
.B(n_8591),
.Y(n_9974)
);

INVx1_ASAP7_75t_L g9975 ( 
.A(n_8200),
.Y(n_9975)
);

INVx1_ASAP7_75t_L g9976 ( 
.A(n_8200),
.Y(n_9976)
);

INVx1_ASAP7_75t_L g9977 ( 
.A(n_8200),
.Y(n_9977)
);

BUFx2_ASAP7_75t_R g9978 ( 
.A(n_8088),
.Y(n_9978)
);

AOI22xp33_ASAP7_75t_L g9979 ( 
.A1(n_8309),
.A2(n_7397),
.B1(n_7426),
.B2(n_7352),
.Y(n_9979)
);

INVx1_ASAP7_75t_SL g9980 ( 
.A(n_9169),
.Y(n_9980)
);

BUFx12f_ASAP7_75t_L g9981 ( 
.A(n_8677),
.Y(n_9981)
);

NOR2xp33_ASAP7_75t_L g9982 ( 
.A(n_7961),
.B(n_8072),
.Y(n_9982)
);

CKINVDCx11_ASAP7_75t_R g9983 ( 
.A(n_8858),
.Y(n_9983)
);

INVx2_ASAP7_75t_L g9984 ( 
.A(n_8789),
.Y(n_9984)
);

INVx1_ASAP7_75t_SL g9985 ( 
.A(n_8298),
.Y(n_9985)
);

INVx1_ASAP7_75t_L g9986 ( 
.A(n_8202),
.Y(n_9986)
);

AOI22xp33_ASAP7_75t_SL g9987 ( 
.A1(n_9118),
.A2(n_7079),
.B1(n_7247),
.B2(n_7246),
.Y(n_9987)
);

INVx1_ASAP7_75t_L g9988 ( 
.A(n_8202),
.Y(n_9988)
);

BUFx6f_ASAP7_75t_L g9989 ( 
.A(n_8797),
.Y(n_9989)
);

INVx1_ASAP7_75t_L g9990 ( 
.A(n_8202),
.Y(n_9990)
);

OAI22xp5_ASAP7_75t_L g9991 ( 
.A1(n_8135),
.A2(n_7432),
.B1(n_7469),
.B2(n_7347),
.Y(n_9991)
);

INVx1_ASAP7_75t_L g9992 ( 
.A(n_8206),
.Y(n_9992)
);

INVx1_ASAP7_75t_L g9993 ( 
.A(n_8206),
.Y(n_9993)
);

INVx2_ASAP7_75t_L g9994 ( 
.A(n_8976),
.Y(n_9994)
);

INVx1_ASAP7_75t_L g9995 ( 
.A(n_8206),
.Y(n_9995)
);

HB1xp67_ASAP7_75t_L g9996 ( 
.A(n_9273),
.Y(n_9996)
);

BUFx2_ASAP7_75t_SL g9997 ( 
.A(n_8851),
.Y(n_9997)
);

BUFx12f_ASAP7_75t_L g9998 ( 
.A(n_8740),
.Y(n_9998)
);

AND2x2_ASAP7_75t_L g9999 ( 
.A(n_7946),
.B(n_6919),
.Y(n_9999)
);

OAI21x1_ASAP7_75t_SL g10000 ( 
.A1(n_8879),
.A2(n_6927),
.B(n_6919),
.Y(n_10000)
);

AOI22xp33_ASAP7_75t_SL g10001 ( 
.A1(n_9118),
.A2(n_8416),
.B1(n_8861),
.B2(n_8871),
.Y(n_10001)
);

CKINVDCx11_ASAP7_75t_R g10002 ( 
.A(n_8858),
.Y(n_10002)
);

INVx2_ASAP7_75t_L g10003 ( 
.A(n_8976),
.Y(n_10003)
);

HB1xp67_ASAP7_75t_L g10004 ( 
.A(n_7979),
.Y(n_10004)
);

BUFx3_ASAP7_75t_L g10005 ( 
.A(n_9221),
.Y(n_10005)
);

HB1xp67_ASAP7_75t_L g10006 ( 
.A(n_7979),
.Y(n_10006)
);

INVx2_ASAP7_75t_L g10007 ( 
.A(n_8976),
.Y(n_10007)
);

OR2x6_ASAP7_75t_L g10008 ( 
.A(n_8837),
.B(n_7109),
.Y(n_10008)
);

OAI21xp5_ASAP7_75t_L g10009 ( 
.A1(n_8406),
.A2(n_7267),
.B(n_7368),
.Y(n_10009)
);

INVx2_ASAP7_75t_L g10010 ( 
.A(n_8983),
.Y(n_10010)
);

OR2x2_ASAP7_75t_L g10011 ( 
.A(n_8484),
.B(n_7702),
.Y(n_10011)
);

INVx1_ASAP7_75t_L g10012 ( 
.A(n_8236),
.Y(n_10012)
);

INVx8_ASAP7_75t_L g10013 ( 
.A(n_9278),
.Y(n_10013)
);

INVx1_ASAP7_75t_L g10014 ( 
.A(n_8236),
.Y(n_10014)
);

OAI21x1_ASAP7_75t_L g10015 ( 
.A1(n_8081),
.A2(n_7862),
.B(n_7850),
.Y(n_10015)
);

INVx3_ASAP7_75t_L g10016 ( 
.A(n_8179),
.Y(n_10016)
);

INVx2_ASAP7_75t_L g10017 ( 
.A(n_8983),
.Y(n_10017)
);

AND2x2_ASAP7_75t_L g10018 ( 
.A(n_7946),
.B(n_6927),
.Y(n_10018)
);

AOI22xp33_ASAP7_75t_L g10019 ( 
.A1(n_8363),
.A2(n_7426),
.B1(n_7435),
.B2(n_7397),
.Y(n_10019)
);

INVx2_ASAP7_75t_L g10020 ( 
.A(n_8983),
.Y(n_10020)
);

INVx2_ASAP7_75t_L g10021 ( 
.A(n_9006),
.Y(n_10021)
);

HB1xp67_ASAP7_75t_L g10022 ( 
.A(n_8016),
.Y(n_10022)
);

BUFx2_ASAP7_75t_L g10023 ( 
.A(n_8933),
.Y(n_10023)
);

INVx2_ASAP7_75t_L g10024 ( 
.A(n_9006),
.Y(n_10024)
);

NAND2xp5_ASAP7_75t_L g10025 ( 
.A(n_8769),
.B(n_7702),
.Y(n_10025)
);

BUFx8_ASAP7_75t_L g10026 ( 
.A(n_8420),
.Y(n_10026)
);

HB1xp67_ASAP7_75t_L g10027 ( 
.A(n_8016),
.Y(n_10027)
);

BUFx2_ASAP7_75t_L g10028 ( 
.A(n_8933),
.Y(n_10028)
);

INVx1_ASAP7_75t_L g10029 ( 
.A(n_8236),
.Y(n_10029)
);

INVx1_ASAP7_75t_L g10030 ( 
.A(n_8239),
.Y(n_10030)
);

AOI22xp33_ASAP7_75t_L g10031 ( 
.A1(n_8371),
.A2(n_7450),
.B1(n_7452),
.B2(n_7435),
.Y(n_10031)
);

BUFx2_ASAP7_75t_L g10032 ( 
.A(n_8933),
.Y(n_10032)
);

CKINVDCx14_ASAP7_75t_R g10033 ( 
.A(n_8602),
.Y(n_10033)
);

CKINVDCx5p33_ASAP7_75t_R g10034 ( 
.A(n_8162),
.Y(n_10034)
);

NOR2xp33_ASAP7_75t_L g10035 ( 
.A(n_7961),
.B(n_7048),
.Y(n_10035)
);

INVx1_ASAP7_75t_L g10036 ( 
.A(n_8239),
.Y(n_10036)
);

OR2x2_ASAP7_75t_L g10037 ( 
.A(n_8484),
.B(n_7702),
.Y(n_10037)
);

BUFx2_ASAP7_75t_L g10038 ( 
.A(n_8933),
.Y(n_10038)
);

CKINVDCx5p33_ASAP7_75t_R g10039 ( 
.A(n_8194),
.Y(n_10039)
);

NOR2xp33_ASAP7_75t_L g10040 ( 
.A(n_7961),
.B(n_7451),
.Y(n_10040)
);

INVx1_ASAP7_75t_L g10041 ( 
.A(n_8239),
.Y(n_10041)
);

BUFx6f_ASAP7_75t_L g10042 ( 
.A(n_8420),
.Y(n_10042)
);

AOI22xp33_ASAP7_75t_L g10043 ( 
.A1(n_8595),
.A2(n_8479),
.B1(n_8861),
.B2(n_9089),
.Y(n_10043)
);

INVx1_ASAP7_75t_L g10044 ( 
.A(n_8248),
.Y(n_10044)
);

AOI21x1_ASAP7_75t_L g10045 ( 
.A1(n_8228),
.A2(n_8057),
.B(n_8271),
.Y(n_10045)
);

AND2x2_ASAP7_75t_L g10046 ( 
.A(n_7946),
.B(n_6927),
.Y(n_10046)
);

AOI22xp33_ASAP7_75t_L g10047 ( 
.A1(n_8595),
.A2(n_7450),
.B1(n_7452),
.B2(n_7435),
.Y(n_10047)
);

INVx4_ASAP7_75t_L g10048 ( 
.A(n_7961),
.Y(n_10048)
);

OA21x2_ASAP7_75t_L g10049 ( 
.A1(n_8081),
.A2(n_7112),
.B(n_7108),
.Y(n_10049)
);

BUFx3_ASAP7_75t_L g10050 ( 
.A(n_9221),
.Y(n_10050)
);

INVx1_ASAP7_75t_L g10051 ( 
.A(n_8248),
.Y(n_10051)
);

NAND2xp5_ASAP7_75t_L g10052 ( 
.A(n_8822),
.B(n_7723),
.Y(n_10052)
);

INVx4_ASAP7_75t_L g10053 ( 
.A(n_8072),
.Y(n_10053)
);

BUFx8_ASAP7_75t_SL g10054 ( 
.A(n_8740),
.Y(n_10054)
);

INVx1_ASAP7_75t_L g10055 ( 
.A(n_8248),
.Y(n_10055)
);

AOI21xp5_ASAP7_75t_L g10056 ( 
.A1(n_8195),
.A2(n_6966),
.B(n_7622),
.Y(n_10056)
);

AOI21x1_ASAP7_75t_L g10057 ( 
.A1(n_8228),
.A2(n_7184),
.B(n_7159),
.Y(n_10057)
);

INVx2_ASAP7_75t_L g10058 ( 
.A(n_9006),
.Y(n_10058)
);

AO21x2_ASAP7_75t_L g10059 ( 
.A1(n_8012),
.A2(n_7166),
.B(n_6965),
.Y(n_10059)
);

BUFx2_ASAP7_75t_R g10060 ( 
.A(n_8298),
.Y(n_10060)
);

BUFx2_ASAP7_75t_L g10061 ( 
.A(n_8933),
.Y(n_10061)
);

INVx1_ASAP7_75t_L g10062 ( 
.A(n_8249),
.Y(n_10062)
);

NAND2xp5_ASAP7_75t_L g10063 ( 
.A(n_8822),
.B(n_7723),
.Y(n_10063)
);

AOI21x1_ASAP7_75t_L g10064 ( 
.A1(n_8057),
.A2(n_7184),
.B(n_7159),
.Y(n_10064)
);

BUFx2_ASAP7_75t_SL g10065 ( 
.A(n_8851),
.Y(n_10065)
);

OAI21xp5_ASAP7_75t_SL g10066 ( 
.A1(n_8406),
.A2(n_7656),
.B(n_6998),
.Y(n_10066)
);

AO21x1_ASAP7_75t_L g10067 ( 
.A1(n_7922),
.A2(n_8234),
.B(n_8284),
.Y(n_10067)
);

BUFx2_ASAP7_75t_SL g10068 ( 
.A(n_8851),
.Y(n_10068)
);

INVx1_ASAP7_75t_L g10069 ( 
.A(n_8249),
.Y(n_10069)
);

INVx6_ASAP7_75t_L g10070 ( 
.A(n_9221),
.Y(n_10070)
);

OAI22xp5_ASAP7_75t_L g10071 ( 
.A1(n_8135),
.A2(n_7469),
.B1(n_7432),
.B2(n_6998),
.Y(n_10071)
);

INVx2_ASAP7_75t_L g10072 ( 
.A(n_9009),
.Y(n_10072)
);

INVx1_ASAP7_75t_SL g10073 ( 
.A(n_9017),
.Y(n_10073)
);

AOI22xp33_ASAP7_75t_L g10074 ( 
.A1(n_8479),
.A2(n_7452),
.B1(n_7466),
.B2(n_7450),
.Y(n_10074)
);

INVx3_ASAP7_75t_L g10075 ( 
.A(n_8179),
.Y(n_10075)
);

INVx2_ASAP7_75t_SL g10076 ( 
.A(n_8425),
.Y(n_10076)
);

INVx2_ASAP7_75t_L g10077 ( 
.A(n_9009),
.Y(n_10077)
);

AOI22xp33_ASAP7_75t_L g10078 ( 
.A1(n_9089),
.A2(n_7468),
.B1(n_7486),
.B2(n_7466),
.Y(n_10078)
);

INVx1_ASAP7_75t_L g10079 ( 
.A(n_8249),
.Y(n_10079)
);

NAND2xp5_ASAP7_75t_L g10080 ( 
.A(n_8928),
.B(n_7723),
.Y(n_10080)
);

INVx2_ASAP7_75t_L g10081 ( 
.A(n_9009),
.Y(n_10081)
);

INVx3_ASAP7_75t_L g10082 ( 
.A(n_8227),
.Y(n_10082)
);

INVx2_ASAP7_75t_L g10083 ( 
.A(n_9011),
.Y(n_10083)
);

INVx2_ASAP7_75t_L g10084 ( 
.A(n_9011),
.Y(n_10084)
);

INVx1_ASAP7_75t_L g10085 ( 
.A(n_8257),
.Y(n_10085)
);

INVx1_ASAP7_75t_L g10086 ( 
.A(n_8257),
.Y(n_10086)
);

OAI22xp5_ASAP7_75t_L g10087 ( 
.A1(n_8005),
.A2(n_7469),
.B1(n_7656),
.B2(n_6939),
.Y(n_10087)
);

INVx2_ASAP7_75t_L g10088 ( 
.A(n_9011),
.Y(n_10088)
);

AOI22xp33_ASAP7_75t_SL g10089 ( 
.A1(n_8871),
.A2(n_7246),
.B1(n_7381),
.B2(n_7247),
.Y(n_10089)
);

AOI22xp33_ASAP7_75t_L g10090 ( 
.A1(n_8005),
.A2(n_7468),
.B1(n_7486),
.B2(n_7466),
.Y(n_10090)
);

INVx1_ASAP7_75t_L g10091 ( 
.A(n_8257),
.Y(n_10091)
);

AOI22xp5_ASAP7_75t_L g10092 ( 
.A1(n_7913),
.A2(n_8156),
.B1(n_8161),
.B2(n_8331),
.Y(n_10092)
);

AOI21x1_ASAP7_75t_L g10093 ( 
.A1(n_8057),
.A2(n_7184),
.B(n_7159),
.Y(n_10093)
);

NAND2xp5_ASAP7_75t_L g10094 ( 
.A(n_8928),
.B(n_7729),
.Y(n_10094)
);

OR2x2_ASAP7_75t_L g10095 ( 
.A(n_8491),
.B(n_7729),
.Y(n_10095)
);

INVx2_ASAP7_75t_L g10096 ( 
.A(n_9018),
.Y(n_10096)
);

NAND2x1p5_ASAP7_75t_L g10097 ( 
.A(n_7992),
.B(n_7780),
.Y(n_10097)
);

NAND2xp5_ASAP7_75t_L g10098 ( 
.A(n_7915),
.B(n_7729),
.Y(n_10098)
);

OR2x2_ASAP7_75t_L g10099 ( 
.A(n_8491),
.B(n_7772),
.Y(n_10099)
);

AND2x4_ASAP7_75t_L g10100 ( 
.A(n_8227),
.B(n_6930),
.Y(n_10100)
);

INVx1_ASAP7_75t_L g10101 ( 
.A(n_8261),
.Y(n_10101)
);

AND2x4_ASAP7_75t_L g10102 ( 
.A(n_8227),
.B(n_7112),
.Y(n_10102)
);

INVx1_ASAP7_75t_L g10103 ( 
.A(n_8261),
.Y(n_10103)
);

INVx6_ASAP7_75t_L g10104 ( 
.A(n_9221),
.Y(n_10104)
);

OAI21x1_ASAP7_75t_L g10105 ( 
.A1(n_8140),
.A2(n_7862),
.B(n_7850),
.Y(n_10105)
);

AOI22xp33_ASAP7_75t_L g10106 ( 
.A1(n_7960),
.A2(n_7486),
.B1(n_7492),
.B2(n_7468),
.Y(n_10106)
);

INVx1_ASAP7_75t_L g10107 ( 
.A(n_8261),
.Y(n_10107)
);

AND2x4_ASAP7_75t_L g10108 ( 
.A(n_8227),
.B(n_7117),
.Y(n_10108)
);

AOI21xp5_ASAP7_75t_L g10109 ( 
.A1(n_8307),
.A2(n_6966),
.B(n_7622),
.Y(n_10109)
);

INVx1_ASAP7_75t_L g10110 ( 
.A(n_8279),
.Y(n_10110)
);

AND2x4_ASAP7_75t_L g10111 ( 
.A(n_8277),
.B(n_7117),
.Y(n_10111)
);

INVx1_ASAP7_75t_L g10112 ( 
.A(n_8279),
.Y(n_10112)
);

NAND2xp5_ASAP7_75t_L g10113 ( 
.A(n_7915),
.B(n_7772),
.Y(n_10113)
);

AND2x2_ASAP7_75t_L g10114 ( 
.A(n_7966),
.B(n_6927),
.Y(n_10114)
);

OAI21x1_ASAP7_75t_SL g10115 ( 
.A1(n_8879),
.A2(n_6935),
.B(n_6933),
.Y(n_10115)
);

OAI221xp5_ASAP7_75t_L g10116 ( 
.A1(n_7909),
.A2(n_7160),
.B1(n_7163),
.B2(n_7157),
.C(n_7117),
.Y(n_10116)
);

INVx1_ASAP7_75t_L g10117 ( 
.A(n_8279),
.Y(n_10117)
);

INVx1_ASAP7_75t_L g10118 ( 
.A(n_8292),
.Y(n_10118)
);

OAI22xp5_ASAP7_75t_L g10119 ( 
.A1(n_8943),
.A2(n_6939),
.B1(n_7013),
.B2(n_7313),
.Y(n_10119)
);

OAI21x1_ASAP7_75t_L g10120 ( 
.A1(n_8140),
.A2(n_8591),
.B(n_7908),
.Y(n_10120)
);

NAND2xp5_ASAP7_75t_L g10121 ( 
.A(n_8812),
.B(n_7772),
.Y(n_10121)
);

AND2x2_ASAP7_75t_L g10122 ( 
.A(n_7966),
.B(n_6933),
.Y(n_10122)
);

INVx3_ASAP7_75t_L g10123 ( 
.A(n_8277),
.Y(n_10123)
);

HB1xp67_ASAP7_75t_L g10124 ( 
.A(n_8064),
.Y(n_10124)
);

OAI21x1_ASAP7_75t_L g10125 ( 
.A1(n_8591),
.A2(n_7862),
.B(n_7850),
.Y(n_10125)
);

BUFx2_ASAP7_75t_L g10126 ( 
.A(n_8933),
.Y(n_10126)
);

INVx2_ASAP7_75t_L g10127 ( 
.A(n_9018),
.Y(n_10127)
);

INVx2_ASAP7_75t_L g10128 ( 
.A(n_9018),
.Y(n_10128)
);

AND2x4_ASAP7_75t_L g10129 ( 
.A(n_8277),
.B(n_7157),
.Y(n_10129)
);

BUFx6f_ASAP7_75t_L g10130 ( 
.A(n_8425),
.Y(n_10130)
);

INVx1_ASAP7_75t_L g10131 ( 
.A(n_8292),
.Y(n_10131)
);

INVx1_ASAP7_75t_L g10132 ( 
.A(n_8292),
.Y(n_10132)
);

INVx2_ASAP7_75t_L g10133 ( 
.A(n_8757),
.Y(n_10133)
);

OAI21xp5_ASAP7_75t_L g10134 ( 
.A1(n_8008),
.A2(n_7558),
.B(n_7523),
.Y(n_10134)
);

OAI22xp5_ASAP7_75t_L g10135 ( 
.A1(n_8943),
.A2(n_7313),
.B1(n_7471),
.B2(n_7447),
.Y(n_10135)
);

OAI21x1_ASAP7_75t_L g10136 ( 
.A1(n_7908),
.A2(n_7862),
.B(n_7850),
.Y(n_10136)
);

AOI22xp33_ASAP7_75t_L g10137 ( 
.A1(n_7960),
.A2(n_7499),
.B1(n_7502),
.B2(n_7492),
.Y(n_10137)
);

BUFx8_ASAP7_75t_L g10138 ( 
.A(n_8425),
.Y(n_10138)
);

AOI22xp33_ASAP7_75t_L g10139 ( 
.A1(n_7976),
.A2(n_7499),
.B1(n_7502),
.B2(n_7492),
.Y(n_10139)
);

NAND2xp5_ASAP7_75t_L g10140 ( 
.A(n_8812),
.B(n_7828),
.Y(n_10140)
);

OAI21x1_ASAP7_75t_L g10141 ( 
.A1(n_7908),
.A2(n_7880),
.B(n_7862),
.Y(n_10141)
);

INVx4_ASAP7_75t_L g10142 ( 
.A(n_8072),
.Y(n_10142)
);

INVx1_ASAP7_75t_L g10143 ( 
.A(n_8294),
.Y(n_10143)
);

INVx2_ASAP7_75t_L g10144 ( 
.A(n_8757),
.Y(n_10144)
);

AND2x4_ASAP7_75t_L g10145 ( 
.A(n_8277),
.B(n_8395),
.Y(n_10145)
);

INVx1_ASAP7_75t_L g10146 ( 
.A(n_8294),
.Y(n_10146)
);

INVx6_ASAP7_75t_L g10147 ( 
.A(n_9221),
.Y(n_10147)
);

OAI22xp5_ASAP7_75t_L g10148 ( 
.A1(n_8446),
.A2(n_7471),
.B1(n_7447),
.B2(n_7576),
.Y(n_10148)
);

INVx1_ASAP7_75t_L g10149 ( 
.A(n_8294),
.Y(n_10149)
);

BUFx2_ASAP7_75t_L g10150 ( 
.A(n_8933),
.Y(n_10150)
);

INVx1_ASAP7_75t_L g10151 ( 
.A(n_8305),
.Y(n_10151)
);

INVx4_ASAP7_75t_L g10152 ( 
.A(n_8072),
.Y(n_10152)
);

INVx2_ASAP7_75t_L g10153 ( 
.A(n_8757),
.Y(n_10153)
);

INVx1_ASAP7_75t_L g10154 ( 
.A(n_8305),
.Y(n_10154)
);

AOI22xp5_ASAP7_75t_L g10155 ( 
.A1(n_7913),
.A2(n_7414),
.B1(n_7017),
.B2(n_7485),
.Y(n_10155)
);

AO21x1_ASAP7_75t_SL g10156 ( 
.A1(n_8284),
.A2(n_7513),
.B(n_7505),
.Y(n_10156)
);

NAND2xp5_ASAP7_75t_SL g10157 ( 
.A(n_8378),
.B(n_7823),
.Y(n_10157)
);

INVx1_ASAP7_75t_L g10158 ( 
.A(n_8305),
.Y(n_10158)
);

AOI22xp5_ASAP7_75t_SL g10159 ( 
.A1(n_8473),
.A2(n_7848),
.B1(n_7876),
.B2(n_7829),
.Y(n_10159)
);

AOI22xp33_ASAP7_75t_L g10160 ( 
.A1(n_7976),
.A2(n_7502),
.B1(n_7536),
.B2(n_7499),
.Y(n_10160)
);

BUFx8_ASAP7_75t_L g10161 ( 
.A(n_8425),
.Y(n_10161)
);

OAI22xp5_ASAP7_75t_L g10162 ( 
.A1(n_8446),
.A2(n_7471),
.B1(n_7596),
.B2(n_7576),
.Y(n_10162)
);

OAI21x1_ASAP7_75t_L g10163 ( 
.A1(n_7908),
.A2(n_7880),
.B(n_7862),
.Y(n_10163)
);

AOI22xp5_ASAP7_75t_L g10164 ( 
.A1(n_8156),
.A2(n_7485),
.B1(n_7732),
.B2(n_7877),
.Y(n_10164)
);

OAI21x1_ASAP7_75t_L g10165 ( 
.A1(n_8819),
.A2(n_7884),
.B(n_7880),
.Y(n_10165)
);

INVx1_ASAP7_75t_L g10166 ( 
.A(n_8306),
.Y(n_10166)
);

OAI22xp5_ASAP7_75t_SL g10167 ( 
.A1(n_8194),
.A2(n_7304),
.B1(n_7360),
.B2(n_7314),
.Y(n_10167)
);

INVx1_ASAP7_75t_L g10168 ( 
.A(n_8306),
.Y(n_10168)
);

NAND2x1p5_ASAP7_75t_L g10169 ( 
.A(n_7992),
.B(n_7780),
.Y(n_10169)
);

INVx2_ASAP7_75t_L g10170 ( 
.A(n_8757),
.Y(n_10170)
);

INVx1_ASAP7_75t_L g10171 ( 
.A(n_8306),
.Y(n_10171)
);

CKINVDCx11_ASAP7_75t_R g10172 ( 
.A(n_9017),
.Y(n_10172)
);

INVx1_ASAP7_75t_L g10173 ( 
.A(n_8310),
.Y(n_10173)
);

NAND2x1p5_ASAP7_75t_L g10174 ( 
.A(n_7992),
.B(n_7780),
.Y(n_10174)
);

INVx4_ASAP7_75t_L g10175 ( 
.A(n_8072),
.Y(n_10175)
);

BUFx2_ASAP7_75t_SL g10176 ( 
.A(n_9312),
.Y(n_10176)
);

NAND2x1p5_ASAP7_75t_L g10177 ( 
.A(n_8115),
.B(n_7780),
.Y(n_10177)
);

INVx1_ASAP7_75t_L g10178 ( 
.A(n_8310),
.Y(n_10178)
);

NAND2xp5_ASAP7_75t_L g10179 ( 
.A(n_8815),
.B(n_7828),
.Y(n_10179)
);

INVx2_ASAP7_75t_L g10180 ( 
.A(n_8757),
.Y(n_10180)
);

INVx1_ASAP7_75t_L g10181 ( 
.A(n_8310),
.Y(n_10181)
);

INVx3_ASAP7_75t_L g10182 ( 
.A(n_8395),
.Y(n_10182)
);

AO21x2_ASAP7_75t_L g10183 ( 
.A1(n_8137),
.A2(n_7317),
.B(n_7264),
.Y(n_10183)
);

AOI22xp33_ASAP7_75t_L g10184 ( 
.A1(n_8130),
.A2(n_7551),
.B1(n_7556),
.B2(n_7536),
.Y(n_10184)
);

OAI22xp33_ASAP7_75t_L g10185 ( 
.A1(n_8587),
.A2(n_7461),
.B1(n_7562),
.B2(n_7293),
.Y(n_10185)
);

AOI22xp33_ASAP7_75t_L g10186 ( 
.A1(n_8130),
.A2(n_7551),
.B1(n_7556),
.B2(n_7536),
.Y(n_10186)
);

AOI22xp33_ASAP7_75t_L g10187 ( 
.A1(n_8876),
.A2(n_7556),
.B1(n_7565),
.B2(n_7551),
.Y(n_10187)
);

AOI21xp5_ASAP7_75t_L g10188 ( 
.A1(n_8037),
.A2(n_7622),
.B(n_7694),
.Y(n_10188)
);

BUFx3_ASAP7_75t_L g10189 ( 
.A(n_8428),
.Y(n_10189)
);

INVx1_ASAP7_75t_L g10190 ( 
.A(n_8312),
.Y(n_10190)
);

INVx1_ASAP7_75t_L g10191 ( 
.A(n_8312),
.Y(n_10191)
);

BUFx2_ASAP7_75t_SL g10192 ( 
.A(n_8428),
.Y(n_10192)
);

AOI21x1_ASAP7_75t_L g10193 ( 
.A1(n_8271),
.A2(n_7192),
.B(n_7184),
.Y(n_10193)
);

NAND2xp5_ASAP7_75t_SL g10194 ( 
.A(n_8378),
.B(n_8635),
.Y(n_10194)
);

AND2x2_ASAP7_75t_L g10195 ( 
.A(n_7966),
.B(n_6933),
.Y(n_10195)
);

CKINVDCx20_ASAP7_75t_R g10196 ( 
.A(n_8318),
.Y(n_10196)
);

INVx1_ASAP7_75t_SL g10197 ( 
.A(n_8318),
.Y(n_10197)
);

INVx1_ASAP7_75t_L g10198 ( 
.A(n_8312),
.Y(n_10198)
);

AOI22xp33_ASAP7_75t_L g10199 ( 
.A1(n_8876),
.A2(n_7591),
.B1(n_7609),
.B2(n_7565),
.Y(n_10199)
);

INVx2_ASAP7_75t_L g10200 ( 
.A(n_8857),
.Y(n_10200)
);

BUFx2_ASAP7_75t_L g10201 ( 
.A(n_8961),
.Y(n_10201)
);

OAI22xp33_ASAP7_75t_SL g10202 ( 
.A1(n_8197),
.A2(n_7461),
.B1(n_7562),
.B2(n_7293),
.Y(n_10202)
);

INVx11_ASAP7_75t_L g10203 ( 
.A(n_8602),
.Y(n_10203)
);

OAI21x1_ASAP7_75t_L g10204 ( 
.A1(n_8819),
.A2(n_7884),
.B(n_7880),
.Y(n_10204)
);

AOI22xp33_ASAP7_75t_L g10205 ( 
.A1(n_8197),
.A2(n_7591),
.B1(n_7609),
.B2(n_7565),
.Y(n_10205)
);

OAI22xp5_ASAP7_75t_L g10206 ( 
.A1(n_8222),
.A2(n_7596),
.B1(n_7610),
.B2(n_7576),
.Y(n_10206)
);

CKINVDCx11_ASAP7_75t_R g10207 ( 
.A(n_8367),
.Y(n_10207)
);

INVx1_ASAP7_75t_L g10208 ( 
.A(n_8321),
.Y(n_10208)
);

AOI22xp33_ASAP7_75t_L g10209 ( 
.A1(n_8583),
.A2(n_7609),
.B1(n_7611),
.B2(n_7591),
.Y(n_10209)
);

BUFx6f_ASAP7_75t_L g10210 ( 
.A(n_8428),
.Y(n_10210)
);

INVx2_ASAP7_75t_L g10211 ( 
.A(n_8857),
.Y(n_10211)
);

AND2x2_ASAP7_75t_L g10212 ( 
.A(n_7981),
.B(n_6933),
.Y(n_10212)
);

AOI21x1_ASAP7_75t_L g10213 ( 
.A1(n_8271),
.A2(n_7215),
.B(n_7192),
.Y(n_10213)
);

INVx2_ASAP7_75t_L g10214 ( 
.A(n_8857),
.Y(n_10214)
);

HB1xp67_ASAP7_75t_L g10215 ( 
.A(n_8064),
.Y(n_10215)
);

INVx2_ASAP7_75t_L g10216 ( 
.A(n_8857),
.Y(n_10216)
);

INVx1_ASAP7_75t_L g10217 ( 
.A(n_8321),
.Y(n_10217)
);

OAI21x1_ASAP7_75t_SL g10218 ( 
.A1(n_8879),
.A2(n_6974),
.B(n_6935),
.Y(n_10218)
);

HB1xp67_ASAP7_75t_L g10219 ( 
.A(n_8106),
.Y(n_10219)
);

INVx2_ASAP7_75t_L g10220 ( 
.A(n_8857),
.Y(n_10220)
);

INVx3_ASAP7_75t_L g10221 ( 
.A(n_8395),
.Y(n_10221)
);

BUFx10_ASAP7_75t_L g10222 ( 
.A(n_9266),
.Y(n_10222)
);

AOI22xp33_ASAP7_75t_L g10223 ( 
.A1(n_8583),
.A2(n_7614),
.B1(n_7661),
.B2(n_7611),
.Y(n_10223)
);

NAND2xp5_ASAP7_75t_L g10224 ( 
.A(n_8815),
.B(n_7828),
.Y(n_10224)
);

NAND2xp5_ASAP7_75t_L g10225 ( 
.A(n_8986),
.B(n_6912),
.Y(n_10225)
);

AND2x4_ASAP7_75t_L g10226 ( 
.A(n_8395),
.B(n_7157),
.Y(n_10226)
);

HB1xp67_ASAP7_75t_SL g10227 ( 
.A(n_9266),
.Y(n_10227)
);

INVx2_ASAP7_75t_L g10228 ( 
.A(n_8857),
.Y(n_10228)
);

INVx2_ASAP7_75t_L g10229 ( 
.A(n_8915),
.Y(n_10229)
);

INVx1_ASAP7_75t_SL g10230 ( 
.A(n_8367),
.Y(n_10230)
);

NAND2xp5_ASAP7_75t_L g10231 ( 
.A(n_8986),
.B(n_6912),
.Y(n_10231)
);

INVx1_ASAP7_75t_L g10232 ( 
.A(n_8321),
.Y(n_10232)
);

CKINVDCx11_ASAP7_75t_R g10233 ( 
.A(n_8380),
.Y(n_10233)
);

HB1xp67_ASAP7_75t_L g10234 ( 
.A(n_8106),
.Y(n_10234)
);

INVx1_ASAP7_75t_L g10235 ( 
.A(n_8326),
.Y(n_10235)
);

AND2x4_ASAP7_75t_L g10236 ( 
.A(n_8402),
.B(n_7160),
.Y(n_10236)
);

HB1xp67_ASAP7_75t_L g10237 ( 
.A(n_8176),
.Y(n_10237)
);

INVx4_ASAP7_75t_L g10238 ( 
.A(n_8072),
.Y(n_10238)
);

OR2x6_ASAP7_75t_L g10239 ( 
.A(n_8086),
.B(n_7109),
.Y(n_10239)
);

OAI21xp5_ASAP7_75t_L g10240 ( 
.A1(n_8008),
.A2(n_7558),
.B(n_7523),
.Y(n_10240)
);

INVx2_ASAP7_75t_L g10241 ( 
.A(n_8915),
.Y(n_10241)
);

AND2x2_ASAP7_75t_L g10242 ( 
.A(n_7981),
.B(n_6935),
.Y(n_10242)
);

INVx5_ASAP7_75t_L g10243 ( 
.A(n_7926),
.Y(n_10243)
);

BUFx8_ASAP7_75t_L g10244 ( 
.A(n_8428),
.Y(n_10244)
);

INVx1_ASAP7_75t_L g10245 ( 
.A(n_8326),
.Y(n_10245)
);

INVx1_ASAP7_75t_L g10246 ( 
.A(n_8326),
.Y(n_10246)
);

AOI21x1_ASAP7_75t_L g10247 ( 
.A1(n_7951),
.A2(n_7215),
.B(n_7192),
.Y(n_10247)
);

NAND2xp5_ASAP7_75t_L g10248 ( 
.A(n_8618),
.B(n_6912),
.Y(n_10248)
);

INVx4_ASAP7_75t_L g10249 ( 
.A(n_8274),
.Y(n_10249)
);

AND2x2_ASAP7_75t_L g10250 ( 
.A(n_7981),
.B(n_6935),
.Y(n_10250)
);

INVx2_ASAP7_75t_L g10251 ( 
.A(n_8915),
.Y(n_10251)
);

BUFx2_ASAP7_75t_L g10252 ( 
.A(n_8961),
.Y(n_10252)
);

CKINVDCx5p33_ASAP7_75t_R g10253 ( 
.A(n_8380),
.Y(n_10253)
);

INVx2_ASAP7_75t_L g10254 ( 
.A(n_8915),
.Y(n_10254)
);

AOI21x1_ASAP7_75t_L g10255 ( 
.A1(n_7951),
.A2(n_7215),
.B(n_7192),
.Y(n_10255)
);

INVx1_ASAP7_75t_L g10256 ( 
.A(n_8335),
.Y(n_10256)
);

AND2x4_ASAP7_75t_L g10257 ( 
.A(n_8402),
.B(n_7160),
.Y(n_10257)
);

INVx2_ASAP7_75t_L g10258 ( 
.A(n_8915),
.Y(n_10258)
);

INVx2_ASAP7_75t_L g10259 ( 
.A(n_8915),
.Y(n_10259)
);

INVx1_ASAP7_75t_L g10260 ( 
.A(n_8335),
.Y(n_10260)
);

BUFx2_ASAP7_75t_L g10261 ( 
.A(n_8364),
.Y(n_10261)
);

HB1xp67_ASAP7_75t_L g10262 ( 
.A(n_8176),
.Y(n_10262)
);

NAND2xp5_ASAP7_75t_L g10263 ( 
.A(n_8544),
.B(n_6912),
.Y(n_10263)
);

INVx3_ASAP7_75t_L g10264 ( 
.A(n_8402),
.Y(n_10264)
);

OA21x2_ASAP7_75t_L g10265 ( 
.A1(n_9016),
.A2(n_8924),
.B(n_8344),
.Y(n_10265)
);

INVx1_ASAP7_75t_L g10266 ( 
.A(n_8335),
.Y(n_10266)
);

INVx1_ASAP7_75t_L g10267 ( 
.A(n_8341),
.Y(n_10267)
);

AND2x2_ASAP7_75t_L g10268 ( 
.A(n_7985),
.B(n_6974),
.Y(n_10268)
);

INVx2_ASAP7_75t_L g10269 ( 
.A(n_8919),
.Y(n_10269)
);

NAND2xp5_ASAP7_75t_L g10270 ( 
.A(n_8544),
.B(n_6936),
.Y(n_10270)
);

NAND2x1p5_ASAP7_75t_L g10271 ( 
.A(n_8115),
.B(n_7780),
.Y(n_10271)
);

OAI22xp5_ASAP7_75t_L g10272 ( 
.A1(n_8222),
.A2(n_7596),
.B1(n_7610),
.B2(n_7576),
.Y(n_10272)
);

CKINVDCx11_ASAP7_75t_R g10273 ( 
.A(n_8390),
.Y(n_10273)
);

AOI22xp5_ASAP7_75t_L g10274 ( 
.A1(n_8331),
.A2(n_7732),
.B1(n_7759),
.B2(n_7753),
.Y(n_10274)
);

INVx1_ASAP7_75t_SL g10275 ( 
.A(n_8390),
.Y(n_10275)
);

INVx1_ASAP7_75t_L g10276 ( 
.A(n_8341),
.Y(n_10276)
);

INVx1_ASAP7_75t_L g10277 ( 
.A(n_8341),
.Y(n_10277)
);

AO21x1_ASAP7_75t_L g10278 ( 
.A1(n_8234),
.A2(n_7869),
.B(n_7856),
.Y(n_10278)
);

INVx1_ASAP7_75t_L g10279 ( 
.A(n_8346),
.Y(n_10279)
);

INVx1_ASAP7_75t_L g10280 ( 
.A(n_8346),
.Y(n_10280)
);

AOI22xp33_ASAP7_75t_L g10281 ( 
.A1(n_8583),
.A2(n_7614),
.B1(n_7661),
.B2(n_7611),
.Y(n_10281)
);

INVx1_ASAP7_75t_L g10282 ( 
.A(n_8346),
.Y(n_10282)
);

INVx1_ASAP7_75t_L g10283 ( 
.A(n_8348),
.Y(n_10283)
);

INVx1_ASAP7_75t_L g10284 ( 
.A(n_8348),
.Y(n_10284)
);

INVx1_ASAP7_75t_L g10285 ( 
.A(n_8348),
.Y(n_10285)
);

INVx1_ASAP7_75t_L g10286 ( 
.A(n_8356),
.Y(n_10286)
);

NAND2xp5_ASAP7_75t_SL g10287 ( 
.A(n_8635),
.B(n_7876),
.Y(n_10287)
);

AOI22xp33_ASAP7_75t_L g10288 ( 
.A1(n_8583),
.A2(n_7661),
.B1(n_7695),
.B2(n_7614),
.Y(n_10288)
);

INVx3_ASAP7_75t_L g10289 ( 
.A(n_8402),
.Y(n_10289)
);

CKINVDCx5p33_ASAP7_75t_R g10290 ( 
.A(n_8674),
.Y(n_10290)
);

OA21x2_ASAP7_75t_L g10291 ( 
.A1(n_9016),
.A2(n_7165),
.B(n_7163),
.Y(n_10291)
);

INVx2_ASAP7_75t_L g10292 ( 
.A(n_8919),
.Y(n_10292)
);

INVx2_ASAP7_75t_L g10293 ( 
.A(n_8919),
.Y(n_10293)
);

INVx1_ASAP7_75t_L g10294 ( 
.A(n_8356),
.Y(n_10294)
);

INVxp67_ASAP7_75t_L g10295 ( 
.A(n_8154),
.Y(n_10295)
);

INVx1_ASAP7_75t_L g10296 ( 
.A(n_8356),
.Y(n_10296)
);

INVx3_ASAP7_75t_L g10297 ( 
.A(n_9055),
.Y(n_10297)
);

HB1xp67_ASAP7_75t_L g10298 ( 
.A(n_8268),
.Y(n_10298)
);

OAI22xp33_ASAP7_75t_L g10299 ( 
.A1(n_8587),
.A2(n_7461),
.B1(n_7562),
.B2(n_7293),
.Y(n_10299)
);

BUFx2_ASAP7_75t_L g10300 ( 
.A(n_8364),
.Y(n_10300)
);

INVx2_ASAP7_75t_L g10301 ( 
.A(n_8919),
.Y(n_10301)
);

OAI22xp33_ASAP7_75t_L g10302 ( 
.A1(n_8350),
.A2(n_7461),
.B1(n_7562),
.B2(n_7293),
.Y(n_10302)
);

INVx1_ASAP7_75t_L g10303 ( 
.A(n_8369),
.Y(n_10303)
);

INVx2_ASAP7_75t_L g10304 ( 
.A(n_8919),
.Y(n_10304)
);

AOI22xp33_ASAP7_75t_L g10305 ( 
.A1(n_8583),
.A2(n_7699),
.B1(n_7718),
.B2(n_7695),
.Y(n_10305)
);

AND2x4_ASAP7_75t_L g10306 ( 
.A(n_8758),
.B(n_7163),
.Y(n_10306)
);

AND2x2_ASAP7_75t_L g10307 ( 
.A(n_7985),
.B(n_6974),
.Y(n_10307)
);

INVx3_ASAP7_75t_L g10308 ( 
.A(n_9055),
.Y(n_10308)
);

INVx2_ASAP7_75t_L g10309 ( 
.A(n_8919),
.Y(n_10309)
);

BUFx3_ASAP7_75t_L g10310 ( 
.A(n_8604),
.Y(n_10310)
);

HB1xp67_ASAP7_75t_L g10311 ( 
.A(n_8268),
.Y(n_10311)
);

INVx1_ASAP7_75t_L g10312 ( 
.A(n_8369),
.Y(n_10312)
);

INVx2_ASAP7_75t_L g10313 ( 
.A(n_8964),
.Y(n_10313)
);

INVx2_ASAP7_75t_L g10314 ( 
.A(n_8964),
.Y(n_10314)
);

INVx1_ASAP7_75t_L g10315 ( 
.A(n_8369),
.Y(n_10315)
);

INVx1_ASAP7_75t_L g10316 ( 
.A(n_8376),
.Y(n_10316)
);

HB1xp67_ASAP7_75t_L g10317 ( 
.A(n_8336),
.Y(n_10317)
);

NAND2xp5_ASAP7_75t_L g10318 ( 
.A(n_8628),
.B(n_6936),
.Y(n_10318)
);

HB1xp67_ASAP7_75t_L g10319 ( 
.A(n_8336),
.Y(n_10319)
);

AOI22xp33_ASAP7_75t_L g10320 ( 
.A1(n_8598),
.A2(n_7699),
.B1(n_7718),
.B2(n_7695),
.Y(n_10320)
);

CKINVDCx20_ASAP7_75t_R g10321 ( 
.A(n_8674),
.Y(n_10321)
);

OR2x2_ASAP7_75t_L g10322 ( 
.A(n_8503),
.B(n_8368),
.Y(n_10322)
);

NAND2xp5_ASAP7_75t_L g10323 ( 
.A(n_8618),
.B(n_6936),
.Y(n_10323)
);

INVx1_ASAP7_75t_L g10324 ( 
.A(n_8376),
.Y(n_10324)
);

INVx1_ASAP7_75t_L g10325 ( 
.A(n_8376),
.Y(n_10325)
);

INVx2_ASAP7_75t_L g10326 ( 
.A(n_8964),
.Y(n_10326)
);

AOI22xp33_ASAP7_75t_L g10327 ( 
.A1(n_8598),
.A2(n_7718),
.B1(n_7727),
.B2(n_7699),
.Y(n_10327)
);

INVx2_ASAP7_75t_L g10328 ( 
.A(n_8964),
.Y(n_10328)
);

INVx1_ASAP7_75t_L g10329 ( 
.A(n_8382),
.Y(n_10329)
);

AOI22xp33_ASAP7_75t_L g10330 ( 
.A1(n_8598),
.A2(n_7751),
.B1(n_7766),
.B2(n_7727),
.Y(n_10330)
);

BUFx2_ASAP7_75t_SL g10331 ( 
.A(n_8604),
.Y(n_10331)
);

INVx2_ASAP7_75t_L g10332 ( 
.A(n_8964),
.Y(n_10332)
);

HB1xp67_ASAP7_75t_L g10333 ( 
.A(n_8464),
.Y(n_10333)
);

INVx1_ASAP7_75t_L g10334 ( 
.A(n_8382),
.Y(n_10334)
);

NAND2xp5_ASAP7_75t_L g10335 ( 
.A(n_8628),
.B(n_6936),
.Y(n_10335)
);

AOI21x1_ASAP7_75t_L g10336 ( 
.A1(n_7951),
.A2(n_7222),
.B(n_7215),
.Y(n_10336)
);

INVx6_ASAP7_75t_L g10337 ( 
.A(n_8274),
.Y(n_10337)
);

INVx1_ASAP7_75t_L g10338 ( 
.A(n_8382),
.Y(n_10338)
);

INVx1_ASAP7_75t_L g10339 ( 
.A(n_8384),
.Y(n_10339)
);

INVx1_ASAP7_75t_L g10340 ( 
.A(n_8384),
.Y(n_10340)
);

INVx1_ASAP7_75t_L g10341 ( 
.A(n_8384),
.Y(n_10341)
);

BUFx6f_ASAP7_75t_L g10342 ( 
.A(n_8604),
.Y(n_10342)
);

INVx1_ASAP7_75t_L g10343 ( 
.A(n_8389),
.Y(n_10343)
);

AND2x2_ASAP7_75t_L g10344 ( 
.A(n_7985),
.B(n_6974),
.Y(n_10344)
);

INVx2_ASAP7_75t_L g10345 ( 
.A(n_8964),
.Y(n_10345)
);

OAI21x1_ASAP7_75t_L g10346 ( 
.A1(n_8045),
.A2(n_7884),
.B(n_7880),
.Y(n_10346)
);

CKINVDCx5p33_ASAP7_75t_R g10347 ( 
.A(n_8217),
.Y(n_10347)
);

BUFx2_ASAP7_75t_L g10348 ( 
.A(n_8364),
.Y(n_10348)
);

AOI22xp33_ASAP7_75t_SL g10349 ( 
.A1(n_8297),
.A2(n_7246),
.B1(n_7381),
.B2(n_7247),
.Y(n_10349)
);

INVx1_ASAP7_75t_L g10350 ( 
.A(n_8389),
.Y(n_10350)
);

INVx2_ASAP7_75t_L g10351 ( 
.A(n_8982),
.Y(n_10351)
);

OR2x2_ASAP7_75t_L g10352 ( 
.A(n_8503),
.B(n_7124),
.Y(n_10352)
);

BUFx6f_ASAP7_75t_SL g10353 ( 
.A(n_8604),
.Y(n_10353)
);

INVx2_ASAP7_75t_L g10354 ( 
.A(n_8982),
.Y(n_10354)
);

INVx2_ASAP7_75t_L g10355 ( 
.A(n_8982),
.Y(n_10355)
);

AOI22xp33_ASAP7_75t_SL g10356 ( 
.A1(n_8297),
.A2(n_7246),
.B1(n_7381),
.B2(n_7247),
.Y(n_10356)
);

INVx1_ASAP7_75t_L g10357 ( 
.A(n_8389),
.Y(n_10357)
);

NAND2x1p5_ASAP7_75t_L g10358 ( 
.A(n_8115),
.B(n_7780),
.Y(n_10358)
);

INVx1_ASAP7_75t_L g10359 ( 
.A(n_8391),
.Y(n_10359)
);

INVx2_ASAP7_75t_L g10360 ( 
.A(n_8982),
.Y(n_10360)
);

INVx1_ASAP7_75t_L g10361 ( 
.A(n_8391),
.Y(n_10361)
);

INVx1_ASAP7_75t_L g10362 ( 
.A(n_8391),
.Y(n_10362)
);

INVx1_ASAP7_75t_L g10363 ( 
.A(n_8393),
.Y(n_10363)
);

CKINVDCx20_ASAP7_75t_R g10364 ( 
.A(n_8831),
.Y(n_10364)
);

INVx6_ASAP7_75t_L g10365 ( 
.A(n_8274),
.Y(n_10365)
);

AND2x2_ASAP7_75t_L g10366 ( 
.A(n_8011),
.B(n_7041),
.Y(n_10366)
);

INVx1_ASAP7_75t_L g10367 ( 
.A(n_8393),
.Y(n_10367)
);

INVx1_ASAP7_75t_L g10368 ( 
.A(n_8393),
.Y(n_10368)
);

INVx1_ASAP7_75t_L g10369 ( 
.A(n_8394),
.Y(n_10369)
);

AO21x1_ASAP7_75t_L g10370 ( 
.A1(n_8457),
.A2(n_7869),
.B(n_7864),
.Y(n_10370)
);

BUFx3_ASAP7_75t_L g10371 ( 
.A(n_8617),
.Y(n_10371)
);

NAND2xp5_ASAP7_75t_L g10372 ( 
.A(n_8154),
.B(n_6997),
.Y(n_10372)
);

INVx2_ASAP7_75t_L g10373 ( 
.A(n_8982),
.Y(n_10373)
);

INVx2_ASAP7_75t_L g10374 ( 
.A(n_8982),
.Y(n_10374)
);

AOI22x1_ASAP7_75t_L g10375 ( 
.A1(n_8274),
.A2(n_7360),
.B1(n_7363),
.B2(n_7314),
.Y(n_10375)
);

INVx1_ASAP7_75t_L g10376 ( 
.A(n_8394),
.Y(n_10376)
);

INVx1_ASAP7_75t_L g10377 ( 
.A(n_8394),
.Y(n_10377)
);

NAND2xp5_ASAP7_75t_L g10378 ( 
.A(n_8191),
.B(n_6997),
.Y(n_10378)
);

AOI22xp33_ASAP7_75t_L g10379 ( 
.A1(n_8598),
.A2(n_7751),
.B1(n_7766),
.B2(n_7727),
.Y(n_10379)
);

HB1xp67_ASAP7_75t_L g10380 ( 
.A(n_8464),
.Y(n_10380)
);

INVx2_ASAP7_75t_L g10381 ( 
.A(n_9001),
.Y(n_10381)
);

OAI22xp33_ASAP7_75t_L g10382 ( 
.A1(n_8350),
.A2(n_7691),
.B1(n_7562),
.B2(n_6920),
.Y(n_10382)
);

INVx3_ASAP7_75t_L g10383 ( 
.A(n_9055),
.Y(n_10383)
);

BUFx2_ASAP7_75t_R g10384 ( 
.A(n_8617),
.Y(n_10384)
);

HB1xp67_ASAP7_75t_L g10385 ( 
.A(n_8647),
.Y(n_10385)
);

AOI22xp33_ASAP7_75t_L g10386 ( 
.A1(n_8598),
.A2(n_7766),
.B1(n_7767),
.B2(n_7751),
.Y(n_10386)
);

BUFx2_ASAP7_75t_L g10387 ( 
.A(n_8364),
.Y(n_10387)
);

OAI22xp5_ASAP7_75t_L g10388 ( 
.A1(n_8342),
.A2(n_7596),
.B1(n_7610),
.B2(n_7576),
.Y(n_10388)
);

INVx1_ASAP7_75t_L g10389 ( 
.A(n_8442),
.Y(n_10389)
);

INVx1_ASAP7_75t_L g10390 ( 
.A(n_8442),
.Y(n_10390)
);

INVx1_ASAP7_75t_L g10391 ( 
.A(n_8442),
.Y(n_10391)
);

INVx2_ASAP7_75t_L g10392 ( 
.A(n_9001),
.Y(n_10392)
);

HB1xp67_ASAP7_75t_L g10393 ( 
.A(n_8647),
.Y(n_10393)
);

NAND2xp5_ASAP7_75t_L g10394 ( 
.A(n_8191),
.B(n_6997),
.Y(n_10394)
);

AOI22xp33_ASAP7_75t_SL g10395 ( 
.A1(n_8115),
.A2(n_7247),
.B1(n_7381),
.B2(n_7043),
.Y(n_10395)
);

AOI21x1_ASAP7_75t_L g10396 ( 
.A1(n_8415),
.A2(n_7224),
.B(n_7222),
.Y(n_10396)
);

BUFx6f_ASAP7_75t_L g10397 ( 
.A(n_8617),
.Y(n_10397)
);

INVx3_ASAP7_75t_L g10398 ( 
.A(n_7926),
.Y(n_10398)
);

INVx2_ASAP7_75t_L g10399 ( 
.A(n_9001),
.Y(n_10399)
);

CKINVDCx20_ASAP7_75t_R g10400 ( 
.A(n_8831),
.Y(n_10400)
);

AND2x2_ASAP7_75t_L g10401 ( 
.A(n_8011),
.B(n_7041),
.Y(n_10401)
);

BUFx2_ASAP7_75t_L g10402 ( 
.A(n_8364),
.Y(n_10402)
);

HB1xp67_ASAP7_75t_L g10403 ( 
.A(n_8654),
.Y(n_10403)
);

OAI22xp5_ASAP7_75t_L g10404 ( 
.A1(n_8342),
.A2(n_7596),
.B1(n_7610),
.B2(n_7576),
.Y(n_10404)
);

AND2x2_ASAP7_75t_L g10405 ( 
.A(n_8011),
.B(n_7041),
.Y(n_10405)
);

BUFx2_ASAP7_75t_L g10406 ( 
.A(n_8364),
.Y(n_10406)
);

OR2x2_ASAP7_75t_L g10407 ( 
.A(n_8368),
.B(n_7124),
.Y(n_10407)
);

BUFx4f_ASAP7_75t_SL g10408 ( 
.A(n_8217),
.Y(n_10408)
);

HB1xp67_ASAP7_75t_L g10409 ( 
.A(n_8654),
.Y(n_10409)
);

INVx6_ASAP7_75t_L g10410 ( 
.A(n_8274),
.Y(n_10410)
);

BUFx4f_ASAP7_75t_SL g10411 ( 
.A(n_8217),
.Y(n_10411)
);

INVx4_ASAP7_75t_L g10412 ( 
.A(n_8274),
.Y(n_10412)
);

INVx6_ASAP7_75t_L g10413 ( 
.A(n_8463),
.Y(n_10413)
);

INVx2_ASAP7_75t_SL g10414 ( 
.A(n_8617),
.Y(n_10414)
);

OA21x2_ASAP7_75t_L g10415 ( 
.A1(n_9016),
.A2(n_7165),
.B(n_7123),
.Y(n_10415)
);

AOI22xp33_ASAP7_75t_L g10416 ( 
.A1(n_8750),
.A2(n_7793),
.B1(n_7808),
.B2(n_7767),
.Y(n_10416)
);

INVx1_ASAP7_75t_L g10417 ( 
.A(n_8482),
.Y(n_10417)
);

INVx1_ASAP7_75t_L g10418 ( 
.A(n_8482),
.Y(n_10418)
);

INVx1_ASAP7_75t_L g10419 ( 
.A(n_8482),
.Y(n_10419)
);

AOI22xp33_ASAP7_75t_L g10420 ( 
.A1(n_8750),
.A2(n_7793),
.B1(n_7808),
.B2(n_7767),
.Y(n_10420)
);

AOI22xp33_ASAP7_75t_L g10421 ( 
.A1(n_8540),
.A2(n_7808),
.B1(n_7838),
.B2(n_7793),
.Y(n_10421)
);

OAI22xp33_ASAP7_75t_L g10422 ( 
.A1(n_8018),
.A2(n_7691),
.B1(n_6920),
.B2(n_7060),
.Y(n_10422)
);

AOI22xp33_ASAP7_75t_SL g10423 ( 
.A1(n_8115),
.A2(n_7247),
.B1(n_7381),
.B2(n_7043),
.Y(n_10423)
);

INVx8_ASAP7_75t_L g10424 ( 
.A(n_9278),
.Y(n_10424)
);

AOI22xp33_ASAP7_75t_L g10425 ( 
.A1(n_8540),
.A2(n_7874),
.B1(n_7881),
.B2(n_7838),
.Y(n_10425)
);

INVx1_ASAP7_75t_L g10426 ( 
.A(n_8487),
.Y(n_10426)
);

AOI21x1_ASAP7_75t_L g10427 ( 
.A1(n_8415),
.A2(n_7224),
.B(n_7222),
.Y(n_10427)
);

OAI22xp5_ASAP7_75t_L g10428 ( 
.A1(n_8419),
.A2(n_7610),
.B1(n_7596),
.B2(n_7564),
.Y(n_10428)
);

OAI21x1_ASAP7_75t_L g10429 ( 
.A1(n_8045),
.A2(n_7884),
.B(n_7880),
.Y(n_10429)
);

INVx1_ASAP7_75t_L g10430 ( 
.A(n_8487),
.Y(n_10430)
);

AOI22xp5_ASAP7_75t_L g10431 ( 
.A1(n_8017),
.A2(n_7753),
.B1(n_7759),
.B2(n_7768),
.Y(n_10431)
);

INVx1_ASAP7_75t_L g10432 ( 
.A(n_8487),
.Y(n_10432)
);

INVx1_ASAP7_75t_L g10433 ( 
.A(n_8498),
.Y(n_10433)
);

CKINVDCx20_ASAP7_75t_R g10434 ( 
.A(n_8323),
.Y(n_10434)
);

INVx1_ASAP7_75t_SL g10435 ( 
.A(n_8419),
.Y(n_10435)
);

AOI22xp33_ASAP7_75t_L g10436 ( 
.A1(n_8017),
.A2(n_7874),
.B1(n_7881),
.B2(n_7838),
.Y(n_10436)
);

AOI22xp33_ASAP7_75t_L g10437 ( 
.A1(n_8243),
.A2(n_7881),
.B1(n_7887),
.B2(n_7874),
.Y(n_10437)
);

INVx2_ASAP7_75t_L g10438 ( 
.A(n_9001),
.Y(n_10438)
);

OA21x2_ASAP7_75t_L g10439 ( 
.A1(n_8924),
.A2(n_7165),
.B(n_7123),
.Y(n_10439)
);

INVx1_ASAP7_75t_L g10440 ( 
.A(n_8498),
.Y(n_10440)
);

BUFx10_ASAP7_75t_L g10441 ( 
.A(n_8087),
.Y(n_10441)
);

INVx1_ASAP7_75t_L g10442 ( 
.A(n_8498),
.Y(n_10442)
);

OAI21x1_ASAP7_75t_L g10443 ( 
.A1(n_8045),
.A2(n_7897),
.B(n_7884),
.Y(n_10443)
);

BUFx6f_ASAP7_75t_L g10444 ( 
.A(n_8633),
.Y(n_10444)
);

INVx2_ASAP7_75t_L g10445 ( 
.A(n_9001),
.Y(n_10445)
);

INVx6_ASAP7_75t_L g10446 ( 
.A(n_8463),
.Y(n_10446)
);

INVx2_ASAP7_75t_L g10447 ( 
.A(n_9001),
.Y(n_10447)
);

OAI22xp5_ASAP7_75t_L g10448 ( 
.A1(n_8610),
.A2(n_7610),
.B1(n_7564),
.B2(n_7571),
.Y(n_10448)
);

INVx1_ASAP7_75t_L g10449 ( 
.A(n_8501),
.Y(n_10449)
);

OAI22xp33_ASAP7_75t_L g10450 ( 
.A1(n_8018),
.A2(n_7691),
.B1(n_6920),
.B2(n_7060),
.Y(n_10450)
);

BUFx3_ASAP7_75t_L g10451 ( 
.A(n_8633),
.Y(n_10451)
);

CKINVDCx20_ASAP7_75t_R g10452 ( 
.A(n_8323),
.Y(n_10452)
);

AOI22xp33_ASAP7_75t_SL g10453 ( 
.A1(n_8115),
.A2(n_7381),
.B1(n_7424),
.B2(n_7043),
.Y(n_10453)
);

INVx1_ASAP7_75t_L g10454 ( 
.A(n_8501),
.Y(n_10454)
);

INVx1_ASAP7_75t_L g10455 ( 
.A(n_8501),
.Y(n_10455)
);

INVx1_ASAP7_75t_L g10456 ( 
.A(n_8504),
.Y(n_10456)
);

INVxp67_ASAP7_75t_L g10457 ( 
.A(n_8241),
.Y(n_10457)
);

INVx1_ASAP7_75t_L g10458 ( 
.A(n_8504),
.Y(n_10458)
);

INVx3_ASAP7_75t_L g10459 ( 
.A(n_7926),
.Y(n_10459)
);

OAI21x1_ASAP7_75t_L g10460 ( 
.A1(n_8066),
.A2(n_7897),
.B(n_7884),
.Y(n_10460)
);

INVx2_ASAP7_75t_L g10461 ( 
.A(n_8979),
.Y(n_10461)
);

BUFx6f_ASAP7_75t_L g10462 ( 
.A(n_8633),
.Y(n_10462)
);

INVx3_ASAP7_75t_L g10463 ( 
.A(n_7926),
.Y(n_10463)
);

NAND2xp5_ASAP7_75t_L g10464 ( 
.A(n_8241),
.B(n_6997),
.Y(n_10464)
);

CKINVDCx5p33_ASAP7_75t_R g10465 ( 
.A(n_8323),
.Y(n_10465)
);

INVx1_ASAP7_75t_L g10466 ( 
.A(n_8504),
.Y(n_10466)
);

OAI21x1_ASAP7_75t_L g10467 ( 
.A1(n_8066),
.A2(n_7897),
.B(n_6937),
.Y(n_10467)
);

INVx1_ASAP7_75t_L g10468 ( 
.A(n_8521),
.Y(n_10468)
);

INVx1_ASAP7_75t_L g10469 ( 
.A(n_8521),
.Y(n_10469)
);

INVx1_ASAP7_75t_L g10470 ( 
.A(n_8521),
.Y(n_10470)
);

INVx1_ASAP7_75t_L g10471 ( 
.A(n_8522),
.Y(n_10471)
);

NAND2x1_ASAP7_75t_L g10472 ( 
.A(n_8231),
.B(n_7482),
.Y(n_10472)
);

NAND2x1p5_ASAP7_75t_L g10473 ( 
.A(n_8044),
.B(n_7780),
.Y(n_10473)
);

NAND2x1p5_ASAP7_75t_L g10474 ( 
.A(n_8044),
.B(n_7795),
.Y(n_10474)
);

BUFx3_ASAP7_75t_L g10475 ( 
.A(n_8633),
.Y(n_10475)
);

AND2x2_ASAP7_75t_L g10476 ( 
.A(n_8047),
.B(n_8157),
.Y(n_10476)
);

INVx6_ASAP7_75t_L g10477 ( 
.A(n_8463),
.Y(n_10477)
);

BUFx6f_ASAP7_75t_L g10478 ( 
.A(n_8684),
.Y(n_10478)
);

OAI21x1_ASAP7_75t_L g10479 ( 
.A1(n_8066),
.A2(n_7897),
.B(n_6937),
.Y(n_10479)
);

AOI22xp33_ASAP7_75t_L g10480 ( 
.A1(n_8243),
.A2(n_7888),
.B1(n_7893),
.B2(n_7887),
.Y(n_10480)
);

INVx1_ASAP7_75t_L g10481 ( 
.A(n_8522),
.Y(n_10481)
);

NAND3xp33_ASAP7_75t_L g10482 ( 
.A(n_7945),
.B(n_7741),
.C(n_7715),
.Y(n_10482)
);

INVx2_ASAP7_75t_L g10483 ( 
.A(n_8979),
.Y(n_10483)
);

OAI21x1_ASAP7_75t_L g10484 ( 
.A1(n_8874),
.A2(n_7897),
.B(n_6937),
.Y(n_10484)
);

CKINVDCx20_ASAP7_75t_R g10485 ( 
.A(n_8496),
.Y(n_10485)
);

OAI21x1_ASAP7_75t_L g10486 ( 
.A1(n_8874),
.A2(n_7897),
.B(n_6937),
.Y(n_10486)
);

INVx2_ASAP7_75t_L g10487 ( 
.A(n_8979),
.Y(n_10487)
);

BUFx6f_ASAP7_75t_L g10488 ( 
.A(n_8684),
.Y(n_10488)
);

CKINVDCx20_ASAP7_75t_R g10489 ( 
.A(n_8496),
.Y(n_10489)
);

NAND2x1p5_ASAP7_75t_L g10490 ( 
.A(n_8044),
.B(n_7795),
.Y(n_10490)
);

AOI21xp5_ASAP7_75t_L g10491 ( 
.A1(n_8037),
.A2(n_7694),
.B(n_7904),
.Y(n_10491)
);

INVx1_ASAP7_75t_L g10492 ( 
.A(n_8522),
.Y(n_10492)
);

AND2x4_ASAP7_75t_L g10493 ( 
.A(n_8758),
.B(n_7143),
.Y(n_10493)
);

INVx1_ASAP7_75t_L g10494 ( 
.A(n_8523),
.Y(n_10494)
);

INVx2_ASAP7_75t_L g10495 ( 
.A(n_8979),
.Y(n_10495)
);

AOI22xp33_ASAP7_75t_L g10496 ( 
.A1(n_9189),
.A2(n_7888),
.B1(n_7893),
.B2(n_7887),
.Y(n_10496)
);

AND2x2_ASAP7_75t_L g10497 ( 
.A(n_8047),
.B(n_7041),
.Y(n_10497)
);

INVxp67_ASAP7_75t_L g10498 ( 
.A(n_8282),
.Y(n_10498)
);

AOI22xp33_ASAP7_75t_SL g10499 ( 
.A1(n_9105),
.A2(n_7424),
.B1(n_7463),
.B2(n_7043),
.Y(n_10499)
);

INVx2_ASAP7_75t_L g10500 ( 
.A(n_8979),
.Y(n_10500)
);

INVx1_ASAP7_75t_L g10501 ( 
.A(n_8523),
.Y(n_10501)
);

INVx2_ASAP7_75t_L g10502 ( 
.A(n_8985),
.Y(n_10502)
);

INVx6_ASAP7_75t_L g10503 ( 
.A(n_8463),
.Y(n_10503)
);

INVx1_ASAP7_75t_L g10504 ( 
.A(n_8523),
.Y(n_10504)
);

CKINVDCx5p33_ASAP7_75t_R g10505 ( 
.A(n_8496),
.Y(n_10505)
);

OAI21x1_ASAP7_75t_L g10506 ( 
.A1(n_8993),
.A2(n_6937),
.B(n_6914),
.Y(n_10506)
);

INVx1_ASAP7_75t_L g10507 ( 
.A(n_8527),
.Y(n_10507)
);

CKINVDCx20_ASAP7_75t_R g10508 ( 
.A(n_8539),
.Y(n_10508)
);

INVx2_ASAP7_75t_L g10509 ( 
.A(n_8985),
.Y(n_10509)
);

INVx1_ASAP7_75t_L g10510 ( 
.A(n_8527),
.Y(n_10510)
);

OAI21x1_ASAP7_75t_L g10511 ( 
.A1(n_8993),
.A2(n_6937),
.B(n_6914),
.Y(n_10511)
);

INVx1_ASAP7_75t_SL g10512 ( 
.A(n_8684),
.Y(n_10512)
);

OAI22xp33_ASAP7_75t_SL g10513 ( 
.A1(n_8921),
.A2(n_7691),
.B1(n_6920),
.B2(n_7060),
.Y(n_10513)
);

AOI21xp5_ASAP7_75t_L g10514 ( 
.A1(n_7909),
.A2(n_7904),
.B(n_7216),
.Y(n_10514)
);

INVx2_ASAP7_75t_L g10515 ( 
.A(n_8985),
.Y(n_10515)
);

HB1xp67_ASAP7_75t_L g10516 ( 
.A(n_8711),
.Y(n_10516)
);

INVx3_ASAP7_75t_L g10517 ( 
.A(n_7926),
.Y(n_10517)
);

AND2x2_ASAP7_75t_L g10518 ( 
.A(n_8047),
.B(n_7058),
.Y(n_10518)
);

INVx11_ASAP7_75t_L g10519 ( 
.A(n_8836),
.Y(n_10519)
);

AOI22xp33_ASAP7_75t_L g10520 ( 
.A1(n_9189),
.A2(n_7893),
.B1(n_7899),
.B2(n_7888),
.Y(n_10520)
);

BUFx2_ASAP7_75t_R g10521 ( 
.A(n_8684),
.Y(n_10521)
);

OAI21x1_ASAP7_75t_L g10522 ( 
.A1(n_8449),
.A2(n_6950),
.B(n_6914),
.Y(n_10522)
);

AOI22xp33_ASAP7_75t_SL g10523 ( 
.A1(n_9105),
.A2(n_7424),
.B1(n_7463),
.B2(n_7043),
.Y(n_10523)
);

INVx1_ASAP7_75t_L g10524 ( 
.A(n_8527),
.Y(n_10524)
);

AOI21x1_ASAP7_75t_L g10525 ( 
.A1(n_8415),
.A2(n_7224),
.B(n_7222),
.Y(n_10525)
);

AOI22xp33_ASAP7_75t_SL g10526 ( 
.A1(n_8044),
.A2(n_7424),
.B1(n_7463),
.B2(n_7043),
.Y(n_10526)
);

HB1xp67_ASAP7_75t_L g10527 ( 
.A(n_8711),
.Y(n_10527)
);

AOI22xp33_ASAP7_75t_SL g10528 ( 
.A1(n_8044),
.A2(n_7424),
.B1(n_7463),
.B2(n_7043),
.Y(n_10528)
);

INVx2_ASAP7_75t_L g10529 ( 
.A(n_8985),
.Y(n_10529)
);

INVx3_ASAP7_75t_L g10530 ( 
.A(n_7926),
.Y(n_10530)
);

INVxp67_ASAP7_75t_SL g10531 ( 
.A(n_9040),
.Y(n_10531)
);

INVx2_ASAP7_75t_L g10532 ( 
.A(n_8985),
.Y(n_10532)
);

INVx2_ASAP7_75t_L g10533 ( 
.A(n_9007),
.Y(n_10533)
);

INVx2_ASAP7_75t_L g10534 ( 
.A(n_9007),
.Y(n_10534)
);

INVx1_ASAP7_75t_L g10535 ( 
.A(n_8542),
.Y(n_10535)
);

INVx1_ASAP7_75t_L g10536 ( 
.A(n_8542),
.Y(n_10536)
);

INVx1_ASAP7_75t_L g10537 ( 
.A(n_8542),
.Y(n_10537)
);

BUFx2_ASAP7_75t_L g10538 ( 
.A(n_8364),
.Y(n_10538)
);

BUFx6f_ASAP7_75t_L g10539 ( 
.A(n_8717),
.Y(n_10539)
);

AND2x4_ASAP7_75t_L g10540 ( 
.A(n_8758),
.B(n_7143),
.Y(n_10540)
);

INVx2_ASAP7_75t_L g10541 ( 
.A(n_9007),
.Y(n_10541)
);

INVx1_ASAP7_75t_L g10542 ( 
.A(n_8568),
.Y(n_10542)
);

INVx1_ASAP7_75t_L g10543 ( 
.A(n_8568),
.Y(n_10543)
);

BUFx4f_ASAP7_75t_L g10544 ( 
.A(n_8539),
.Y(n_10544)
);

OAI22xp33_ASAP7_75t_L g10545 ( 
.A1(n_8530),
.A2(n_7691),
.B1(n_6920),
.B2(n_7060),
.Y(n_10545)
);

INVx3_ASAP7_75t_L g10546 ( 
.A(n_8026),
.Y(n_10546)
);

INVx1_ASAP7_75t_L g10547 ( 
.A(n_8568),
.Y(n_10547)
);

INVxp67_ASAP7_75t_SL g10548 ( 
.A(n_9040),
.Y(n_10548)
);

AO21x2_ASAP7_75t_L g10549 ( 
.A1(n_8137),
.A2(n_7317),
.B(n_7264),
.Y(n_10549)
);

INVx1_ASAP7_75t_L g10550 ( 
.A(n_8584),
.Y(n_10550)
);

AOI22xp33_ASAP7_75t_L g10551 ( 
.A1(n_8616),
.A2(n_7899),
.B1(n_6922),
.B2(n_6945),
.Y(n_10551)
);

HB1xp67_ASAP7_75t_L g10552 ( 
.A(n_8770),
.Y(n_10552)
);

INVx3_ASAP7_75t_L g10553 ( 
.A(n_8026),
.Y(n_10553)
);

AOI22xp33_ASAP7_75t_L g10554 ( 
.A1(n_8616),
.A2(n_7899),
.B1(n_6922),
.B2(n_6945),
.Y(n_10554)
);

AND2x2_ASAP7_75t_L g10555 ( 
.A(n_8157),
.B(n_7058),
.Y(n_10555)
);

INVx1_ASAP7_75t_L g10556 ( 
.A(n_8584),
.Y(n_10556)
);

OAI22xp33_ASAP7_75t_L g10557 ( 
.A1(n_8530),
.A2(n_8454),
.B1(n_8810),
.B2(n_8505),
.Y(n_10557)
);

INVx1_ASAP7_75t_L g10558 ( 
.A(n_8584),
.Y(n_10558)
);

BUFx3_ASAP7_75t_L g10559 ( 
.A(n_8717),
.Y(n_10559)
);

INVx1_ASAP7_75t_L g10560 ( 
.A(n_8614),
.Y(n_10560)
);

AND2x2_ASAP7_75t_L g10561 ( 
.A(n_8157),
.B(n_7058),
.Y(n_10561)
);

INVx1_ASAP7_75t_L g10562 ( 
.A(n_8614),
.Y(n_10562)
);

INVx2_ASAP7_75t_L g10563 ( 
.A(n_9007),
.Y(n_10563)
);

INVx1_ASAP7_75t_L g10564 ( 
.A(n_8614),
.Y(n_10564)
);

INVx2_ASAP7_75t_L g10565 ( 
.A(n_9007),
.Y(n_10565)
);

OA21x2_ASAP7_75t_L g10566 ( 
.A1(n_8924),
.A2(n_7123),
.B(n_7111),
.Y(n_10566)
);

BUFx16f_ASAP7_75t_R g10567 ( 
.A(n_8539),
.Y(n_10567)
);

AOI22xp33_ASAP7_75t_L g10568 ( 
.A1(n_8345),
.A2(n_8535),
.B1(n_8506),
.B2(n_8463),
.Y(n_10568)
);

AND2x2_ASAP7_75t_L g10569 ( 
.A(n_8168),
.B(n_7058),
.Y(n_10569)
);

AOI22xp5_ASAP7_75t_L g10570 ( 
.A1(n_8911),
.A2(n_7768),
.B1(n_7451),
.B2(n_7102),
.Y(n_10570)
);

AOI22xp33_ASAP7_75t_L g10571 ( 
.A1(n_8345),
.A2(n_6922),
.B1(n_6945),
.B2(n_6938),
.Y(n_10571)
);

HB1xp67_ASAP7_75t_L g10572 ( 
.A(n_8770),
.Y(n_10572)
);

INVx2_ASAP7_75t_SL g10573 ( 
.A(n_8717),
.Y(n_10573)
);

NAND2xp5_ASAP7_75t_SL g10574 ( 
.A(n_8463),
.B(n_7493),
.Y(n_10574)
);

INVx1_ASAP7_75t_L g10575 ( 
.A(n_8619),
.Y(n_10575)
);

AO21x1_ASAP7_75t_L g10576 ( 
.A1(n_8457),
.A2(n_7869),
.B(n_7864),
.Y(n_10576)
);

AO21x2_ASAP7_75t_L g10577 ( 
.A1(n_8352),
.A2(n_7390),
.B(n_7348),
.Y(n_10577)
);

INVx1_ASAP7_75t_L g10578 ( 
.A(n_8619),
.Y(n_10578)
);

INVx3_ASAP7_75t_L g10579 ( 
.A(n_8026),
.Y(n_10579)
);

AOI22xp33_ASAP7_75t_L g10580 ( 
.A1(n_8535),
.A2(n_6922),
.B1(n_6945),
.B2(n_6938),
.Y(n_10580)
);

INVx1_ASAP7_75t_L g10581 ( 
.A(n_8619),
.Y(n_10581)
);

AOI22xp33_ASAP7_75t_L g10582 ( 
.A1(n_8506),
.A2(n_6922),
.B1(n_6945),
.B2(n_6938),
.Y(n_10582)
);

NAND2xp5_ASAP7_75t_L g10583 ( 
.A(n_8921),
.B(n_7039),
.Y(n_10583)
);

INVx1_ASAP7_75t_L g10584 ( 
.A(n_8625),
.Y(n_10584)
);

OAI22xp33_ASAP7_75t_L g10585 ( 
.A1(n_8454),
.A2(n_7060),
.B1(n_6775),
.B2(n_7258),
.Y(n_10585)
);

INVx1_ASAP7_75t_L g10586 ( 
.A(n_8625),
.Y(n_10586)
);

INVx2_ASAP7_75t_L g10587 ( 
.A(n_9020),
.Y(n_10587)
);

NAND2xp5_ASAP7_75t_L g10588 ( 
.A(n_9083),
.B(n_7039),
.Y(n_10588)
);

INVx2_ASAP7_75t_L g10589 ( 
.A(n_9020),
.Y(n_10589)
);

CKINVDCx6p67_ASAP7_75t_R g10590 ( 
.A(n_8606),
.Y(n_10590)
);

INVx2_ASAP7_75t_SL g10591 ( 
.A(n_8717),
.Y(n_10591)
);

OAI21x1_ASAP7_75t_L g10592 ( 
.A1(n_8449),
.A2(n_6950),
.B(n_6914),
.Y(n_10592)
);

INVx5_ASAP7_75t_L g10593 ( 
.A(n_8026),
.Y(n_10593)
);

OAI22xp5_ASAP7_75t_L g10594 ( 
.A1(n_8610),
.A2(n_7571),
.B1(n_7578),
.B2(n_7560),
.Y(n_10594)
);

AOI21x1_ASAP7_75t_L g10595 ( 
.A1(n_8246),
.A2(n_7226),
.B(n_7224),
.Y(n_10595)
);

INVx1_ASAP7_75t_L g10596 ( 
.A(n_8625),
.Y(n_10596)
);

INVx1_ASAP7_75t_L g10597 ( 
.A(n_8634),
.Y(n_10597)
);

INVx2_ASAP7_75t_L g10598 ( 
.A(n_9020),
.Y(n_10598)
);

INVx2_ASAP7_75t_L g10599 ( 
.A(n_9020),
.Y(n_10599)
);

INVx1_ASAP7_75t_L g10600 ( 
.A(n_8634),
.Y(n_10600)
);

NAND2xp5_ASAP7_75t_L g10601 ( 
.A(n_9083),
.B(n_7039),
.Y(n_10601)
);

INVx3_ASAP7_75t_L g10602 ( 
.A(n_8026),
.Y(n_10602)
);

INVx1_ASAP7_75t_L g10603 ( 
.A(n_8634),
.Y(n_10603)
);

OAI21xp5_ASAP7_75t_L g10604 ( 
.A1(n_8438),
.A2(n_7320),
.B(n_7319),
.Y(n_10604)
);

AND2x4_ASAP7_75t_L g10605 ( 
.A(n_8758),
.B(n_7143),
.Y(n_10605)
);

INVx1_ASAP7_75t_L g10606 ( 
.A(n_8642),
.Y(n_10606)
);

INVx1_ASAP7_75t_L g10607 ( 
.A(n_8642),
.Y(n_10607)
);

OR2x2_ASAP7_75t_L g10608 ( 
.A(n_8401),
.B(n_7124),
.Y(n_10608)
);

BUFx3_ASAP7_75t_L g10609 ( 
.A(n_8744),
.Y(n_10609)
);

CKINVDCx20_ASAP7_75t_R g10610 ( 
.A(n_8606),
.Y(n_10610)
);

INVx1_ASAP7_75t_SL g10611 ( 
.A(n_8744),
.Y(n_10611)
);

OAI21x1_ASAP7_75t_L g10612 ( 
.A1(n_8449),
.A2(n_6950),
.B(n_6914),
.Y(n_10612)
);

OR2x6_ASAP7_75t_L g10613 ( 
.A(n_8086),
.B(n_7109),
.Y(n_10613)
);

INVx1_ASAP7_75t_L g10614 ( 
.A(n_8642),
.Y(n_10614)
);

INVx1_ASAP7_75t_L g10615 ( 
.A(n_8648),
.Y(n_10615)
);

INVx1_ASAP7_75t_L g10616 ( 
.A(n_8648),
.Y(n_10616)
);

INVx1_ASAP7_75t_L g10617 ( 
.A(n_8648),
.Y(n_10617)
);

AND2x2_ASAP7_75t_L g10618 ( 
.A(n_8168),
.B(n_7077),
.Y(n_10618)
);

INVx2_ASAP7_75t_L g10619 ( 
.A(n_9020),
.Y(n_10619)
);

INVx1_ASAP7_75t_L g10620 ( 
.A(n_8649),
.Y(n_10620)
);

INVx1_ASAP7_75t_L g10621 ( 
.A(n_8649),
.Y(n_10621)
);

INVx2_ASAP7_75t_SL g10622 ( 
.A(n_8744),
.Y(n_10622)
);

INVx1_ASAP7_75t_L g10623 ( 
.A(n_8649),
.Y(n_10623)
);

BUFx6f_ASAP7_75t_L g10624 ( 
.A(n_8744),
.Y(n_10624)
);

INVx3_ASAP7_75t_L g10625 ( 
.A(n_8026),
.Y(n_10625)
);

BUFx2_ASAP7_75t_R g10626 ( 
.A(n_8753),
.Y(n_10626)
);

INVx1_ASAP7_75t_L g10627 ( 
.A(n_8664),
.Y(n_10627)
);

CKINVDCx16_ASAP7_75t_R g10628 ( 
.A(n_8753),
.Y(n_10628)
);

INVx3_ASAP7_75t_L g10629 ( 
.A(n_8026),
.Y(n_10629)
);

INVx1_ASAP7_75t_L g10630 ( 
.A(n_8664),
.Y(n_10630)
);

BUFx3_ASAP7_75t_L g10631 ( 
.A(n_8753),
.Y(n_10631)
);

AOI22xp33_ASAP7_75t_L g10632 ( 
.A1(n_8506),
.A2(n_6922),
.B1(n_6945),
.B2(n_6938),
.Y(n_10632)
);

OAI21xp5_ASAP7_75t_L g10633 ( 
.A1(n_8438),
.A2(n_7320),
.B(n_7319),
.Y(n_10633)
);

INVx1_ASAP7_75t_SL g10634 ( 
.A(n_8753),
.Y(n_10634)
);

INVx2_ASAP7_75t_L g10635 ( 
.A(n_9077),
.Y(n_10635)
);

AOI21x1_ASAP7_75t_L g10636 ( 
.A1(n_8246),
.A2(n_7230),
.B(n_7226),
.Y(n_10636)
);

AOI22xp33_ASAP7_75t_SL g10637 ( 
.A1(n_8044),
.A2(n_7424),
.B1(n_7463),
.B2(n_7043),
.Y(n_10637)
);

INVx2_ASAP7_75t_L g10638 ( 
.A(n_9077),
.Y(n_10638)
);

INVx1_ASAP7_75t_L g10639 ( 
.A(n_8664),
.Y(n_10639)
);

INVx2_ASAP7_75t_SL g10640 ( 
.A(n_8756),
.Y(n_10640)
);

BUFx3_ASAP7_75t_L g10641 ( 
.A(n_8756),
.Y(n_10641)
);

INVx2_ASAP7_75t_L g10642 ( 
.A(n_9077),
.Y(n_10642)
);

INVx1_ASAP7_75t_L g10643 ( 
.A(n_8687),
.Y(n_10643)
);

OAI22xp5_ASAP7_75t_L g10644 ( 
.A1(n_8810),
.A2(n_7578),
.B1(n_7580),
.B2(n_7560),
.Y(n_10644)
);

INVxp67_ASAP7_75t_SL g10645 ( 
.A(n_9040),
.Y(n_10645)
);

AO21x1_ASAP7_75t_SL g10646 ( 
.A1(n_9190),
.A2(n_7580),
.B(n_7715),
.Y(n_10646)
);

CKINVDCx5p33_ASAP7_75t_R g10647 ( 
.A(n_8606),
.Y(n_10647)
);

AOI22xp33_ASAP7_75t_L g10648 ( 
.A1(n_8506),
.A2(n_6938),
.B1(n_6991),
.B2(n_6948),
.Y(n_10648)
);

INVx1_ASAP7_75t_L g10649 ( 
.A(n_8687),
.Y(n_10649)
);

INVx2_ASAP7_75t_L g10650 ( 
.A(n_9077),
.Y(n_10650)
);

NAND2x1p5_ASAP7_75t_L g10651 ( 
.A(n_8758),
.B(n_7795),
.Y(n_10651)
);

INVx1_ASAP7_75t_L g10652 ( 
.A(n_8687),
.Y(n_10652)
);

INVx1_ASAP7_75t_L g10653 ( 
.A(n_8690),
.Y(n_10653)
);

INVx2_ASAP7_75t_L g10654 ( 
.A(n_9077),
.Y(n_10654)
);

NAND2xp5_ASAP7_75t_L g10655 ( 
.A(n_9224),
.B(n_7039),
.Y(n_10655)
);

OAI21x1_ASAP7_75t_L g10656 ( 
.A1(n_8855),
.A2(n_6950),
.B(n_6914),
.Y(n_10656)
);

INVx1_ASAP7_75t_L g10657 ( 
.A(n_8690),
.Y(n_10657)
);

INVx1_ASAP7_75t_L g10658 ( 
.A(n_8690),
.Y(n_10658)
);

HB1xp67_ASAP7_75t_L g10659 ( 
.A(n_8867),
.Y(n_10659)
);

BUFx10_ASAP7_75t_L g10660 ( 
.A(n_8087),
.Y(n_10660)
);

AOI22xp33_ASAP7_75t_L g10661 ( 
.A1(n_8506),
.A2(n_6938),
.B1(n_6991),
.B2(n_6948),
.Y(n_10661)
);

INVx1_ASAP7_75t_L g10662 ( 
.A(n_8697),
.Y(n_10662)
);

AOI22xp5_ASAP7_75t_L g10663 ( 
.A1(n_8911),
.A2(n_7102),
.B1(n_7784),
.B2(n_7510),
.Y(n_10663)
);

OAI21x1_ASAP7_75t_L g10664 ( 
.A1(n_8855),
.A2(n_6957),
.B(n_6950),
.Y(n_10664)
);

INVx3_ASAP7_75t_L g10665 ( 
.A(n_8026),
.Y(n_10665)
);

AO21x1_ASAP7_75t_L g10666 ( 
.A1(n_8453),
.A2(n_7547),
.B(n_7095),
.Y(n_10666)
);

INVx6_ASAP7_75t_L g10667 ( 
.A(n_8506),
.Y(n_10667)
);

INVx1_ASAP7_75t_SL g10668 ( 
.A(n_8756),
.Y(n_10668)
);

OAI21x1_ASAP7_75t_L g10669 ( 
.A1(n_8855),
.A2(n_6957),
.B(n_6950),
.Y(n_10669)
);

OR2x2_ASAP7_75t_L g10670 ( 
.A(n_8401),
.B(n_7124),
.Y(n_10670)
);

AOI22xp33_ASAP7_75t_L g10671 ( 
.A1(n_8685),
.A2(n_6948),
.B1(n_6996),
.B2(n_6991),
.Y(n_10671)
);

AND2x2_ASAP7_75t_L g10672 ( 
.A(n_8168),
.B(n_7077),
.Y(n_10672)
);

INVxp33_ASAP7_75t_L g10673 ( 
.A(n_8836),
.Y(n_10673)
);

INVx1_ASAP7_75t_L g10674 ( 
.A(n_8697),
.Y(n_10674)
);

INVx1_ASAP7_75t_L g10675 ( 
.A(n_8697),
.Y(n_10675)
);

INVx1_ASAP7_75t_L g10676 ( 
.A(n_8703),
.Y(n_10676)
);

AOI22xp33_ASAP7_75t_L g10677 ( 
.A1(n_8685),
.A2(n_6948),
.B1(n_6996),
.B2(n_6991),
.Y(n_10677)
);

INVx1_ASAP7_75t_L g10678 ( 
.A(n_8703),
.Y(n_10678)
);

INVx1_ASAP7_75t_L g10679 ( 
.A(n_8703),
.Y(n_10679)
);

INVx1_ASAP7_75t_L g10680 ( 
.A(n_8733),
.Y(n_10680)
);

BUFx6f_ASAP7_75t_L g10681 ( 
.A(n_8756),
.Y(n_10681)
);

OAI22xp5_ASAP7_75t_L g10682 ( 
.A1(n_8529),
.A2(n_7424),
.B1(n_7463),
.B2(n_7582),
.Y(n_10682)
);

INVx2_ASAP7_75t_L g10683 ( 
.A(n_9080),
.Y(n_10683)
);

INVx1_ASAP7_75t_L g10684 ( 
.A(n_8733),
.Y(n_10684)
);

INVx2_ASAP7_75t_L g10685 ( 
.A(n_9080),
.Y(n_10685)
);

HB1xp67_ASAP7_75t_L g10686 ( 
.A(n_8867),
.Y(n_10686)
);

INVx1_ASAP7_75t_L g10687 ( 
.A(n_8733),
.Y(n_10687)
);

INVx1_ASAP7_75t_L g10688 ( 
.A(n_8742),
.Y(n_10688)
);

INVx1_ASAP7_75t_L g10689 ( 
.A(n_8742),
.Y(n_10689)
);

CKINVDCx20_ASAP7_75t_R g10690 ( 
.A(n_8888),
.Y(n_10690)
);

AOI22xp33_ASAP7_75t_L g10691 ( 
.A1(n_8685),
.A2(n_8594),
.B1(n_8155),
.B2(n_8429),
.Y(n_10691)
);

HB1xp67_ASAP7_75t_L g10692 ( 
.A(n_8991),
.Y(n_10692)
);

INVx1_ASAP7_75t_L g10693 ( 
.A(n_8742),
.Y(n_10693)
);

INVx2_ASAP7_75t_L g10694 ( 
.A(n_9080),
.Y(n_10694)
);

AOI22xp33_ASAP7_75t_L g10695 ( 
.A1(n_8685),
.A2(n_6948),
.B1(n_6996),
.B2(n_6991),
.Y(n_10695)
);

HB1xp67_ASAP7_75t_L g10696 ( 
.A(n_8991),
.Y(n_10696)
);

OA21x2_ASAP7_75t_L g10697 ( 
.A1(n_8924),
.A2(n_7126),
.B(n_7111),
.Y(n_10697)
);

INVx2_ASAP7_75t_L g10698 ( 
.A(n_9080),
.Y(n_10698)
);

BUFx12f_ASAP7_75t_L g10699 ( 
.A(n_8685),
.Y(n_10699)
);

AOI22xp33_ASAP7_75t_SL g10700 ( 
.A1(n_8407),
.A2(n_7424),
.B1(n_7463),
.B2(n_7440),
.Y(n_10700)
);

INVx2_ASAP7_75t_L g10701 ( 
.A(n_9080),
.Y(n_10701)
);

AND2x2_ASAP7_75t_L g10702 ( 
.A(n_8187),
.B(n_7077),
.Y(n_10702)
);

OAI21xp33_ASAP7_75t_SL g10703 ( 
.A1(n_8056),
.A2(n_7114),
.B(n_7077),
.Y(n_10703)
);

INVx2_ASAP7_75t_L g10704 ( 
.A(n_9165),
.Y(n_10704)
);

INVx2_ASAP7_75t_L g10705 ( 
.A(n_9165),
.Y(n_10705)
);

CKINVDCx5p33_ASAP7_75t_R g10706 ( 
.A(n_8888),
.Y(n_10706)
);

AOI22xp33_ASAP7_75t_L g10707 ( 
.A1(n_8685),
.A2(n_6948),
.B1(n_6996),
.B2(n_6991),
.Y(n_10707)
);

INVx1_ASAP7_75t_L g10708 ( 
.A(n_8761),
.Y(n_10708)
);

BUFx3_ASAP7_75t_L g10709 ( 
.A(n_8780),
.Y(n_10709)
);

INVx1_ASAP7_75t_L g10710 ( 
.A(n_8761),
.Y(n_10710)
);

INVx1_ASAP7_75t_L g10711 ( 
.A(n_8761),
.Y(n_10711)
);

AND2x2_ASAP7_75t_L g10712 ( 
.A(n_8187),
.B(n_7114),
.Y(n_10712)
);

AOI22xp5_ASAP7_75t_L g10713 ( 
.A1(n_8429),
.A2(n_7102),
.B1(n_7784),
.B2(n_7510),
.Y(n_10713)
);

INVx2_ASAP7_75t_L g10714 ( 
.A(n_9165),
.Y(n_10714)
);

AOI22xp5_ASAP7_75t_L g10715 ( 
.A1(n_7945),
.A2(n_7784),
.B1(n_7463),
.B2(n_7495),
.Y(n_10715)
);

HB1xp67_ASAP7_75t_L g10716 ( 
.A(n_9019),
.Y(n_10716)
);

BUFx2_ASAP7_75t_L g10717 ( 
.A(n_8364),
.Y(n_10717)
);

OAI22xp5_ASAP7_75t_SL g10718 ( 
.A1(n_8662),
.A2(n_7363),
.B1(n_7495),
.B2(n_7493),
.Y(n_10718)
);

BUFx2_ASAP7_75t_L g10719 ( 
.A(n_8364),
.Y(n_10719)
);

NAND2x1p5_ASAP7_75t_L g10720 ( 
.A(n_8758),
.B(n_7795),
.Y(n_10720)
);

NAND2xp5_ASAP7_75t_L g10721 ( 
.A(n_9224),
.B(n_7056),
.Y(n_10721)
);

HB1xp67_ASAP7_75t_L g10722 ( 
.A(n_9019),
.Y(n_10722)
);

NOR2x1_ASAP7_75t_R g10723 ( 
.A(n_8780),
.B(n_8842),
.Y(n_10723)
);

BUFx3_ASAP7_75t_L g10724 ( 
.A(n_9668),
.Y(n_10724)
);

BUFx6f_ASAP7_75t_L g10725 ( 
.A(n_9419),
.Y(n_10725)
);

INVx1_ASAP7_75t_L g10726 ( 
.A(n_9313),
.Y(n_10726)
);

INVx2_ASAP7_75t_L g10727 ( 
.A(n_10476),
.Y(n_10727)
);

BUFx2_ASAP7_75t_L g10728 ( 
.A(n_9419),
.Y(n_10728)
);

NAND2xp5_ASAP7_75t_L g10729 ( 
.A(n_9542),
.B(n_8028),
.Y(n_10729)
);

INVx1_ASAP7_75t_L g10730 ( 
.A(n_9313),
.Y(n_10730)
);

BUFx6f_ASAP7_75t_L g10731 ( 
.A(n_9419),
.Y(n_10731)
);

AOI22xp33_ASAP7_75t_L g10732 ( 
.A1(n_9340),
.A2(n_8351),
.B1(n_7973),
.B2(n_8225),
.Y(n_10732)
);

INVx1_ASAP7_75t_L g10733 ( 
.A(n_9322),
.Y(n_10733)
);

INVx3_ASAP7_75t_L g10734 ( 
.A(n_9719),
.Y(n_10734)
);

HB1xp67_ASAP7_75t_L g10735 ( 
.A(n_9451),
.Y(n_10735)
);

INVx2_ASAP7_75t_L g10736 ( 
.A(n_10476),
.Y(n_10736)
);

INVx1_ASAP7_75t_L g10737 ( 
.A(n_9322),
.Y(n_10737)
);

AND2x2_ASAP7_75t_L g10738 ( 
.A(n_9379),
.B(n_8187),
.Y(n_10738)
);

BUFx2_ASAP7_75t_L g10739 ( 
.A(n_9583),
.Y(n_10739)
);

HB1xp67_ASAP7_75t_L g10740 ( 
.A(n_9462),
.Y(n_10740)
);

INVx1_ASAP7_75t_L g10741 ( 
.A(n_9372),
.Y(n_10741)
);

INVx2_ASAP7_75t_L g10742 ( 
.A(n_10396),
.Y(n_10742)
);

INVxp67_ASAP7_75t_L g10743 ( 
.A(n_9496),
.Y(n_10743)
);

OR2x2_ASAP7_75t_L g10744 ( 
.A(n_10025),
.B(n_7935),
.Y(n_10744)
);

INVx2_ASAP7_75t_L g10745 ( 
.A(n_10396),
.Y(n_10745)
);

NAND2xp33_ASAP7_75t_L g10746 ( 
.A(n_9314),
.B(n_9195),
.Y(n_10746)
);

INVx2_ASAP7_75t_L g10747 ( 
.A(n_10427),
.Y(n_10747)
);

AND2x2_ASAP7_75t_L g10748 ( 
.A(n_9379),
.B(n_8780),
.Y(n_10748)
);

INVx1_ASAP7_75t_L g10749 ( 
.A(n_9365),
.Y(n_10749)
);

INVx1_ASAP7_75t_L g10750 ( 
.A(n_9365),
.Y(n_10750)
);

INVx2_ASAP7_75t_L g10751 ( 
.A(n_10427),
.Y(n_10751)
);

INVx2_ASAP7_75t_SL g10752 ( 
.A(n_9898),
.Y(n_10752)
);

INVx1_ASAP7_75t_L g10753 ( 
.A(n_9366),
.Y(n_10753)
);

AND2x4_ASAP7_75t_L g10754 ( 
.A(n_9593),
.B(n_8758),
.Y(n_10754)
);

OAI21x1_ASAP7_75t_L g10755 ( 
.A1(n_10525),
.A2(n_9213),
.B(n_8875),
.Y(n_10755)
);

AOI21xp5_ASAP7_75t_L g10756 ( 
.A1(n_9602),
.A2(n_10194),
.B(n_9335),
.Y(n_10756)
);

INVx3_ASAP7_75t_L g10757 ( 
.A(n_9719),
.Y(n_10757)
);

BUFx2_ASAP7_75t_SL g10758 ( 
.A(n_9341),
.Y(n_10758)
);

BUFx2_ASAP7_75t_L g10759 ( 
.A(n_9583),
.Y(n_10759)
);

HB1xp67_ASAP7_75t_L g10760 ( 
.A(n_9843),
.Y(n_10760)
);

NAND2xp5_ASAP7_75t_L g10761 ( 
.A(n_9596),
.B(n_8028),
.Y(n_10761)
);

OAI22xp5_ASAP7_75t_L g10762 ( 
.A1(n_9559),
.A2(n_8791),
.B1(n_8692),
.B2(n_8529),
.Y(n_10762)
);

BUFx3_ASAP7_75t_L g10763 ( 
.A(n_9668),
.Y(n_10763)
);

INVx1_ASAP7_75t_SL g10764 ( 
.A(n_9745),
.Y(n_10764)
);

AOI22xp33_ASAP7_75t_L g10765 ( 
.A1(n_9358),
.A2(n_8351),
.B1(n_7973),
.B2(n_8225),
.Y(n_10765)
);

INVx1_ASAP7_75t_L g10766 ( 
.A(n_9342),
.Y(n_10766)
);

OR2x2_ASAP7_75t_L g10767 ( 
.A(n_10322),
.B(n_7935),
.Y(n_10767)
);

INVx1_ASAP7_75t_L g10768 ( 
.A(n_9342),
.Y(n_10768)
);

BUFx3_ASAP7_75t_L g10769 ( 
.A(n_9634),
.Y(n_10769)
);

INVx4_ASAP7_75t_L g10770 ( 
.A(n_9341),
.Y(n_10770)
);

INVx2_ASAP7_75t_L g10771 ( 
.A(n_10525),
.Y(n_10771)
);

INVx2_ASAP7_75t_L g10772 ( 
.A(n_9887),
.Y(n_10772)
);

INVx2_ASAP7_75t_L g10773 ( 
.A(n_9887),
.Y(n_10773)
);

AO21x2_ASAP7_75t_L g10774 ( 
.A1(n_9856),
.A2(n_8352),
.B(n_8056),
.Y(n_10774)
);

OR2x2_ASAP7_75t_L g10775 ( 
.A(n_10322),
.B(n_7963),
.Y(n_10775)
);

OAI21x1_ASAP7_75t_L g10776 ( 
.A1(n_10125),
.A2(n_10592),
.B(n_10522),
.Y(n_10776)
);

INVx3_ASAP7_75t_L g10777 ( 
.A(n_9719),
.Y(n_10777)
);

INVx2_ASAP7_75t_L g10778 ( 
.A(n_9887),
.Y(n_10778)
);

NAND2x1p5_ASAP7_75t_L g10779 ( 
.A(n_9719),
.B(n_8262),
.Y(n_10779)
);

INVx1_ASAP7_75t_L g10780 ( 
.A(n_9359),
.Y(n_10780)
);

INVx1_ASAP7_75t_L g10781 ( 
.A(n_9359),
.Y(n_10781)
);

INVx1_ASAP7_75t_L g10782 ( 
.A(n_9452),
.Y(n_10782)
);

OAI21x1_ASAP7_75t_L g10783 ( 
.A1(n_10125),
.A2(n_9213),
.B(n_8875),
.Y(n_10783)
);

INVx2_ASAP7_75t_L g10784 ( 
.A(n_9893),
.Y(n_10784)
);

OR2x2_ASAP7_75t_L g10785 ( 
.A(n_10011),
.B(n_10037),
.Y(n_10785)
);

OR2x2_ASAP7_75t_L g10786 ( 
.A(n_10011),
.B(n_7963),
.Y(n_10786)
);

INVx1_ASAP7_75t_L g10787 ( 
.A(n_9452),
.Y(n_10787)
);

OAI21xp5_ASAP7_75t_L g10788 ( 
.A1(n_9864),
.A2(n_7950),
.B(n_8136),
.Y(n_10788)
);

HB1xp67_ASAP7_75t_L g10789 ( 
.A(n_9849),
.Y(n_10789)
);

HB1xp67_ASAP7_75t_L g10790 ( 
.A(n_9854),
.Y(n_10790)
);

INVx1_ASAP7_75t_L g10791 ( 
.A(n_9453),
.Y(n_10791)
);

INVx2_ASAP7_75t_L g10792 ( 
.A(n_9893),
.Y(n_10792)
);

INVxp67_ASAP7_75t_L g10793 ( 
.A(n_9496),
.Y(n_10793)
);

AND2x2_ASAP7_75t_L g10794 ( 
.A(n_9387),
.B(n_8780),
.Y(n_10794)
);

BUFx3_ASAP7_75t_L g10795 ( 
.A(n_9853),
.Y(n_10795)
);

INVx1_ASAP7_75t_L g10796 ( 
.A(n_9453),
.Y(n_10796)
);

OR2x2_ASAP7_75t_L g10797 ( 
.A(n_10095),
.B(n_8003),
.Y(n_10797)
);

BUFx2_ASAP7_75t_L g10798 ( 
.A(n_9583),
.Y(n_10798)
);

OR2x6_ASAP7_75t_L g10799 ( 
.A(n_9997),
.B(n_9278),
.Y(n_10799)
);

INVxp67_ASAP7_75t_L g10800 ( 
.A(n_9768),
.Y(n_10800)
);

INVx3_ASAP7_75t_SL g10801 ( 
.A(n_9355),
.Y(n_10801)
);

HB1xp67_ASAP7_75t_L g10802 ( 
.A(n_9996),
.Y(n_10802)
);

INVx2_ASAP7_75t_L g10803 ( 
.A(n_9893),
.Y(n_10803)
);

INVx2_ASAP7_75t_L g10804 ( 
.A(n_9894),
.Y(n_10804)
);

BUFx3_ASAP7_75t_L g10805 ( 
.A(n_9853),
.Y(n_10805)
);

NAND2xp5_ASAP7_75t_L g10806 ( 
.A(n_9844),
.B(n_8051),
.Y(n_10806)
);

AND2x2_ASAP7_75t_L g10807 ( 
.A(n_9387),
.B(n_8100),
.Y(n_10807)
);

INVx1_ASAP7_75t_L g10808 ( 
.A(n_9403),
.Y(n_10808)
);

INVx2_ASAP7_75t_SL g10809 ( 
.A(n_9898),
.Y(n_10809)
);

INVx1_ASAP7_75t_L g10810 ( 
.A(n_9403),
.Y(n_10810)
);

HB1xp67_ASAP7_75t_L g10811 ( 
.A(n_10004),
.Y(n_10811)
);

INVx2_ASAP7_75t_L g10812 ( 
.A(n_9894),
.Y(n_10812)
);

OR2x2_ASAP7_75t_L g10813 ( 
.A(n_10037),
.B(n_8003),
.Y(n_10813)
);

INVx2_ASAP7_75t_L g10814 ( 
.A(n_9894),
.Y(n_10814)
);

HB1xp67_ASAP7_75t_L g10815 ( 
.A(n_10006),
.Y(n_10815)
);

INVx1_ASAP7_75t_L g10816 ( 
.A(n_9456),
.Y(n_10816)
);

INVx1_ASAP7_75t_L g10817 ( 
.A(n_9456),
.Y(n_10817)
);

OR2x2_ASAP7_75t_L g10818 ( 
.A(n_10099),
.B(n_8022),
.Y(n_10818)
);

INVx2_ASAP7_75t_L g10819 ( 
.A(n_9895),
.Y(n_10819)
);

INVx1_ASAP7_75t_L g10820 ( 
.A(n_9466),
.Y(n_10820)
);

INVxp67_ASAP7_75t_R g10821 ( 
.A(n_9839),
.Y(n_10821)
);

AND2x2_ASAP7_75t_L g10822 ( 
.A(n_9400),
.B(n_8100),
.Y(n_10822)
);

INVx1_ASAP7_75t_L g10823 ( 
.A(n_9466),
.Y(n_10823)
);

OR2x6_ASAP7_75t_L g10824 ( 
.A(n_9997),
.B(n_9278),
.Y(n_10824)
);

INVx2_ASAP7_75t_L g10825 ( 
.A(n_9895),
.Y(n_10825)
);

INVx2_ASAP7_75t_L g10826 ( 
.A(n_9895),
.Y(n_10826)
);

INVx1_ASAP7_75t_L g10827 ( 
.A(n_9475),
.Y(n_10827)
);

OAI21x1_ASAP7_75t_L g10828 ( 
.A1(n_10522),
.A2(n_9213),
.B(n_8875),
.Y(n_10828)
);

BUFx2_ASAP7_75t_L g10829 ( 
.A(n_9583),
.Y(n_10829)
);

INVx3_ASAP7_75t_L g10830 ( 
.A(n_9719),
.Y(n_10830)
);

INVx1_ASAP7_75t_L g10831 ( 
.A(n_9475),
.Y(n_10831)
);

BUFx12f_ASAP7_75t_L g10832 ( 
.A(n_9317),
.Y(n_10832)
);

BUFx2_ASAP7_75t_SL g10833 ( 
.A(n_9341),
.Y(n_10833)
);

INVx2_ASAP7_75t_L g10834 ( 
.A(n_9897),
.Y(n_10834)
);

INVx1_ASAP7_75t_L g10835 ( 
.A(n_9476),
.Y(n_10835)
);

INVx1_ASAP7_75t_L g10836 ( 
.A(n_9476),
.Y(n_10836)
);

AND2x2_ASAP7_75t_L g10837 ( 
.A(n_9400),
.B(n_8100),
.Y(n_10837)
);

INVx1_ASAP7_75t_L g10838 ( 
.A(n_9405),
.Y(n_10838)
);

INVx1_ASAP7_75t_L g10839 ( 
.A(n_9405),
.Y(n_10839)
);

CKINVDCx5p33_ASAP7_75t_R g10840 ( 
.A(n_9828),
.Y(n_10840)
);

HB1xp67_ASAP7_75t_L g10841 ( 
.A(n_10022),
.Y(n_10841)
);

AOI211xp5_ASAP7_75t_L g10842 ( 
.A1(n_9491),
.A2(n_8328),
.B(n_8515),
.C(n_7950),
.Y(n_10842)
);

HB1xp67_ASAP7_75t_L g10843 ( 
.A(n_10027),
.Y(n_10843)
);

HB1xp67_ASAP7_75t_L g10844 ( 
.A(n_10124),
.Y(n_10844)
);

OAI22xp5_ASAP7_75t_L g10845 ( 
.A1(n_9559),
.A2(n_8791),
.B1(n_8692),
.B2(n_8771),
.Y(n_10845)
);

INVx2_ASAP7_75t_L g10846 ( 
.A(n_9897),
.Y(n_10846)
);

HB1xp67_ASAP7_75t_SL g10847 ( 
.A(n_9464),
.Y(n_10847)
);

HB1xp67_ASAP7_75t_L g10848 ( 
.A(n_10215),
.Y(n_10848)
);

AND2x4_ASAP7_75t_L g10849 ( 
.A(n_9593),
.B(n_8758),
.Y(n_10849)
);

NAND2xp5_ASAP7_75t_L g10850 ( 
.A(n_9383),
.B(n_8051),
.Y(n_10850)
);

INVx2_ASAP7_75t_L g10851 ( 
.A(n_9897),
.Y(n_10851)
);

OAI21x1_ASAP7_75t_L g10852 ( 
.A1(n_10592),
.A2(n_8553),
.B(n_8547),
.Y(n_10852)
);

INVx2_ASAP7_75t_L g10853 ( 
.A(n_9901),
.Y(n_10853)
);

INVx1_ASAP7_75t_L g10854 ( 
.A(n_9388),
.Y(n_10854)
);

INVx1_ASAP7_75t_L g10855 ( 
.A(n_9388),
.Y(n_10855)
);

INVx1_ASAP7_75t_L g10856 ( 
.A(n_9389),
.Y(n_10856)
);

INVx1_ASAP7_75t_L g10857 ( 
.A(n_9389),
.Y(n_10857)
);

INVx2_ASAP7_75t_L g10858 ( 
.A(n_9901),
.Y(n_10858)
);

INVx1_ASAP7_75t_L g10859 ( 
.A(n_9398),
.Y(n_10859)
);

BUFx3_ASAP7_75t_L g10860 ( 
.A(n_9853),
.Y(n_10860)
);

AOI22xp33_ASAP7_75t_L g10861 ( 
.A1(n_9358),
.A2(n_9867),
.B1(n_9524),
.B2(n_10092),
.Y(n_10861)
);

AND2x2_ASAP7_75t_L g10862 ( 
.A(n_10628),
.B(n_8104),
.Y(n_10862)
);

CKINVDCx5p33_ASAP7_75t_R g10863 ( 
.A(n_10054),
.Y(n_10863)
);

AOI22xp33_ASAP7_75t_SL g10864 ( 
.A1(n_9375),
.A2(n_7970),
.B1(n_9173),
.B2(n_8352),
.Y(n_10864)
);

INVx1_ASAP7_75t_L g10865 ( 
.A(n_9391),
.Y(n_10865)
);

INVx1_ASAP7_75t_L g10866 ( 
.A(n_9391),
.Y(n_10866)
);

AND2x2_ASAP7_75t_L g10867 ( 
.A(n_10628),
.B(n_8104),
.Y(n_10867)
);

INVx1_ASAP7_75t_L g10868 ( 
.A(n_9444),
.Y(n_10868)
);

INVx2_ASAP7_75t_L g10869 ( 
.A(n_9901),
.Y(n_10869)
);

INVx2_ASAP7_75t_L g10870 ( 
.A(n_9905),
.Y(n_10870)
);

OAI21x1_ASAP7_75t_L g10871 ( 
.A1(n_10612),
.A2(n_8553),
.B(n_8547),
.Y(n_10871)
);

BUFx2_ASAP7_75t_L g10872 ( 
.A(n_9317),
.Y(n_10872)
);

INVx1_ASAP7_75t_L g10873 ( 
.A(n_9444),
.Y(n_10873)
);

INVx2_ASAP7_75t_L g10874 ( 
.A(n_9905),
.Y(n_10874)
);

OR2x2_ASAP7_75t_L g10875 ( 
.A(n_10095),
.B(n_8022),
.Y(n_10875)
);

BUFx2_ASAP7_75t_L g10876 ( 
.A(n_9317),
.Y(n_10876)
);

OAI21x1_ASAP7_75t_L g10877 ( 
.A1(n_10612),
.A2(n_8553),
.B(n_8547),
.Y(n_10877)
);

AND2x2_ASAP7_75t_L g10878 ( 
.A(n_9414),
.B(n_8104),
.Y(n_10878)
);

AND2x4_ASAP7_75t_L g10879 ( 
.A(n_9623),
.B(n_9414),
.Y(n_10879)
);

INVx1_ASAP7_75t_L g10880 ( 
.A(n_9486),
.Y(n_10880)
);

AND2x6_ASAP7_75t_L g10881 ( 
.A(n_9317),
.B(n_8842),
.Y(n_10881)
);

AND2x2_ASAP7_75t_L g10882 ( 
.A(n_9414),
.B(n_8141),
.Y(n_10882)
);

OA21x2_ASAP7_75t_L g10883 ( 
.A1(n_10370),
.A2(n_7964),
.B(n_7955),
.Y(n_10883)
);

OAI21x1_ASAP7_75t_L g10884 ( 
.A1(n_10656),
.A2(n_8553),
.B(n_8547),
.Y(n_10884)
);

HB1xp67_ASAP7_75t_L g10885 ( 
.A(n_10219),
.Y(n_10885)
);

INVx2_ASAP7_75t_L g10886 ( 
.A(n_9905),
.Y(n_10886)
);

AND2x2_ASAP7_75t_L g10887 ( 
.A(n_9414),
.B(n_8141),
.Y(n_10887)
);

NAND2xp5_ASAP7_75t_L g10888 ( 
.A(n_10295),
.B(n_8282),
.Y(n_10888)
);

INVx2_ASAP7_75t_L g10889 ( 
.A(n_9908),
.Y(n_10889)
);

OR2x2_ASAP7_75t_L g10890 ( 
.A(n_10099),
.B(n_8423),
.Y(n_10890)
);

INVx2_ASAP7_75t_L g10891 ( 
.A(n_9908),
.Y(n_10891)
);

HB1xp67_ASAP7_75t_L g10892 ( 
.A(n_10234),
.Y(n_10892)
);

INVx2_ASAP7_75t_L g10893 ( 
.A(n_9908),
.Y(n_10893)
);

INVx2_ASAP7_75t_L g10894 ( 
.A(n_9911),
.Y(n_10894)
);

INVx2_ASAP7_75t_L g10895 ( 
.A(n_9911),
.Y(n_10895)
);

AND2x2_ASAP7_75t_L g10896 ( 
.A(n_9447),
.B(n_8141),
.Y(n_10896)
);

INVx1_ASAP7_75t_L g10897 ( 
.A(n_9446),
.Y(n_10897)
);

INVx3_ASAP7_75t_L g10898 ( 
.A(n_9719),
.Y(n_10898)
);

INVx3_ASAP7_75t_L g10899 ( 
.A(n_9808),
.Y(n_10899)
);

INVx2_ASAP7_75t_L g10900 ( 
.A(n_9911),
.Y(n_10900)
);

AO21x1_ASAP7_75t_SL g10901 ( 
.A1(n_9571),
.A2(n_9190),
.B(n_8942),
.Y(n_10901)
);

INVx2_ASAP7_75t_L g10902 ( 
.A(n_9915),
.Y(n_10902)
);

AOI31xp67_ASAP7_75t_L g10903 ( 
.A1(n_10287),
.A2(n_9173),
.A3(n_7930),
.B(n_7953),
.Y(n_10903)
);

BUFx3_ASAP7_75t_L g10904 ( 
.A(n_9916),
.Y(n_10904)
);

INVx2_ASAP7_75t_SL g10905 ( 
.A(n_9898),
.Y(n_10905)
);

OR2x2_ASAP7_75t_L g10906 ( 
.A(n_9508),
.B(n_8423),
.Y(n_10906)
);

AND2x2_ASAP7_75t_L g10907 ( 
.A(n_9447),
.B(n_8842),
.Y(n_10907)
);

INVx2_ASAP7_75t_L g10908 ( 
.A(n_9915),
.Y(n_10908)
);

INVx1_ASAP7_75t_L g10909 ( 
.A(n_9446),
.Y(n_10909)
);

INVx1_ASAP7_75t_L g10910 ( 
.A(n_9459),
.Y(n_10910)
);

CKINVDCx20_ASAP7_75t_R g10911 ( 
.A(n_9983),
.Y(n_10911)
);

BUFx2_ASAP7_75t_L g10912 ( 
.A(n_9317),
.Y(n_10912)
);

INVx3_ASAP7_75t_L g10913 ( 
.A(n_9808),
.Y(n_10913)
);

INVx1_ASAP7_75t_L g10914 ( 
.A(n_9459),
.Y(n_10914)
);

INVx1_ASAP7_75t_L g10915 ( 
.A(n_9481),
.Y(n_10915)
);

INVx1_ASAP7_75t_L g10916 ( 
.A(n_9481),
.Y(n_10916)
);

CKINVDCx20_ASAP7_75t_R g10917 ( 
.A(n_10002),
.Y(n_10917)
);

INVx2_ASAP7_75t_L g10918 ( 
.A(n_9915),
.Y(n_10918)
);

INVx2_ASAP7_75t_L g10919 ( 
.A(n_9918),
.Y(n_10919)
);

OAI21x1_ASAP7_75t_L g10920 ( 
.A1(n_10656),
.A2(n_8561),
.B(n_8405),
.Y(n_10920)
);

INVx1_ASAP7_75t_L g10921 ( 
.A(n_9752),
.Y(n_10921)
);

INVx1_ASAP7_75t_SL g10922 ( 
.A(n_9869),
.Y(n_10922)
);

AND2x4_ASAP7_75t_L g10923 ( 
.A(n_9623),
.B(n_8758),
.Y(n_10923)
);

INVx2_ASAP7_75t_L g10924 ( 
.A(n_9918),
.Y(n_10924)
);

INVx1_ASAP7_75t_L g10925 ( 
.A(n_9671),
.Y(n_10925)
);

INVx1_ASAP7_75t_L g10926 ( 
.A(n_9671),
.Y(n_10926)
);

INVx1_ASAP7_75t_L g10927 ( 
.A(n_9688),
.Y(n_10927)
);

AND2x2_ASAP7_75t_L g10928 ( 
.A(n_9447),
.B(n_8842),
.Y(n_10928)
);

INVx3_ASAP7_75t_L g10929 ( 
.A(n_9808),
.Y(n_10929)
);

NOR2xp33_ASAP7_75t_L g10930 ( 
.A(n_9733),
.B(n_8599),
.Y(n_10930)
);

AND2x2_ASAP7_75t_L g10931 ( 
.A(n_9447),
.B(n_8907),
.Y(n_10931)
);

INVx2_ASAP7_75t_L g10932 ( 
.A(n_9918),
.Y(n_10932)
);

OAI21xp5_ASAP7_75t_L g10933 ( 
.A1(n_9872),
.A2(n_8136),
.B(n_8929),
.Y(n_10933)
);

NOR2xp33_ASAP7_75t_L g10934 ( 
.A(n_9404),
.B(n_9317),
.Y(n_10934)
);

OR2x2_ASAP7_75t_L g10935 ( 
.A(n_9508),
.B(n_9928),
.Y(n_10935)
);

INVx1_ASAP7_75t_L g10936 ( 
.A(n_9344),
.Y(n_10936)
);

AO31x2_ASAP7_75t_L g10937 ( 
.A1(n_9963),
.A2(n_8328),
.A3(n_8669),
.B(n_8772),
.Y(n_10937)
);

OAI21xp5_ASAP7_75t_L g10938 ( 
.A1(n_10482),
.A2(n_9966),
.B(n_10001),
.Y(n_10938)
);

INVx1_ASAP7_75t_L g10939 ( 
.A(n_9344),
.Y(n_10939)
);

INVx1_ASAP7_75t_L g10940 ( 
.A(n_9372),
.Y(n_10940)
);

INVx1_ASAP7_75t_L g10941 ( 
.A(n_9440),
.Y(n_10941)
);

HB1xp67_ASAP7_75t_L g10942 ( 
.A(n_10237),
.Y(n_10942)
);

AND2x2_ASAP7_75t_L g10943 ( 
.A(n_9712),
.B(n_8907),
.Y(n_10943)
);

INVx2_ASAP7_75t_L g10944 ( 
.A(n_9923),
.Y(n_10944)
);

INVx2_ASAP7_75t_L g10945 ( 
.A(n_9923),
.Y(n_10945)
);

INVx1_ASAP7_75t_L g10946 ( 
.A(n_9440),
.Y(n_10946)
);

INVx1_ASAP7_75t_L g10947 ( 
.A(n_9441),
.Y(n_10947)
);

INVx1_ASAP7_75t_L g10948 ( 
.A(n_9441),
.Y(n_10948)
);

INVx2_ASAP7_75t_L g10949 ( 
.A(n_9923),
.Y(n_10949)
);

INVx3_ASAP7_75t_L g10950 ( 
.A(n_9808),
.Y(n_10950)
);

BUFx2_ASAP7_75t_SL g10951 ( 
.A(n_9341),
.Y(n_10951)
);

INVx1_ASAP7_75t_L g10952 ( 
.A(n_9479),
.Y(n_10952)
);

OAI21x1_ASAP7_75t_L g10953 ( 
.A1(n_10664),
.A2(n_8561),
.B(n_8405),
.Y(n_10953)
);

OAI21x1_ASAP7_75t_L g10954 ( 
.A1(n_10664),
.A2(n_8561),
.B(n_8405),
.Y(n_10954)
);

AND2x2_ASAP7_75t_L g10955 ( 
.A(n_9712),
.B(n_8907),
.Y(n_10955)
);

OAI21xp5_ASAP7_75t_L g10956 ( 
.A1(n_10092),
.A2(n_8929),
.B(n_8536),
.Y(n_10956)
);

OA21x2_ASAP7_75t_L g10957 ( 
.A1(n_10370),
.A2(n_7964),
.B(n_7955),
.Y(n_10957)
);

BUFx4f_ASAP7_75t_L g10958 ( 
.A(n_9320),
.Y(n_10958)
);

INVx3_ASAP7_75t_L g10959 ( 
.A(n_9808),
.Y(n_10959)
);

INVx11_ASAP7_75t_L g10960 ( 
.A(n_9751),
.Y(n_10960)
);

BUFx6f_ASAP7_75t_L g10961 ( 
.A(n_9395),
.Y(n_10961)
);

INVx1_ASAP7_75t_L g10962 ( 
.A(n_9479),
.Y(n_10962)
);

INVx1_ASAP7_75t_L g10963 ( 
.A(n_9489),
.Y(n_10963)
);

INVx2_ASAP7_75t_L g10964 ( 
.A(n_9930),
.Y(n_10964)
);

OAI22xp5_ASAP7_75t_L g10965 ( 
.A1(n_10043),
.A2(n_9371),
.B1(n_9945),
.B2(n_9938),
.Y(n_10965)
);

BUFx2_ASAP7_75t_L g10966 ( 
.A(n_9320),
.Y(n_10966)
);

INVx1_ASAP7_75t_L g10967 ( 
.A(n_9407),
.Y(n_10967)
);

OAI21xp5_ASAP7_75t_L g10968 ( 
.A1(n_10009),
.A2(n_8536),
.B(n_8517),
.Y(n_10968)
);

INVx1_ASAP7_75t_L g10969 ( 
.A(n_9407),
.Y(n_10969)
);

OAI21x1_ASAP7_75t_L g10970 ( 
.A1(n_10669),
.A2(n_8561),
.B(n_8387),
.Y(n_10970)
);

INVx2_ASAP7_75t_L g10971 ( 
.A(n_9930),
.Y(n_10971)
);

AND2x4_ASAP7_75t_L g10972 ( 
.A(n_9712),
.B(n_8764),
.Y(n_10972)
);

INVx1_ASAP7_75t_L g10973 ( 
.A(n_9408),
.Y(n_10973)
);

BUFx2_ASAP7_75t_L g10974 ( 
.A(n_9320),
.Y(n_10974)
);

INVx1_ASAP7_75t_L g10975 ( 
.A(n_9408),
.Y(n_10975)
);

AND2x2_ASAP7_75t_L g10976 ( 
.A(n_9712),
.B(n_8907),
.Y(n_10976)
);

INVx2_ASAP7_75t_L g10977 ( 
.A(n_9930),
.Y(n_10977)
);

OA21x2_ASAP7_75t_L g10978 ( 
.A1(n_10576),
.A2(n_7964),
.B(n_7955),
.Y(n_10978)
);

AND2x2_ASAP7_75t_L g10979 ( 
.A(n_10145),
.B(n_10435),
.Y(n_10979)
);

AND2x2_ASAP7_75t_SL g10980 ( 
.A(n_9404),
.B(n_8262),
.Y(n_10980)
);

AND2x2_ASAP7_75t_L g10981 ( 
.A(n_9912),
.B(n_7990),
.Y(n_10981)
);

INVx1_ASAP7_75t_L g10982 ( 
.A(n_9449),
.Y(n_10982)
);

INVx1_ASAP7_75t_L g10983 ( 
.A(n_9449),
.Y(n_10983)
);

OAI21xp33_ASAP7_75t_L g10984 ( 
.A1(n_10274),
.A2(n_8344),
.B(n_8517),
.Y(n_10984)
);

HB1xp67_ASAP7_75t_L g10985 ( 
.A(n_10262),
.Y(n_10985)
);

AND2x2_ASAP7_75t_L g10986 ( 
.A(n_10145),
.B(n_8917),
.Y(n_10986)
);

OAI21x1_ASAP7_75t_L g10987 ( 
.A1(n_10669),
.A2(n_8387),
.B(n_9041),
.Y(n_10987)
);

OAI21x1_ASAP7_75t_L g10988 ( 
.A1(n_9974),
.A2(n_8387),
.B(n_9041),
.Y(n_10988)
);

OAI21x1_ASAP7_75t_L g10989 ( 
.A1(n_9974),
.A2(n_9041),
.B(n_8467),
.Y(n_10989)
);

HB1xp67_ASAP7_75t_L g10990 ( 
.A(n_10298),
.Y(n_10990)
);

AND2x4_ASAP7_75t_L g10991 ( 
.A(n_10145),
.B(n_8764),
.Y(n_10991)
);

BUFx2_ASAP7_75t_L g10992 ( 
.A(n_9320),
.Y(n_10992)
);

AND2x2_ASAP7_75t_L g10993 ( 
.A(n_10145),
.B(n_8917),
.Y(n_10993)
);

INVx2_ASAP7_75t_SL g10994 ( 
.A(n_9898),
.Y(n_10994)
);

INVx2_ASAP7_75t_L g10995 ( 
.A(n_9951),
.Y(n_10995)
);

INVx1_ASAP7_75t_L g10996 ( 
.A(n_9474),
.Y(n_10996)
);

AO21x2_ASAP7_75t_L g10997 ( 
.A1(n_9856),
.A2(n_8669),
.B(n_8328),
.Y(n_10997)
);

INVx2_ASAP7_75t_L g10998 ( 
.A(n_9951),
.Y(n_10998)
);

INVx2_ASAP7_75t_L g10999 ( 
.A(n_9951),
.Y(n_10999)
);

INVx1_ASAP7_75t_L g11000 ( 
.A(n_9474),
.Y(n_11000)
);

INVx2_ASAP7_75t_L g11001 ( 
.A(n_9954),
.Y(n_11001)
);

AND2x4_ASAP7_75t_L g11002 ( 
.A(n_9912),
.B(n_8764),
.Y(n_11002)
);

INVx3_ASAP7_75t_L g11003 ( 
.A(n_9808),
.Y(n_11003)
);

INVx2_ASAP7_75t_L g11004 ( 
.A(n_9954),
.Y(n_11004)
);

INVx3_ASAP7_75t_L g11005 ( 
.A(n_10243),
.Y(n_11005)
);

INVx2_ASAP7_75t_SL g11006 ( 
.A(n_9961),
.Y(n_11006)
);

INVx1_ASAP7_75t_L g11007 ( 
.A(n_9497),
.Y(n_11007)
);

INVx1_ASAP7_75t_L g11008 ( 
.A(n_9497),
.Y(n_11008)
);

AND2x2_ASAP7_75t_L g11009 ( 
.A(n_9436),
.B(n_8917),
.Y(n_11009)
);

AOI22xp33_ASAP7_75t_L g11010 ( 
.A1(n_9963),
.A2(n_7973),
.B1(n_8558),
.B2(n_8407),
.Y(n_11010)
);

BUFx6f_ASAP7_75t_L g11011 ( 
.A(n_9395),
.Y(n_11011)
);

INVx2_ASAP7_75t_L g11012 ( 
.A(n_9954),
.Y(n_11012)
);

INVx1_ASAP7_75t_L g11013 ( 
.A(n_9498),
.Y(n_11013)
);

AND2x2_ASAP7_75t_L g11014 ( 
.A(n_9436),
.B(n_8917),
.Y(n_11014)
);

INVx1_ASAP7_75t_L g11015 ( 
.A(n_9498),
.Y(n_11015)
);

AND2x2_ASAP7_75t_L g11016 ( 
.A(n_9436),
.B(n_8956),
.Y(n_11016)
);

INVx2_ASAP7_75t_L g11017 ( 
.A(n_9958),
.Y(n_11017)
);

AND2x4_ASAP7_75t_L g11018 ( 
.A(n_10243),
.B(n_8764),
.Y(n_11018)
);

CKINVDCx5p33_ASAP7_75t_R g11019 ( 
.A(n_9420),
.Y(n_11019)
);

INVx2_ASAP7_75t_L g11020 ( 
.A(n_9958),
.Y(n_11020)
);

INVx2_ASAP7_75t_L g11021 ( 
.A(n_9958),
.Y(n_11021)
);

INVx2_ASAP7_75t_L g11022 ( 
.A(n_9970),
.Y(n_11022)
);

INVx3_ASAP7_75t_L g11023 ( 
.A(n_10243),
.Y(n_11023)
);

INVx1_ASAP7_75t_L g11024 ( 
.A(n_9454),
.Y(n_11024)
);

INVx2_ASAP7_75t_L g11025 ( 
.A(n_9970),
.Y(n_11025)
);

INVx1_ASAP7_75t_L g11026 ( 
.A(n_9454),
.Y(n_11026)
);

INVx2_ASAP7_75t_L g11027 ( 
.A(n_9970),
.Y(n_11027)
);

INVx1_ASAP7_75t_L g11028 ( 
.A(n_9489),
.Y(n_11028)
);

BUFx3_ASAP7_75t_L g11029 ( 
.A(n_9916),
.Y(n_11029)
);

NOR2xp33_ASAP7_75t_L g11030 ( 
.A(n_9320),
.B(n_8599),
.Y(n_11030)
);

OAI21xp5_ASAP7_75t_L g11031 ( 
.A1(n_10134),
.A2(n_8256),
.B(n_8278),
.Y(n_11031)
);

INVx1_ASAP7_75t_L g11032 ( 
.A(n_9519),
.Y(n_11032)
);

INVx1_ASAP7_75t_L g11033 ( 
.A(n_9519),
.Y(n_11033)
);

INVx1_ASAP7_75t_L g11034 ( 
.A(n_9537),
.Y(n_11034)
);

HB1xp67_ASAP7_75t_L g11035 ( 
.A(n_10311),
.Y(n_11035)
);

INVx2_ASAP7_75t_L g11036 ( 
.A(n_9984),
.Y(n_11036)
);

INVx2_ASAP7_75t_SL g11037 ( 
.A(n_9961),
.Y(n_11037)
);

BUFx3_ASAP7_75t_L g11038 ( 
.A(n_9916),
.Y(n_11038)
);

INVx1_ASAP7_75t_L g11039 ( 
.A(n_9537),
.Y(n_11039)
);

NAND2x1p5_ASAP7_75t_L g11040 ( 
.A(n_10243),
.B(n_8764),
.Y(n_11040)
);

BUFx3_ASAP7_75t_L g11041 ( 
.A(n_9998),
.Y(n_11041)
);

BUFx3_ASAP7_75t_L g11042 ( 
.A(n_9998),
.Y(n_11042)
);

OR2x6_ASAP7_75t_L g11043 ( 
.A(n_10065),
.B(n_9278),
.Y(n_11043)
);

NOR2xp33_ASAP7_75t_L g11044 ( 
.A(n_9320),
.B(n_8956),
.Y(n_11044)
);

AND2x2_ASAP7_75t_L g11045 ( 
.A(n_9436),
.B(n_8956),
.Y(n_11045)
);

OAI21x1_ASAP7_75t_L g11046 ( 
.A1(n_10120),
.A2(n_8467),
.B(n_8887),
.Y(n_11046)
);

INVx2_ASAP7_75t_L g11047 ( 
.A(n_9984),
.Y(n_11047)
);

INVx2_ASAP7_75t_L g11048 ( 
.A(n_9984),
.Y(n_11048)
);

HB1xp67_ASAP7_75t_L g11049 ( 
.A(n_10317),
.Y(n_11049)
);

INVx1_ASAP7_75t_L g11050 ( 
.A(n_9385),
.Y(n_11050)
);

NAND2xp5_ASAP7_75t_L g11051 ( 
.A(n_10457),
.B(n_9309),
.Y(n_11051)
);

OR2x2_ASAP7_75t_L g11052 ( 
.A(n_9928),
.B(n_8474),
.Y(n_11052)
);

NAND2xp5_ASAP7_75t_L g11053 ( 
.A(n_9595),
.B(n_9309),
.Y(n_11053)
);

AOI21xp33_ASAP7_75t_SL g11054 ( 
.A1(n_10157),
.A2(n_9275),
.B(n_9195),
.Y(n_11054)
);

AND2x2_ASAP7_75t_L g11055 ( 
.A(n_9535),
.B(n_8956),
.Y(n_11055)
);

AOI22xp5_ASAP7_75t_SL g11056 ( 
.A1(n_9375),
.A2(n_9005),
.B1(n_9149),
.B2(n_9056),
.Y(n_11056)
);

AO21x1_ASAP7_75t_L g11057 ( 
.A1(n_10531),
.A2(n_9155),
.B(n_8787),
.Y(n_11057)
);

BUFx6f_ASAP7_75t_L g11058 ( 
.A(n_9395),
.Y(n_11058)
);

INVx2_ASAP7_75t_L g11059 ( 
.A(n_10595),
.Y(n_11059)
);

INVx1_ASAP7_75t_L g11060 ( 
.A(n_9398),
.Y(n_11060)
);

OR2x2_ASAP7_75t_L g11061 ( 
.A(n_10098),
.B(n_8474),
.Y(n_11061)
);

INVx1_ASAP7_75t_L g11062 ( 
.A(n_9413),
.Y(n_11062)
);

INVx2_ASAP7_75t_SL g11063 ( 
.A(n_9961),
.Y(n_11063)
);

INVx1_ASAP7_75t_L g11064 ( 
.A(n_9413),
.Y(n_11064)
);

INVx2_ASAP7_75t_L g11065 ( 
.A(n_10595),
.Y(n_11065)
);

INVx2_ASAP7_75t_L g11066 ( 
.A(n_10636),
.Y(n_11066)
);

OAI21x1_ASAP7_75t_L g11067 ( 
.A1(n_10120),
.A2(n_8467),
.B(n_8887),
.Y(n_11067)
);

CKINVDCx12_ASAP7_75t_R g11068 ( 
.A(n_9943),
.Y(n_11068)
);

OAI21x1_ASAP7_75t_L g11069 ( 
.A1(n_10636),
.A2(n_8897),
.B(n_8887),
.Y(n_11069)
);

INVx1_ASAP7_75t_L g11070 ( 
.A(n_9433),
.Y(n_11070)
);

OAI21x1_ASAP7_75t_L g11071 ( 
.A1(n_9370),
.A2(n_8897),
.B(n_8887),
.Y(n_11071)
);

INVx1_ASAP7_75t_L g11072 ( 
.A(n_9433),
.Y(n_11072)
);

BUFx3_ASAP7_75t_L g11073 ( 
.A(n_9998),
.Y(n_11073)
);

BUFx2_ASAP7_75t_L g11074 ( 
.A(n_9331),
.Y(n_11074)
);

INVx1_ASAP7_75t_L g11075 ( 
.A(n_9448),
.Y(n_11075)
);

INVx2_ASAP7_75t_L g11076 ( 
.A(n_10133),
.Y(n_11076)
);

OAI22xp5_ASAP7_75t_L g11077 ( 
.A1(n_9455),
.A2(n_8771),
.B1(n_8450),
.B2(n_8621),
.Y(n_11077)
);

BUFx3_ASAP7_75t_L g11078 ( 
.A(n_9751),
.Y(n_11078)
);

INVx2_ASAP7_75t_L g11079 ( 
.A(n_10133),
.Y(n_11079)
);

NOR2xp33_ASAP7_75t_L g11080 ( 
.A(n_9331),
.B(n_9005),
.Y(n_11080)
);

OAI22xp5_ASAP7_75t_L g11081 ( 
.A1(n_9873),
.A2(n_8450),
.B1(n_8621),
.B2(n_8505),
.Y(n_11081)
);

INVx1_ASAP7_75t_L g11082 ( 
.A(n_9448),
.Y(n_11082)
);

INVx1_ASAP7_75t_L g11083 ( 
.A(n_9547),
.Y(n_11083)
);

BUFx3_ASAP7_75t_L g11084 ( 
.A(n_9866),
.Y(n_11084)
);

INVx1_ASAP7_75t_L g11085 ( 
.A(n_9547),
.Y(n_11085)
);

INVx3_ASAP7_75t_L g11086 ( 
.A(n_10243),
.Y(n_11086)
);

NOR2xp33_ASAP7_75t_L g11087 ( 
.A(n_9331),
.B(n_9357),
.Y(n_11087)
);

BUFx2_ASAP7_75t_L g11088 ( 
.A(n_9331),
.Y(n_11088)
);

NAND2xp5_ASAP7_75t_L g11089 ( 
.A(n_10113),
.B(n_9546),
.Y(n_11089)
);

OR2x2_ASAP7_75t_L g11090 ( 
.A(n_10248),
.B(n_8474),
.Y(n_11090)
);

NAND2xp5_ASAP7_75t_L g11091 ( 
.A(n_9612),
.B(n_8128),
.Y(n_11091)
);

INVx3_ASAP7_75t_L g11092 ( 
.A(n_10243),
.Y(n_11092)
);

INVx1_ASAP7_75t_L g11093 ( 
.A(n_9549),
.Y(n_11093)
);

OAI22xp5_ASAP7_75t_L g11094 ( 
.A1(n_9315),
.A2(n_8865),
.B1(n_8712),
.B2(n_8811),
.Y(n_11094)
);

INVx3_ASAP7_75t_L g11095 ( 
.A(n_10593),
.Y(n_11095)
);

OAI21x1_ASAP7_75t_L g11096 ( 
.A1(n_9370),
.A2(n_8901),
.B(n_8897),
.Y(n_11096)
);

INVx2_ASAP7_75t_L g11097 ( 
.A(n_10133),
.Y(n_11097)
);

INVx1_ASAP7_75t_L g11098 ( 
.A(n_9366),
.Y(n_11098)
);

OAI21x1_ASAP7_75t_L g11099 ( 
.A1(n_9461),
.A2(n_8901),
.B(n_8897),
.Y(n_11099)
);

INVx1_ASAP7_75t_L g11100 ( 
.A(n_9367),
.Y(n_11100)
);

INVx2_ASAP7_75t_L g11101 ( 
.A(n_10144),
.Y(n_11101)
);

HB1xp67_ASAP7_75t_L g11102 ( 
.A(n_10319),
.Y(n_11102)
);

AND2x2_ASAP7_75t_L g11103 ( 
.A(n_9535),
.B(n_9005),
.Y(n_11103)
);

INVx1_ASAP7_75t_L g11104 ( 
.A(n_9367),
.Y(n_11104)
);

AOI21x1_ASAP7_75t_L g11105 ( 
.A1(n_9503),
.A2(n_8971),
.B(n_8914),
.Y(n_11105)
);

INVx1_ASAP7_75t_L g11106 ( 
.A(n_9495),
.Y(n_11106)
);

NAND2xp5_ASAP7_75t_L g11107 ( 
.A(n_9399),
.B(n_8128),
.Y(n_11107)
);

INVx2_ASAP7_75t_L g11108 ( 
.A(n_10144),
.Y(n_11108)
);

INVx1_ASAP7_75t_L g11109 ( 
.A(n_9430),
.Y(n_11109)
);

INVx2_ASAP7_75t_L g11110 ( 
.A(n_10144),
.Y(n_11110)
);

INVx2_ASAP7_75t_L g11111 ( 
.A(n_10153),
.Y(n_11111)
);

INVx1_ASAP7_75t_L g11112 ( 
.A(n_9430),
.Y(n_11112)
);

INVx1_ASAP7_75t_L g11113 ( 
.A(n_9431),
.Y(n_11113)
);

NOR2xp33_ASAP7_75t_L g11114 ( 
.A(n_9331),
.B(n_9005),
.Y(n_11114)
);

INVx1_ASAP7_75t_L g11115 ( 
.A(n_9431),
.Y(n_11115)
);

INVx1_ASAP7_75t_L g11116 ( 
.A(n_9536),
.Y(n_11116)
);

BUFx2_ASAP7_75t_L g11117 ( 
.A(n_9331),
.Y(n_11117)
);

INVx1_ASAP7_75t_L g11118 ( 
.A(n_9337),
.Y(n_11118)
);

BUFx6f_ASAP7_75t_L g11119 ( 
.A(n_9395),
.Y(n_11119)
);

INVx1_ASAP7_75t_L g11120 ( 
.A(n_9337),
.Y(n_11120)
);

INVx2_ASAP7_75t_L g11121 ( 
.A(n_10153),
.Y(n_11121)
);

OA21x2_ASAP7_75t_L g11122 ( 
.A1(n_10576),
.A2(n_7964),
.B(n_7955),
.Y(n_11122)
);

AO21x2_ASAP7_75t_L g11123 ( 
.A1(n_10548),
.A2(n_8669),
.B(n_8231),
.Y(n_11123)
);

NOR2xp33_ASAP7_75t_L g11124 ( 
.A(n_9357),
.B(n_9056),
.Y(n_11124)
);

INVx1_ASAP7_75t_L g11125 ( 
.A(n_9631),
.Y(n_11125)
);

OR2x2_ASAP7_75t_L g11126 ( 
.A(n_10263),
.B(n_8474),
.Y(n_11126)
);

AND2x2_ASAP7_75t_L g11127 ( 
.A(n_9535),
.B(n_9056),
.Y(n_11127)
);

AOI221xp5_ASAP7_75t_L g11128 ( 
.A1(n_10278),
.A2(n_8848),
.B1(n_8453),
.B2(n_8950),
.C(n_8835),
.Y(n_11128)
);

INVx1_ASAP7_75t_L g11129 ( 
.A(n_9631),
.Y(n_11129)
);

AND2x2_ASAP7_75t_L g11130 ( 
.A(n_9535),
.B(n_9056),
.Y(n_11130)
);

HB1xp67_ASAP7_75t_L g11131 ( 
.A(n_10333),
.Y(n_11131)
);

CKINVDCx14_ASAP7_75t_R g11132 ( 
.A(n_10033),
.Y(n_11132)
);

INVx3_ASAP7_75t_L g11133 ( 
.A(n_10593),
.Y(n_11133)
);

OAI21x1_ASAP7_75t_L g11134 ( 
.A1(n_9461),
.A2(n_8908),
.B(n_8901),
.Y(n_11134)
);

NAND2x1_ASAP7_75t_L g11135 ( 
.A(n_10000),
.B(n_10115),
.Y(n_11135)
);

INVx1_ASAP7_75t_L g11136 ( 
.A(n_9522),
.Y(n_11136)
);

INVx1_ASAP7_75t_L g11137 ( 
.A(n_9522),
.Y(n_11137)
);

BUFx3_ASAP7_75t_L g11138 ( 
.A(n_9866),
.Y(n_11138)
);

INVx2_ASAP7_75t_L g11139 ( 
.A(n_10153),
.Y(n_11139)
);

AND2x2_ASAP7_75t_L g11140 ( 
.A(n_9776),
.B(n_9149),
.Y(n_11140)
);

NAND2x1p5_ASAP7_75t_L g11141 ( 
.A(n_10593),
.B(n_8764),
.Y(n_11141)
);

INVx1_ASAP7_75t_L g11142 ( 
.A(n_9532),
.Y(n_11142)
);

OAI21x1_ASAP7_75t_L g11143 ( 
.A1(n_9592),
.A2(n_8908),
.B(n_8901),
.Y(n_11143)
);

CKINVDCx8_ASAP7_75t_R g11144 ( 
.A(n_10176),
.Y(n_11144)
);

HB1xp67_ASAP7_75t_L g11145 ( 
.A(n_10380),
.Y(n_11145)
);

INVx1_ASAP7_75t_L g11146 ( 
.A(n_9532),
.Y(n_11146)
);

OR2x6_ASAP7_75t_L g11147 ( 
.A(n_10065),
.B(n_9278),
.Y(n_11147)
);

INVx1_ASAP7_75t_L g11148 ( 
.A(n_9609),
.Y(n_11148)
);

NAND2xp5_ASAP7_75t_L g11149 ( 
.A(n_9334),
.B(n_8144),
.Y(n_11149)
);

INVx1_ASAP7_75t_L g11150 ( 
.A(n_9385),
.Y(n_11150)
);

INVx2_ASAP7_75t_L g11151 ( 
.A(n_10170),
.Y(n_11151)
);

HB1xp67_ASAP7_75t_L g11152 ( 
.A(n_10385),
.Y(n_11152)
);

INVx2_ASAP7_75t_SL g11153 ( 
.A(n_9961),
.Y(n_11153)
);

INVx1_ASAP7_75t_L g11154 ( 
.A(n_9438),
.Y(n_11154)
);

INVx1_ASAP7_75t_L g11155 ( 
.A(n_9438),
.Y(n_11155)
);

INVx1_ASAP7_75t_L g11156 ( 
.A(n_9486),
.Y(n_11156)
);

INVx3_ASAP7_75t_L g11157 ( 
.A(n_10593),
.Y(n_11157)
);

AND2x4_ASAP7_75t_L g11158 ( 
.A(n_10593),
.B(n_8764),
.Y(n_11158)
);

INVx1_ASAP7_75t_L g11159 ( 
.A(n_9509),
.Y(n_11159)
);

INVx2_ASAP7_75t_L g11160 ( 
.A(n_10170),
.Y(n_11160)
);

BUFx2_ASAP7_75t_L g11161 ( 
.A(n_9357),
.Y(n_11161)
);

INVx2_ASAP7_75t_SL g11162 ( 
.A(n_10222),
.Y(n_11162)
);

INVx1_ASAP7_75t_L g11163 ( 
.A(n_9509),
.Y(n_11163)
);

INVx1_ASAP7_75t_L g11164 ( 
.A(n_9597),
.Y(n_11164)
);

INVx3_ASAP7_75t_L g11165 ( 
.A(n_10593),
.Y(n_11165)
);

INVx1_ASAP7_75t_L g11166 ( 
.A(n_9597),
.Y(n_11166)
);

INVx1_ASAP7_75t_L g11167 ( 
.A(n_9635),
.Y(n_11167)
);

INVx2_ASAP7_75t_SL g11168 ( 
.A(n_10222),
.Y(n_11168)
);

OAI21x1_ASAP7_75t_L g11169 ( 
.A1(n_9592),
.A2(n_8927),
.B(n_8908),
.Y(n_11169)
);

INVx1_ASAP7_75t_L g11170 ( 
.A(n_9636),
.Y(n_11170)
);

AOI21xp33_ASAP7_75t_L g11171 ( 
.A1(n_9876),
.A2(n_8787),
.B(n_8659),
.Y(n_11171)
);

AND2x2_ASAP7_75t_L g11172 ( 
.A(n_9776),
.B(n_9149),
.Y(n_11172)
);

INVx2_ASAP7_75t_L g11173 ( 
.A(n_10170),
.Y(n_11173)
);

INVx3_ASAP7_75t_L g11174 ( 
.A(n_10651),
.Y(n_11174)
);

AOI22xp5_ASAP7_75t_L g11175 ( 
.A1(n_9316),
.A2(n_8605),
.B1(n_8594),
.B2(n_9148),
.Y(n_11175)
);

INVx1_ASAP7_75t_L g11176 ( 
.A(n_9578),
.Y(n_11176)
);

INVx4_ASAP7_75t_L g11177 ( 
.A(n_9341),
.Y(n_11177)
);

NAND2xp5_ASAP7_75t_L g11178 ( 
.A(n_9368),
.B(n_8144),
.Y(n_11178)
);

INVx1_ASAP7_75t_L g11179 ( 
.A(n_9579),
.Y(n_11179)
);

AND2x2_ASAP7_75t_L g11180 ( 
.A(n_9776),
.B(n_9149),
.Y(n_11180)
);

HB1xp67_ASAP7_75t_L g11181 ( 
.A(n_10393),
.Y(n_11181)
);

BUFx2_ASAP7_75t_L g11182 ( 
.A(n_9357),
.Y(n_11182)
);

AOI21xp5_ASAP7_75t_L g11183 ( 
.A1(n_10557),
.A2(n_8515),
.B(n_8869),
.Y(n_11183)
);

AND2x2_ASAP7_75t_L g11184 ( 
.A(n_9776),
.B(n_9270),
.Y(n_11184)
);

INVx1_ASAP7_75t_L g11185 ( 
.A(n_9579),
.Y(n_11185)
);

INVx1_ASAP7_75t_L g11186 ( 
.A(n_9639),
.Y(n_11186)
);

NAND2xp5_ASAP7_75t_L g11187 ( 
.A(n_9835),
.B(n_8158),
.Y(n_11187)
);

INVx3_ASAP7_75t_L g11188 ( 
.A(n_10651),
.Y(n_11188)
);

OAI22xp5_ASAP7_75t_SL g11189 ( 
.A1(n_10364),
.A2(n_7784),
.B1(n_7517),
.B2(n_7785),
.Y(n_11189)
);

INVx3_ASAP7_75t_L g11190 ( 
.A(n_10651),
.Y(n_11190)
);

HB1xp67_ASAP7_75t_SL g11191 ( 
.A(n_9892),
.Y(n_11191)
);

INVx2_ASAP7_75t_L g11192 ( 
.A(n_10180),
.Y(n_11192)
);

INVx1_ASAP7_75t_L g11193 ( 
.A(n_9639),
.Y(n_11193)
);

OA21x2_ASAP7_75t_L g11194 ( 
.A1(n_10645),
.A2(n_7993),
.B(n_7983),
.Y(n_11194)
);

NOR2xp33_ASAP7_75t_L g11195 ( 
.A(n_9357),
.B(n_9270),
.Y(n_11195)
);

INVx1_ASAP7_75t_L g11196 ( 
.A(n_9656),
.Y(n_11196)
);

OAI21x1_ASAP7_75t_L g11197 ( 
.A1(n_9655),
.A2(n_8927),
.B(n_8908),
.Y(n_11197)
);

INVx1_ASAP7_75t_L g11198 ( 
.A(n_9656),
.Y(n_11198)
);

BUFx2_ASAP7_75t_L g11199 ( 
.A(n_9357),
.Y(n_11199)
);

INVx1_ASAP7_75t_L g11200 ( 
.A(n_9362),
.Y(n_11200)
);

INVx1_ASAP7_75t_L g11201 ( 
.A(n_9362),
.Y(n_11201)
);

AO21x2_ASAP7_75t_L g11202 ( 
.A1(n_9876),
.A2(n_8231),
.B(n_9155),
.Y(n_11202)
);

INVx3_ASAP7_75t_L g11203 ( 
.A(n_10720),
.Y(n_11203)
);

HB1xp67_ASAP7_75t_L g11204 ( 
.A(n_10403),
.Y(n_11204)
);

INVx2_ASAP7_75t_L g11205 ( 
.A(n_10180),
.Y(n_11205)
);

BUFx12f_ASAP7_75t_L g11206 ( 
.A(n_9432),
.Y(n_11206)
);

INVx1_ASAP7_75t_L g11207 ( 
.A(n_9380),
.Y(n_11207)
);

INVx4_ASAP7_75t_L g11208 ( 
.A(n_9341),
.Y(n_11208)
);

INVx3_ASAP7_75t_L g11209 ( 
.A(n_10720),
.Y(n_11209)
);

INVx1_ASAP7_75t_L g11210 ( 
.A(n_9423),
.Y(n_11210)
);

INVx1_ASAP7_75t_L g11211 ( 
.A(n_9423),
.Y(n_11211)
);

INVxp33_ASAP7_75t_L g11212 ( 
.A(n_9943),
.Y(n_11212)
);

INVx1_ASAP7_75t_L g11213 ( 
.A(n_9517),
.Y(n_11213)
);

INVx2_ASAP7_75t_L g11214 ( 
.A(n_10180),
.Y(n_11214)
);

OAI21xp5_ASAP7_75t_L g11215 ( 
.A1(n_10240),
.A2(n_8256),
.B(n_8278),
.Y(n_11215)
);

BUFx2_ASAP7_75t_L g11216 ( 
.A(n_9919),
.Y(n_11216)
);

AND2x4_ASAP7_75t_L g11217 ( 
.A(n_9339),
.B(n_8764),
.Y(n_11217)
);

INVx1_ASAP7_75t_L g11218 ( 
.A(n_9517),
.Y(n_11218)
);

AO21x1_ASAP7_75t_SL g11219 ( 
.A1(n_9577),
.A2(n_10715),
.B(n_10164),
.Y(n_11219)
);

BUFx2_ASAP7_75t_L g11220 ( 
.A(n_9919),
.Y(n_11220)
);

INVx1_ASAP7_75t_L g11221 ( 
.A(n_9578),
.Y(n_11221)
);

INVx1_ASAP7_75t_L g11222 ( 
.A(n_9657),
.Y(n_11222)
);

INVx2_ASAP7_75t_L g11223 ( 
.A(n_10247),
.Y(n_11223)
);

BUFx2_ASAP7_75t_L g11224 ( 
.A(n_9919),
.Y(n_11224)
);

CKINVDCx11_ASAP7_75t_R g11225 ( 
.A(n_10567),
.Y(n_11225)
);

AND2x2_ASAP7_75t_L g11226 ( 
.A(n_9802),
.B(n_9270),
.Y(n_11226)
);

INVx2_ASAP7_75t_L g11227 ( 
.A(n_10247),
.Y(n_11227)
);

AOI21x1_ASAP7_75t_L g11228 ( 
.A1(n_9503),
.A2(n_10045),
.B(n_10201),
.Y(n_11228)
);

INVx3_ASAP7_75t_L g11229 ( 
.A(n_10720),
.Y(n_11229)
);

INVx1_ASAP7_75t_L g11230 ( 
.A(n_9581),
.Y(n_11230)
);

INVx2_ASAP7_75t_SL g11231 ( 
.A(n_10222),
.Y(n_11231)
);

INVxp67_ASAP7_75t_SL g11232 ( 
.A(n_9605),
.Y(n_11232)
);

AO21x2_ASAP7_75t_L g11233 ( 
.A1(n_10666),
.A2(n_8534),
.B(n_8260),
.Y(n_11233)
);

INVx1_ASAP7_75t_L g11234 ( 
.A(n_9581),
.Y(n_11234)
);

INVx1_ASAP7_75t_L g11235 ( 
.A(n_9582),
.Y(n_11235)
);

HB1xp67_ASAP7_75t_L g11236 ( 
.A(n_10409),
.Y(n_11236)
);

CKINVDCx5p33_ASAP7_75t_R g11237 ( 
.A(n_9755),
.Y(n_11237)
);

INVx3_ASAP7_75t_L g11238 ( 
.A(n_10472),
.Y(n_11238)
);

INVx2_ASAP7_75t_SL g11239 ( 
.A(n_10222),
.Y(n_11239)
);

INVx1_ASAP7_75t_SL g11240 ( 
.A(n_9978),
.Y(n_11240)
);

AND2x2_ASAP7_75t_L g11241 ( 
.A(n_9802),
.B(n_9270),
.Y(n_11241)
);

INVx1_ASAP7_75t_L g11242 ( 
.A(n_9582),
.Y(n_11242)
);

INVx1_ASAP7_75t_L g11243 ( 
.A(n_9635),
.Y(n_11243)
);

INVx1_ASAP7_75t_L g11244 ( 
.A(n_9636),
.Y(n_11244)
);

INVx2_ASAP7_75t_L g11245 ( 
.A(n_10255),
.Y(n_11245)
);

INVx1_ASAP7_75t_L g11246 ( 
.A(n_9697),
.Y(n_11246)
);

BUFx2_ASAP7_75t_L g11247 ( 
.A(n_9919),
.Y(n_11247)
);

BUFx3_ASAP7_75t_L g11248 ( 
.A(n_9981),
.Y(n_11248)
);

INVx1_ASAP7_75t_L g11249 ( 
.A(n_9697),
.Y(n_11249)
);

INVx1_ASAP7_75t_L g11250 ( 
.A(n_9732),
.Y(n_11250)
);

INVx2_ASAP7_75t_L g11251 ( 
.A(n_10255),
.Y(n_11251)
);

INVx1_ASAP7_75t_L g11252 ( 
.A(n_9732),
.Y(n_11252)
);

INVx2_ASAP7_75t_L g11253 ( 
.A(n_10336),
.Y(n_11253)
);

INVx2_ASAP7_75t_L g11254 ( 
.A(n_10336),
.Y(n_11254)
);

AOI21x1_ASAP7_75t_L g11255 ( 
.A1(n_10045),
.A2(n_8971),
.B(n_8914),
.Y(n_11255)
);

AND2x2_ASAP7_75t_L g11256 ( 
.A(n_9802),
.B(n_9200),
.Y(n_11256)
);

INVx2_ASAP7_75t_L g11257 ( 
.A(n_10183),
.Y(n_11257)
);

BUFx2_ASAP7_75t_L g11258 ( 
.A(n_10026),
.Y(n_11258)
);

INVx3_ASAP7_75t_L g11259 ( 
.A(n_10472),
.Y(n_11259)
);

INVx2_ASAP7_75t_L g11260 ( 
.A(n_10183),
.Y(n_11260)
);

INVx1_ASAP7_75t_L g11261 ( 
.A(n_9752),
.Y(n_11261)
);

INVx1_ASAP7_75t_L g11262 ( 
.A(n_9753),
.Y(n_11262)
);

INVx1_ASAP7_75t_L g11263 ( 
.A(n_9753),
.Y(n_11263)
);

OA21x2_ASAP7_75t_L g11264 ( 
.A1(n_9378),
.A2(n_7993),
.B(n_7983),
.Y(n_11264)
);

BUFx3_ASAP7_75t_L g11265 ( 
.A(n_9981),
.Y(n_11265)
);

INVx1_ASAP7_75t_L g11266 ( 
.A(n_9771),
.Y(n_11266)
);

INVx1_ASAP7_75t_SL g11267 ( 
.A(n_9699),
.Y(n_11267)
);

INVx3_ASAP7_75t_L g11268 ( 
.A(n_10493),
.Y(n_11268)
);

AO21x2_ASAP7_75t_L g11269 ( 
.A1(n_10666),
.A2(n_8534),
.B(n_8260),
.Y(n_11269)
);

BUFx6f_ASAP7_75t_L g11270 ( 
.A(n_9395),
.Y(n_11270)
);

AND2x2_ASAP7_75t_L g11271 ( 
.A(n_9802),
.B(n_9200),
.Y(n_11271)
);

INVx1_ASAP7_75t_L g11272 ( 
.A(n_9756),
.Y(n_11272)
);

INVx1_ASAP7_75t_L g11273 ( 
.A(n_9756),
.Y(n_11273)
);

NOR2x1_ASAP7_75t_SL g11274 ( 
.A(n_9784),
.B(n_9277),
.Y(n_11274)
);

INVx1_ASAP7_75t_L g11275 ( 
.A(n_9757),
.Y(n_11275)
);

INVx3_ASAP7_75t_L g11276 ( 
.A(n_10493),
.Y(n_11276)
);

BUFx2_ASAP7_75t_L g11277 ( 
.A(n_10026),
.Y(n_11277)
);

INVx2_ASAP7_75t_SL g11278 ( 
.A(n_10203),
.Y(n_11278)
);

INVx1_ASAP7_75t_L g11279 ( 
.A(n_9757),
.Y(n_11279)
);

INVx2_ASAP7_75t_L g11280 ( 
.A(n_10183),
.Y(n_11280)
);

INVx2_ASAP7_75t_L g11281 ( 
.A(n_10549),
.Y(n_11281)
);

INVx2_ASAP7_75t_L g11282 ( 
.A(n_10549),
.Y(n_11282)
);

INVx1_ASAP7_75t_L g11283 ( 
.A(n_9825),
.Y(n_11283)
);

OAI21x1_ASAP7_75t_L g11284 ( 
.A1(n_9655),
.A2(n_8927),
.B(n_8582),
.Y(n_11284)
);

INVx1_ASAP7_75t_SL g11285 ( 
.A(n_9739),
.Y(n_11285)
);

INVx1_ASAP7_75t_L g11286 ( 
.A(n_9717),
.Y(n_11286)
);

HB1xp67_ASAP7_75t_L g11287 ( 
.A(n_10516),
.Y(n_11287)
);

INVx2_ASAP7_75t_L g11288 ( 
.A(n_10549),
.Y(n_11288)
);

INVx2_ASAP7_75t_L g11289 ( 
.A(n_9738),
.Y(n_11289)
);

INVx1_ASAP7_75t_L g11290 ( 
.A(n_9717),
.Y(n_11290)
);

CKINVDCx20_ASAP7_75t_R g11291 ( 
.A(n_10172),
.Y(n_11291)
);

OR2x2_ASAP7_75t_L g11292 ( 
.A(n_10270),
.B(n_8474),
.Y(n_11292)
);

OAI21x1_ASAP7_75t_L g11293 ( 
.A1(n_9779),
.A2(n_8927),
.B(n_8582),
.Y(n_11293)
);

NAND2xp5_ASAP7_75t_L g11294 ( 
.A(n_9868),
.B(n_8158),
.Y(n_11294)
);

INVx2_ASAP7_75t_L g11295 ( 
.A(n_9738),
.Y(n_11295)
);

INVx3_ASAP7_75t_L g11296 ( 
.A(n_10493),
.Y(n_11296)
);

INVx1_ASAP7_75t_L g11297 ( 
.A(n_9737),
.Y(n_11297)
);

INVx1_ASAP7_75t_L g11298 ( 
.A(n_9737),
.Y(n_11298)
);

BUFx2_ASAP7_75t_L g11299 ( 
.A(n_10026),
.Y(n_11299)
);

INVx2_ASAP7_75t_L g11300 ( 
.A(n_9804),
.Y(n_11300)
);

INVx2_ASAP7_75t_L g11301 ( 
.A(n_9804),
.Y(n_11301)
);

INVx2_ASAP7_75t_L g11302 ( 
.A(n_9832),
.Y(n_11302)
);

INVx2_ASAP7_75t_L g11303 ( 
.A(n_9832),
.Y(n_11303)
);

OAI22xp5_ASAP7_75t_SL g11304 ( 
.A1(n_10400),
.A2(n_7517),
.B1(n_7785),
.B2(n_6730),
.Y(n_11304)
);

INVx2_ASAP7_75t_L g11305 ( 
.A(n_10057),
.Y(n_11305)
);

INVx1_ASAP7_75t_L g11306 ( 
.A(n_9740),
.Y(n_11306)
);

INVx1_ASAP7_75t_L g11307 ( 
.A(n_9740),
.Y(n_11307)
);

OAI22xp5_ASAP7_75t_SL g11308 ( 
.A1(n_9343),
.A2(n_7785),
.B1(n_6730),
.B2(n_6677),
.Y(n_11308)
);

OAI21xp5_ASAP7_75t_L g11309 ( 
.A1(n_10715),
.A2(n_8256),
.B(n_8865),
.Y(n_11309)
);

NAND2x1p5_ASAP7_75t_L g11310 ( 
.A(n_10188),
.B(n_8764),
.Y(n_11310)
);

INVx1_ASAP7_75t_L g11311 ( 
.A(n_9772),
.Y(n_11311)
);

OR2x2_ASAP7_75t_L g11312 ( 
.A(n_10318),
.B(n_8474),
.Y(n_11312)
);

BUFx2_ASAP7_75t_L g11313 ( 
.A(n_10026),
.Y(n_11313)
);

INVx3_ASAP7_75t_L g11314 ( 
.A(n_10493),
.Y(n_11314)
);

HB1xp67_ASAP7_75t_L g11315 ( 
.A(n_10527),
.Y(n_11315)
);

INVx1_ASAP7_75t_L g11316 ( 
.A(n_9772),
.Y(n_11316)
);

HB1xp67_ASAP7_75t_L g11317 ( 
.A(n_10552),
.Y(n_11317)
);

OAI22xp33_ASAP7_75t_L g11318 ( 
.A1(n_9541),
.A2(n_9236),
.B1(n_8558),
.B2(n_8570),
.Y(n_11318)
);

BUFx6f_ASAP7_75t_L g11319 ( 
.A(n_9395),
.Y(n_11319)
);

NOR2xp33_ASAP7_75t_L g11320 ( 
.A(n_9343),
.B(n_8888),
.Y(n_11320)
);

BUFx2_ASAP7_75t_L g11321 ( 
.A(n_10138),
.Y(n_11321)
);

NAND2xp5_ASAP7_75t_L g11322 ( 
.A(n_10052),
.B(n_8165),
.Y(n_11322)
);

OAI21x1_ASAP7_75t_L g11323 ( 
.A1(n_9779),
.A2(n_8582),
.B(n_8565),
.Y(n_11323)
);

INVx1_ASAP7_75t_L g11324 ( 
.A(n_9657),
.Y(n_11324)
);

INVx2_ASAP7_75t_L g11325 ( 
.A(n_10057),
.Y(n_11325)
);

AND2x4_ASAP7_75t_L g11326 ( 
.A(n_9339),
.B(n_8788),
.Y(n_11326)
);

INVx1_ASAP7_75t_L g11327 ( 
.A(n_9666),
.Y(n_11327)
);

INVx1_ASAP7_75t_L g11328 ( 
.A(n_9666),
.Y(n_11328)
);

INVx4_ASAP7_75t_L g11329 ( 
.A(n_9416),
.Y(n_11329)
);

INVx1_ASAP7_75t_L g11330 ( 
.A(n_9667),
.Y(n_11330)
);

BUFx3_ASAP7_75t_L g11331 ( 
.A(n_9355),
.Y(n_11331)
);

INVx1_ASAP7_75t_L g11332 ( 
.A(n_9609),
.Y(n_11332)
);

BUFx2_ASAP7_75t_L g11333 ( 
.A(n_10138),
.Y(n_11333)
);

INVxp67_ASAP7_75t_SL g11334 ( 
.A(n_9480),
.Y(n_11334)
);

NAND2x1_ASAP7_75t_L g11335 ( 
.A(n_10000),
.B(n_8260),
.Y(n_11335)
);

INVx1_ASAP7_75t_L g11336 ( 
.A(n_9573),
.Y(n_11336)
);

INVx2_ASAP7_75t_L g11337 ( 
.A(n_9319),
.Y(n_11337)
);

BUFx2_ASAP7_75t_L g11338 ( 
.A(n_10138),
.Y(n_11338)
);

INVx2_ASAP7_75t_L g11339 ( 
.A(n_9319),
.Y(n_11339)
);

INVx2_ASAP7_75t_L g11340 ( 
.A(n_9329),
.Y(n_11340)
);

HB1xp67_ASAP7_75t_L g11341 ( 
.A(n_10572),
.Y(n_11341)
);

INVx2_ASAP7_75t_L g11342 ( 
.A(n_9329),
.Y(n_11342)
);

OAI21x1_ASAP7_75t_L g11343 ( 
.A1(n_9826),
.A2(n_8582),
.B(n_8565),
.Y(n_11343)
);

INVx1_ASAP7_75t_L g11344 ( 
.A(n_9549),
.Y(n_11344)
);

BUFx2_ASAP7_75t_L g11345 ( 
.A(n_10138),
.Y(n_11345)
);

AND2x2_ASAP7_75t_L g11346 ( 
.A(n_9831),
.B(n_9240),
.Y(n_11346)
);

INVx2_ASAP7_75t_L g11347 ( 
.A(n_9380),
.Y(n_11347)
);

OAI21x1_ASAP7_75t_L g11348 ( 
.A1(n_9826),
.A2(n_8585),
.B(n_8565),
.Y(n_11348)
);

INVx2_ASAP7_75t_L g11349 ( 
.A(n_9495),
.Y(n_11349)
);

INVx3_ASAP7_75t_L g11350 ( 
.A(n_10540),
.Y(n_11350)
);

OAI21x1_ASAP7_75t_L g11351 ( 
.A1(n_10473),
.A2(n_10490),
.B(n_10474),
.Y(n_11351)
);

INVx1_ASAP7_75t_L g11352 ( 
.A(n_9667),
.Y(n_11352)
);

INVx2_ASAP7_75t_L g11353 ( 
.A(n_9526),
.Y(n_11353)
);

BUFx3_ASAP7_75t_L g11354 ( 
.A(n_9858),
.Y(n_11354)
);

INVx2_ASAP7_75t_L g11355 ( 
.A(n_9526),
.Y(n_11355)
);

INVx1_ASAP7_75t_L g11356 ( 
.A(n_9618),
.Y(n_11356)
);

AOI221xp5_ASAP7_75t_L g11357 ( 
.A1(n_10278),
.A2(n_8848),
.B1(n_8950),
.B2(n_8835),
.C(n_8611),
.Y(n_11357)
);

INVx1_ASAP7_75t_L g11358 ( 
.A(n_9618),
.Y(n_11358)
);

BUFx2_ASAP7_75t_L g11359 ( 
.A(n_10161),
.Y(n_11359)
);

OAI21x1_ASAP7_75t_L g11360 ( 
.A1(n_10473),
.A2(n_8585),
.B(n_8565),
.Y(n_11360)
);

INVx2_ASAP7_75t_L g11361 ( 
.A(n_9536),
.Y(n_11361)
);

OR2x2_ASAP7_75t_L g11362 ( 
.A(n_10323),
.B(n_8474),
.Y(n_11362)
);

NOR2xp67_ASAP7_75t_L g11363 ( 
.A(n_10703),
.B(n_9168),
.Y(n_11363)
);

AO21x2_ASAP7_75t_L g11364 ( 
.A1(n_10115),
.A2(n_8458),
.B(n_8300),
.Y(n_11364)
);

OAI21x1_ASAP7_75t_L g11365 ( 
.A1(n_10473),
.A2(n_10490),
.B(n_10474),
.Y(n_11365)
);

INVx1_ASAP7_75t_L g11366 ( 
.A(n_9726),
.Y(n_11366)
);

OAI21x1_ASAP7_75t_L g11367 ( 
.A1(n_10474),
.A2(n_8586),
.B(n_8585),
.Y(n_11367)
);

INVx2_ASAP7_75t_L g11368 ( 
.A(n_9573),
.Y(n_11368)
);

INVx1_ASAP7_75t_L g11369 ( 
.A(n_9643),
.Y(n_11369)
);

OAI22x1_ASAP7_75t_L g11370 ( 
.A1(n_10663),
.A2(n_9214),
.B1(n_9275),
.B2(n_9195),
.Y(n_11370)
);

INVxp67_ASAP7_75t_L g11371 ( 
.A(n_9768),
.Y(n_11371)
);

INVx1_ASAP7_75t_L g11372 ( 
.A(n_9643),
.Y(n_11372)
);

BUFx2_ASAP7_75t_L g11373 ( 
.A(n_10161),
.Y(n_11373)
);

INVx2_ASAP7_75t_L g11374 ( 
.A(n_9574),
.Y(n_11374)
);

AND2x2_ASAP7_75t_L g11375 ( 
.A(n_9831),
.B(n_9240),
.Y(n_11375)
);

OAI21x1_ASAP7_75t_L g11376 ( 
.A1(n_10490),
.A2(n_8586),
.B(n_8585),
.Y(n_11376)
);

HB1xp67_ASAP7_75t_L g11377 ( 
.A(n_10659),
.Y(n_11377)
);

INVx1_ASAP7_75t_L g11378 ( 
.A(n_9691),
.Y(n_11378)
);

INVx2_ASAP7_75t_L g11379 ( 
.A(n_9574),
.Y(n_11379)
);

INVx2_ASAP7_75t_L g11380 ( 
.A(n_9575),
.Y(n_11380)
);

NAND2xp5_ASAP7_75t_L g11381 ( 
.A(n_10063),
.B(n_8165),
.Y(n_11381)
);

INVx2_ASAP7_75t_L g11382 ( 
.A(n_9575),
.Y(n_11382)
);

INVx1_ASAP7_75t_L g11383 ( 
.A(n_9624),
.Y(n_11383)
);

AOI22xp33_ASAP7_75t_L g11384 ( 
.A1(n_10067),
.A2(n_7973),
.B1(n_8407),
.B2(n_8458),
.Y(n_11384)
);

INVx2_ASAP7_75t_L g11385 ( 
.A(n_9624),
.Y(n_11385)
);

INVx2_ASAP7_75t_L g11386 ( 
.A(n_9627),
.Y(n_11386)
);

BUFx2_ASAP7_75t_L g11387 ( 
.A(n_10161),
.Y(n_11387)
);

INVx1_ASAP7_75t_L g11388 ( 
.A(n_9713),
.Y(n_11388)
);

AND2x2_ASAP7_75t_L g11389 ( 
.A(n_9831),
.B(n_9244),
.Y(n_11389)
);

INVx1_ASAP7_75t_L g11390 ( 
.A(n_9713),
.Y(n_11390)
);

INVx1_ASAP7_75t_L g11391 ( 
.A(n_9846),
.Y(n_11391)
);

INVx3_ASAP7_75t_L g11392 ( 
.A(n_10540),
.Y(n_11392)
);

CKINVDCx5p33_ASAP7_75t_R g11393 ( 
.A(n_9513),
.Y(n_11393)
);

AND2x2_ASAP7_75t_L g11394 ( 
.A(n_9831),
.B(n_9244),
.Y(n_11394)
);

INVx1_ASAP7_75t_L g11395 ( 
.A(n_9659),
.Y(n_11395)
);

AOI211x1_ASAP7_75t_L g11396 ( 
.A1(n_9613),
.A2(n_9277),
.B(n_8772),
.C(n_8942),
.Y(n_11396)
);

INVx1_ASAP7_75t_L g11397 ( 
.A(n_9659),
.Y(n_11397)
);

AND2x4_ASAP7_75t_L g11398 ( 
.A(n_9339),
.B(n_8788),
.Y(n_11398)
);

INVx1_ASAP7_75t_L g11399 ( 
.A(n_9627),
.Y(n_11399)
);

AND2x4_ASAP7_75t_L g11400 ( 
.A(n_9384),
.B(n_8788),
.Y(n_11400)
);

OAI21x1_ASAP7_75t_L g11401 ( 
.A1(n_9669),
.A2(n_8593),
.B(n_8586),
.Y(n_11401)
);

AND2x2_ASAP7_75t_L g11402 ( 
.A(n_9949),
.B(n_8229),
.Y(n_11402)
);

NAND2xp5_ASAP7_75t_L g11403 ( 
.A(n_10080),
.B(n_8192),
.Y(n_11403)
);

AO31x2_ASAP7_75t_L g11404 ( 
.A1(n_10067),
.A2(n_8772),
.A3(n_8612),
.B(n_8566),
.Y(n_11404)
);

AOI22xp33_ASAP7_75t_SL g11405 ( 
.A1(n_10135),
.A2(n_7970),
.B1(n_8077),
.B2(n_8458),
.Y(n_11405)
);

HB1xp67_ASAP7_75t_L g11406 ( 
.A(n_10686),
.Y(n_11406)
);

OAI21x1_ASAP7_75t_L g11407 ( 
.A1(n_9669),
.A2(n_8593),
.B(n_8586),
.Y(n_11407)
);

NAND2xp5_ASAP7_75t_L g11408 ( 
.A(n_10094),
.B(n_8192),
.Y(n_11408)
);

HB1xp67_ASAP7_75t_L g11409 ( 
.A(n_10692),
.Y(n_11409)
);

NAND2xp5_ASAP7_75t_L g11410 ( 
.A(n_10121),
.B(n_8207),
.Y(n_11410)
);

OAI21x1_ASAP7_75t_L g11411 ( 
.A1(n_9669),
.A2(n_8601),
.B(n_8593),
.Y(n_11411)
);

OR2x2_ASAP7_75t_L g11412 ( 
.A(n_10335),
.B(n_8474),
.Y(n_11412)
);

INVx2_ASAP7_75t_SL g11413 ( 
.A(n_10203),
.Y(n_11413)
);

HB1xp67_ASAP7_75t_L g11414 ( 
.A(n_10696),
.Y(n_11414)
);

INVx2_ASAP7_75t_SL g11415 ( 
.A(n_9858),
.Y(n_11415)
);

BUFx3_ASAP7_75t_L g11416 ( 
.A(n_9858),
.Y(n_11416)
);

INVx2_ASAP7_75t_L g11417 ( 
.A(n_9651),
.Y(n_11417)
);

NOR2xp33_ASAP7_75t_SL g11418 ( 
.A(n_10060),
.B(n_8984),
.Y(n_11418)
);

INVx3_ASAP7_75t_L g11419 ( 
.A(n_10540),
.Y(n_11419)
);

INVx1_ASAP7_75t_L g11420 ( 
.A(n_9691),
.Y(n_11420)
);

HB1xp67_ASAP7_75t_L g11421 ( 
.A(n_10716),
.Y(n_11421)
);

INVx1_ASAP7_75t_L g11422 ( 
.A(n_9692),
.Y(n_11422)
);

CKINVDCx6p67_ASAP7_75t_R g11423 ( 
.A(n_9610),
.Y(n_11423)
);

AOI22xp33_ASAP7_75t_L g11424 ( 
.A1(n_9421),
.A2(n_7973),
.B1(n_8524),
.B2(n_7970),
.Y(n_11424)
);

INVx2_ASAP7_75t_L g11425 ( 
.A(n_9651),
.Y(n_11425)
);

INVx1_ASAP7_75t_L g11426 ( 
.A(n_9695),
.Y(n_11426)
);

INVx2_ASAP7_75t_L g11427 ( 
.A(n_9660),
.Y(n_11427)
);

INVx1_ASAP7_75t_L g11428 ( 
.A(n_9695),
.Y(n_11428)
);

INVx2_ASAP7_75t_L g11429 ( 
.A(n_9660),
.Y(n_11429)
);

INVx1_ASAP7_75t_SL g11430 ( 
.A(n_9543),
.Y(n_11430)
);

AND2x2_ASAP7_75t_L g11431 ( 
.A(n_9949),
.B(n_8229),
.Y(n_11431)
);

INVx1_ASAP7_75t_L g11432 ( 
.A(n_9688),
.Y(n_11432)
);

AND2x2_ASAP7_75t_L g11433 ( 
.A(n_9949),
.B(n_9973),
.Y(n_11433)
);

INVx2_ASAP7_75t_L g11434 ( 
.A(n_9676),
.Y(n_11434)
);

INVx1_ASAP7_75t_L g11435 ( 
.A(n_9777),
.Y(n_11435)
);

INVx1_ASAP7_75t_L g11436 ( 
.A(n_9777),
.Y(n_11436)
);

BUFx6f_ASAP7_75t_L g11437 ( 
.A(n_9416),
.Y(n_11437)
);

INVx1_ASAP7_75t_L g11438 ( 
.A(n_9822),
.Y(n_11438)
);

INVx2_ASAP7_75t_L g11439 ( 
.A(n_9676),
.Y(n_11439)
);

OAI21x1_ASAP7_75t_L g11440 ( 
.A1(n_9708),
.A2(n_8601),
.B(n_8593),
.Y(n_11440)
);

BUFx2_ASAP7_75t_L g11441 ( 
.A(n_10161),
.Y(n_11441)
);

INVx1_ASAP7_75t_L g11442 ( 
.A(n_9788),
.Y(n_11442)
);

AND2x2_ASAP7_75t_L g11443 ( 
.A(n_9949),
.B(n_8229),
.Y(n_11443)
);

INVx1_ASAP7_75t_L g11444 ( 
.A(n_9788),
.Y(n_11444)
);

INVx3_ASAP7_75t_L g11445 ( 
.A(n_10540),
.Y(n_11445)
);

BUFx3_ASAP7_75t_L g11446 ( 
.A(n_9858),
.Y(n_11446)
);

BUFx3_ASAP7_75t_L g11447 ( 
.A(n_9416),
.Y(n_11447)
);

INVx2_ASAP7_75t_L g11448 ( 
.A(n_9692),
.Y(n_11448)
);

INVx1_ASAP7_75t_L g11449 ( 
.A(n_9711),
.Y(n_11449)
);

INVx2_ASAP7_75t_L g11450 ( 
.A(n_9693),
.Y(n_11450)
);

INVx3_ASAP7_75t_L g11451 ( 
.A(n_10605),
.Y(n_11451)
);

INVx2_ASAP7_75t_L g11452 ( 
.A(n_9693),
.Y(n_11452)
);

HB1xp67_ASAP7_75t_L g11453 ( 
.A(n_10722),
.Y(n_11453)
);

INVx1_ASAP7_75t_L g11454 ( 
.A(n_9886),
.Y(n_11454)
);

INVx2_ASAP7_75t_L g11455 ( 
.A(n_9696),
.Y(n_11455)
);

BUFx2_ASAP7_75t_L g11456 ( 
.A(n_10244),
.Y(n_11456)
);

HB1xp67_ASAP7_75t_L g11457 ( 
.A(n_9494),
.Y(n_11457)
);

INVx1_ASAP7_75t_L g11458 ( 
.A(n_9771),
.Y(n_11458)
);

NAND2xp5_ASAP7_75t_L g11459 ( 
.A(n_10140),
.B(n_8207),
.Y(n_11459)
);

INVx1_ASAP7_75t_L g11460 ( 
.A(n_9830),
.Y(n_11460)
);

AOI22xp33_ASAP7_75t_L g11461 ( 
.A1(n_9613),
.A2(n_8524),
.B1(n_7970),
.B2(n_9185),
.Y(n_11461)
);

INVxp67_ASAP7_75t_SL g11462 ( 
.A(n_9518),
.Y(n_11462)
);

INVx1_ASAP7_75t_L g11463 ( 
.A(n_9775),
.Y(n_11463)
);

BUFx3_ASAP7_75t_L g11464 ( 
.A(n_9416),
.Y(n_11464)
);

OAI21x1_ASAP7_75t_L g11465 ( 
.A1(n_9708),
.A2(n_8603),
.B(n_8601),
.Y(n_11465)
);

BUFx3_ASAP7_75t_L g11466 ( 
.A(n_9416),
.Y(n_11466)
);

BUFx6f_ASAP7_75t_SL g11467 ( 
.A(n_9416),
.Y(n_11467)
);

AO21x2_ASAP7_75t_L g11468 ( 
.A1(n_10218),
.A2(n_8300),
.B(n_8801),
.Y(n_11468)
);

AOI22xp33_ASAP7_75t_L g11469 ( 
.A1(n_9652),
.A2(n_7970),
.B1(n_9185),
.B2(n_8611),
.Y(n_11469)
);

INVx4_ASAP7_75t_SL g11470 ( 
.A(n_9434),
.Y(n_11470)
);

HB1xp67_ASAP7_75t_L g11471 ( 
.A(n_9630),
.Y(n_11471)
);

INVx1_ASAP7_75t_L g11472 ( 
.A(n_9946),
.Y(n_11472)
);

INVx2_ASAP7_75t_L g11473 ( 
.A(n_9696),
.Y(n_11473)
);

INVx1_ASAP7_75t_L g11474 ( 
.A(n_9790),
.Y(n_11474)
);

NAND2xp5_ASAP7_75t_L g11475 ( 
.A(n_10179),
.B(n_8502),
.Y(n_11475)
);

HB1xp67_ASAP7_75t_L g11476 ( 
.A(n_9640),
.Y(n_11476)
);

AO21x2_ASAP7_75t_L g11477 ( 
.A1(n_10218),
.A2(n_8300),
.B(n_8801),
.Y(n_11477)
);

INVx2_ASAP7_75t_L g11478 ( 
.A(n_9711),
.Y(n_11478)
);

AND2x4_ASAP7_75t_L g11479 ( 
.A(n_9384),
.B(n_8788),
.Y(n_11479)
);

AND2x2_ASAP7_75t_L g11480 ( 
.A(n_9973),
.B(n_8362),
.Y(n_11480)
);

INVx1_ASAP7_75t_L g11481 ( 
.A(n_9792),
.Y(n_11481)
);

BUFx2_ASAP7_75t_L g11482 ( 
.A(n_10244),
.Y(n_11482)
);

INVx2_ASAP7_75t_L g11483 ( 
.A(n_9726),
.Y(n_11483)
);

BUFx3_ASAP7_75t_L g11484 ( 
.A(n_9434),
.Y(n_11484)
);

INVx1_ASAP7_75t_L g11485 ( 
.A(n_9830),
.Y(n_11485)
);

INVx1_ASAP7_75t_L g11486 ( 
.A(n_9870),
.Y(n_11486)
);

INVx1_ASAP7_75t_L g11487 ( 
.A(n_9870),
.Y(n_11487)
);

NAND2xp5_ASAP7_75t_L g11488 ( 
.A(n_10224),
.B(n_8502),
.Y(n_11488)
);

INVx1_ASAP7_75t_L g11489 ( 
.A(n_9871),
.Y(n_11489)
);

NAND2x1p5_ASAP7_75t_L g11490 ( 
.A(n_10201),
.B(n_8788),
.Y(n_11490)
);

HB1xp67_ASAP7_75t_L g11491 ( 
.A(n_9649),
.Y(n_11491)
);

INVx1_ASAP7_75t_L g11492 ( 
.A(n_9736),
.Y(n_11492)
);

INVx1_ASAP7_75t_L g11493 ( 
.A(n_9736),
.Y(n_11493)
);

INVx1_ASAP7_75t_L g11494 ( 
.A(n_9775),
.Y(n_11494)
);

INVx2_ASAP7_75t_SL g11495 ( 
.A(n_9434),
.Y(n_11495)
);

AOI21xp5_ASAP7_75t_L g11496 ( 
.A1(n_10056),
.A2(n_8869),
.B(n_8541),
.Y(n_11496)
);

INVx2_ASAP7_75t_L g11497 ( 
.A(n_9728),
.Y(n_11497)
);

INVx1_ASAP7_75t_L g11498 ( 
.A(n_9815),
.Y(n_11498)
);

OR2x2_ASAP7_75t_L g11499 ( 
.A(n_10352),
.B(n_8474),
.Y(n_11499)
);

INVx2_ASAP7_75t_L g11500 ( 
.A(n_9728),
.Y(n_11500)
);

AND2x2_ASAP7_75t_L g11501 ( 
.A(n_9973),
.B(n_8362),
.Y(n_11501)
);

OA21x2_ASAP7_75t_L g11502 ( 
.A1(n_9378),
.A2(n_7993),
.B(n_7983),
.Y(n_11502)
);

INVx1_ASAP7_75t_L g11503 ( 
.A(n_9790),
.Y(n_11503)
);

INVx2_ASAP7_75t_L g11504 ( 
.A(n_9792),
.Y(n_11504)
);

AO21x2_ASAP7_75t_L g11505 ( 
.A1(n_9652),
.A2(n_10109),
.B(n_9397),
.Y(n_11505)
);

BUFx12f_ASAP7_75t_L g11506 ( 
.A(n_9663),
.Y(n_11506)
);

INVx2_ASAP7_75t_L g11507 ( 
.A(n_9798),
.Y(n_11507)
);

INVx2_ASAP7_75t_SL g11508 ( 
.A(n_9434),
.Y(n_11508)
);

INVx2_ASAP7_75t_L g11509 ( 
.A(n_9798),
.Y(n_11509)
);

AO21x1_ASAP7_75t_SL g11510 ( 
.A1(n_10164),
.A2(n_9236),
.B(n_9142),
.Y(n_11510)
);

AOI221x1_ASAP7_75t_L g11511 ( 
.A1(n_9807),
.A2(n_8538),
.B1(n_9023),
.B2(n_9032),
.C(n_8636),
.Y(n_11511)
);

OAI21xp5_ASAP7_75t_L g11512 ( 
.A1(n_9680),
.A2(n_8256),
.B(n_8267),
.Y(n_11512)
);

INVx2_ASAP7_75t_L g11513 ( 
.A(n_9803),
.Y(n_11513)
);

OA21x2_ASAP7_75t_L g11514 ( 
.A1(n_9642),
.A2(n_7993),
.B(n_7983),
.Y(n_11514)
);

INVx2_ASAP7_75t_L g11515 ( 
.A(n_9803),
.Y(n_11515)
);

INVx1_ASAP7_75t_L g11516 ( 
.A(n_9838),
.Y(n_11516)
);

HB1xp67_ASAP7_75t_L g11517 ( 
.A(n_9677),
.Y(n_11517)
);

INVx1_ASAP7_75t_L g11518 ( 
.A(n_9825),
.Y(n_11518)
);

OAI21xp5_ASAP7_75t_L g11519 ( 
.A1(n_9468),
.A2(n_8267),
.B(n_8171),
.Y(n_11519)
);

OAI21x1_ASAP7_75t_L g11520 ( 
.A1(n_9708),
.A2(n_8603),
.B(n_8601),
.Y(n_11520)
);

INVx1_ASAP7_75t_L g11521 ( 
.A(n_9811),
.Y(n_11521)
);

NAND2xp5_ASAP7_75t_L g11522 ( 
.A(n_9932),
.B(n_8783),
.Y(n_11522)
);

AND2x4_ASAP7_75t_L g11523 ( 
.A(n_9384),
.B(n_8788),
.Y(n_11523)
);

INVx1_ASAP7_75t_L g11524 ( 
.A(n_9857),
.Y(n_11524)
);

INVx1_ASAP7_75t_L g11525 ( 
.A(n_9857),
.Y(n_11525)
);

INVx1_ASAP7_75t_L g11526 ( 
.A(n_9859),
.Y(n_11526)
);

INVx2_ASAP7_75t_L g11527 ( 
.A(n_9811),
.Y(n_11527)
);

AND2x2_ASAP7_75t_L g11528 ( 
.A(n_9973),
.B(n_8362),
.Y(n_11528)
);

INVx2_ASAP7_75t_L g11529 ( 
.A(n_9813),
.Y(n_11529)
);

INVx3_ASAP7_75t_L g11530 ( 
.A(n_10605),
.Y(n_11530)
);

CKINVDCx5p33_ASAP7_75t_R g11531 ( 
.A(n_9529),
.Y(n_11531)
);

INVx1_ASAP7_75t_L g11532 ( 
.A(n_9822),
.Y(n_11532)
);

INVx1_ASAP7_75t_L g11533 ( 
.A(n_9838),
.Y(n_11533)
);

INVx2_ASAP7_75t_L g11534 ( 
.A(n_9813),
.Y(n_11534)
);

INVx1_ASAP7_75t_L g11535 ( 
.A(n_9815),
.Y(n_11535)
);

INVx2_ASAP7_75t_L g11536 ( 
.A(n_9840),
.Y(n_11536)
);

INVx1_ASAP7_75t_L g11537 ( 
.A(n_9871),
.Y(n_11537)
);

INVx1_ASAP7_75t_L g11538 ( 
.A(n_9883),
.Y(n_11538)
);

INVx1_ASAP7_75t_L g11539 ( 
.A(n_9883),
.Y(n_11539)
);

AO21x2_ASAP7_75t_L g11540 ( 
.A1(n_9397),
.A2(n_8801),
.B(n_8246),
.Y(n_11540)
);

AO31x2_ASAP7_75t_L g11541 ( 
.A1(n_10048),
.A2(n_8612),
.A3(n_8778),
.B(n_8566),
.Y(n_11541)
);

OAI21x1_ASAP7_75t_L g11542 ( 
.A1(n_9940),
.A2(n_8607),
.B(n_8603),
.Y(n_11542)
);

INVx1_ASAP7_75t_L g11543 ( 
.A(n_9948),
.Y(n_11543)
);

INVx3_ASAP7_75t_L g11544 ( 
.A(n_10605),
.Y(n_11544)
);

INVx1_ASAP7_75t_L g11545 ( 
.A(n_9948),
.Y(n_11545)
);

AND2x4_ASAP7_75t_L g11546 ( 
.A(n_9429),
.B(n_8788),
.Y(n_11546)
);

INVx2_ASAP7_75t_SL g11547 ( 
.A(n_9434),
.Y(n_11547)
);

INVx2_ASAP7_75t_L g11548 ( 
.A(n_9840),
.Y(n_11548)
);

INVx1_ASAP7_75t_L g11549 ( 
.A(n_9859),
.Y(n_11549)
);

INVx2_ASAP7_75t_L g11550 ( 
.A(n_9846),
.Y(n_11550)
);

INVx1_ASAP7_75t_L g11551 ( 
.A(n_9879),
.Y(n_11551)
);

AND2x6_ASAP7_75t_L g11552 ( 
.A(n_9434),
.B(n_8693),
.Y(n_11552)
);

INVx1_ASAP7_75t_L g11553 ( 
.A(n_9933),
.Y(n_11553)
);

BUFx2_ASAP7_75t_L g11554 ( 
.A(n_10244),
.Y(n_11554)
);

HB1xp67_ASAP7_75t_L g11555 ( 
.A(n_9758),
.Y(n_11555)
);

INVx1_ASAP7_75t_SL g11556 ( 
.A(n_9604),
.Y(n_11556)
);

INVx1_ASAP7_75t_L g11557 ( 
.A(n_9882),
.Y(n_11557)
);

AND2x2_ASAP7_75t_L g11558 ( 
.A(n_10100),
.B(n_10512),
.Y(n_11558)
);

INVx1_ASAP7_75t_L g11559 ( 
.A(n_9882),
.Y(n_11559)
);

AND2x2_ASAP7_75t_L g11560 ( 
.A(n_10100),
.B(n_8373),
.Y(n_11560)
);

OAI21x1_ASAP7_75t_L g11561 ( 
.A1(n_9940),
.A2(n_8607),
.B(n_8603),
.Y(n_11561)
);

AND2x2_ASAP7_75t_L g11562 ( 
.A(n_10100),
.B(n_8373),
.Y(n_11562)
);

HB1xp67_ASAP7_75t_L g11563 ( 
.A(n_9787),
.Y(n_11563)
);

INVx2_ASAP7_75t_L g11564 ( 
.A(n_9851),
.Y(n_11564)
);

AND2x4_ASAP7_75t_L g11565 ( 
.A(n_9429),
.B(n_8788),
.Y(n_11565)
);

HB1xp67_ASAP7_75t_L g11566 ( 
.A(n_9821),
.Y(n_11566)
);

INVx2_ASAP7_75t_SL g11567 ( 
.A(n_9472),
.Y(n_11567)
);

INVx2_ASAP7_75t_L g11568 ( 
.A(n_9851),
.Y(n_11568)
);

INVx2_ASAP7_75t_L g11569 ( 
.A(n_9879),
.Y(n_11569)
);

INVx1_ASAP7_75t_L g11570 ( 
.A(n_9904),
.Y(n_11570)
);

INVx2_ASAP7_75t_L g11571 ( 
.A(n_9881),
.Y(n_11571)
);

OR2x2_ASAP7_75t_L g11572 ( 
.A(n_10352),
.B(n_9250),
.Y(n_11572)
);

HB1xp67_ASAP7_75t_L g11573 ( 
.A(n_9881),
.Y(n_11573)
);

INVx2_ASAP7_75t_L g11574 ( 
.A(n_9886),
.Y(n_11574)
);

INVx2_ASAP7_75t_L g11575 ( 
.A(n_9904),
.Y(n_11575)
);

INVx1_ASAP7_75t_L g11576 ( 
.A(n_9909),
.Y(n_11576)
);

INVx3_ASAP7_75t_L g11577 ( 
.A(n_10605),
.Y(n_11577)
);

AND2x4_ASAP7_75t_L g11578 ( 
.A(n_9429),
.B(n_8788),
.Y(n_11578)
);

OAI21x1_ASAP7_75t_L g11579 ( 
.A1(n_9940),
.A2(n_8622),
.B(n_8607),
.Y(n_11579)
);

AO21x2_ASAP7_75t_L g11580 ( 
.A1(n_10577),
.A2(n_8801),
.B(n_8372),
.Y(n_11580)
);

INVx2_ASAP7_75t_L g11581 ( 
.A(n_9909),
.Y(n_11581)
);

BUFx3_ASAP7_75t_L g11582 ( 
.A(n_9472),
.Y(n_11582)
);

INVx1_ASAP7_75t_L g11583 ( 
.A(n_9952),
.Y(n_11583)
);

AND2x2_ASAP7_75t_L g11584 ( 
.A(n_10100),
.B(n_8373),
.Y(n_11584)
);

HB1xp67_ASAP7_75t_L g11585 ( 
.A(n_9914),
.Y(n_11585)
);

INVx2_ASAP7_75t_SL g11586 ( 
.A(n_9472),
.Y(n_11586)
);

INVx1_ASAP7_75t_L g11587 ( 
.A(n_9952),
.Y(n_11587)
);

OAI21x1_ASAP7_75t_L g11588 ( 
.A1(n_10097),
.A2(n_8622),
.B(n_8607),
.Y(n_11588)
);

INVx1_ASAP7_75t_L g11589 ( 
.A(n_9977),
.Y(n_11589)
);

INVx2_ASAP7_75t_L g11590 ( 
.A(n_9914),
.Y(n_11590)
);

HB1xp67_ASAP7_75t_L g11591 ( 
.A(n_9917),
.Y(n_11591)
);

INVx2_ASAP7_75t_L g11592 ( 
.A(n_9917),
.Y(n_11592)
);

AO21x2_ASAP7_75t_L g11593 ( 
.A1(n_10577),
.A2(n_8801),
.B(n_8372),
.Y(n_11593)
);

INVx1_ASAP7_75t_L g11594 ( 
.A(n_10029),
.Y(n_11594)
);

INVx1_ASAP7_75t_L g11595 ( 
.A(n_10029),
.Y(n_11595)
);

INVxp67_ASAP7_75t_L g11596 ( 
.A(n_10384),
.Y(n_11596)
);

INVxp67_ASAP7_75t_L g11597 ( 
.A(n_10521),
.Y(n_11597)
);

AOI21x1_ASAP7_75t_L g11598 ( 
.A1(n_10252),
.A2(n_8994),
.B(n_8027),
.Y(n_11598)
);

AO31x2_ASAP7_75t_L g11599 ( 
.A1(n_10048),
.A2(n_8612),
.A3(n_8778),
.B(n_8566),
.Y(n_11599)
);

AND2x2_ASAP7_75t_L g11600 ( 
.A(n_10611),
.B(n_8411),
.Y(n_11600)
);

AND2x2_ASAP7_75t_L g11601 ( 
.A(n_10634),
.B(n_8411),
.Y(n_11601)
);

INVx1_ASAP7_75t_L g11602 ( 
.A(n_10030),
.Y(n_11602)
);

INVx1_ASAP7_75t_L g11603 ( 
.A(n_10030),
.Y(n_11603)
);

AND2x2_ASAP7_75t_L g11604 ( 
.A(n_10668),
.B(n_8411),
.Y(n_11604)
);

NAND2xp5_ASAP7_75t_L g11605 ( 
.A(n_9690),
.B(n_8783),
.Y(n_11605)
);

INVx1_ASAP7_75t_L g11606 ( 
.A(n_9969),
.Y(n_11606)
);

NAND2xp5_ASAP7_75t_L g11607 ( 
.A(n_9730),
.B(n_9010),
.Y(n_11607)
);

AOI22xp5_ASAP7_75t_SL g11608 ( 
.A1(n_10673),
.A2(n_7590),
.B1(n_7650),
.B2(n_7567),
.Y(n_11608)
);

CKINVDCx5p33_ASAP7_75t_R g11609 ( 
.A(n_10207),
.Y(n_11609)
);

INVx1_ASAP7_75t_L g11610 ( 
.A(n_9933),
.Y(n_11610)
);

NAND2xp5_ASAP7_75t_L g11611 ( 
.A(n_9778),
.B(n_9010),
.Y(n_11611)
);

INVx1_ASAP7_75t_L g11612 ( 
.A(n_9975),
.Y(n_11612)
);

INVx2_ASAP7_75t_L g11613 ( 
.A(n_9924),
.Y(n_11613)
);

INVx1_ASAP7_75t_L g11614 ( 
.A(n_9975),
.Y(n_11614)
);

BUFx3_ASAP7_75t_L g11615 ( 
.A(n_9472),
.Y(n_11615)
);

HB1xp67_ASAP7_75t_L g11616 ( 
.A(n_9924),
.Y(n_11616)
);

INVx1_ASAP7_75t_L g11617 ( 
.A(n_9936),
.Y(n_11617)
);

AOI22xp33_ASAP7_75t_SL g11618 ( 
.A1(n_10148),
.A2(n_7970),
.B1(n_8077),
.B2(n_9171),
.Y(n_11618)
);

HB1xp67_ASAP7_75t_L g11619 ( 
.A(n_9936),
.Y(n_11619)
);

AOI22xp5_ASAP7_75t_L g11620 ( 
.A1(n_10594),
.A2(n_8605),
.B1(n_9148),
.B2(n_9181),
.Y(n_11620)
);

INVx3_ASAP7_75t_L g11621 ( 
.A(n_9472),
.Y(n_11621)
);

INVx1_ASAP7_75t_L g11622 ( 
.A(n_9990),
.Y(n_11622)
);

OAI21x1_ASAP7_75t_L g11623 ( 
.A1(n_10097),
.A2(n_10174),
.B(n_10169),
.Y(n_11623)
);

INVx1_ASAP7_75t_L g11624 ( 
.A(n_9990),
.Y(n_11624)
);

INVx1_ASAP7_75t_L g11625 ( 
.A(n_10041),
.Y(n_11625)
);

CKINVDCx14_ASAP7_75t_R g11626 ( 
.A(n_10233),
.Y(n_11626)
);

INVx1_ASAP7_75t_L g11627 ( 
.A(n_10041),
.Y(n_11627)
);

AND2x2_ASAP7_75t_L g11628 ( 
.A(n_9350),
.B(n_8480),
.Y(n_11628)
);

CKINVDCx6p67_ASAP7_75t_R g11629 ( 
.A(n_9472),
.Y(n_11629)
);

INVx2_ASAP7_75t_L g11630 ( 
.A(n_9946),
.Y(n_11630)
);

AND2x2_ASAP7_75t_L g11631 ( 
.A(n_9350),
.B(n_8480),
.Y(n_11631)
);

HB1xp67_ASAP7_75t_L g11632 ( 
.A(n_9950),
.Y(n_11632)
);

CKINVDCx6p67_ASAP7_75t_R g11633 ( 
.A(n_9558),
.Y(n_11633)
);

INVx1_ASAP7_75t_L g11634 ( 
.A(n_9993),
.Y(n_11634)
);

INVx2_ASAP7_75t_L g11635 ( 
.A(n_9950),
.Y(n_11635)
);

INVx1_ASAP7_75t_SL g11636 ( 
.A(n_10273),
.Y(n_11636)
);

OAI21x1_ASAP7_75t_L g11637 ( 
.A1(n_10097),
.A2(n_8627),
.B(n_8622),
.Y(n_11637)
);

BUFx2_ASAP7_75t_L g11638 ( 
.A(n_10244),
.Y(n_11638)
);

INVx1_ASAP7_75t_L g11639 ( 
.A(n_9969),
.Y(n_11639)
);

INVx1_ASAP7_75t_L g11640 ( 
.A(n_9986),
.Y(n_11640)
);

INVx1_ASAP7_75t_L g11641 ( 
.A(n_9986),
.Y(n_11641)
);

HB1xp67_ASAP7_75t_L g11642 ( 
.A(n_9955),
.Y(n_11642)
);

INVx2_ASAP7_75t_SL g11643 ( 
.A(n_10441),
.Y(n_11643)
);

INVx1_ASAP7_75t_L g11644 ( 
.A(n_10014),
.Y(n_11644)
);

AND2x2_ASAP7_75t_L g11645 ( 
.A(n_9350),
.B(n_8480),
.Y(n_11645)
);

INVx2_ASAP7_75t_L g11646 ( 
.A(n_9955),
.Y(n_11646)
);

BUFx3_ASAP7_75t_L g11647 ( 
.A(n_10434),
.Y(n_11647)
);

INVx2_ASAP7_75t_SL g11648 ( 
.A(n_10441),
.Y(n_11648)
);

INVx1_ASAP7_75t_L g11649 ( 
.A(n_9988),
.Y(n_11649)
);

AND2x2_ASAP7_75t_L g11650 ( 
.A(n_9350),
.B(n_9251),
.Y(n_11650)
);

INVx1_ASAP7_75t_L g11651 ( 
.A(n_9976),
.Y(n_11651)
);

INVx2_ASAP7_75t_L g11652 ( 
.A(n_9964),
.Y(n_11652)
);

INVx1_ASAP7_75t_L g11653 ( 
.A(n_9976),
.Y(n_11653)
);

CKINVDCx20_ASAP7_75t_R g11654 ( 
.A(n_9880),
.Y(n_11654)
);

INVx1_ASAP7_75t_L g11655 ( 
.A(n_9992),
.Y(n_11655)
);

NAND2xp5_ASAP7_75t_L g11656 ( 
.A(n_10604),
.B(n_9052),
.Y(n_11656)
);

INVx2_ASAP7_75t_L g11657 ( 
.A(n_9964),
.Y(n_11657)
);

BUFx3_ASAP7_75t_L g11658 ( 
.A(n_10452),
.Y(n_11658)
);

INVx1_ASAP7_75t_L g11659 ( 
.A(n_9993),
.Y(n_11659)
);

INVx3_ASAP7_75t_L g11660 ( 
.A(n_10297),
.Y(n_11660)
);

OA21x2_ASAP7_75t_L g11661 ( 
.A1(n_9642),
.A2(n_8204),
.B(n_8203),
.Y(n_11661)
);

INVx4_ASAP7_75t_L g11662 ( 
.A(n_9343),
.Y(n_11662)
);

AO21x2_ASAP7_75t_L g11663 ( 
.A1(n_10577),
.A2(n_8372),
.B(n_8160),
.Y(n_11663)
);

OR2x6_ASAP7_75t_L g11664 ( 
.A(n_10068),
.B(n_7971),
.Y(n_11664)
);

INVx1_ASAP7_75t_L g11665 ( 
.A(n_9995),
.Y(n_11665)
);

INVx2_ASAP7_75t_L g11666 ( 
.A(n_9967),
.Y(n_11666)
);

BUFx6f_ASAP7_75t_L g11667 ( 
.A(n_9343),
.Y(n_11667)
);

AND2x2_ASAP7_75t_L g11668 ( 
.A(n_9354),
.B(n_9251),
.Y(n_11668)
);

INVx2_ASAP7_75t_L g11669 ( 
.A(n_9967),
.Y(n_11669)
);

OR2x2_ASAP7_75t_L g11670 ( 
.A(n_10407),
.B(n_10608),
.Y(n_11670)
);

INVx1_ASAP7_75t_L g11671 ( 
.A(n_10091),
.Y(n_11671)
);

AND2x2_ASAP7_75t_L g11672 ( 
.A(n_9354),
.B(n_9260),
.Y(n_11672)
);

INVx2_ASAP7_75t_L g11673 ( 
.A(n_9977),
.Y(n_11673)
);

INVx1_ASAP7_75t_L g11674 ( 
.A(n_9988),
.Y(n_11674)
);

INVx1_ASAP7_75t_L g11675 ( 
.A(n_10085),
.Y(n_11675)
);

INVx1_ASAP7_75t_L g11676 ( 
.A(n_10085),
.Y(n_11676)
);

BUFx2_ASAP7_75t_L g11677 ( 
.A(n_10723),
.Y(n_11677)
);

OAI21xp5_ASAP7_75t_L g11678 ( 
.A1(n_10066),
.A2(n_8267),
.B(n_8171),
.Y(n_11678)
);

AND2x2_ASAP7_75t_L g11679 ( 
.A(n_9354),
.B(n_9260),
.Y(n_11679)
);

OAI21x1_ASAP7_75t_L g11680 ( 
.A1(n_10169),
.A2(n_10174),
.B(n_10177),
.Y(n_11680)
);

BUFx3_ASAP7_75t_L g11681 ( 
.A(n_10485),
.Y(n_11681)
);

OA21x2_ASAP7_75t_L g11682 ( 
.A1(n_10461),
.A2(n_8204),
.B(n_8203),
.Y(n_11682)
);

INVx2_ASAP7_75t_L g11683 ( 
.A(n_9992),
.Y(n_11683)
);

INVx2_ASAP7_75t_SL g11684 ( 
.A(n_10441),
.Y(n_11684)
);

INVx2_ASAP7_75t_L g11685 ( 
.A(n_9995),
.Y(n_11685)
);

OR2x6_ASAP7_75t_L g11686 ( 
.A(n_10068),
.B(n_7971),
.Y(n_11686)
);

INVx2_ASAP7_75t_L g11687 ( 
.A(n_10012),
.Y(n_11687)
);

INVx3_ASAP7_75t_L g11688 ( 
.A(n_10297),
.Y(n_11688)
);

INVx2_ASAP7_75t_L g11689 ( 
.A(n_10012),
.Y(n_11689)
);

HB1xp67_ASAP7_75t_L g11690 ( 
.A(n_10014),
.Y(n_11690)
);

INVx2_ASAP7_75t_L g11691 ( 
.A(n_10036),
.Y(n_11691)
);

NAND2xp5_ASAP7_75t_L g11692 ( 
.A(n_10633),
.B(n_9052),
.Y(n_11692)
);

AND2x2_ASAP7_75t_L g11693 ( 
.A(n_9354),
.B(n_9364),
.Y(n_11693)
);

INVx3_ASAP7_75t_L g11694 ( 
.A(n_10297),
.Y(n_11694)
);

AND2x4_ASAP7_75t_L g11695 ( 
.A(n_9533),
.B(n_8881),
.Y(n_11695)
);

OAI21x1_ASAP7_75t_L g11696 ( 
.A1(n_10169),
.A2(n_8627),
.B(n_8622),
.Y(n_11696)
);

INVx1_ASAP7_75t_L g11697 ( 
.A(n_10062),
.Y(n_11697)
);

AND2x2_ASAP7_75t_L g11698 ( 
.A(n_9364),
.B(n_9263),
.Y(n_11698)
);

INVx1_ASAP7_75t_L g11699 ( 
.A(n_10062),
.Y(n_11699)
);

INVx1_ASAP7_75t_L g11700 ( 
.A(n_10086),
.Y(n_11700)
);

INVx1_ASAP7_75t_L g11701 ( 
.A(n_10086),
.Y(n_11701)
);

HB1xp67_ASAP7_75t_L g11702 ( 
.A(n_10036),
.Y(n_11702)
);

INVx4_ASAP7_75t_L g11703 ( 
.A(n_10519),
.Y(n_11703)
);

INVx2_ASAP7_75t_L g11704 ( 
.A(n_10044),
.Y(n_11704)
);

HB1xp67_ASAP7_75t_L g11705 ( 
.A(n_10044),
.Y(n_11705)
);

INVxp67_ASAP7_75t_L g11706 ( 
.A(n_10626),
.Y(n_11706)
);

INVx1_ASAP7_75t_SL g11707 ( 
.A(n_10227),
.Y(n_11707)
);

INVx2_ASAP7_75t_L g11708 ( 
.A(n_10051),
.Y(n_11708)
);

INVx1_ASAP7_75t_L g11709 ( 
.A(n_10051),
.Y(n_11709)
);

AO21x2_ASAP7_75t_L g11710 ( 
.A1(n_9927),
.A2(n_8372),
.B(n_8160),
.Y(n_11710)
);

AND2x2_ASAP7_75t_L g11711 ( 
.A(n_9364),
.B(n_9263),
.Y(n_11711)
);

BUFx3_ASAP7_75t_L g11712 ( 
.A(n_10489),
.Y(n_11712)
);

OAI21x1_ASAP7_75t_L g11713 ( 
.A1(n_10174),
.A2(n_8630),
.B(n_8627),
.Y(n_11713)
);

INVx1_ASAP7_75t_L g11714 ( 
.A(n_10079),
.Y(n_11714)
);

INVx1_ASAP7_75t_L g11715 ( 
.A(n_10079),
.Y(n_11715)
);

AOI22xp33_ASAP7_75t_L g11716 ( 
.A1(n_9731),
.A2(n_8571),
.B1(n_8570),
.B2(n_9145),
.Y(n_11716)
);

BUFx2_ASAP7_75t_L g11717 ( 
.A(n_10723),
.Y(n_11717)
);

INVx1_ASAP7_75t_L g11718 ( 
.A(n_10091),
.Y(n_11718)
);

BUFx3_ASAP7_75t_L g11719 ( 
.A(n_10508),
.Y(n_11719)
);

OAI21x1_ASAP7_75t_L g11720 ( 
.A1(n_10177),
.A2(n_8630),
.B(n_8627),
.Y(n_11720)
);

INVx2_ASAP7_75t_SL g11721 ( 
.A(n_10441),
.Y(n_11721)
);

BUFx3_ASAP7_75t_L g11722 ( 
.A(n_10610),
.Y(n_11722)
);

INVx1_ASAP7_75t_L g11723 ( 
.A(n_10107),
.Y(n_11723)
);

CKINVDCx5p33_ASAP7_75t_R g11724 ( 
.A(n_9321),
.Y(n_11724)
);

INVxp67_ASAP7_75t_SL g11725 ( 
.A(n_9807),
.Y(n_11725)
);

INVx2_ASAP7_75t_L g11726 ( 
.A(n_10055),
.Y(n_11726)
);

INVx3_ASAP7_75t_L g11727 ( 
.A(n_10297),
.Y(n_11727)
);

INVx2_ASAP7_75t_L g11728 ( 
.A(n_10055),
.Y(n_11728)
);

CKINVDCx5p33_ASAP7_75t_R g11729 ( 
.A(n_10176),
.Y(n_11729)
);

INVx2_ASAP7_75t_L g11730 ( 
.A(n_10069),
.Y(n_11730)
);

INVx2_ASAP7_75t_L g11731 ( 
.A(n_10069),
.Y(n_11731)
);

AND2x2_ASAP7_75t_L g11732 ( 
.A(n_9364),
.B(n_7990),
.Y(n_11732)
);

INVx1_ASAP7_75t_L g11733 ( 
.A(n_10151),
.Y(n_11733)
);

INVx2_ASAP7_75t_L g11734 ( 
.A(n_10101),
.Y(n_11734)
);

BUFx3_ASAP7_75t_L g11735 ( 
.A(n_10690),
.Y(n_11735)
);

INVx1_ASAP7_75t_L g11736 ( 
.A(n_10151),
.Y(n_11736)
);

BUFx3_ASAP7_75t_L g11737 ( 
.A(n_9558),
.Y(n_11737)
);

NAND2x1p5_ASAP7_75t_L g11738 ( 
.A(n_10252),
.B(n_8881),
.Y(n_11738)
);

HB1xp67_ASAP7_75t_L g11739 ( 
.A(n_10101),
.Y(n_11739)
);

INVx2_ASAP7_75t_L g11740 ( 
.A(n_10103),
.Y(n_11740)
);

INVx1_ASAP7_75t_L g11741 ( 
.A(n_10117),
.Y(n_11741)
);

INVx1_ASAP7_75t_L g11742 ( 
.A(n_10117),
.Y(n_11742)
);

OA21x2_ASAP7_75t_L g11743 ( 
.A1(n_10461),
.A2(n_8204),
.B(n_8203),
.Y(n_11743)
);

INVx1_ASAP7_75t_L g11744 ( 
.A(n_10118),
.Y(n_11744)
);

INVx2_ASAP7_75t_SL g11745 ( 
.A(n_10660),
.Y(n_11745)
);

AND2x2_ASAP7_75t_L g11746 ( 
.A(n_9386),
.B(n_7990),
.Y(n_11746)
);

INVx1_ASAP7_75t_L g11747 ( 
.A(n_10118),
.Y(n_11747)
);

INVx2_ASAP7_75t_L g11748 ( 
.A(n_10103),
.Y(n_11748)
);

INVx2_ASAP7_75t_L g11749 ( 
.A(n_10107),
.Y(n_11749)
);

BUFx4f_ASAP7_75t_SL g11750 ( 
.A(n_9902),
.Y(n_11750)
);

AOI22xp33_ASAP7_75t_L g11751 ( 
.A1(n_9731),
.A2(n_8571),
.B1(n_9145),
.B2(n_8518),
.Y(n_11751)
);

INVx1_ASAP7_75t_L g11752 ( 
.A(n_10198),
.Y(n_11752)
);

INVx2_ASAP7_75t_L g11753 ( 
.A(n_10110),
.Y(n_11753)
);

INVx1_ASAP7_75t_L g11754 ( 
.A(n_10198),
.Y(n_11754)
);

OAI21xp5_ASAP7_75t_L g11755 ( 
.A1(n_9527),
.A2(n_8267),
.B(n_8171),
.Y(n_11755)
);

INVx1_ASAP7_75t_L g11756 ( 
.A(n_10112),
.Y(n_11756)
);

INVx1_ASAP7_75t_L g11757 ( 
.A(n_10112),
.Y(n_11757)
);

INVx2_ASAP7_75t_L g11758 ( 
.A(n_10110),
.Y(n_11758)
);

INVx1_ASAP7_75t_L g11759 ( 
.A(n_10143),
.Y(n_11759)
);

AND2x2_ASAP7_75t_L g11760 ( 
.A(n_9386),
.B(n_8027),
.Y(n_11760)
);

INVx2_ASAP7_75t_L g11761 ( 
.A(n_10131),
.Y(n_11761)
);

INVx1_ASAP7_75t_L g11762 ( 
.A(n_10143),
.Y(n_11762)
);

INVx2_ASAP7_75t_L g11763 ( 
.A(n_10131),
.Y(n_11763)
);

INVx2_ASAP7_75t_L g11764 ( 
.A(n_10132),
.Y(n_11764)
);

AOI21x1_ASAP7_75t_L g11765 ( 
.A1(n_9706),
.A2(n_8994),
.B(n_8058),
.Y(n_11765)
);

INVx1_ASAP7_75t_L g11766 ( 
.A(n_10171),
.Y(n_11766)
);

INVx1_ASAP7_75t_L g11767 ( 
.A(n_10171),
.Y(n_11767)
);

HB1xp67_ASAP7_75t_SL g11768 ( 
.A(n_9878),
.Y(n_11768)
);

AND2x2_ASAP7_75t_L g11769 ( 
.A(n_9386),
.B(n_9484),
.Y(n_11769)
);

AOI22xp33_ASAP7_75t_L g11770 ( 
.A1(n_9791),
.A2(n_8518),
.B1(n_8288),
.B2(n_8455),
.Y(n_11770)
);

INVx4_ASAP7_75t_L g11771 ( 
.A(n_10519),
.Y(n_11771)
);

AOI21xp5_ASAP7_75t_SL g11772 ( 
.A1(n_9530),
.A2(n_8984),
.B(n_8538),
.Y(n_11772)
);

NOR2xp33_ASAP7_75t_L g11773 ( 
.A(n_9349),
.B(n_7785),
.Y(n_11773)
);

OAI21x1_ASAP7_75t_L g11774 ( 
.A1(n_10177),
.A2(n_8631),
.B(n_8630),
.Y(n_11774)
);

INVx2_ASAP7_75t_L g11775 ( 
.A(n_10132),
.Y(n_11775)
);

INVx1_ASAP7_75t_L g11776 ( 
.A(n_10154),
.Y(n_11776)
);

INVx1_ASAP7_75t_L g11777 ( 
.A(n_10154),
.Y(n_11777)
);

INVx1_ASAP7_75t_L g11778 ( 
.A(n_10166),
.Y(n_11778)
);

INVx3_ASAP7_75t_L g11779 ( 
.A(n_10308),
.Y(n_11779)
);

INVx1_ASAP7_75t_L g11780 ( 
.A(n_10166),
.Y(n_11780)
);

INVx1_ASAP7_75t_L g11781 ( 
.A(n_10284),
.Y(n_11781)
);

CKINVDCx20_ASAP7_75t_R g11782 ( 
.A(n_10196),
.Y(n_11782)
);

OA21x2_ASAP7_75t_L g11783 ( 
.A1(n_10461),
.A2(n_7962),
.B(n_7959),
.Y(n_11783)
);

INVx3_ASAP7_75t_L g11784 ( 
.A(n_10308),
.Y(n_11784)
);

INVx1_ASAP7_75t_L g11785 ( 
.A(n_10208),
.Y(n_11785)
);

AOI21xp33_ASAP7_75t_L g11786 ( 
.A1(n_10202),
.A2(n_8659),
.B(n_8333),
.Y(n_11786)
);

AND2x4_ASAP7_75t_L g11787 ( 
.A(n_9533),
.B(n_8881),
.Y(n_11787)
);

INVx1_ASAP7_75t_L g11788 ( 
.A(n_10208),
.Y(n_11788)
);

INVx1_ASAP7_75t_L g11789 ( 
.A(n_10245),
.Y(n_11789)
);

HB1xp67_ASAP7_75t_L g11790 ( 
.A(n_10146),
.Y(n_11790)
);

INVx2_ASAP7_75t_L g11791 ( 
.A(n_10146),
.Y(n_11791)
);

INVx1_ASAP7_75t_L g11792 ( 
.A(n_10168),
.Y(n_11792)
);

INVx2_ASAP7_75t_L g11793 ( 
.A(n_10149),
.Y(n_11793)
);

OAI21x1_ASAP7_75t_L g11794 ( 
.A1(n_10271),
.A2(n_8631),
.B(n_8630),
.Y(n_11794)
);

NAND2xp5_ASAP7_75t_L g11795 ( 
.A(n_9959),
.B(n_8712),
.Y(n_11795)
);

INVx1_ASAP7_75t_L g11796 ( 
.A(n_10158),
.Y(n_11796)
);

OAI21x1_ASAP7_75t_L g11797 ( 
.A1(n_10271),
.A2(n_8637),
.B(n_8631),
.Y(n_11797)
);

INVx1_ASAP7_75t_L g11798 ( 
.A(n_10158),
.Y(n_11798)
);

AND2x4_ASAP7_75t_L g11799 ( 
.A(n_9533),
.B(n_8881),
.Y(n_11799)
);

INVx2_ASAP7_75t_L g11800 ( 
.A(n_10149),
.Y(n_11800)
);

OAI221xp5_ASAP7_75t_L g11801 ( 
.A1(n_9907),
.A2(n_9168),
.B1(n_9214),
.B2(n_9294),
.C(n_9283),
.Y(n_11801)
);

INVx4_ASAP7_75t_L g11802 ( 
.A(n_9601),
.Y(n_11802)
);

INVx1_ASAP7_75t_L g11803 ( 
.A(n_10284),
.Y(n_11803)
);

INVx1_ASAP7_75t_L g11804 ( 
.A(n_10285),
.Y(n_11804)
);

BUFx3_ASAP7_75t_L g11805 ( 
.A(n_9402),
.Y(n_11805)
);

OAI22xp5_ASAP7_75t_L g11806 ( 
.A1(n_9424),
.A2(n_8811),
.B1(n_8729),
.B2(n_9286),
.Y(n_11806)
);

INVx1_ASAP7_75t_L g11807 ( 
.A(n_10245),
.Y(n_11807)
);

INVx2_ASAP7_75t_L g11808 ( 
.A(n_10168),
.Y(n_11808)
);

AND2x4_ASAP7_75t_L g11809 ( 
.A(n_9560),
.B(n_8881),
.Y(n_11809)
);

BUFx3_ASAP7_75t_L g11810 ( 
.A(n_9417),
.Y(n_11810)
);

INVx1_ASAP7_75t_L g11811 ( 
.A(n_10173),
.Y(n_11811)
);

INVx1_ASAP7_75t_L g11812 ( 
.A(n_10173),
.Y(n_11812)
);

INVx2_ASAP7_75t_L g11813 ( 
.A(n_10178),
.Y(n_11813)
);

INVx1_ASAP7_75t_L g11814 ( 
.A(n_10282),
.Y(n_11814)
);

INVx1_ASAP7_75t_L g11815 ( 
.A(n_10282),
.Y(n_11815)
);

HB1xp67_ASAP7_75t_L g11816 ( 
.A(n_10178),
.Y(n_11816)
);

INVx1_ASAP7_75t_L g11817 ( 
.A(n_10190),
.Y(n_11817)
);

INVx1_ASAP7_75t_L g11818 ( 
.A(n_10190),
.Y(n_11818)
);

BUFx6f_ASAP7_75t_L g11819 ( 
.A(n_9501),
.Y(n_11819)
);

INVx2_ASAP7_75t_L g11820 ( 
.A(n_10181),
.Y(n_11820)
);

INVx1_ASAP7_75t_L g11821 ( 
.A(n_10191),
.Y(n_11821)
);

INVx2_ASAP7_75t_L g11822 ( 
.A(n_10181),
.Y(n_11822)
);

INVx1_ASAP7_75t_L g11823 ( 
.A(n_10256),
.Y(n_11823)
);

INVx1_ASAP7_75t_L g11824 ( 
.A(n_10256),
.Y(n_11824)
);

INVx2_ASAP7_75t_SL g11825 ( 
.A(n_10660),
.Y(n_11825)
);

INVx2_ASAP7_75t_SL g11826 ( 
.A(n_10660),
.Y(n_11826)
);

NAND3xp33_ASAP7_75t_L g11827 ( 
.A(n_10274),
.B(n_8077),
.C(n_8759),
.Y(n_11827)
);

NAND3xp33_ASAP7_75t_L g11828 ( 
.A(n_10713),
.B(n_8077),
.C(n_8759),
.Y(n_11828)
);

INVx1_ASAP7_75t_L g11829 ( 
.A(n_10267),
.Y(n_11829)
);

INVx1_ASAP7_75t_L g11830 ( 
.A(n_10267),
.Y(n_11830)
);

AND2x2_ASAP7_75t_L g11831 ( 
.A(n_9386),
.B(n_8027),
.Y(n_11831)
);

INVx1_ASAP7_75t_L g11832 ( 
.A(n_10217),
.Y(n_11832)
);

AND2x2_ASAP7_75t_L g11833 ( 
.A(n_9484),
.B(n_8058),
.Y(n_11833)
);

BUFx2_ASAP7_75t_L g11834 ( 
.A(n_10590),
.Y(n_11834)
);

INVx4_ASAP7_75t_L g11835 ( 
.A(n_9601),
.Y(n_11835)
);

INVx1_ASAP7_75t_L g11836 ( 
.A(n_10246),
.Y(n_11836)
);

INVx2_ASAP7_75t_L g11837 ( 
.A(n_10191),
.Y(n_11837)
);

NAND2x1p5_ASAP7_75t_L g11838 ( 
.A(n_9723),
.B(n_8881),
.Y(n_11838)
);

INVx1_ASAP7_75t_L g11839 ( 
.A(n_10232),
.Y(n_11839)
);

INVx1_ASAP7_75t_L g11840 ( 
.A(n_10232),
.Y(n_11840)
);

INVx2_ASAP7_75t_L g11841 ( 
.A(n_10217),
.Y(n_11841)
);

NAND2xp5_ASAP7_75t_L g11842 ( 
.A(n_9972),
.B(n_8729),
.Y(n_11842)
);

NAND2xp5_ASAP7_75t_L g11843 ( 
.A(n_9412),
.B(n_9469),
.Y(n_11843)
);

AND2x2_ASAP7_75t_L g11844 ( 
.A(n_9484),
.B(n_8058),
.Y(n_11844)
);

INVx2_ASAP7_75t_L g11845 ( 
.A(n_10235),
.Y(n_11845)
);

BUFx2_ASAP7_75t_L g11846 ( 
.A(n_10590),
.Y(n_11846)
);

BUFx6f_ASAP7_75t_L g11847 ( 
.A(n_9501),
.Y(n_11847)
);

INVx2_ASAP7_75t_L g11848 ( 
.A(n_10235),
.Y(n_11848)
);

INVx3_ASAP7_75t_L g11849 ( 
.A(n_10308),
.Y(n_11849)
);

INVx2_ASAP7_75t_L g11850 ( 
.A(n_10246),
.Y(n_11850)
);

INVxp67_ASAP7_75t_L g11851 ( 
.A(n_9796),
.Y(n_11851)
);

INVx1_ASAP7_75t_L g11852 ( 
.A(n_10283),
.Y(n_11852)
);

BUFx2_ASAP7_75t_SL g11853 ( 
.A(n_9373),
.Y(n_11853)
);

AND2x2_ASAP7_75t_L g11854 ( 
.A(n_9484),
.B(n_8146),
.Y(n_11854)
);

INVx1_ASAP7_75t_L g11855 ( 
.A(n_10286),
.Y(n_11855)
);

INVx3_ASAP7_75t_L g11856 ( 
.A(n_10308),
.Y(n_11856)
);

BUFx3_ASAP7_75t_L g11857 ( 
.A(n_9896),
.Y(n_11857)
);

NAND2xp5_ASAP7_75t_L g11858 ( 
.A(n_9590),
.B(n_8755),
.Y(n_11858)
);

INVx1_ASAP7_75t_L g11859 ( 
.A(n_10277),
.Y(n_11859)
);

INVx3_ASAP7_75t_L g11860 ( 
.A(n_10383),
.Y(n_11860)
);

INVx3_ASAP7_75t_L g11861 ( 
.A(n_10383),
.Y(n_11861)
);

INVx2_ASAP7_75t_SL g11862 ( 
.A(n_10660),
.Y(n_11862)
);

INVx1_ASAP7_75t_L g11863 ( 
.A(n_10277),
.Y(n_11863)
);

BUFx2_ASAP7_75t_L g11864 ( 
.A(n_10699),
.Y(n_11864)
);

OA21x2_ASAP7_75t_L g11865 ( 
.A1(n_10483),
.A2(n_7962),
.B(n_7959),
.Y(n_11865)
);

INVx2_ASAP7_75t_L g11866 ( 
.A(n_10260),
.Y(n_11866)
);

INVx1_ASAP7_75t_L g11867 ( 
.A(n_10279),
.Y(n_11867)
);

BUFx8_ASAP7_75t_SL g11868 ( 
.A(n_10347),
.Y(n_11868)
);

INVx2_ASAP7_75t_L g11869 ( 
.A(n_10260),
.Y(n_11869)
);

INVx1_ASAP7_75t_L g11870 ( 
.A(n_10266),
.Y(n_11870)
);

INVx2_ASAP7_75t_L g11871 ( 
.A(n_10266),
.Y(n_11871)
);

OAI21x1_ASAP7_75t_L g11872 ( 
.A1(n_10271),
.A2(n_8637),
.B(n_8631),
.Y(n_11872)
);

INVx1_ASAP7_75t_L g11873 ( 
.A(n_10283),
.Y(n_11873)
);

AND2x4_ASAP7_75t_L g11874 ( 
.A(n_9560),
.B(n_8881),
.Y(n_11874)
);

INVx2_ASAP7_75t_SL g11875 ( 
.A(n_10042),
.Y(n_11875)
);

INVx2_ASAP7_75t_SL g11876 ( 
.A(n_10042),
.Y(n_11876)
);

OAI21x1_ASAP7_75t_L g11877 ( 
.A1(n_10358),
.A2(n_8638),
.B(n_8637),
.Y(n_11877)
);

OAI21x1_ASAP7_75t_L g11878 ( 
.A1(n_10358),
.A2(n_8638),
.B(n_8637),
.Y(n_11878)
);

INVx1_ASAP7_75t_L g11879 ( 
.A(n_10285),
.Y(n_11879)
);

OAI21xp5_ASAP7_75t_L g11880 ( 
.A1(n_10119),
.A2(n_8339),
.B(n_8223),
.Y(n_11880)
);

AND2x2_ASAP7_75t_L g11881 ( 
.A(n_9555),
.B(n_8146),
.Y(n_11881)
);

INVx2_ASAP7_75t_L g11882 ( 
.A(n_10276),
.Y(n_11882)
);

AND2x4_ASAP7_75t_L g11883 ( 
.A(n_9560),
.B(n_9606),
.Y(n_11883)
);

INVx2_ASAP7_75t_L g11884 ( 
.A(n_10276),
.Y(n_11884)
);

OAI22xp33_ASAP7_75t_L g11885 ( 
.A1(n_9541),
.A2(n_9204),
.B1(n_8930),
.B2(n_9142),
.Y(n_11885)
);

INVx1_ASAP7_75t_L g11886 ( 
.A(n_10312),
.Y(n_11886)
);

OAI21x1_ASAP7_75t_L g11887 ( 
.A1(n_10358),
.A2(n_8638),
.B(n_8782),
.Y(n_11887)
);

INVx2_ASAP7_75t_SL g11888 ( 
.A(n_10042),
.Y(n_11888)
);

OA21x2_ASAP7_75t_L g11889 ( 
.A1(n_10483),
.A2(n_7962),
.B(n_7959),
.Y(n_11889)
);

INVx2_ASAP7_75t_L g11890 ( 
.A(n_10279),
.Y(n_11890)
);

INVx1_ASAP7_75t_L g11891 ( 
.A(n_10303),
.Y(n_11891)
);

AND2x2_ASAP7_75t_L g11892 ( 
.A(n_9555),
.B(n_8146),
.Y(n_11892)
);

NOR2xp33_ASAP7_75t_L g11893 ( 
.A(n_9356),
.B(n_9311),
.Y(n_11893)
);

INVx5_ASAP7_75t_L g11894 ( 
.A(n_9501),
.Y(n_11894)
);

AND2x2_ASAP7_75t_L g11895 ( 
.A(n_9555),
.B(n_8211),
.Y(n_11895)
);

INVxp67_ASAP7_75t_L g11896 ( 
.A(n_9796),
.Y(n_11896)
);

INVx1_ASAP7_75t_L g11897 ( 
.A(n_10294),
.Y(n_11897)
);

INVx1_ASAP7_75t_L g11898 ( 
.A(n_10294),
.Y(n_11898)
);

INVx2_ASAP7_75t_L g11899 ( 
.A(n_10280),
.Y(n_11899)
);

INVx2_ASAP7_75t_L g11900 ( 
.A(n_10280),
.Y(n_11900)
);

INVx2_ASAP7_75t_L g11901 ( 
.A(n_10286),
.Y(n_11901)
);

INVx2_ASAP7_75t_L g11902 ( 
.A(n_10296),
.Y(n_11902)
);

NAND2xp5_ASAP7_75t_L g11903 ( 
.A(n_9670),
.B(n_8755),
.Y(n_11903)
);

INVx2_ASAP7_75t_L g11904 ( 
.A(n_10296),
.Y(n_11904)
);

INVx1_ASAP7_75t_L g11905 ( 
.A(n_10312),
.Y(n_11905)
);

INVx2_ASAP7_75t_L g11906 ( 
.A(n_10303),
.Y(n_11906)
);

AND2x2_ASAP7_75t_L g11907 ( 
.A(n_9555),
.B(n_8211),
.Y(n_11907)
);

INVx2_ASAP7_75t_L g11908 ( 
.A(n_10315),
.Y(n_11908)
);

INVx1_ASAP7_75t_L g11909 ( 
.A(n_10315),
.Y(n_11909)
);

INVx2_ASAP7_75t_L g11910 ( 
.A(n_10316),
.Y(n_11910)
);

INVx1_ASAP7_75t_L g11911 ( 
.A(n_10316),
.Y(n_11911)
);

NAND2xp5_ASAP7_75t_L g11912 ( 
.A(n_9947),
.B(n_8854),
.Y(n_11912)
);

INVx1_ASAP7_75t_L g11913 ( 
.A(n_10361),
.Y(n_11913)
);

INVx3_ASAP7_75t_L g11914 ( 
.A(n_10383),
.Y(n_11914)
);

INVx1_ASAP7_75t_L g11915 ( 
.A(n_10361),
.Y(n_11915)
);

OR2x2_ASAP7_75t_L g11916 ( 
.A(n_10407),
.B(n_9250),
.Y(n_11916)
);

INVx1_ASAP7_75t_L g11917 ( 
.A(n_10362),
.Y(n_11917)
);

AND2x2_ASAP7_75t_L g11918 ( 
.A(n_9564),
.B(n_8211),
.Y(n_11918)
);

HB1xp67_ASAP7_75t_L g11919 ( 
.A(n_10324),
.Y(n_11919)
);

OR2x2_ASAP7_75t_L g11920 ( 
.A(n_10608),
.B(n_9088),
.Y(n_11920)
);

INVx1_ASAP7_75t_L g11921 ( 
.A(n_10362),
.Y(n_11921)
);

OAI21xp5_ASAP7_75t_L g11922 ( 
.A1(n_10514),
.A2(n_8339),
.B(n_8223),
.Y(n_11922)
);

AND2x2_ASAP7_75t_L g11923 ( 
.A(n_9564),
.B(n_8218),
.Y(n_11923)
);

INVx3_ASAP7_75t_L g11924 ( 
.A(n_10383),
.Y(n_11924)
);

INVx1_ASAP7_75t_L g11925 ( 
.A(n_10363),
.Y(n_11925)
);

INVx2_ASAP7_75t_L g11926 ( 
.A(n_10324),
.Y(n_11926)
);

OR2x2_ASAP7_75t_L g11927 ( 
.A(n_10670),
.B(n_9088),
.Y(n_11927)
);

INVx1_ASAP7_75t_L g11928 ( 
.A(n_10343),
.Y(n_11928)
);

AND2x2_ASAP7_75t_L g11929 ( 
.A(n_9564),
.B(n_8218),
.Y(n_11929)
);

BUFx12f_ASAP7_75t_L g11930 ( 
.A(n_10465),
.Y(n_11930)
);

BUFx6f_ASAP7_75t_L g11931 ( 
.A(n_9501),
.Y(n_11931)
);

AOI22xp33_ASAP7_75t_SL g11932 ( 
.A1(n_10965),
.A2(n_10116),
.B1(n_9377),
.B2(n_9784),
.Y(n_11932)
);

AOI22xp33_ASAP7_75t_L g11933 ( 
.A1(n_10956),
.A2(n_10646),
.B1(n_9539),
.B2(n_9675),
.Y(n_11933)
);

AND2x2_ASAP7_75t_L g11934 ( 
.A(n_10748),
.B(n_9654),
.Y(n_11934)
);

AOI22xp33_ASAP7_75t_L g11935 ( 
.A1(n_10933),
.A2(n_10646),
.B1(n_10156),
.B2(n_9551),
.Y(n_11935)
);

INVx1_ASAP7_75t_L g11936 ( 
.A(n_10735),
.Y(n_11936)
);

OAI222xp33_ASAP7_75t_L g11937 ( 
.A1(n_10732),
.A2(n_10713),
.B1(n_9921),
.B2(n_9346),
.C1(n_10090),
.C2(n_9903),
.Y(n_11937)
);

OR2x2_ASAP7_75t_L g11938 ( 
.A(n_10761),
.B(n_10670),
.Y(n_11938)
);

AOI22xp33_ASAP7_75t_L g11939 ( 
.A1(n_10980),
.A2(n_10156),
.B1(n_10356),
.B2(n_10349),
.Y(n_11939)
);

AOI22xp33_ASAP7_75t_SL g11940 ( 
.A1(n_10980),
.A2(n_9377),
.B1(n_10087),
.B2(n_10202),
.Y(n_11940)
);

OAI22xp5_ASAP7_75t_L g11941 ( 
.A1(n_11010),
.A2(n_9458),
.B1(n_9900),
.B2(n_9477),
.Y(n_11941)
);

AOI21xp5_ASAP7_75t_SL g11942 ( 
.A1(n_11467),
.A2(n_9530),
.B(n_10353),
.Y(n_11942)
);

OAI221xp5_ASAP7_75t_L g11943 ( 
.A1(n_10765),
.A2(n_10031),
.B1(n_10019),
.B2(n_9965),
.C(n_9829),
.Y(n_11943)
);

OAI22xp33_ASAP7_75t_L g11944 ( 
.A1(n_11175),
.A2(n_9900),
.B1(n_10663),
.B2(n_10431),
.Y(n_11944)
);

HB1xp67_ASAP7_75t_L g11945 ( 
.A(n_11457),
.Y(n_11945)
);

BUFx2_ASAP7_75t_L g11946 ( 
.A(n_11132),
.Y(n_11946)
);

NAND2xp5_ASAP7_75t_L g11947 ( 
.A(n_10861),
.B(n_9422),
.Y(n_11947)
);

AND2x2_ASAP7_75t_L g11948 ( 
.A(n_10794),
.B(n_9654),
.Y(n_11948)
);

AND2x2_ASAP7_75t_L g11949 ( 
.A(n_11433),
.B(n_9684),
.Y(n_11949)
);

INVx1_ASAP7_75t_L g11950 ( 
.A(n_10735),
.Y(n_11950)
);

INVx2_ASAP7_75t_L g11951 ( 
.A(n_10872),
.Y(n_11951)
);

AOI22xp33_ASAP7_75t_L g11952 ( 
.A1(n_11081),
.A2(n_9333),
.B1(n_9591),
.B2(n_9506),
.Y(n_11952)
);

NAND2xp5_ASAP7_75t_L g11953 ( 
.A(n_10861),
.B(n_9487),
.Y(n_11953)
);

AOI222xp33_ASAP7_75t_L g11954 ( 
.A1(n_10938),
.A2(n_10644),
.B1(n_10074),
.B2(n_9600),
.C1(n_9599),
.C2(n_10071),
.Y(n_11954)
);

OAI22xp5_ASAP7_75t_L g11955 ( 
.A1(n_11010),
.A2(n_9427),
.B1(n_9720),
.B2(n_10691),
.Y(n_11955)
);

AOI222xp33_ASAP7_75t_L g11956 ( 
.A1(n_11357),
.A2(n_9842),
.B1(n_9572),
.B2(n_9899),
.C1(n_9587),
.C2(n_9465),
.Y(n_11956)
);

O2A1O1Ixp33_ASAP7_75t_L g11957 ( 
.A1(n_11171),
.A2(n_10302),
.B(n_10382),
.C(n_9769),
.Y(n_11957)
);

AOI22xp33_ASAP7_75t_L g11958 ( 
.A1(n_11031),
.A2(n_9411),
.B1(n_9506),
.B2(n_9318),
.Y(n_11958)
);

OR2x2_ASAP7_75t_L g11959 ( 
.A(n_10806),
.B(n_9361),
.Y(n_11959)
);

INVx2_ASAP7_75t_L g11960 ( 
.A(n_10876),
.Y(n_11960)
);

AOI22xp5_ASAP7_75t_L g11961 ( 
.A1(n_11077),
.A2(n_9710),
.B1(n_10718),
.B2(n_9720),
.Y(n_11961)
);

AOI21xp33_ASAP7_75t_L g11962 ( 
.A1(n_10765),
.A2(n_9506),
.B(n_9411),
.Y(n_11962)
);

OAI22xp33_ASAP7_75t_L g11963 ( 
.A1(n_11620),
.A2(n_10431),
.B1(n_9570),
.B2(n_10155),
.Y(n_11963)
);

AOI22xp33_ASAP7_75t_L g11964 ( 
.A1(n_11215),
.A2(n_9506),
.B1(n_9411),
.B2(n_10499),
.Y(n_11964)
);

OAI211xp5_ASAP7_75t_L g11965 ( 
.A1(n_10732),
.A2(n_10570),
.B(n_10137),
.C(n_10139),
.Y(n_11965)
);

AND2x2_ASAP7_75t_L g11966 ( 
.A(n_10743),
.B(n_9684),
.Y(n_11966)
);

AOI22xp33_ASAP7_75t_L g11967 ( 
.A1(n_11318),
.A2(n_9506),
.B1(n_9411),
.B2(n_10523),
.Y(n_11967)
);

OAI22xp33_ASAP7_75t_L g11968 ( 
.A1(n_11183),
.A2(n_9570),
.B1(n_10155),
.B2(n_9628),
.Y(n_11968)
);

NOR2x1_ASAP7_75t_SL g11969 ( 
.A(n_10774),
.B(n_9411),
.Y(n_11969)
);

OAI22xp5_ASAP7_75t_L g11970 ( 
.A1(n_11716),
.A2(n_9628),
.B1(n_10570),
.B2(n_9979),
.Y(n_11970)
);

AOI22xp33_ASAP7_75t_SL g11971 ( 
.A1(n_10788),
.A2(n_9710),
.B1(n_10159),
.B2(n_10162),
.Y(n_11971)
);

OAI211xp5_ASAP7_75t_L g11972 ( 
.A1(n_11751),
.A2(n_10106),
.B(n_10160),
.C(n_10568),
.Y(n_11972)
);

AOI22xp33_ASAP7_75t_L g11973 ( 
.A1(n_11318),
.A2(n_11716),
.B1(n_10984),
.B2(n_10968),
.Y(n_11973)
);

INVx2_ASAP7_75t_SL g11974 ( 
.A(n_10960),
.Y(n_11974)
);

NAND2xp5_ASAP7_75t_L g11975 ( 
.A(n_11089),
.B(n_9548),
.Y(n_11975)
);

INVx1_ASAP7_75t_L g11976 ( 
.A(n_10740),
.Y(n_11976)
);

INVx1_ASAP7_75t_L g11977 ( 
.A(n_10740),
.Y(n_11977)
);

AND2x2_ASAP7_75t_L g11978 ( 
.A(n_10793),
.B(n_10189),
.Y(n_11978)
);

OAI221xp5_ASAP7_75t_L g11979 ( 
.A1(n_11424),
.A2(n_10700),
.B1(n_10526),
.B2(n_10637),
.C(n_10528),
.Y(n_11979)
);

AOI221xp5_ASAP7_75t_L g11980 ( 
.A1(n_11424),
.A2(n_11461),
.B1(n_11770),
.B2(n_11469),
.C(n_11751),
.Y(n_11980)
);

INVx5_ASAP7_75t_SL g11981 ( 
.A(n_11423),
.Y(n_11981)
);

INVx2_ASAP7_75t_L g11982 ( 
.A(n_10912),
.Y(n_11982)
);

INVx2_ASAP7_75t_L g11983 ( 
.A(n_10966),
.Y(n_11983)
);

INVx1_ASAP7_75t_L g11984 ( 
.A(n_11585),
.Y(n_11984)
);

AOI22xp33_ASAP7_75t_L g11985 ( 
.A1(n_10845),
.A2(n_9500),
.B1(n_9515),
.B2(n_9505),
.Y(n_11985)
);

NAND4xp25_ASAP7_75t_L g11986 ( 
.A(n_10756),
.B(n_9701),
.C(n_9700),
.D(n_10159),
.Y(n_11986)
);

BUFx6f_ASAP7_75t_L g11987 ( 
.A(n_10725),
.Y(n_11987)
);

AOI22xp33_ASAP7_75t_L g11988 ( 
.A1(n_10762),
.A2(n_9563),
.B1(n_9648),
.B2(n_9637),
.Y(n_11988)
);

A2O1A1Ixp33_ASAP7_75t_L g11989 ( 
.A1(n_10842),
.A2(n_10491),
.B(n_10703),
.C(n_9741),
.Y(n_11989)
);

OA21x2_ASAP7_75t_L g11990 ( 
.A1(n_11511),
.A2(n_9741),
.B(n_9706),
.Y(n_11990)
);

OAI22xp33_ASAP7_75t_L g11991 ( 
.A1(n_10779),
.A2(n_9324),
.B1(n_9336),
.B2(n_10448),
.Y(n_11991)
);

AND2x2_ASAP7_75t_L g11992 ( 
.A(n_10800),
.B(n_10189),
.Y(n_11992)
);

INVx1_ASAP7_75t_L g11993 ( 
.A(n_11591),
.Y(n_11993)
);

AND2x4_ASAP7_75t_L g11994 ( 
.A(n_11415),
.B(n_10189),
.Y(n_11994)
);

NOR2xp67_ASAP7_75t_L g11995 ( 
.A(n_11496),
.B(n_9564),
.Y(n_11995)
);

AOI22xp33_ASAP7_75t_L g11996 ( 
.A1(n_11827),
.A2(n_9662),
.B1(n_9463),
.B2(n_9471),
.Y(n_11996)
);

INVx2_ASAP7_75t_L g11997 ( 
.A(n_10974),
.Y(n_11997)
);

AOI211xp5_ASAP7_75t_L g11998 ( 
.A1(n_11212),
.A2(n_9944),
.B(n_10718),
.C(n_10299),
.Y(n_11998)
);

INVx2_ASAP7_75t_L g11999 ( 
.A(n_10992),
.Y(n_11999)
);

AOI22xp33_ASAP7_75t_SL g12000 ( 
.A1(n_11725),
.A2(n_9646),
.B1(n_9797),
.B2(n_9793),
.Y(n_12000)
);

OAI21xp33_ASAP7_75t_L g12001 ( 
.A1(n_11461),
.A2(n_11469),
.B(n_11770),
.Y(n_12001)
);

AOI22xp33_ASAP7_75t_L g12002 ( 
.A1(n_11219),
.A2(n_9330),
.B1(n_9744),
.B2(n_9742),
.Y(n_12002)
);

AOI22xp33_ASAP7_75t_L g12003 ( 
.A1(n_10746),
.A2(n_10395),
.B1(n_10423),
.B2(n_9661),
.Y(n_12003)
);

INVx2_ASAP7_75t_L g12004 ( 
.A(n_11074),
.Y(n_12004)
);

NAND2xp5_ASAP7_75t_L g12005 ( 
.A(n_10729),
.B(n_10498),
.Y(n_12005)
);

AND2x2_ASAP7_75t_L g12006 ( 
.A(n_11371),
.B(n_10310),
.Y(n_12006)
);

AND2x4_ASAP7_75t_L g12007 ( 
.A(n_11415),
.B(n_10310),
.Y(n_12007)
);

NAND2xp5_ASAP7_75t_L g12008 ( 
.A(n_11903),
.B(n_9764),
.Y(n_12008)
);

AND2x2_ASAP7_75t_L g12009 ( 
.A(n_10979),
.B(n_10310),
.Y(n_12009)
);

OAI221xp5_ASAP7_75t_SL g12010 ( 
.A1(n_11384),
.A2(n_10186),
.B1(n_10184),
.B2(n_10223),
.C(n_10209),
.Y(n_12010)
);

OR2x6_ASAP7_75t_L g12011 ( 
.A(n_11206),
.B(n_9499),
.Y(n_12011)
);

AOI22xp33_ASAP7_75t_L g12012 ( 
.A1(n_10746),
.A2(n_9783),
.B1(n_9698),
.B2(n_9633),
.Y(n_12012)
);

AOI21xp33_ASAP7_75t_L g12013 ( 
.A1(n_11212),
.A2(n_9336),
.B(n_9324),
.Y(n_12013)
);

AND2x2_ASAP7_75t_L g12014 ( 
.A(n_10907),
.B(n_10371),
.Y(n_12014)
);

INVx1_ASAP7_75t_L g12015 ( 
.A(n_11573),
.Y(n_12015)
);

AO21x2_ASAP7_75t_L g12016 ( 
.A1(n_11505),
.A2(n_10059),
.B(n_9927),
.Y(n_12016)
);

OAI221xp5_ASAP7_75t_L g12017 ( 
.A1(n_11384),
.A2(n_10288),
.B1(n_10320),
.B2(n_10305),
.C(n_10281),
.Y(n_12017)
);

OR2x2_ASAP7_75t_L g12018 ( 
.A(n_10888),
.B(n_9361),
.Y(n_12018)
);

AOI22xp33_ASAP7_75t_L g12019 ( 
.A1(n_11510),
.A2(n_9616),
.B1(n_9557),
.B2(n_9584),
.Y(n_12019)
);

AOI33xp33_ASAP7_75t_L g12020 ( 
.A1(n_11618),
.A2(n_10386),
.A3(n_10330),
.B1(n_10379),
.B2(n_10327),
.B3(n_10437),
.Y(n_12020)
);

NAND2xp5_ASAP7_75t_L g12021 ( 
.A(n_11091),
.B(n_11656),
.Y(n_12021)
);

AND2x2_ASAP7_75t_SL g12022 ( 
.A(n_11418),
.B(n_9723),
.Y(n_12022)
);

AOI22xp33_ASAP7_75t_L g12023 ( 
.A1(n_11405),
.A2(n_9557),
.B1(n_9584),
.B2(n_9501),
.Y(n_12023)
);

AND2x2_ASAP7_75t_L g12024 ( 
.A(n_10928),
.B(n_10371),
.Y(n_12024)
);

INVxp67_ASAP7_75t_L g12025 ( 
.A(n_11191),
.Y(n_12025)
);

AOI22xp33_ASAP7_75t_L g12026 ( 
.A1(n_11505),
.A2(n_9557),
.B1(n_9584),
.B2(n_9501),
.Y(n_12026)
);

AOI222xp33_ASAP7_75t_L g12027 ( 
.A1(n_11128),
.A2(n_10480),
.B1(n_9953),
.B2(n_9925),
.C1(n_9797),
.C2(n_9805),
.Y(n_12027)
);

CKINVDCx20_ASAP7_75t_R g12028 ( 
.A(n_10911),
.Y(n_12028)
);

OAI22xp5_ASAP7_75t_L g12029 ( 
.A1(n_10779),
.A2(n_9502),
.B1(n_9694),
.B2(n_9679),
.Y(n_12029)
);

AOI22xp33_ASAP7_75t_L g12030 ( 
.A1(n_11828),
.A2(n_9584),
.B1(n_9761),
.B2(n_9557),
.Y(n_12030)
);

AOI22xp33_ASAP7_75t_L g12031 ( 
.A1(n_11094),
.A2(n_9584),
.B1(n_9761),
.B2(n_9557),
.Y(n_12031)
);

OAI221xp5_ASAP7_75t_L g12032 ( 
.A1(n_10864),
.A2(n_10453),
.B1(n_10205),
.B2(n_9934),
.C(n_9931),
.Y(n_12032)
);

OAI221xp5_ASAP7_75t_L g12033 ( 
.A1(n_11512),
.A2(n_10078),
.B1(n_10187),
.B2(n_10199),
.C(n_9565),
.Y(n_12033)
);

AND2x2_ASAP7_75t_L g12034 ( 
.A(n_10931),
.B(n_10371),
.Y(n_12034)
);

OAI22xp33_ASAP7_75t_L g12035 ( 
.A1(n_11692),
.A2(n_9324),
.B1(n_9336),
.B2(n_9991),
.Y(n_12035)
);

OAI22xp5_ASAP7_75t_L g12036 ( 
.A1(n_11396),
.A2(n_11144),
.B1(n_11896),
.B2(n_11851),
.Y(n_12036)
);

NAND2xp5_ASAP7_75t_L g12037 ( 
.A(n_11795),
.B(n_9764),
.Y(n_12037)
);

AND2x2_ASAP7_75t_L g12038 ( 
.A(n_10943),
.B(n_10955),
.Y(n_12038)
);

INVx2_ASAP7_75t_SL g12039 ( 
.A(n_10769),
.Y(n_12039)
);

NAND2xp5_ASAP7_75t_L g12040 ( 
.A(n_11842),
.B(n_11053),
.Y(n_12040)
);

INVx2_ASAP7_75t_L g12041 ( 
.A(n_11088),
.Y(n_12041)
);

AND2x2_ASAP7_75t_L g12042 ( 
.A(n_10976),
.B(n_10451),
.Y(n_12042)
);

BUFx4f_ASAP7_75t_SL g12043 ( 
.A(n_10911),
.Y(n_12043)
);

AOI21xp33_ASAP7_75t_L g12044 ( 
.A1(n_11056),
.A2(n_9336),
.B(n_9324),
.Y(n_12044)
);

INVx1_ASAP7_75t_L g12045 ( 
.A(n_11573),
.Y(n_12045)
);

AND2x4_ASAP7_75t_L g12046 ( 
.A(n_10879),
.B(n_10451),
.Y(n_12046)
);

OAI22xp5_ASAP7_75t_L g12047 ( 
.A1(n_11144),
.A2(n_9987),
.B1(n_9819),
.B2(n_9817),
.Y(n_12047)
);

OAI22xp33_ASAP7_75t_L g12048 ( 
.A1(n_11363),
.A2(n_9324),
.B1(n_9336),
.B2(n_9765),
.Y(n_12048)
);

NAND2xp5_ASAP7_75t_L g12049 ( 
.A(n_11858),
.B(n_9786),
.Y(n_12049)
);

OR2x2_ASAP7_75t_L g12050 ( 
.A(n_11843),
.B(n_10225),
.Y(n_12050)
);

AOI222xp33_ASAP7_75t_L g12051 ( 
.A1(n_11806),
.A2(n_9863),
.B1(n_9793),
.B2(n_9888),
.C1(n_9885),
.C2(n_9805),
.Y(n_12051)
);

AOI221xp5_ASAP7_75t_L g12052 ( 
.A1(n_11885),
.A2(n_9888),
.B1(n_9926),
.B2(n_9885),
.C(n_9863),
.Y(n_12052)
);

NAND2xp5_ASAP7_75t_L g12053 ( 
.A(n_11607),
.B(n_9786),
.Y(n_12053)
);

OAI221xp5_ASAP7_75t_L g12054 ( 
.A1(n_11309),
.A2(n_11880),
.B1(n_11678),
.B2(n_11755),
.C(n_11786),
.Y(n_12054)
);

NAND2xp5_ASAP7_75t_L g12055 ( 
.A(n_11611),
.B(n_9836),
.Y(n_12055)
);

NAND2xp5_ASAP7_75t_L g12056 ( 
.A(n_11232),
.B(n_9836),
.Y(n_12056)
);

INVx1_ASAP7_75t_L g12057 ( 
.A(n_11585),
.Y(n_12057)
);

AO221x1_ASAP7_75t_L g12058 ( 
.A1(n_11885),
.A2(n_10185),
.B1(n_10682),
.B2(n_10545),
.C(n_9942),
.Y(n_12058)
);

CKINVDCx5p33_ASAP7_75t_R g12059 ( 
.A(n_11237),
.Y(n_12059)
);

OAI21x1_ASAP7_75t_L g12060 ( 
.A1(n_11105),
.A2(n_9678),
.B(n_9428),
.Y(n_12060)
);

NAND2xp5_ASAP7_75t_L g12061 ( 
.A(n_11522),
.B(n_9884),
.Y(n_12061)
);

OAI22xp5_ASAP7_75t_L g12062 ( 
.A1(n_11132),
.A2(n_9816),
.B1(n_10047),
.B2(n_9749),
.Y(n_12062)
);

NAND2xp5_ASAP7_75t_SL g12063 ( 
.A(n_11054),
.B(n_9723),
.Y(n_12063)
);

AOI22xp33_ASAP7_75t_L g12064 ( 
.A1(n_10901),
.A2(n_9584),
.B1(n_9761),
.B2(n_9557),
.Y(n_12064)
);

OR2x2_ASAP7_75t_L g12065 ( 
.A(n_10850),
.B(n_10231),
.Y(n_12065)
);

INVx1_ASAP7_75t_L g12066 ( 
.A(n_11619),
.Y(n_12066)
);

OAI22xp33_ASAP7_75t_L g12067 ( 
.A1(n_11801),
.A2(n_9619),
.B1(n_8713),
.B2(n_8930),
.Y(n_12067)
);

INVx2_ASAP7_75t_SL g12068 ( 
.A(n_10769),
.Y(n_12068)
);

AND2x4_ASAP7_75t_L g12069 ( 
.A(n_10879),
.B(n_10451),
.Y(n_12069)
);

NOR2xp33_ASAP7_75t_L g12070 ( 
.A(n_10801),
.B(n_9935),
.Y(n_12070)
);

AOI22xp33_ASAP7_75t_L g12071 ( 
.A1(n_11225),
.A2(n_9818),
.B1(n_9824),
.B2(n_9761),
.Y(n_12071)
);

OAI22xp5_ASAP7_75t_L g12072 ( 
.A1(n_11596),
.A2(n_9780),
.B1(n_10089),
.B2(n_9567),
.Y(n_12072)
);

AOI22xp33_ASAP7_75t_L g12073 ( 
.A1(n_11225),
.A2(n_9818),
.B1(n_9824),
.B2(n_9761),
.Y(n_12073)
);

AOI21xp33_ASAP7_75t_SL g12074 ( 
.A1(n_10801),
.A2(n_10167),
.B(n_9839),
.Y(n_12074)
);

BUFx3_ASAP7_75t_L g12075 ( 
.A(n_10917),
.Y(n_12075)
);

AOI22xp33_ASAP7_75t_L g12076 ( 
.A1(n_11057),
.A2(n_9818),
.B1(n_9824),
.B2(n_9761),
.Y(n_12076)
);

AOI21xp33_ASAP7_75t_L g12077 ( 
.A1(n_11370),
.A2(n_10934),
.B(n_11540),
.Y(n_12077)
);

AOI22xp33_ASAP7_75t_L g12078 ( 
.A1(n_10934),
.A2(n_9824),
.B1(n_9890),
.B2(n_9818),
.Y(n_12078)
);

AOI22xp33_ASAP7_75t_SL g12079 ( 
.A1(n_11274),
.A2(n_9941),
.B1(n_9942),
.B2(n_9926),
.Y(n_12079)
);

OAI211xp5_ASAP7_75t_L g12080 ( 
.A1(n_11922),
.A2(n_10023),
.B(n_10028),
.C(n_9941),
.Y(n_12080)
);

OAI211xp5_ASAP7_75t_SL g12081 ( 
.A1(n_11519),
.A2(n_10073),
.B(n_10230),
.C(n_10197),
.Y(n_12081)
);

CKINVDCx20_ASAP7_75t_R g12082 ( 
.A(n_10917),
.Y(n_12082)
);

OAI22xp5_ASAP7_75t_L g12083 ( 
.A1(n_11597),
.A2(n_9735),
.B1(n_10420),
.B2(n_10416),
.Y(n_12083)
);

OA21x2_ASAP7_75t_L g12084 ( 
.A1(n_11228),
.A2(n_11260),
.B(n_11257),
.Y(n_12084)
);

AND2x2_ASAP7_75t_L g12085 ( 
.A(n_10986),
.B(n_10475),
.Y(n_12085)
);

BUFx8_ASAP7_75t_L g12086 ( 
.A(n_11206),
.Y(n_12086)
);

AOI221xp5_ASAP7_75t_L g12087 ( 
.A1(n_11370),
.A2(n_10032),
.B1(n_10038),
.B2(n_10028),
.C(n_10023),
.Y(n_12087)
);

A2O1A1Ixp33_ASAP7_75t_L g12088 ( 
.A1(n_10958),
.A2(n_10038),
.B(n_10061),
.C(n_10032),
.Y(n_12088)
);

AOI22xp33_ASAP7_75t_SL g12089 ( 
.A1(n_11677),
.A2(n_10126),
.B1(n_10150),
.B2(n_10061),
.Y(n_12089)
);

OAI22xp5_ASAP7_75t_L g12090 ( 
.A1(n_11706),
.A2(n_9812),
.B1(n_9794),
.B2(n_10436),
.Y(n_12090)
);

INVx1_ASAP7_75t_L g12091 ( 
.A(n_11616),
.Y(n_12091)
);

NAND3xp33_ASAP7_75t_L g12092 ( 
.A(n_11087),
.B(n_8077),
.C(n_10048),
.Y(n_12092)
);

OAI211xp5_ASAP7_75t_SL g12093 ( 
.A1(n_10930),
.A2(n_10275),
.B(n_9327),
.C(n_10574),
.Y(n_12093)
);

INVx1_ASAP7_75t_L g12094 ( 
.A(n_11616),
.Y(n_12094)
);

CKINVDCx5p33_ASAP7_75t_R g12095 ( 
.A(n_11237),
.Y(n_12095)
);

AOI221xp5_ASAP7_75t_L g12096 ( 
.A1(n_11540),
.A2(n_10150),
.B1(n_10126),
.B2(n_10300),
.C(n_10261),
.Y(n_12096)
);

INVx2_ASAP7_75t_SL g12097 ( 
.A(n_10958),
.Y(n_12097)
);

INVx4_ASAP7_75t_SL g12098 ( 
.A(n_10832),
.Y(n_12098)
);

AOI22xp33_ASAP7_75t_L g12099 ( 
.A1(n_10728),
.A2(n_9824),
.B1(n_9890),
.B2(n_9818),
.Y(n_12099)
);

AOI22xp33_ASAP7_75t_L g12100 ( 
.A1(n_11864),
.A2(n_9824),
.B1(n_9890),
.B2(n_9818),
.Y(n_12100)
);

AOI222xp33_ASAP7_75t_L g12101 ( 
.A1(n_10930),
.A2(n_10348),
.B1(n_10261),
.B2(n_10402),
.C1(n_10387),
.C2(n_10300),
.Y(n_12101)
);

AND2x2_ASAP7_75t_L g12102 ( 
.A(n_10993),
.B(n_10475),
.Y(n_12102)
);

AOI22xp33_ASAP7_75t_L g12103 ( 
.A1(n_11331),
.A2(n_10759),
.B1(n_10798),
.B2(n_10739),
.Y(n_12103)
);

AOI222xp33_ASAP7_75t_L g12104 ( 
.A1(n_11189),
.A2(n_10402),
.B1(n_10348),
.B2(n_10538),
.C1(n_10406),
.C2(n_10387),
.Y(n_12104)
);

OAI211xp5_ASAP7_75t_L g12105 ( 
.A1(n_11717),
.A2(n_10406),
.B(n_10717),
.C(n_10538),
.Y(n_12105)
);

AOI22xp33_ASAP7_75t_SL g12106 ( 
.A1(n_11626),
.A2(n_8077),
.B1(n_10719),
.B2(n_10717),
.Y(n_12106)
);

AOI222xp33_ASAP7_75t_L g12107 ( 
.A1(n_11117),
.A2(n_10719),
.B1(n_8710),
.B2(n_10554),
.C1(n_10551),
.C2(n_8850),
.Y(n_12107)
);

AND2x2_ASAP7_75t_L g12108 ( 
.A(n_10862),
.B(n_10475),
.Y(n_12108)
);

OAI22xp33_ASAP7_75t_L g12109 ( 
.A1(n_10821),
.A2(n_9619),
.B1(n_8713),
.B2(n_9644),
.Y(n_12109)
);

OAI211xp5_ASAP7_75t_L g12110 ( 
.A1(n_11772),
.A2(n_10425),
.B(n_10421),
.C(n_10496),
.Y(n_12110)
);

AO21x2_ASAP7_75t_L g12111 ( 
.A1(n_11257),
.A2(n_10059),
.B(n_9927),
.Y(n_12111)
);

AND2x2_ASAP7_75t_L g12112 ( 
.A(n_10867),
.B(n_11009),
.Y(n_12112)
);

INVx1_ASAP7_75t_L g12113 ( 
.A(n_11642),
.Y(n_12113)
);

AND2x4_ASAP7_75t_L g12114 ( 
.A(n_10879),
.B(n_10559),
.Y(n_12114)
);

OA21x2_ASAP7_75t_L g12115 ( 
.A1(n_11260),
.A2(n_10487),
.B(n_10483),
.Y(n_12115)
);

OAI221xp5_ASAP7_75t_L g12116 ( 
.A1(n_11087),
.A2(n_9982),
.B1(n_9707),
.B2(n_9703),
.C(n_10580),
.Y(n_12116)
);

AND2x4_ASAP7_75t_L g12117 ( 
.A(n_11354),
.B(n_10559),
.Y(n_12117)
);

OAI21xp33_ASAP7_75t_L g12118 ( 
.A1(n_11090),
.A2(n_10571),
.B(n_10520),
.Y(n_12118)
);

OAI22xp5_ASAP7_75t_L g12119 ( 
.A1(n_11729),
.A2(n_9286),
.B1(n_9799),
.B2(n_9723),
.Y(n_12119)
);

OAI22xp33_ASAP7_75t_L g12120 ( 
.A1(n_11126),
.A2(n_9619),
.B1(n_9644),
.B2(n_10042),
.Y(n_12120)
);

OAI22xp33_ASAP7_75t_L g12121 ( 
.A1(n_11292),
.A2(n_9619),
.B1(n_9644),
.B2(n_10042),
.Y(n_12121)
);

AOI22xp33_ASAP7_75t_L g12122 ( 
.A1(n_11331),
.A2(n_9922),
.B1(n_9989),
.B2(n_9890),
.Y(n_12122)
);

AND2x2_ASAP7_75t_L g12123 ( 
.A(n_11014),
.B(n_10559),
.Y(n_12123)
);

AOI22xp33_ASAP7_75t_SL g12124 ( 
.A1(n_11626),
.A2(n_7912),
.B1(n_7956),
.B2(n_7949),
.Y(n_12124)
);

AOI22xp33_ASAP7_75t_L g12125 ( 
.A1(n_10829),
.A2(n_9922),
.B1(n_9989),
.B2(n_9890),
.Y(n_12125)
);

AOI22xp33_ASAP7_75t_L g12126 ( 
.A1(n_11161),
.A2(n_11182),
.B1(n_11199),
.B2(n_11737),
.Y(n_12126)
);

BUFx4f_ASAP7_75t_SL g12127 ( 
.A(n_11291),
.Y(n_12127)
);

NAND2xp5_ASAP7_75t_L g12128 ( 
.A(n_11605),
.B(n_9884),
.Y(n_12128)
);

AO21x1_ASAP7_75t_L g12129 ( 
.A1(n_11490),
.A2(n_10513),
.B(n_9626),
.Y(n_12129)
);

BUFx2_ASAP7_75t_L g12130 ( 
.A(n_11930),
.Y(n_12130)
);

BUFx6f_ASAP7_75t_L g12131 ( 
.A(n_10725),
.Y(n_12131)
);

AOI22xp33_ASAP7_75t_L g12132 ( 
.A1(n_11737),
.A2(n_9922),
.B1(n_9989),
.B2(n_9890),
.Y(n_12132)
);

AOI221xp5_ASAP7_75t_L g12133 ( 
.A1(n_11312),
.A2(n_9538),
.B1(n_9392),
.B2(n_9351),
.C(n_8710),
.Y(n_12133)
);

INVx3_ASAP7_75t_L g12134 ( 
.A(n_11002),
.Y(n_12134)
);

INVx3_ASAP7_75t_L g12135 ( 
.A(n_11002),
.Y(n_12135)
);

AOI22xp33_ASAP7_75t_L g12136 ( 
.A1(n_11883),
.A2(n_11216),
.B1(n_11224),
.B2(n_11220),
.Y(n_12136)
);

OR2x2_ASAP7_75t_L g12137 ( 
.A(n_11051),
.B(n_10588),
.Y(n_12137)
);

OAI211xp5_ASAP7_75t_L g12138 ( 
.A1(n_11772),
.A2(n_7928),
.B(n_8103),
.C(n_7980),
.Y(n_12138)
);

AND2x2_ASAP7_75t_L g12139 ( 
.A(n_11016),
.B(n_10609),
.Y(n_12139)
);

OAI221xp5_ASAP7_75t_L g12140 ( 
.A1(n_10958),
.A2(n_10613),
.B1(n_10239),
.B2(n_10365),
.C(n_10410),
.Y(n_12140)
);

AOI22xp33_ASAP7_75t_L g12141 ( 
.A1(n_11883),
.A2(n_9989),
.B1(n_9922),
.B2(n_10337),
.Y(n_12141)
);

OAI22xp5_ASAP7_75t_L g12142 ( 
.A1(n_11729),
.A2(n_10544),
.B1(n_9799),
.B2(n_9781),
.Y(n_12142)
);

OAI211xp5_ASAP7_75t_L g12143 ( 
.A1(n_11362),
.A2(n_7928),
.B(n_8103),
.C(n_7980),
.Y(n_12143)
);

AOI222xp33_ASAP7_75t_L g12144 ( 
.A1(n_11506),
.A2(n_8850),
.B1(n_9110),
.B2(n_8880),
.C1(n_9718),
.C2(n_8884),
.Y(n_12144)
);

INVx2_ASAP7_75t_L g12145 ( 
.A(n_11268),
.Y(n_12145)
);

OAI21xp5_ASAP7_75t_L g12146 ( 
.A1(n_10903),
.A2(n_10513),
.B(n_8339),
.Y(n_12146)
);

INVx1_ASAP7_75t_L g12147 ( 
.A(n_11739),
.Y(n_12147)
);

AND2x2_ASAP7_75t_L g12148 ( 
.A(n_11045),
.B(n_10609),
.Y(n_12148)
);

AOI22xp33_ASAP7_75t_L g12149 ( 
.A1(n_11883),
.A2(n_9989),
.B1(n_9922),
.B2(n_10337),
.Y(n_12149)
);

OAI21xp5_ASAP7_75t_L g12150 ( 
.A1(n_11030),
.A2(n_8223),
.B(n_8259),
.Y(n_12150)
);

INVx1_ASAP7_75t_L g12151 ( 
.A(n_11642),
.Y(n_12151)
);

INVx2_ASAP7_75t_SL g12152 ( 
.A(n_10840),
.Y(n_12152)
);

AOI22xp33_ASAP7_75t_L g12153 ( 
.A1(n_11247),
.A2(n_9989),
.B1(n_9922),
.B2(n_10337),
.Y(n_12153)
);

NOR2xp33_ASAP7_75t_L g12154 ( 
.A(n_11423),
.B(n_9985),
.Y(n_12154)
);

AOI211xp5_ASAP7_75t_L g12155 ( 
.A1(n_11030),
.A2(n_11080),
.B(n_11114),
.C(n_11044),
.Y(n_12155)
);

AOI221xp5_ASAP7_75t_L g12156 ( 
.A1(n_11412),
.A2(n_9392),
.B1(n_9538),
.B2(n_9351),
.C(n_10059),
.Y(n_12156)
);

OAI22xp5_ASAP7_75t_L g12157 ( 
.A1(n_10847),
.A2(n_11633),
.B1(n_10799),
.B2(n_11043),
.Y(n_12157)
);

OAI22xp5_ASAP7_75t_L g12158 ( 
.A1(n_11633),
.A2(n_10544),
.B1(n_9799),
.B2(n_9850),
.Y(n_12158)
);

OAI221xp5_ASAP7_75t_L g12159 ( 
.A1(n_11044),
.A2(n_10613),
.B1(n_10239),
.B2(n_10365),
.C(n_10410),
.Y(n_12159)
);

NOR2xp33_ASAP7_75t_L g12160 ( 
.A(n_11506),
.B(n_9561),
.Y(n_12160)
);

INVx3_ASAP7_75t_L g12161 ( 
.A(n_11002),
.Y(n_12161)
);

AOI21xp5_ASAP7_75t_L g12162 ( 
.A1(n_11304),
.A2(n_11707),
.B(n_10544),
.Y(n_12162)
);

AOI22xp5_ASAP7_75t_L g12163 ( 
.A1(n_11068),
.A2(n_10353),
.B1(n_9181),
.B2(n_10130),
.Y(n_12163)
);

AOI221xp5_ASAP7_75t_L g12164 ( 
.A1(n_11334),
.A2(n_9392),
.B1(n_9538),
.B2(n_9351),
.C(n_8160),
.Y(n_12164)
);

OAI22xp5_ASAP7_75t_L g12165 ( 
.A1(n_10799),
.A2(n_10544),
.B1(n_9799),
.B2(n_9789),
.Y(n_12165)
);

NOR2x1_ASAP7_75t_L g12166 ( 
.A(n_11354),
.B(n_10609),
.Y(n_12166)
);

INVx2_ASAP7_75t_L g12167 ( 
.A(n_11268),
.Y(n_12167)
);

AOI221xp5_ASAP7_75t_L g12168 ( 
.A1(n_11462),
.A2(n_8160),
.B1(n_8966),
.B2(n_9013),
.C(n_8541),
.Y(n_12168)
);

AOI222xp33_ASAP7_75t_L g12169 ( 
.A1(n_10832),
.A2(n_9110),
.B1(n_8880),
.B2(n_8884),
.C1(n_8825),
.C2(n_8799),
.Y(n_12169)
);

AOI22xp33_ASAP7_75t_L g12170 ( 
.A1(n_11258),
.A2(n_10365),
.B1(n_10410),
.B2(n_10337),
.Y(n_12170)
);

AND2x2_ASAP7_75t_L g12171 ( 
.A(n_11055),
.B(n_10631),
.Y(n_12171)
);

OAI22xp5_ASAP7_75t_L g12172 ( 
.A1(n_10799),
.A2(n_11043),
.B1(n_11147),
.B2(n_10824),
.Y(n_12172)
);

NAND2xp5_ASAP7_75t_L g12173 ( 
.A(n_11912),
.B(n_9910),
.Y(n_12173)
);

CKINVDCx20_ASAP7_75t_R g12174 ( 
.A(n_11291),
.Y(n_12174)
);

NOR2x1_ASAP7_75t_SL g12175 ( 
.A(n_10774),
.B(n_9619),
.Y(n_12175)
);

AOI22xp33_ASAP7_75t_L g12176 ( 
.A1(n_11277),
.A2(n_10410),
.B1(n_10413),
.B2(n_10365),
.Y(n_12176)
);

OAI221xp5_ASAP7_75t_L g12177 ( 
.A1(n_11080),
.A2(n_10613),
.B1(n_10239),
.B2(n_10446),
.C(n_10477),
.Y(n_12177)
);

AO21x2_ASAP7_75t_L g12178 ( 
.A1(n_11280),
.A2(n_10495),
.B(n_10487),
.Y(n_12178)
);

HB1xp67_ASAP7_75t_L g12179 ( 
.A(n_11457),
.Y(n_12179)
);

INVx1_ASAP7_75t_L g12180 ( 
.A(n_11591),
.Y(n_12180)
);

AOI22xp33_ASAP7_75t_SL g12181 ( 
.A1(n_11202),
.A2(n_7912),
.B1(n_7956),
.B2(n_7949),
.Y(n_12181)
);

AOI221xp5_ASAP7_75t_L g12182 ( 
.A1(n_11061),
.A2(n_11667),
.B1(n_11202),
.B2(n_11124),
.C(n_11195),
.Y(n_12182)
);

NAND3xp33_ASAP7_75t_L g12183 ( 
.A(n_11667),
.B(n_10053),
.C(n_10048),
.Y(n_12183)
);

BUFx2_ASAP7_75t_L g12184 ( 
.A(n_11930),
.Y(n_12184)
);

INVx8_ASAP7_75t_L g12185 ( 
.A(n_10725),
.Y(n_12185)
);

AOI22xp5_ASAP7_75t_L g12186 ( 
.A1(n_11068),
.A2(n_10353),
.B1(n_10130),
.B2(n_10210),
.Y(n_12186)
);

BUFx3_ASAP7_75t_L g12187 ( 
.A(n_11857),
.Y(n_12187)
);

OAI211xp5_ASAP7_75t_SL g12188 ( 
.A1(n_11114),
.A2(n_11195),
.B(n_11124),
.C(n_11430),
.Y(n_12188)
);

OAI211xp5_ASAP7_75t_SL g12189 ( 
.A1(n_11556),
.A2(n_9724),
.B(n_9382),
.C(n_9937),
.Y(n_12189)
);

OAI211xp5_ASAP7_75t_L g12190 ( 
.A1(n_10883),
.A2(n_7928),
.B(n_8103),
.C(n_7980),
.Y(n_12190)
);

AND2x2_ASAP7_75t_L g12191 ( 
.A(n_11103),
.B(n_10631),
.Y(n_12191)
);

NOR2x1_ASAP7_75t_SL g12192 ( 
.A(n_11364),
.B(n_11664),
.Y(n_12192)
);

AOI22xp5_ASAP7_75t_L g12193 ( 
.A1(n_11467),
.A2(n_10353),
.B1(n_10130),
.B2(n_10210),
.Y(n_12193)
);

INVx3_ASAP7_75t_L g12194 ( 
.A(n_11040),
.Y(n_12194)
);

AOI22xp33_ASAP7_75t_L g12195 ( 
.A1(n_11299),
.A2(n_10446),
.B1(n_10477),
.B2(n_10413),
.Y(n_12195)
);

NAND2xp5_ASAP7_75t_L g12196 ( 
.A(n_11107),
.B(n_9910),
.Y(n_12196)
);

OAI22xp33_ASAP7_75t_L g12197 ( 
.A1(n_10824),
.A2(n_9644),
.B1(n_10130),
.B2(n_10042),
.Y(n_12197)
);

AND2x2_ASAP7_75t_L g12198 ( 
.A(n_11127),
.B(n_10631),
.Y(n_12198)
);

NAND3xp33_ASAP7_75t_L g12199 ( 
.A(n_11667),
.B(n_10142),
.C(n_10053),
.Y(n_12199)
);

NAND2xp5_ASAP7_75t_L g12200 ( 
.A(n_11475),
.B(n_10076),
.Y(n_12200)
);

AOI22xp33_ASAP7_75t_L g12201 ( 
.A1(n_11313),
.A2(n_10446),
.B1(n_10477),
.B2(n_10413),
.Y(n_12201)
);

AOI22xp33_ASAP7_75t_L g12202 ( 
.A1(n_11321),
.A2(n_11338),
.B1(n_11345),
.B2(n_11333),
.Y(n_12202)
);

AOI22xp33_ASAP7_75t_SL g12203 ( 
.A1(n_11359),
.A2(n_7912),
.B1(n_7956),
.B2(n_7949),
.Y(n_12203)
);

A2O1A1Ixp33_ASAP7_75t_L g12204 ( 
.A1(n_11608),
.A2(n_8623),
.B(n_8947),
.C(n_8555),
.Y(n_12204)
);

HB1xp67_ASAP7_75t_L g12205 ( 
.A(n_11471),
.Y(n_12205)
);

INVx2_ASAP7_75t_L g12206 ( 
.A(n_11268),
.Y(n_12206)
);

AOI22xp33_ASAP7_75t_L g12207 ( 
.A1(n_11373),
.A2(n_10446),
.B1(n_10477),
.B2(n_10413),
.Y(n_12207)
);

AOI22xp33_ASAP7_75t_L g12208 ( 
.A1(n_11387),
.A2(n_10667),
.B1(n_10503),
.B2(n_9390),
.Y(n_12208)
);

OAI211xp5_ASAP7_75t_L g12209 ( 
.A1(n_10883),
.A2(n_7928),
.B(n_8103),
.C(n_7980),
.Y(n_12209)
);

AOI22xp33_ASAP7_75t_L g12210 ( 
.A1(n_11441),
.A2(n_10667),
.B1(n_10503),
.B2(n_9390),
.Y(n_12210)
);

AOI221xp5_ASAP7_75t_L g12211 ( 
.A1(n_11667),
.A2(n_11662),
.B1(n_11476),
.B2(n_11517),
.C(n_11491),
.Y(n_12211)
);

OAI321xp33_ASAP7_75t_L g12212 ( 
.A1(n_11490),
.A2(n_10613),
.A3(n_10239),
.B1(n_10422),
.B2(n_10450),
.C(n_10585),
.Y(n_12212)
);

OAI211xp5_ASAP7_75t_L g12213 ( 
.A1(n_10883),
.A2(n_7928),
.B(n_8103),
.C(n_7980),
.Y(n_12213)
);

INVx1_ASAP7_75t_L g12214 ( 
.A(n_11705),
.Y(n_12214)
);

AOI221xp5_ASAP7_75t_L g12215 ( 
.A1(n_11662),
.A2(n_8160),
.B1(n_8966),
.B2(n_9013),
.C(n_8049),
.Y(n_12215)
);

BUFx4f_ASAP7_75t_SL g12216 ( 
.A(n_11654),
.Y(n_12216)
);

OR2x2_ASAP7_75t_L g12217 ( 
.A(n_10744),
.B(n_10601),
.Y(n_12217)
);

OAI22xp33_ASAP7_75t_L g12218 ( 
.A1(n_10824),
.A2(n_9644),
.B1(n_10210),
.B2(n_10130),
.Y(n_12218)
);

OAI22xp5_ASAP7_75t_L g12219 ( 
.A1(n_11043),
.A2(n_8948),
.B1(n_9483),
.B2(n_9390),
.Y(n_12219)
);

AOI21xp5_ASAP7_75t_L g12220 ( 
.A1(n_11308),
.A2(n_9760),
.B(n_9000),
.Y(n_12220)
);

AND2x2_ASAP7_75t_L g12221 ( 
.A(n_11130),
.B(n_10641),
.Y(n_12221)
);

AOI22xp33_ASAP7_75t_SL g12222 ( 
.A1(n_11456),
.A2(n_7912),
.B1(n_7956),
.B2(n_7949),
.Y(n_12222)
);

AOI221xp5_ASAP7_75t_L g12223 ( 
.A1(n_11662),
.A2(n_8049),
.B1(n_8947),
.B2(n_8962),
.C(n_9008),
.Y(n_12223)
);

CKINVDCx5p33_ASAP7_75t_R g12224 ( 
.A(n_11609),
.Y(n_12224)
);

INVx6_ASAP7_75t_L g12225 ( 
.A(n_11703),
.Y(n_12225)
);

AOI22xp33_ASAP7_75t_SL g12226 ( 
.A1(n_11482),
.A2(n_7912),
.B1(n_7956),
.B2(n_7949),
.Y(n_12226)
);

AOI222xp33_ASAP7_75t_SL g12227 ( 
.A1(n_10881),
.A2(n_10167),
.B1(n_9980),
.B2(n_9435),
.C1(n_9325),
.C2(n_9457),
.Y(n_12227)
);

AOI22xp33_ASAP7_75t_L g12228 ( 
.A1(n_11554),
.A2(n_10667),
.B1(n_10503),
.B2(n_9483),
.Y(n_12228)
);

INVx2_ASAP7_75t_L g12229 ( 
.A(n_11276),
.Y(n_12229)
);

AOI22xp33_ASAP7_75t_L g12230 ( 
.A1(n_11638),
.A2(n_10667),
.B1(n_10503),
.B2(n_9483),
.Y(n_12230)
);

AND2x2_ASAP7_75t_L g12231 ( 
.A(n_11140),
.B(n_10641),
.Y(n_12231)
);

AOI22xp33_ASAP7_75t_L g12232 ( 
.A1(n_10725),
.A2(n_10731),
.B1(n_10805),
.B2(n_10795),
.Y(n_12232)
);

AOI221xp5_ASAP7_75t_L g12233 ( 
.A1(n_11471),
.A2(n_8049),
.B1(n_8962),
.B2(n_9008),
.C(n_9000),
.Y(n_12233)
);

NAND2xp5_ASAP7_75t_L g12234 ( 
.A(n_11488),
.B(n_10076),
.Y(n_12234)
);

OAI22xp33_ASAP7_75t_L g12235 ( 
.A1(n_11147),
.A2(n_10210),
.B1(n_10342),
.B2(n_10130),
.Y(n_12235)
);

OAI22xp5_ASAP7_75t_L g12236 ( 
.A1(n_11147),
.A2(n_8948),
.B1(n_9483),
.B2(n_9390),
.Y(n_12236)
);

OAI211xp5_ASAP7_75t_SL g12237 ( 
.A1(n_10764),
.A2(n_9709),
.B(n_10573),
.C(n_10414),
.Y(n_12237)
);

CKINVDCx20_ASAP7_75t_R g12238 ( 
.A(n_11654),
.Y(n_12238)
);

AND2x2_ASAP7_75t_L g12239 ( 
.A(n_11172),
.B(n_11180),
.Y(n_12239)
);

NAND2xp5_ASAP7_75t_L g12240 ( 
.A(n_11149),
.B(n_10414),
.Y(n_12240)
);

NAND2xp5_ASAP7_75t_L g12241 ( 
.A(n_11178),
.B(n_10573),
.Y(n_12241)
);

OAI31xp33_ASAP7_75t_SL g12242 ( 
.A1(n_11320),
.A2(n_9275),
.A3(n_10375),
.B(n_9214),
.Y(n_12242)
);

OAI22xp33_ASAP7_75t_L g12243 ( 
.A1(n_11499),
.A2(n_10210),
.B1(n_10397),
.B2(n_10342),
.Y(n_12243)
);

INVx4_ASAP7_75t_L g12244 ( 
.A(n_10731),
.Y(n_12244)
);

AND2x2_ASAP7_75t_L g12245 ( 
.A(n_11184),
.B(n_10641),
.Y(n_12245)
);

OAI22xp5_ASAP7_75t_L g12246 ( 
.A1(n_10752),
.A2(n_9514),
.B1(n_9727),
.B2(n_9889),
.Y(n_12246)
);

OA21x2_ASAP7_75t_L g12247 ( 
.A1(n_11280),
.A2(n_10495),
.B(n_10487),
.Y(n_12247)
);

INVx2_ASAP7_75t_L g12248 ( 
.A(n_11276),
.Y(n_12248)
);

OAI22xp5_ASAP7_75t_L g12249 ( 
.A1(n_10752),
.A2(n_9889),
.B1(n_10070),
.B2(n_9913),
.Y(n_12249)
);

NAND2xp33_ASAP7_75t_L g12250 ( 
.A(n_10840),
.B(n_10375),
.Y(n_12250)
);

AOI22x1_ASAP7_75t_L g12251 ( 
.A1(n_11703),
.A2(n_10331),
.B1(n_10192),
.B2(n_10142),
.Y(n_12251)
);

AOI21xp5_ASAP7_75t_L g12252 ( 
.A1(n_11636),
.A2(n_8596),
.B(n_10035),
.Y(n_12252)
);

OAI22xp5_ASAP7_75t_L g12253 ( 
.A1(n_10809),
.A2(n_9889),
.B1(n_10070),
.B2(n_9913),
.Y(n_12253)
);

AOI22xp5_ASAP7_75t_L g12254 ( 
.A1(n_11467),
.A2(n_10210),
.B1(n_10397),
.B2(n_10342),
.Y(n_12254)
);

NOR2x1_ASAP7_75t_L g12255 ( 
.A(n_11416),
.B(n_11446),
.Y(n_12255)
);

AND2x2_ASAP7_75t_L g12256 ( 
.A(n_11226),
.B(n_10709),
.Y(n_12256)
);

NOR2xp33_ASAP7_75t_L g12257 ( 
.A(n_10922),
.B(n_10505),
.Y(n_12257)
);

AOI22xp33_ASAP7_75t_L g12258 ( 
.A1(n_10731),
.A2(n_10142),
.B1(n_10152),
.B2(n_10053),
.Y(n_12258)
);

BUFx3_ASAP7_75t_L g12259 ( 
.A(n_11857),
.Y(n_12259)
);

OAI22xp33_ASAP7_75t_L g12260 ( 
.A1(n_11052),
.A2(n_10397),
.B1(n_10444),
.B2(n_10342),
.Y(n_12260)
);

AOI22xp33_ASAP7_75t_L g12261 ( 
.A1(n_10731),
.A2(n_10142),
.B1(n_10152),
.B2(n_10053),
.Y(n_12261)
);

NOR2xp33_ASAP7_75t_L g12262 ( 
.A(n_11240),
.B(n_10647),
.Y(n_12262)
);

AOI221xp5_ASAP7_75t_L g12263 ( 
.A1(n_11476),
.A2(n_8049),
.B1(n_8623),
.B2(n_8636),
.C(n_9121),
.Y(n_12263)
);

AOI21xp5_ASAP7_75t_L g12264 ( 
.A1(n_11320),
.A2(n_8596),
.B(n_10040),
.Y(n_12264)
);

OAI21x1_ASAP7_75t_L g12265 ( 
.A1(n_11738),
.A2(n_9678),
.B(n_9428),
.Y(n_12265)
);

INVx2_ASAP7_75t_L g12266 ( 
.A(n_11276),
.Y(n_12266)
);

AOI21xp5_ASAP7_75t_L g12267 ( 
.A1(n_11609),
.A2(n_9664),
.B(n_9499),
.Y(n_12267)
);

NAND2xp5_ASAP7_75t_SL g12268 ( 
.A(n_11894),
.B(n_10342),
.Y(n_12268)
);

INVx2_ASAP7_75t_L g12269 ( 
.A(n_11296),
.Y(n_12269)
);

OAI22xp33_ASAP7_75t_L g12270 ( 
.A1(n_11738),
.A2(n_10397),
.B1(n_10444),
.B2(n_10342),
.Y(n_12270)
);

OAI22xp5_ASAP7_75t_L g12271 ( 
.A1(n_10809),
.A2(n_9889),
.B1(n_10070),
.B2(n_9913),
.Y(n_12271)
);

OAI22xp5_ASAP7_75t_L g12272 ( 
.A1(n_10905),
.A2(n_11006),
.B1(n_11037),
.B2(n_10994),
.Y(n_12272)
);

AOI22xp33_ASAP7_75t_L g12273 ( 
.A1(n_10795),
.A2(n_10175),
.B1(n_10238),
.B2(n_10152),
.Y(n_12273)
);

OAI22xp33_ASAP7_75t_L g12274 ( 
.A1(n_11894),
.A2(n_10397),
.B1(n_10462),
.B2(n_10444),
.Y(n_12274)
);

INVx1_ASAP7_75t_L g12275 ( 
.A(n_11619),
.Y(n_12275)
);

AOI22xp33_ASAP7_75t_L g12276 ( 
.A1(n_10805),
.A2(n_10175),
.B1(n_10238),
.B2(n_10152),
.Y(n_12276)
);

AOI22xp33_ASAP7_75t_L g12277 ( 
.A1(n_10860),
.A2(n_10238),
.B1(n_10249),
.B2(n_10175),
.Y(n_12277)
);

INVx3_ASAP7_75t_L g12278 ( 
.A(n_11040),
.Y(n_12278)
);

HB1xp67_ASAP7_75t_L g12279 ( 
.A(n_11491),
.Y(n_12279)
);

OR2x6_ASAP7_75t_L g12280 ( 
.A(n_11703),
.B(n_9499),
.Y(n_12280)
);

AOI22xp33_ASAP7_75t_L g12281 ( 
.A1(n_10860),
.A2(n_10238),
.B1(n_10249),
.B2(n_10175),
.Y(n_12281)
);

AND2x2_ASAP7_75t_L g12282 ( 
.A(n_11241),
.B(n_10709),
.Y(n_12282)
);

INVx2_ASAP7_75t_SL g12283 ( 
.A(n_10863),
.Y(n_12283)
);

OAI22xp33_ASAP7_75t_L g12284 ( 
.A1(n_11894),
.A2(n_10397),
.B1(n_10462),
.B2(n_10444),
.Y(n_12284)
);

INVx1_ASAP7_75t_L g12285 ( 
.A(n_11702),
.Y(n_12285)
);

INVx1_ASAP7_75t_L g12286 ( 
.A(n_11702),
.Y(n_12286)
);

INVx1_ASAP7_75t_L g12287 ( 
.A(n_11816),
.Y(n_12287)
);

NAND3xp33_ASAP7_75t_L g12288 ( 
.A(n_10957),
.B(n_10412),
.C(n_10249),
.Y(n_12288)
);

OAI22xp33_ASAP7_75t_L g12289 ( 
.A1(n_11894),
.A2(n_10462),
.B1(n_10478),
.B2(n_10444),
.Y(n_12289)
);

INVx1_ASAP7_75t_L g12290 ( 
.A(n_11816),
.Y(n_12290)
);

AOI22xp33_ASAP7_75t_L g12291 ( 
.A1(n_10904),
.A2(n_10412),
.B1(n_10249),
.B2(n_10070),
.Y(n_12291)
);

INVx2_ASAP7_75t_L g12292 ( 
.A(n_11296),
.Y(n_12292)
);

AND2x2_ASAP7_75t_L g12293 ( 
.A(n_11558),
.B(n_11256),
.Y(n_12293)
);

NAND2xp5_ASAP7_75t_L g12294 ( 
.A(n_11187),
.B(n_10591),
.Y(n_12294)
);

HB1xp67_ASAP7_75t_L g12295 ( 
.A(n_11517),
.Y(n_12295)
);

INVx1_ASAP7_75t_L g12296 ( 
.A(n_11632),
.Y(n_12296)
);

AND2x2_ASAP7_75t_L g12297 ( 
.A(n_11271),
.B(n_10709),
.Y(n_12297)
);

INVx2_ASAP7_75t_L g12298 ( 
.A(n_11296),
.Y(n_12298)
);

AOI22xp33_ASAP7_75t_L g12299 ( 
.A1(n_10904),
.A2(n_10412),
.B1(n_10104),
.B2(n_10147),
.Y(n_12299)
);

OAI221xp5_ASAP7_75t_L g12300 ( 
.A1(n_11310),
.A2(n_10613),
.B1(n_10239),
.B2(n_9360),
.C(n_9435),
.Y(n_12300)
);

AOI22xp33_ASAP7_75t_L g12301 ( 
.A1(n_11029),
.A2(n_10412),
.B1(n_10104),
.B2(n_10147),
.Y(n_12301)
);

BUFx6f_ASAP7_75t_L g12302 ( 
.A(n_10724),
.Y(n_12302)
);

A2O1A1Ixp33_ASAP7_75t_L g12303 ( 
.A1(n_11267),
.A2(n_8555),
.B(n_8592),
.C(n_8870),
.Y(n_12303)
);

AND2x2_ASAP7_75t_L g12304 ( 
.A(n_11346),
.B(n_10192),
.Y(n_12304)
);

AOI22xp33_ASAP7_75t_L g12305 ( 
.A1(n_11029),
.A2(n_11038),
.B1(n_11042),
.B2(n_11041),
.Y(n_12305)
);

AOI22xp33_ASAP7_75t_SL g12306 ( 
.A1(n_10997),
.A2(n_7912),
.B1(n_7956),
.B2(n_7949),
.Y(n_12306)
);

AOI22xp33_ASAP7_75t_L g12307 ( 
.A1(n_11038),
.A2(n_10104),
.B1(n_10147),
.B2(n_9913),
.Y(n_12307)
);

AOI22xp33_ASAP7_75t_L g12308 ( 
.A1(n_11041),
.A2(n_10147),
.B1(n_10104),
.B2(n_10699),
.Y(n_12308)
);

AO21x2_ASAP7_75t_L g12309 ( 
.A1(n_11281),
.A2(n_10500),
.B(n_10495),
.Y(n_12309)
);

NAND2xp5_ASAP7_75t_L g12310 ( 
.A(n_11294),
.B(n_10591),
.Y(n_12310)
);

INVx1_ASAP7_75t_L g12311 ( 
.A(n_11632),
.Y(n_12311)
);

AOI21xp33_ASAP7_75t_SL g12312 ( 
.A1(n_10863),
.A2(n_10706),
.B(n_10039),
.Y(n_12312)
);

OR2x2_ASAP7_75t_L g12313 ( 
.A(n_10890),
.B(n_10655),
.Y(n_12313)
);

INVx1_ASAP7_75t_L g12314 ( 
.A(n_11690),
.Y(n_12314)
);

BUFx4f_ASAP7_75t_SL g12315 ( 
.A(n_11782),
.Y(n_12315)
);

AOI22xp33_ASAP7_75t_L g12316 ( 
.A1(n_11042),
.A2(n_11073),
.B1(n_11771),
.B2(n_10881),
.Y(n_12316)
);

AOI22xp33_ASAP7_75t_SL g12317 ( 
.A1(n_10997),
.A2(n_9855),
.B1(n_9848),
.B2(n_9171),
.Y(n_12317)
);

INVx3_ASAP7_75t_L g12318 ( 
.A(n_11141),
.Y(n_12318)
);

AND2x2_ASAP7_75t_L g12319 ( 
.A(n_11375),
.B(n_10331),
.Y(n_12319)
);

AOI221xp5_ASAP7_75t_L g12320 ( 
.A1(n_11555),
.A2(n_8049),
.B1(n_9121),
.B2(n_9023),
.C(n_8372),
.Y(n_12320)
);

AND2x2_ASAP7_75t_L g12321 ( 
.A(n_11389),
.B(n_10444),
.Y(n_12321)
);

AOI22xp33_ASAP7_75t_L g12322 ( 
.A1(n_11073),
.A2(n_10699),
.B1(n_9607),
.B2(n_9606),
.Y(n_12322)
);

AOI22xp33_ASAP7_75t_L g12323 ( 
.A1(n_11771),
.A2(n_9607),
.B1(n_9606),
.B2(n_10206),
.Y(n_12323)
);

OAI33xp33_ASAP7_75t_L g12324 ( 
.A1(n_10726),
.A2(n_8923),
.A3(n_8854),
.B1(n_8826),
.B2(n_10329),
.B3(n_10325),
.Y(n_12324)
);

INVx1_ASAP7_75t_L g12325 ( 
.A(n_11690),
.Y(n_12325)
);

BUFx6f_ASAP7_75t_L g12326 ( 
.A(n_10724),
.Y(n_12326)
);

AOI221xp5_ASAP7_75t_L g12327 ( 
.A1(n_11555),
.A2(n_8188),
.B1(n_9029),
.B2(n_8988),
.C(n_9122),
.Y(n_12327)
);

A2O1A1Ixp33_ASAP7_75t_L g12328 ( 
.A1(n_11285),
.A2(n_8592),
.B(n_8870),
.C(n_8259),
.Y(n_12328)
);

AOI22xp33_ASAP7_75t_L g12329 ( 
.A1(n_11771),
.A2(n_9607),
.B1(n_10272),
.B2(n_9762),
.Y(n_12329)
);

OAI21xp5_ASAP7_75t_SL g12330 ( 
.A1(n_11834),
.A2(n_10404),
.B(n_10388),
.Y(n_12330)
);

AOI22xp5_ASAP7_75t_L g12331 ( 
.A1(n_10881),
.A2(n_10478),
.B1(n_10488),
.B2(n_10462),
.Y(n_12331)
);

HB1xp67_ASAP7_75t_L g12332 ( 
.A(n_11563),
.Y(n_12332)
);

AOI22xp33_ASAP7_75t_L g12333 ( 
.A1(n_10881),
.A2(n_9762),
.B1(n_9766),
.B2(n_9686),
.Y(n_12333)
);

OAI22xp5_ASAP7_75t_L g12334 ( 
.A1(n_10905),
.A2(n_8968),
.B1(n_8662),
.B2(n_8730),
.Y(n_12334)
);

INVx1_ASAP7_75t_L g12335 ( 
.A(n_11739),
.Y(n_12335)
);

OAI22xp5_ASAP7_75t_L g12336 ( 
.A1(n_10994),
.A2(n_8968),
.B1(n_8700),
.B2(n_8730),
.Y(n_12336)
);

BUFx12f_ASAP7_75t_L g12337 ( 
.A(n_11019),
.Y(n_12337)
);

INVx1_ASAP7_75t_L g12338 ( 
.A(n_11919),
.Y(n_12338)
);

OAI22xp5_ASAP7_75t_L g12339 ( 
.A1(n_11006),
.A2(n_8700),
.B1(n_8970),
.B2(n_9116),
.Y(n_12339)
);

AOI22xp33_ASAP7_75t_L g12340 ( 
.A1(n_10881),
.A2(n_9762),
.B1(n_9766),
.B2(n_9686),
.Y(n_12340)
);

INVx1_ASAP7_75t_L g12341 ( 
.A(n_11705),
.Y(n_12341)
);

NOR4xp25_ASAP7_75t_L g12342 ( 
.A(n_11495),
.B(n_10640),
.C(n_10622),
.D(n_8988),
.Y(n_12342)
);

OA21x2_ASAP7_75t_L g12343 ( 
.A1(n_11281),
.A2(n_10502),
.B(n_10500),
.Y(n_12343)
);

OAI221xp5_ASAP7_75t_L g12344 ( 
.A1(n_11310),
.A2(n_9360),
.B1(n_9457),
.B2(n_9353),
.C(n_9325),
.Y(n_12344)
);

AND2x2_ASAP7_75t_L g12345 ( 
.A(n_11394),
.B(n_10462),
.Y(n_12345)
);

OA21x2_ASAP7_75t_L g12346 ( 
.A1(n_11282),
.A2(n_10502),
.B(n_10500),
.Y(n_12346)
);

INVx1_ASAP7_75t_L g12347 ( 
.A(n_11790),
.Y(n_12347)
);

INVx2_ASAP7_75t_L g12348 ( 
.A(n_11314),
.Y(n_12348)
);

OAI21x1_ASAP7_75t_L g12349 ( 
.A1(n_11598),
.A2(n_10204),
.B(n_10165),
.Y(n_12349)
);

AOI22xp33_ASAP7_75t_L g12350 ( 
.A1(n_11846),
.A2(n_9766),
.B1(n_9801),
.B2(n_9686),
.Y(n_12350)
);

BUFx2_ASAP7_75t_L g12351 ( 
.A(n_11868),
.Y(n_12351)
);

AOI22xp33_ASAP7_75t_L g12352 ( 
.A1(n_11819),
.A2(n_9806),
.B1(n_9810),
.B2(n_9801),
.Y(n_12352)
);

AOI33xp33_ASAP7_75t_L g12353 ( 
.A1(n_11495),
.A2(n_8455),
.A3(n_9248),
.B1(n_9116),
.B2(n_9039),
.B3(n_9111),
.Y(n_12353)
);

AND2x2_ASAP7_75t_L g12354 ( 
.A(n_11650),
.B(n_11668),
.Y(n_12354)
);

AND2x4_ASAP7_75t_L g12355 ( 
.A(n_11416),
.B(n_9499),
.Y(n_12355)
);

AOI222xp33_ASAP7_75t_L g12356 ( 
.A1(n_11750),
.A2(n_8825),
.B1(n_8799),
.B2(n_8560),
.C1(n_8906),
.C2(n_8926),
.Y(n_12356)
);

AOI22xp33_ASAP7_75t_L g12357 ( 
.A1(n_11819),
.A2(n_9806),
.B1(n_9810),
.B2(n_9801),
.Y(n_12357)
);

AOI221xp5_ASAP7_75t_L g12358 ( 
.A1(n_11563),
.A2(n_8188),
.B1(n_9029),
.B2(n_9122),
.C(n_9032),
.Y(n_12358)
);

AOI22xp33_ASAP7_75t_L g12359 ( 
.A1(n_11819),
.A2(n_9810),
.B1(n_9861),
.B2(n_9806),
.Y(n_12359)
);

INVx1_ASAP7_75t_L g12360 ( 
.A(n_11790),
.Y(n_12360)
);

AOI22xp33_ASAP7_75t_L g12361 ( 
.A1(n_11819),
.A2(n_9862),
.B1(n_9891),
.B2(n_9861),
.Y(n_12361)
);

AND2x2_ASAP7_75t_L g12362 ( 
.A(n_11672),
.B(n_10462),
.Y(n_12362)
);

AOI22xp5_ASAP7_75t_L g12363 ( 
.A1(n_11893),
.A2(n_10488),
.B1(n_10539),
.B2(n_10478),
.Y(n_12363)
);

AOI22xp33_ASAP7_75t_SL g12364 ( 
.A1(n_11446),
.A2(n_9855),
.B1(n_9848),
.B2(n_9171),
.Y(n_12364)
);

OAI22xp5_ASAP7_75t_L g12365 ( 
.A1(n_11037),
.A2(n_8970),
.B1(n_9248),
.B2(n_9442),
.Y(n_12365)
);

AOI222xp33_ASAP7_75t_L g12366 ( 
.A1(n_11750),
.A2(n_8560),
.B1(n_8906),
.B2(n_8926),
.C1(n_8155),
.C2(n_8719),
.Y(n_12366)
);

AND2x2_ASAP7_75t_L g12367 ( 
.A(n_11679),
.B(n_10478),
.Y(n_12367)
);

AOI22xp33_ASAP7_75t_L g12368 ( 
.A1(n_11847),
.A2(n_9861),
.B1(n_9891),
.B2(n_9862),
.Y(n_12368)
);

NOR2xp33_ASAP7_75t_L g12369 ( 
.A(n_10763),
.B(n_9632),
.Y(n_12369)
);

INVx1_ASAP7_75t_L g12370 ( 
.A(n_11919),
.Y(n_12370)
);

AOI33xp33_ASAP7_75t_L g12371 ( 
.A1(n_11508),
.A2(n_9039),
.A3(n_9111),
.B1(n_9144),
.B2(n_8990),
.B3(n_9133),
.Y(n_12371)
);

OAI22xp33_ASAP7_75t_L g12372 ( 
.A1(n_11664),
.A2(n_10488),
.B1(n_10539),
.B2(n_10478),
.Y(n_12372)
);

AOI22xp33_ASAP7_75t_L g12373 ( 
.A1(n_11847),
.A2(n_9862),
.B1(n_9920),
.B2(n_9891),
.Y(n_12373)
);

OAI22xp5_ASAP7_75t_L g12374 ( 
.A1(n_11063),
.A2(n_9442),
.B1(n_8922),
.B2(n_9294),
.Y(n_12374)
);

OAI211xp5_ASAP7_75t_L g12375 ( 
.A1(n_10957),
.A2(n_7980),
.B(n_8103),
.C(n_7928),
.Y(n_12375)
);

AOI22xp33_ASAP7_75t_L g12376 ( 
.A1(n_11847),
.A2(n_9920),
.B1(n_10005),
.B2(n_9957),
.Y(n_12376)
);

AND2x2_ASAP7_75t_L g12377 ( 
.A(n_11698),
.B(n_10478),
.Y(n_12377)
);

OAI22xp5_ASAP7_75t_L g12378 ( 
.A1(n_11063),
.A2(n_9442),
.B1(n_8922),
.B2(n_9283),
.Y(n_12378)
);

OAI211xp5_ASAP7_75t_L g12379 ( 
.A1(n_10957),
.A2(n_8125),
.B(n_8734),
.C(n_8151),
.Y(n_12379)
);

OAI22xp33_ASAP7_75t_L g12380 ( 
.A1(n_11664),
.A2(n_10539),
.B1(n_10624),
.B2(n_10488),
.Y(n_12380)
);

INVxp67_ASAP7_75t_L g12381 ( 
.A(n_11893),
.Y(n_12381)
);

OAI22xp5_ASAP7_75t_L g12382 ( 
.A1(n_11153),
.A2(n_11168),
.B1(n_11231),
.B2(n_11162),
.Y(n_12382)
);

AOI22xp33_ASAP7_75t_L g12383 ( 
.A1(n_11847),
.A2(n_9920),
.B1(n_10005),
.B2(n_9957),
.Y(n_12383)
);

OAI21x1_ASAP7_75t_L g12384 ( 
.A1(n_11141),
.A2(n_11680),
.B(n_11365),
.Y(n_12384)
);

INVx3_ASAP7_75t_L g12385 ( 
.A(n_11018),
.Y(n_12385)
);

AOI22xp33_ASAP7_75t_L g12386 ( 
.A1(n_11931),
.A2(n_9957),
.B1(n_10050),
.B2(n_10005),
.Y(n_12386)
);

NAND3xp33_ASAP7_75t_L g12387 ( 
.A(n_10978),
.B(n_8288),
.C(n_8151),
.Y(n_12387)
);

AOI22xp33_ASAP7_75t_SL g12388 ( 
.A1(n_11153),
.A2(n_9855),
.B1(n_9848),
.B2(n_9171),
.Y(n_12388)
);

OAI22xp5_ASAP7_75t_L g12389 ( 
.A1(n_11162),
.A2(n_9442),
.B1(n_8937),
.B2(n_9632),
.Y(n_12389)
);

AND2x2_ASAP7_75t_L g12390 ( 
.A(n_11711),
.B(n_10488),
.Y(n_12390)
);

OAI211xp5_ASAP7_75t_SL g12391 ( 
.A1(n_11621),
.A2(n_10640),
.B(n_10622),
.C(n_10398),
.Y(n_12391)
);

OA21x2_ASAP7_75t_L g12392 ( 
.A1(n_11282),
.A2(n_10509),
.B(n_10502),
.Y(n_12392)
);

OA21x2_ASAP7_75t_L g12393 ( 
.A1(n_11288),
.A2(n_10515),
.B(n_10509),
.Y(n_12393)
);

OAI221xp5_ASAP7_75t_L g12394 ( 
.A1(n_11168),
.A2(n_9556),
.B1(n_9353),
.B2(n_9664),
.C(n_10582),
.Y(n_12394)
);

OA21x2_ASAP7_75t_L g12395 ( 
.A1(n_11288),
.A2(n_10515),
.B(n_10509),
.Y(n_12395)
);

INVx2_ASAP7_75t_L g12396 ( 
.A(n_11314),
.Y(n_12396)
);

AND2x2_ASAP7_75t_L g12397 ( 
.A(n_10878),
.B(n_10488),
.Y(n_12397)
);

CKINVDCx5p33_ASAP7_75t_R g12398 ( 
.A(n_11868),
.Y(n_12398)
);

AOI22xp33_ASAP7_75t_L g12399 ( 
.A1(n_11931),
.A2(n_10050),
.B1(n_9171),
.B2(n_10539),
.Y(n_12399)
);

OAI22xp5_ASAP7_75t_L g12400 ( 
.A1(n_11231),
.A2(n_9442),
.B1(n_8937),
.B2(n_10539),
.Y(n_12400)
);

OAI22xp5_ASAP7_75t_L g12401 ( 
.A1(n_11239),
.A2(n_10539),
.B1(n_10681),
.B2(n_10624),
.Y(n_12401)
);

AND2x2_ASAP7_75t_L g12402 ( 
.A(n_10882),
.B(n_10624),
.Y(n_12402)
);

OAI22xp5_ASAP7_75t_L g12403 ( 
.A1(n_11239),
.A2(n_10624),
.B1(n_10681),
.B2(n_9311),
.Y(n_12403)
);

AOI22xp33_ASAP7_75t_L g12404 ( 
.A1(n_11931),
.A2(n_10050),
.B1(n_9171),
.B2(n_10624),
.Y(n_12404)
);

INVx3_ASAP7_75t_L g12405 ( 
.A(n_11018),
.Y(n_12405)
);

AND2x2_ASAP7_75t_L g12406 ( 
.A(n_10887),
.B(n_10624),
.Y(n_12406)
);

INVx4_ASAP7_75t_SL g12407 ( 
.A(n_10763),
.Y(n_12407)
);

NAND2xp5_ASAP7_75t_L g12408 ( 
.A(n_11508),
.B(n_11547),
.Y(n_12408)
);

INVx1_ASAP7_75t_L g12409 ( 
.A(n_10760),
.Y(n_12409)
);

HB1xp67_ASAP7_75t_L g12410 ( 
.A(n_11566),
.Y(n_12410)
);

AOI22xp33_ASAP7_75t_L g12411 ( 
.A1(n_11931),
.A2(n_10681),
.B1(n_9664),
.B2(n_9714),
.Y(n_12411)
);

OAI22xp5_ASAP7_75t_L g12412 ( 
.A1(n_11629),
.A2(n_10681),
.B1(n_9311),
.B2(n_10411),
.Y(n_12412)
);

INVx1_ASAP7_75t_L g12413 ( 
.A(n_10760),
.Y(n_12413)
);

BUFx6f_ASAP7_75t_L g12414 ( 
.A(n_11078),
.Y(n_12414)
);

INVxp67_ASAP7_75t_SL g12415 ( 
.A(n_11566),
.Y(n_12415)
);

INVx3_ASAP7_75t_L g12416 ( 
.A(n_11018),
.Y(n_12416)
);

AND2x4_ASAP7_75t_L g12417 ( 
.A(n_11547),
.B(n_9664),
.Y(n_12417)
);

OR2x2_ASAP7_75t_L g12418 ( 
.A(n_10906),
.B(n_10721),
.Y(n_12418)
);

INVx1_ASAP7_75t_L g12419 ( 
.A(n_10789),
.Y(n_12419)
);

INVx1_ASAP7_75t_L g12420 ( 
.A(n_10789),
.Y(n_12420)
);

OAI22xp5_ASAP7_75t_L g12421 ( 
.A1(n_11629),
.A2(n_10681),
.B1(n_10408),
.B2(n_10648),
.Y(n_12421)
);

AOI22xp33_ASAP7_75t_L g12422 ( 
.A1(n_11447),
.A2(n_10681),
.B1(n_9714),
.B2(n_10428),
.Y(n_12422)
);

BUFx3_ASAP7_75t_L g12423 ( 
.A(n_11805),
.Y(n_12423)
);

BUFx2_ASAP7_75t_L g12424 ( 
.A(n_11078),
.Y(n_12424)
);

AOI22xp33_ASAP7_75t_L g12425 ( 
.A1(n_11447),
.A2(n_9714),
.B1(n_10008),
.B2(n_9877),
.Y(n_12425)
);

BUFx6f_ASAP7_75t_L g12426 ( 
.A(n_11084),
.Y(n_12426)
);

OAI211xp5_ASAP7_75t_SL g12427 ( 
.A1(n_11621),
.A2(n_10398),
.B(n_10463),
.C(n_10459),
.Y(n_12427)
);

AND2x4_ASAP7_75t_L g12428 ( 
.A(n_11567),
.B(n_9714),
.Y(n_12428)
);

AOI22xp33_ASAP7_75t_L g12429 ( 
.A1(n_11464),
.A2(n_10008),
.B1(n_9877),
.B2(n_8288),
.Y(n_12429)
);

AOI22xp33_ASAP7_75t_L g12430 ( 
.A1(n_11464),
.A2(n_11484),
.B1(n_11582),
.B2(n_11466),
.Y(n_12430)
);

OAI22xp5_ASAP7_75t_L g12431 ( 
.A1(n_11773),
.A2(n_10661),
.B1(n_10671),
.B2(n_10632),
.Y(n_12431)
);

INVx1_ASAP7_75t_L g12432 ( 
.A(n_10790),
.Y(n_12432)
);

OAI22xp5_ASAP7_75t_L g12433 ( 
.A1(n_11773),
.A2(n_10695),
.B1(n_10707),
.B2(n_10677),
.Y(n_12433)
);

BUFx4f_ASAP7_75t_SL g12434 ( 
.A(n_11782),
.Y(n_12434)
);

AOI22xp33_ASAP7_75t_L g12435 ( 
.A1(n_11466),
.A2(n_10008),
.B1(n_9877),
.B2(n_8288),
.Y(n_12435)
);

AOI22xp33_ASAP7_75t_L g12436 ( 
.A1(n_11484),
.A2(n_10008),
.B1(n_9877),
.B2(n_8288),
.Y(n_12436)
);

OAI221xp5_ASAP7_75t_SL g12437 ( 
.A1(n_11686),
.A2(n_10008),
.B1(n_9877),
.B2(n_9243),
.C(n_9144),
.Y(n_12437)
);

AND2x4_ASAP7_75t_L g12438 ( 
.A(n_11567),
.B(n_9328),
.Y(n_12438)
);

AND2x4_ASAP7_75t_L g12439 ( 
.A(n_11586),
.B(n_9328),
.Y(n_12439)
);

INVx2_ASAP7_75t_L g12440 ( 
.A(n_11314),
.Y(n_12440)
);

BUFx3_ASAP7_75t_L g12441 ( 
.A(n_11805),
.Y(n_12441)
);

AOI22xp33_ASAP7_75t_L g12442 ( 
.A1(n_11582),
.A2(n_8288),
.B1(n_9556),
.B2(n_9285),
.Y(n_12442)
);

BUFx2_ASAP7_75t_R g12443 ( 
.A(n_11019),
.Y(n_12443)
);

AOI22xp33_ASAP7_75t_SL g12444 ( 
.A1(n_11853),
.A2(n_7940),
.B1(n_7943),
.B2(n_8188),
.Y(n_12444)
);

OAI22xp5_ASAP7_75t_L g12445 ( 
.A1(n_11322),
.A2(n_9243),
.B1(n_8990),
.B2(n_9418),
.Y(n_12445)
);

INVx2_ASAP7_75t_L g12446 ( 
.A(n_11350),
.Y(n_12446)
);

INVx1_ASAP7_75t_L g12447 ( 
.A(n_10790),
.Y(n_12447)
);

BUFx2_ASAP7_75t_L g12448 ( 
.A(n_11084),
.Y(n_12448)
);

AND2x2_ASAP7_75t_L g12449 ( 
.A(n_10896),
.B(n_9580),
.Y(n_12449)
);

AOI221xp5_ASAP7_75t_L g12450 ( 
.A1(n_10802),
.A2(n_8188),
.B1(n_9032),
.B2(n_8185),
.C(n_9256),
.Y(n_12450)
);

AOI22xp5_ASAP7_75t_L g12451 ( 
.A1(n_11586),
.A2(n_9285),
.B1(n_9256),
.B2(n_9208),
.Y(n_12451)
);

INVx1_ASAP7_75t_L g12452 ( 
.A(n_10802),
.Y(n_12452)
);

INVx1_ASAP7_75t_L g12453 ( 
.A(n_10811),
.Y(n_12453)
);

OR2x2_ASAP7_75t_L g12454 ( 
.A(n_10767),
.B(n_10583),
.Y(n_12454)
);

AOI222xp33_ASAP7_75t_L g12455 ( 
.A1(n_11647),
.A2(n_8719),
.B1(n_8938),
.B2(n_8974),
.C1(n_9101),
.C2(n_9004),
.Y(n_12455)
);

AND2x2_ASAP7_75t_L g12456 ( 
.A(n_11402),
.B(n_9580),
.Y(n_12456)
);

AND2x2_ASAP7_75t_L g12457 ( 
.A(n_11431),
.B(n_9580),
.Y(n_12457)
);

OA21x2_ASAP7_75t_L g12458 ( 
.A1(n_10776),
.A2(n_10529),
.B(n_10515),
.Y(n_12458)
);

OAI221xp5_ASAP7_75t_L g12459 ( 
.A1(n_11329),
.A2(n_9512),
.B1(n_9534),
.B2(n_9490),
.C(n_9439),
.Y(n_12459)
);

AND2x4_ASAP7_75t_L g12460 ( 
.A(n_11621),
.B(n_9418),
.Y(n_12460)
);

AO21x2_ASAP7_75t_L g12461 ( 
.A1(n_11580),
.A2(n_10532),
.B(n_10529),
.Y(n_12461)
);

AOI221xp5_ASAP7_75t_L g12462 ( 
.A1(n_10811),
.A2(n_8188),
.B1(n_8185),
.B2(n_8250),
.C(n_9101),
.Y(n_12462)
);

AOI22xp33_ASAP7_75t_L g12463 ( 
.A1(n_11615),
.A2(n_8333),
.B1(n_8327),
.B2(n_10102),
.Y(n_12463)
);

AOI221xp5_ASAP7_75t_L g12464 ( 
.A1(n_10815),
.A2(n_8185),
.B1(n_8250),
.B2(n_8923),
.C(n_9004),
.Y(n_12464)
);

OAI22xp33_ASAP7_75t_L g12465 ( 
.A1(n_11686),
.A2(n_9204),
.B1(n_8266),
.B2(n_8182),
.Y(n_12465)
);

OAI221xp5_ASAP7_75t_L g12466 ( 
.A1(n_11329),
.A2(n_9512),
.B1(n_9534),
.B2(n_9490),
.C(n_9439),
.Y(n_12466)
);

AOI22xp33_ASAP7_75t_L g12467 ( 
.A1(n_11615),
.A2(n_8333),
.B1(n_8327),
.B2(n_10102),
.Y(n_12467)
);

INVx2_ASAP7_75t_L g12468 ( 
.A(n_11350),
.Y(n_12468)
);

AOI22xp33_ASAP7_75t_L g12469 ( 
.A1(n_10961),
.A2(n_8327),
.B1(n_10108),
.B2(n_10102),
.Y(n_12469)
);

HB1xp67_ASAP7_75t_L g12470 ( 
.A(n_10815),
.Y(n_12470)
);

NOR2xp67_ASAP7_75t_L g12471 ( 
.A(n_10734),
.B(n_9580),
.Y(n_12471)
);

HB1xp67_ASAP7_75t_L g12472 ( 
.A(n_10841),
.Y(n_12472)
);

INVx1_ASAP7_75t_L g12473 ( 
.A(n_10841),
.Y(n_12473)
);

OAI22xp33_ASAP7_75t_L g12474 ( 
.A1(n_11686),
.A2(n_9204),
.B1(n_8266),
.B2(n_8182),
.Y(n_12474)
);

INVx1_ASAP7_75t_L g12475 ( 
.A(n_10843),
.Y(n_12475)
);

BUFx6f_ASAP7_75t_L g12476 ( 
.A(n_11138),
.Y(n_12476)
);

OAI21xp33_ASAP7_75t_L g12477 ( 
.A1(n_11381),
.A2(n_9117),
.B(n_9192),
.Y(n_12477)
);

HB1xp67_ASAP7_75t_L g12478 ( 
.A(n_10843),
.Y(n_12478)
);

AND2x2_ASAP7_75t_L g12479 ( 
.A(n_11443),
.B(n_9620),
.Y(n_12479)
);

AOI22xp33_ASAP7_75t_L g12480 ( 
.A1(n_10961),
.A2(n_10108),
.B1(n_10111),
.B2(n_10102),
.Y(n_12480)
);

NAND3xp33_ASAP7_75t_L g12481 ( 
.A(n_10978),
.B(n_8151),
.C(n_8125),
.Y(n_12481)
);

AOI22xp33_ASAP7_75t_SL g12482 ( 
.A1(n_11647),
.A2(n_7940),
.B1(n_7943),
.B2(n_8125),
.Y(n_12482)
);

INVx2_ASAP7_75t_L g12483 ( 
.A(n_11350),
.Y(n_12483)
);

HB1xp67_ASAP7_75t_L g12484 ( 
.A(n_10844),
.Y(n_12484)
);

OAI21xp5_ASAP7_75t_L g12485 ( 
.A1(n_11838),
.A2(n_8259),
.B(n_8170),
.Y(n_12485)
);

NAND2xp5_ASAP7_75t_L g12486 ( 
.A(n_11403),
.B(n_9042),
.Y(n_12486)
);

OAI211xp5_ASAP7_75t_L g12487 ( 
.A1(n_10978),
.A2(n_8125),
.B(n_8734),
.C(n_8151),
.Y(n_12487)
);

AND2x2_ASAP7_75t_L g12488 ( 
.A(n_11480),
.B(n_9620),
.Y(n_12488)
);

AND2x2_ASAP7_75t_L g12489 ( 
.A(n_11501),
.B(n_9620),
.Y(n_12489)
);

OAI211xp5_ASAP7_75t_L g12490 ( 
.A1(n_11122),
.A2(n_8125),
.B(n_8734),
.C(n_8151),
.Y(n_12490)
);

OAI22xp5_ASAP7_75t_SL g12491 ( 
.A1(n_11278),
.A2(n_10321),
.B1(n_9554),
.B2(n_9608),
.Y(n_12491)
);

INVx1_ASAP7_75t_L g12492 ( 
.A(n_10844),
.Y(n_12492)
);

INVx1_ASAP7_75t_L g12493 ( 
.A(n_10848),
.Y(n_12493)
);

INVx1_ASAP7_75t_L g12494 ( 
.A(n_10848),
.Y(n_12494)
);

AND2x2_ASAP7_75t_L g12495 ( 
.A(n_11528),
.B(n_9620),
.Y(n_12495)
);

AOI21xp5_ASAP7_75t_L g12496 ( 
.A1(n_11278),
.A2(n_10013),
.B(n_9820),
.Y(n_12496)
);

NOR2xp33_ASAP7_75t_L g12497 ( 
.A(n_11138),
.B(n_10034),
.Y(n_12497)
);

NAND2xp5_ASAP7_75t_L g12498 ( 
.A(n_11408),
.B(n_9042),
.Y(n_12498)
);

AOI22xp33_ASAP7_75t_L g12499 ( 
.A1(n_10961),
.A2(n_10111),
.B1(n_10129),
.B2(n_10108),
.Y(n_12499)
);

BUFx4f_ASAP7_75t_SL g12500 ( 
.A(n_11810),
.Y(n_12500)
);

AO31x2_ASAP7_75t_L g12501 ( 
.A1(n_11329),
.A2(n_10532),
.A3(n_10533),
.B(n_10529),
.Y(n_12501)
);

INVx1_ASAP7_75t_L g12502 ( 
.A(n_10885),
.Y(n_12502)
);

AOI21xp33_ASAP7_75t_L g12503 ( 
.A1(n_11643),
.A2(n_8518),
.B(n_8250),
.Y(n_12503)
);

A2O1A1Ixp33_ASAP7_75t_L g12504 ( 
.A1(n_11248),
.A2(n_8259),
.B(n_9235),
.C(n_8675),
.Y(n_12504)
);

AOI22xp33_ASAP7_75t_L g12505 ( 
.A1(n_10961),
.A2(n_10111),
.B1(n_10129),
.B2(n_10108),
.Y(n_12505)
);

AND2x2_ASAP7_75t_L g12506 ( 
.A(n_11560),
.B(n_9629),
.Y(n_12506)
);

AND2x2_ASAP7_75t_L g12507 ( 
.A(n_11562),
.B(n_9629),
.Y(n_12507)
);

AOI22xp33_ASAP7_75t_L g12508 ( 
.A1(n_11011),
.A2(n_10129),
.B1(n_10226),
.B2(n_10111),
.Y(n_12508)
);

AOI221xp5_ASAP7_75t_L g12509 ( 
.A1(n_10885),
.A2(n_10942),
.B1(n_10990),
.B2(n_10985),
.C(n_10892),
.Y(n_12509)
);

INVx2_ASAP7_75t_L g12510 ( 
.A(n_11392),
.Y(n_12510)
);

AOI22xp33_ASAP7_75t_L g12511 ( 
.A1(n_11011),
.A2(n_10226),
.B1(n_10236),
.B2(n_10129),
.Y(n_12511)
);

AOI21xp5_ASAP7_75t_L g12512 ( 
.A1(n_11413),
.A2(n_10013),
.B(n_9820),
.Y(n_12512)
);

AOI22xp33_ASAP7_75t_L g12513 ( 
.A1(n_11011),
.A2(n_10236),
.B1(n_10257),
.B2(n_10226),
.Y(n_12513)
);

INVx1_ASAP7_75t_L g12514 ( 
.A(n_10892),
.Y(n_12514)
);

NAND3xp33_ASAP7_75t_L g12515 ( 
.A(n_11122),
.B(n_8151),
.C(n_8125),
.Y(n_12515)
);

OAI222xp33_ASAP7_75t_L g12516 ( 
.A1(n_11838),
.A2(n_8266),
.B1(n_8675),
.B2(n_9512),
.C1(n_9490),
.C2(n_9439),
.Y(n_12516)
);

AND2x4_ASAP7_75t_L g12517 ( 
.A(n_11875),
.B(n_9426),
.Y(n_12517)
);

OR2x2_ASAP7_75t_L g12518 ( 
.A(n_10775),
.B(n_10785),
.Y(n_12518)
);

AOI22xp5_ASAP7_75t_L g12519 ( 
.A1(n_11413),
.A2(n_9208),
.B1(n_8589),
.B2(n_9426),
.Y(n_12519)
);

AOI22xp33_ASAP7_75t_L g12520 ( 
.A1(n_11011),
.A2(n_11119),
.B1(n_11270),
.B2(n_11058),
.Y(n_12520)
);

AOI22xp33_ASAP7_75t_L g12521 ( 
.A1(n_11058),
.A2(n_10236),
.B1(n_10257),
.B2(n_10226),
.Y(n_12521)
);

OAI22xp5_ASAP7_75t_L g12522 ( 
.A1(n_11410),
.A2(n_9510),
.B1(n_9615),
.B2(n_9576),
.Y(n_12522)
);

NAND2xp5_ASAP7_75t_L g12523 ( 
.A(n_11459),
.B(n_9119),
.Y(n_12523)
);

OAI21xp5_ASAP7_75t_L g12524 ( 
.A1(n_10989),
.A2(n_8170),
.B(n_8357),
.Y(n_12524)
);

NAND2xp5_ASAP7_75t_L g12525 ( 
.A(n_11600),
.B(n_9119),
.Y(n_12525)
);

OAI21xp33_ASAP7_75t_L g12526 ( 
.A1(n_10935),
.A2(n_9117),
.B(n_9192),
.Y(n_12526)
);

AOI22xp5_ASAP7_75t_L g12527 ( 
.A1(n_11058),
.A2(n_11119),
.B1(n_11319),
.B2(n_11270),
.Y(n_12527)
);

AOI22xp33_ASAP7_75t_L g12528 ( 
.A1(n_11058),
.A2(n_10257),
.B1(n_10236),
.B2(n_9146),
.Y(n_12528)
);

OAI22xp5_ASAP7_75t_L g12529 ( 
.A1(n_11658),
.A2(n_9510),
.B1(n_9615),
.B2(n_9576),
.Y(n_12529)
);

INVxp67_ASAP7_75t_L g12530 ( 
.A(n_11768),
.Y(n_12530)
);

OAI22xp5_ASAP7_75t_L g12531 ( 
.A1(n_11658),
.A2(n_9641),
.B1(n_9650),
.B2(n_9645),
.Y(n_12531)
);

AOI22xp33_ASAP7_75t_L g12532 ( 
.A1(n_11119),
.A2(n_10257),
.B1(n_9146),
.B2(n_10013),
.Y(n_12532)
);

AOI22xp33_ASAP7_75t_L g12533 ( 
.A1(n_11119),
.A2(n_9146),
.B1(n_10013),
.B2(n_9820),
.Y(n_12533)
);

OAI33xp33_ASAP7_75t_L g12534 ( 
.A1(n_10730),
.A2(n_10749),
.A3(n_10737),
.B1(n_10750),
.B2(n_10741),
.B3(n_10733),
.Y(n_12534)
);

AOI22xp5_ASAP7_75t_SL g12535 ( 
.A1(n_11552),
.A2(n_9437),
.B1(n_10290),
.B2(n_10253),
.Y(n_12535)
);

AOI22xp5_ASAP7_75t_L g12536 ( 
.A1(n_11270),
.A2(n_8589),
.B1(n_9645),
.B2(n_9641),
.Y(n_12536)
);

AOI22xp33_ASAP7_75t_L g12537 ( 
.A1(n_11270),
.A2(n_10013),
.B1(n_10424),
.B2(n_9820),
.Y(n_12537)
);

AOI22xp33_ASAP7_75t_L g12538 ( 
.A1(n_11319),
.A2(n_11437),
.B1(n_11265),
.B2(n_11248),
.Y(n_12538)
);

BUFx4f_ASAP7_75t_SL g12539 ( 
.A(n_11810),
.Y(n_12539)
);

OA21x2_ASAP7_75t_L g12540 ( 
.A1(n_10776),
.A2(n_10533),
.B(n_10532),
.Y(n_12540)
);

INVx1_ASAP7_75t_L g12541 ( 
.A(n_10942),
.Y(n_12541)
);

AOI21xp5_ASAP7_75t_L g12542 ( 
.A1(n_11233),
.A2(n_10424),
.B(n_9820),
.Y(n_12542)
);

AND2x2_ASAP7_75t_L g12543 ( 
.A(n_11584),
.B(n_9629),
.Y(n_12543)
);

AOI22xp33_ASAP7_75t_L g12544 ( 
.A1(n_11319),
.A2(n_11437),
.B1(n_11265),
.B2(n_11552),
.Y(n_12544)
);

AOI22xp33_ASAP7_75t_L g12545 ( 
.A1(n_11319),
.A2(n_10424),
.B1(n_9650),
.B2(n_9704),
.Y(n_12545)
);

OAI22xp5_ASAP7_75t_L g12546 ( 
.A1(n_11681),
.A2(n_9674),
.B1(n_9721),
.B2(n_9704),
.Y(n_12546)
);

INVx2_ASAP7_75t_SL g12547 ( 
.A(n_11393),
.Y(n_12547)
);

AOI211xp5_ASAP7_75t_L g12548 ( 
.A1(n_11437),
.A2(n_8170),
.B(n_8163),
.C(n_7994),
.Y(n_12548)
);

AOI221xp5_ASAP7_75t_L g12549 ( 
.A1(n_10985),
.A2(n_8185),
.B1(n_8250),
.B2(n_8826),
.C(n_8938),
.Y(n_12549)
);

INVx1_ASAP7_75t_L g12550 ( 
.A(n_10990),
.Y(n_12550)
);

OAI21x1_ASAP7_75t_L g12551 ( 
.A1(n_11680),
.A2(n_10204),
.B(n_10165),
.Y(n_12551)
);

INVx1_ASAP7_75t_L g12552 ( 
.A(n_11035),
.Y(n_12552)
);

HB1xp67_ASAP7_75t_L g12553 ( 
.A(n_11035),
.Y(n_12553)
);

AOI221xp5_ASAP7_75t_L g12554 ( 
.A1(n_11049),
.A2(n_8185),
.B1(n_8250),
.B2(n_8974),
.C(n_8518),
.Y(n_12554)
);

AND2x2_ASAP7_75t_L g12555 ( 
.A(n_11601),
.B(n_9629),
.Y(n_12555)
);

NAND2xp5_ASAP7_75t_L g12556 ( 
.A(n_11604),
.B(n_9094),
.Y(n_12556)
);

OAI22xp5_ASAP7_75t_L g12557 ( 
.A1(n_11681),
.A2(n_9674),
.B1(n_9746),
.B2(n_9721),
.Y(n_12557)
);

AOI21xp5_ASAP7_75t_L g12558 ( 
.A1(n_11233),
.A2(n_10424),
.B(n_8997),
.Y(n_12558)
);

OAI222xp33_ASAP7_75t_L g12559 ( 
.A1(n_11875),
.A2(n_9534),
.B1(n_9621),
.B2(n_9550),
.C1(n_8182),
.C2(n_8212),
.Y(n_12559)
);

NAND2xp5_ASAP7_75t_L g12560 ( 
.A(n_11437),
.B(n_9094),
.Y(n_12560)
);

NAND2xp5_ASAP7_75t_L g12561 ( 
.A(n_11888),
.B(n_9279),
.Y(n_12561)
);

INVx1_ASAP7_75t_L g12562 ( 
.A(n_11049),
.Y(n_12562)
);

OR2x2_ASAP7_75t_L g12563 ( 
.A(n_10786),
.B(n_10372),
.Y(n_12563)
);

INVx2_ASAP7_75t_L g12564 ( 
.A(n_11392),
.Y(n_12564)
);

OAI31xp33_ASAP7_75t_SL g12565 ( 
.A1(n_10981),
.A2(n_10306),
.A3(n_8845),
.B(n_8090),
.Y(n_12565)
);

AOI22xp33_ASAP7_75t_L g12566 ( 
.A1(n_11552),
.A2(n_10424),
.B1(n_9746),
.B2(n_8734),
.Y(n_12566)
);

AOI22xp33_ASAP7_75t_L g12567 ( 
.A1(n_11552),
.A2(n_8734),
.B1(n_9722),
.B2(n_9665),
.Y(n_12567)
);

INVx2_ASAP7_75t_L g12568 ( 
.A(n_11392),
.Y(n_12568)
);

OAI221xp5_ASAP7_75t_SL g12569 ( 
.A1(n_10981),
.A2(n_8997),
.B1(n_9281),
.B2(n_8212),
.C(n_8030),
.Y(n_12569)
);

OAI21x1_ASAP7_75t_L g12570 ( 
.A1(n_11351),
.A2(n_10459),
.B(n_10398),
.Y(n_12570)
);

AOI22xp33_ASAP7_75t_L g12571 ( 
.A1(n_11552),
.A2(n_8734),
.B1(n_9722),
.B2(n_9665),
.Y(n_12571)
);

INVx1_ASAP7_75t_L g12572 ( 
.A(n_11102),
.Y(n_12572)
);

AOI21xp5_ASAP7_75t_SL g12573 ( 
.A1(n_10770),
.A2(n_8778),
.B(n_7590),
.Y(n_12573)
);

OAI211xp5_ASAP7_75t_L g12574 ( 
.A1(n_11122),
.A2(n_9183),
.B(n_10697),
.C(n_10566),
.Y(n_12574)
);

AOI21xp5_ASAP7_75t_L g12575 ( 
.A1(n_11269),
.A2(n_8849),
.B(n_8784),
.Y(n_12575)
);

INVx2_ASAP7_75t_L g12576 ( 
.A(n_11419),
.Y(n_12576)
);

AOI22xp33_ASAP7_75t_L g12577 ( 
.A1(n_11802),
.A2(n_9665),
.B1(n_9734),
.B2(n_9722),
.Y(n_12577)
);

OAI211xp5_ASAP7_75t_L g12578 ( 
.A1(n_11181),
.A2(n_9183),
.B(n_10697),
.C(n_10566),
.Y(n_12578)
);

INVx1_ASAP7_75t_L g12579 ( 
.A(n_11102),
.Y(n_12579)
);

AND2x2_ASAP7_75t_L g12580 ( 
.A(n_10738),
.B(n_10807),
.Y(n_12580)
);

AOI21xp5_ASAP7_75t_SL g12581 ( 
.A1(n_10770),
.A2(n_7650),
.B(n_7567),
.Y(n_12581)
);

INVx1_ASAP7_75t_L g12582 ( 
.A(n_11131),
.Y(n_12582)
);

AOI222xp33_ASAP7_75t_L g12583 ( 
.A1(n_11712),
.A2(n_8272),
.B1(n_8632),
.B2(n_8071),
.C1(n_8098),
.C2(n_8101),
.Y(n_12583)
);

OAI22xp5_ASAP7_75t_SL g12584 ( 
.A1(n_11802),
.A2(n_6730),
.B1(n_6677),
.B2(n_7658),
.Y(n_12584)
);

AOI22xp33_ASAP7_75t_L g12585 ( 
.A1(n_11802),
.A2(n_11835),
.B1(n_11719),
.B2(n_11722),
.Y(n_12585)
);

OAI21xp33_ASAP7_75t_L g12586 ( 
.A1(n_11670),
.A2(n_7994),
.B(n_9281),
.Y(n_12586)
);

NAND2xp5_ASAP7_75t_L g12587 ( 
.A(n_11876),
.B(n_9279),
.Y(n_12587)
);

AOI22xp33_ASAP7_75t_L g12588 ( 
.A1(n_11835),
.A2(n_9665),
.B1(n_9734),
.B2(n_9722),
.Y(n_12588)
);

AOI22xp33_ASAP7_75t_L g12589 ( 
.A1(n_11835),
.A2(n_9734),
.B1(n_9767),
.B2(n_9754),
.Y(n_12589)
);

NAND2x1_ASAP7_75t_L g12590 ( 
.A(n_11238),
.B(n_9734),
.Y(n_12590)
);

BUFx2_ASAP7_75t_L g12591 ( 
.A(n_11712),
.Y(n_12591)
);

AOI221xp5_ASAP7_75t_L g12592 ( 
.A1(n_11131),
.A2(n_8518),
.B1(n_8497),
.B2(n_8489),
.C(n_8488),
.Y(n_12592)
);

AOI222xp33_ASAP7_75t_L g12593 ( 
.A1(n_11719),
.A2(n_8272),
.B1(n_8632),
.B2(n_8071),
.C1(n_8090),
.C2(n_8101),
.Y(n_12593)
);

NOR2x1_ASAP7_75t_SL g12594 ( 
.A(n_11364),
.B(n_8030),
.Y(n_12594)
);

AOI22xp33_ASAP7_75t_SL g12595 ( 
.A1(n_11722),
.A2(n_7940),
.B1(n_7943),
.B2(n_9183),
.Y(n_12595)
);

INVx1_ASAP7_75t_L g12596 ( 
.A(n_11145),
.Y(n_12596)
);

INVx1_ASAP7_75t_L g12597 ( 
.A(n_11145),
.Y(n_12597)
);

AOI22xp33_ASAP7_75t_L g12598 ( 
.A1(n_11735),
.A2(n_9754),
.B1(n_9785),
.B2(n_9767),
.Y(n_12598)
);

AOI22xp33_ASAP7_75t_SL g12599 ( 
.A1(n_11735),
.A2(n_7940),
.B1(n_7943),
.B2(n_9183),
.Y(n_12599)
);

AOI22xp5_ASAP7_75t_L g12600 ( 
.A1(n_10758),
.A2(n_7003),
.B1(n_7040),
.B2(n_6999),
.Y(n_12600)
);

AO21x2_ASAP7_75t_L g12601 ( 
.A1(n_11580),
.A2(n_10534),
.B(n_10533),
.Y(n_12601)
);

INVx2_ASAP7_75t_L g12602 ( 
.A(n_11419),
.Y(n_12602)
);

OA21x2_ASAP7_75t_L g12603 ( 
.A1(n_11351),
.A2(n_10541),
.B(n_10534),
.Y(n_12603)
);

INVx1_ASAP7_75t_L g12604 ( 
.A(n_11152),
.Y(n_12604)
);

AOI22xp33_ASAP7_75t_L g12605 ( 
.A1(n_10833),
.A2(n_9754),
.B1(n_9785),
.B2(n_9767),
.Y(n_12605)
);

BUFx6f_ASAP7_75t_L g12606 ( 
.A(n_11393),
.Y(n_12606)
);

INVx2_ASAP7_75t_L g12607 ( 
.A(n_11419),
.Y(n_12607)
);

AOI222xp33_ASAP7_75t_L g12608 ( 
.A1(n_11152),
.A2(n_8272),
.B1(n_8071),
.B2(n_8090),
.C1(n_8101),
.C2(n_8099),
.Y(n_12608)
);

OAI21x1_ASAP7_75t_L g12609 ( 
.A1(n_11365),
.A2(n_10459),
.B(n_10398),
.Y(n_12609)
);

OAI22xp5_ASAP7_75t_L g12610 ( 
.A1(n_11643),
.A2(n_8693),
.B1(n_9767),
.B2(n_9754),
.Y(n_12610)
);

AND2x2_ASAP7_75t_L g12611 ( 
.A(n_10822),
.B(n_9785),
.Y(n_12611)
);

INVx1_ASAP7_75t_L g12612 ( 
.A(n_11181),
.Y(n_12612)
);

NAND2xp5_ASAP7_75t_L g12613 ( 
.A(n_11876),
.B(n_11888),
.Y(n_12613)
);

CKINVDCx20_ASAP7_75t_R g12614 ( 
.A(n_11724),
.Y(n_12614)
);

AND2x4_ASAP7_75t_SL g12615 ( 
.A(n_10770),
.B(n_7734),
.Y(n_12615)
);

AOI22xp33_ASAP7_75t_L g12616 ( 
.A1(n_10951),
.A2(n_9785),
.B1(n_10016),
.B2(n_9971),
.Y(n_12616)
);

AOI221xp5_ASAP7_75t_L g12617 ( 
.A1(n_11204),
.A2(n_8497),
.B1(n_8489),
.B2(n_8488),
.C(n_9264),
.Y(n_12617)
);

AND2x2_ASAP7_75t_L g12618 ( 
.A(n_10837),
.B(n_9971),
.Y(n_12618)
);

OAI21xp5_ASAP7_75t_L g12619 ( 
.A1(n_10989),
.A2(n_10849),
.B(n_10754),
.Y(n_12619)
);

INVx1_ASAP7_75t_L g12620 ( 
.A(n_11204),
.Y(n_12620)
);

OAI221xp5_ASAP7_75t_SL g12621 ( 
.A1(n_11236),
.A2(n_8212),
.B1(n_8030),
.B2(n_9264),
.C(n_8784),
.Y(n_12621)
);

INVx2_ASAP7_75t_L g12622 ( 
.A(n_11445),
.Y(n_12622)
);

AOI22xp33_ASAP7_75t_L g12623 ( 
.A1(n_11177),
.A2(n_9971),
.B1(n_10075),
.B2(n_10016),
.Y(n_12623)
);

AOI22xp33_ASAP7_75t_L g12624 ( 
.A1(n_11177),
.A2(n_11208),
.B1(n_11326),
.B2(n_11217),
.Y(n_12624)
);

OAI22xp5_ASAP7_75t_L g12625 ( 
.A1(n_11648),
.A2(n_8693),
.B1(n_10016),
.B2(n_9971),
.Y(n_12625)
);

AOI22xp33_ASAP7_75t_L g12626 ( 
.A1(n_11177),
.A2(n_10016),
.B1(n_10082),
.B2(n_10075),
.Y(n_12626)
);

AOI221xp5_ASAP7_75t_L g12627 ( 
.A1(n_11236),
.A2(n_8497),
.B1(n_8489),
.B2(n_8488),
.C(n_9323),
.Y(n_12627)
);

OR2x2_ASAP7_75t_L g12628 ( 
.A(n_10797),
.B(n_10378),
.Y(n_12628)
);

AND2x2_ASAP7_75t_L g12629 ( 
.A(n_11217),
.B(n_11326),
.Y(n_12629)
);

CKINVDCx5p33_ASAP7_75t_R g12630 ( 
.A(n_11724),
.Y(n_12630)
);

AOI22xp33_ASAP7_75t_L g12631 ( 
.A1(n_11208),
.A2(n_10075),
.B1(n_10123),
.B2(n_10082),
.Y(n_12631)
);

NAND2xp5_ASAP7_75t_L g12632 ( 
.A(n_11287),
.B(n_9310),
.Y(n_12632)
);

OAI22xp33_ASAP7_75t_L g12633 ( 
.A1(n_11648),
.A2(n_8849),
.B1(n_10082),
.B2(n_10075),
.Y(n_12633)
);

AND2x4_ASAP7_75t_L g12634 ( 
.A(n_11470),
.B(n_9929),
.Y(n_12634)
);

INVx1_ASAP7_75t_SL g12635 ( 
.A(n_11531),
.Y(n_12635)
);

AOI22xp33_ASAP7_75t_L g12636 ( 
.A1(n_11208),
.A2(n_11326),
.B1(n_11398),
.B2(n_11217),
.Y(n_12636)
);

INVx1_ASAP7_75t_L g12637 ( 
.A(n_11287),
.Y(n_12637)
);

INVx2_ASAP7_75t_L g12638 ( 
.A(n_11445),
.Y(n_12638)
);

CKINVDCx5p33_ASAP7_75t_R g12639 ( 
.A(n_11531),
.Y(n_12639)
);

OAI22xp5_ASAP7_75t_L g12640 ( 
.A1(n_11684),
.A2(n_8693),
.B1(n_10123),
.B2(n_10082),
.Y(n_12640)
);

NAND2xp5_ASAP7_75t_L g12641 ( 
.A(n_11315),
.B(n_9310),
.Y(n_12641)
);

NAND2xp5_ASAP7_75t_L g12642 ( 
.A(n_11315),
.B(n_8724),
.Y(n_12642)
);

A2O1A1Ixp33_ASAP7_75t_SL g12643 ( 
.A1(n_10734),
.A2(n_10459),
.B(n_10517),
.C(n_10463),
.Y(n_12643)
);

AND2x2_ASAP7_75t_L g12644 ( 
.A(n_11398),
.B(n_10123),
.Y(n_12644)
);

AND2x4_ASAP7_75t_L g12645 ( 
.A(n_11470),
.B(n_9929),
.Y(n_12645)
);

AOI21xp5_ASAP7_75t_L g12646 ( 
.A1(n_11269),
.A2(n_11593),
.B(n_11663),
.Y(n_12646)
);

AOI221xp5_ASAP7_75t_L g12647 ( 
.A1(n_11317),
.A2(n_8497),
.B1(n_8489),
.B2(n_8488),
.C(n_9323),
.Y(n_12647)
);

BUFx3_ASAP7_75t_L g12648 ( 
.A(n_11398),
.Y(n_12648)
);

AOI21xp5_ASAP7_75t_L g12649 ( 
.A1(n_11593),
.A2(n_8849),
.B(n_8680),
.Y(n_12649)
);

BUFx3_ASAP7_75t_L g12650 ( 
.A(n_11400),
.Y(n_12650)
);

AND2x2_ASAP7_75t_L g12651 ( 
.A(n_11400),
.B(n_10123),
.Y(n_12651)
);

CKINVDCx5p33_ASAP7_75t_R g12652 ( 
.A(n_11470),
.Y(n_12652)
);

OAI22xp5_ASAP7_75t_SL g12653 ( 
.A1(n_11684),
.A2(n_7669),
.B1(n_7721),
.B2(n_7658),
.Y(n_12653)
);

AOI22xp33_ASAP7_75t_L g12654 ( 
.A1(n_11400),
.A2(n_10182),
.B1(n_10264),
.B2(n_10221),
.Y(n_12654)
);

HB1xp67_ASAP7_75t_L g12655 ( 
.A(n_11317),
.Y(n_12655)
);

AOI221xp5_ASAP7_75t_L g12656 ( 
.A1(n_11341),
.A2(n_8497),
.B1(n_8489),
.B2(n_8488),
.C(n_9323),
.Y(n_12656)
);

OAI22xp5_ASAP7_75t_L g12657 ( 
.A1(n_11721),
.A2(n_8693),
.B1(n_10221),
.B2(n_10182),
.Y(n_12657)
);

OAI321xp33_ASAP7_75t_L g12658 ( 
.A1(n_11765),
.A2(n_9550),
.A3(n_9621),
.B1(n_10064),
.B2(n_10093),
.C(n_8332),
.Y(n_12658)
);

OAI22xp33_ASAP7_75t_L g12659 ( 
.A1(n_11721),
.A2(n_10221),
.B1(n_10264),
.B2(n_10182),
.Y(n_12659)
);

AOI22xp5_ASAP7_75t_L g12660 ( 
.A1(n_11479),
.A2(n_7003),
.B1(n_7040),
.B2(n_6999),
.Y(n_12660)
);

OR2x2_ASAP7_75t_L g12661 ( 
.A(n_10813),
.B(n_10394),
.Y(n_12661)
);

AOI22xp33_ASAP7_75t_L g12662 ( 
.A1(n_11479),
.A2(n_10182),
.B1(n_10264),
.B2(n_10221),
.Y(n_12662)
);

AND2x2_ASAP7_75t_L g12663 ( 
.A(n_11479),
.B(n_10264),
.Y(n_12663)
);

INVx3_ASAP7_75t_L g12664 ( 
.A(n_11158),
.Y(n_12664)
);

INVx1_ASAP7_75t_L g12665 ( 
.A(n_11341),
.Y(n_12665)
);

NAND2xp5_ASAP7_75t_L g12666 ( 
.A(n_11377),
.B(n_8724),
.Y(n_12666)
);

INVx1_ASAP7_75t_SL g12667 ( 
.A(n_11523),
.Y(n_12667)
);

INVx3_ASAP7_75t_L g12668 ( 
.A(n_11158),
.Y(n_12668)
);

NAND3xp33_ASAP7_75t_L g12669 ( 
.A(n_11377),
.B(n_8408),
.C(n_8358),
.Y(n_12669)
);

AOI22xp33_ASAP7_75t_L g12670 ( 
.A1(n_11523),
.A2(n_10289),
.B1(n_9183),
.B2(n_7948),
.Y(n_12670)
);

AOI22xp33_ASAP7_75t_L g12671 ( 
.A1(n_11523),
.A2(n_10289),
.B1(n_9183),
.B2(n_7948),
.Y(n_12671)
);

INVx1_ASAP7_75t_L g12672 ( 
.A(n_11406),
.Y(n_12672)
);

AND2x2_ASAP7_75t_L g12673 ( 
.A(n_11546),
.B(n_10289),
.Y(n_12673)
);

AND2x4_ASAP7_75t_L g12674 ( 
.A(n_10972),
.B(n_10289),
.Y(n_12674)
);

AOI22xp5_ASAP7_75t_L g12675 ( 
.A1(n_11546),
.A2(n_7003),
.B1(n_7040),
.B2(n_6999),
.Y(n_12675)
);

AOI22xp33_ASAP7_75t_L g12676 ( 
.A1(n_11546),
.A2(n_7948),
.B1(n_7914),
.B2(n_6999),
.Y(n_12676)
);

INVx2_ASAP7_75t_L g12677 ( 
.A(n_11445),
.Y(n_12677)
);

HB1xp67_ASAP7_75t_L g12678 ( 
.A(n_11406),
.Y(n_12678)
);

OAI22xp33_ASAP7_75t_L g12679 ( 
.A1(n_11745),
.A2(n_8965),
.B1(n_9074),
.B2(n_8813),
.Y(n_12679)
);

HB1xp67_ASAP7_75t_L g12680 ( 
.A(n_11409),
.Y(n_12680)
);

OR2x2_ASAP7_75t_L g12681 ( 
.A(n_10818),
.B(n_10464),
.Y(n_12681)
);

AOI22xp33_ASAP7_75t_L g12682 ( 
.A1(n_11565),
.A2(n_7948),
.B1(n_7914),
.B2(n_6999),
.Y(n_12682)
);

INVx3_ASAP7_75t_L g12683 ( 
.A(n_11158),
.Y(n_12683)
);

NAND2xp5_ASAP7_75t_L g12684 ( 
.A(n_11409),
.B(n_8213),
.Y(n_12684)
);

OR2x2_ASAP7_75t_L g12685 ( 
.A(n_10875),
.B(n_9135),
.Y(n_12685)
);

AOI21xp5_ASAP7_75t_L g12686 ( 
.A1(n_11663),
.A2(n_8680),
.B(n_8676),
.Y(n_12686)
);

OAI222xp33_ASAP7_75t_L g12687 ( 
.A1(n_11745),
.A2(n_9550),
.B1(n_9621),
.B2(n_8218),
.C1(n_8846),
.C2(n_8443),
.Y(n_12687)
);

INVx2_ASAP7_75t_L g12688 ( 
.A(n_11451),
.Y(n_12688)
);

INVx1_ASAP7_75t_SL g12689 ( 
.A(n_11565),
.Y(n_12689)
);

AOI221xp5_ASAP7_75t_L g12690 ( 
.A1(n_11414),
.A2(n_9326),
.B1(n_9348),
.B2(n_9338),
.C(n_9332),
.Y(n_12690)
);

AOI22xp33_ASAP7_75t_L g12691 ( 
.A1(n_11565),
.A2(n_7948),
.B1(n_7914),
.B2(n_6999),
.Y(n_12691)
);

AOI22xp33_ASAP7_75t_L g12692 ( 
.A1(n_11578),
.A2(n_11787),
.B1(n_11799),
.B2(n_11695),
.Y(n_12692)
);

INVx2_ASAP7_75t_L g12693 ( 
.A(n_11451),
.Y(n_12693)
);

BUFx3_ASAP7_75t_L g12694 ( 
.A(n_11578),
.Y(n_12694)
);

INVx2_ASAP7_75t_L g12695 ( 
.A(n_11451),
.Y(n_12695)
);

AOI22xp33_ASAP7_75t_L g12696 ( 
.A1(n_11578),
.A2(n_7948),
.B1(n_7914),
.B2(n_7003),
.Y(n_12696)
);

NOR2xp33_ASAP7_75t_L g12697 ( 
.A(n_11825),
.B(n_7669),
.Y(n_12697)
);

CKINVDCx20_ASAP7_75t_R g12698 ( 
.A(n_11825),
.Y(n_12698)
);

BUFx4f_ASAP7_75t_L g12699 ( 
.A(n_11695),
.Y(n_12699)
);

OAI221xp5_ASAP7_75t_L g12700 ( 
.A1(n_11826),
.A2(n_9235),
.B1(n_8119),
.B2(n_10697),
.C(n_10566),
.Y(n_12700)
);

NAND2xp5_ASAP7_75t_L g12701 ( 
.A(n_11414),
.B(n_8213),
.Y(n_12701)
);

AND2x2_ASAP7_75t_L g12702 ( 
.A(n_11695),
.B(n_9406),
.Y(n_12702)
);

AOI22xp33_ASAP7_75t_L g12703 ( 
.A1(n_11787),
.A2(n_7914),
.B1(n_7003),
.B2(n_7045),
.Y(n_12703)
);

NOR2xp33_ASAP7_75t_L g12704 ( 
.A(n_11826),
.B(n_7721),
.Y(n_12704)
);

AOI22xp33_ASAP7_75t_SL g12705 ( 
.A1(n_11123),
.A2(n_7940),
.B1(n_7943),
.B2(n_8357),
.Y(n_12705)
);

AND2x2_ASAP7_75t_L g12706 ( 
.A(n_11787),
.B(n_9406),
.Y(n_12706)
);

INVx1_ASAP7_75t_L g12707 ( 
.A(n_11421),
.Y(n_12707)
);

OAI31xp33_ASAP7_75t_SL g12708 ( 
.A1(n_11799),
.A2(n_10306),
.A3(n_8845),
.B(n_8098),
.Y(n_12708)
);

OAI22xp33_ASAP7_75t_L g12709 ( 
.A1(n_11862),
.A2(n_8965),
.B1(n_9074),
.B2(n_8813),
.Y(n_12709)
);

AOI221xp5_ASAP7_75t_L g12710 ( 
.A1(n_11421),
.A2(n_9332),
.B1(n_9348),
.B2(n_9338),
.C(n_9326),
.Y(n_12710)
);

INVx1_ASAP7_75t_L g12711 ( 
.A(n_11453),
.Y(n_12711)
);

AND2x6_ASAP7_75t_SL g12712 ( 
.A(n_11799),
.B(n_11809),
.Y(n_12712)
);

AND2x4_ASAP7_75t_L g12713 ( 
.A(n_10972),
.B(n_10991),
.Y(n_12713)
);

AOI22xp33_ASAP7_75t_SL g12714 ( 
.A1(n_11123),
.A2(n_7940),
.B1(n_7943),
.B2(n_8357),
.Y(n_12714)
);

CKINVDCx11_ASAP7_75t_R g12715 ( 
.A(n_11809),
.Y(n_12715)
);

OAI211xp5_ASAP7_75t_L g12716 ( 
.A1(n_11453),
.A2(n_10697),
.B(n_10566),
.C(n_10265),
.Y(n_12716)
);

AOI22xp33_ASAP7_75t_SL g12717 ( 
.A1(n_11710),
.A2(n_8360),
.B1(n_9114),
.B2(n_9092),
.Y(n_12717)
);

OAI211xp5_ASAP7_75t_L g12718 ( 
.A1(n_11194),
.A2(n_10265),
.B(n_8408),
.C(n_10439),
.Y(n_12718)
);

OAI21xp33_ASAP7_75t_L g12719 ( 
.A1(n_11862),
.A2(n_7994),
.B(n_8098),
.Y(n_12719)
);

INVx1_ASAP7_75t_L g12720 ( 
.A(n_10753),
.Y(n_12720)
);

BUFx2_ASAP7_75t_L g12721 ( 
.A(n_10754),
.Y(n_12721)
);

AOI22xp33_ASAP7_75t_L g12722 ( 
.A1(n_11809),
.A2(n_7914),
.B1(n_7003),
.B2(n_7045),
.Y(n_12722)
);

INVx5_ASAP7_75t_SL g12723 ( 
.A(n_11874),
.Y(n_12723)
);

OAI22xp5_ASAP7_75t_L g12724 ( 
.A1(n_10727),
.A2(n_8693),
.B1(n_8661),
.B2(n_8296),
.Y(n_12724)
);

NAND2xp5_ASAP7_75t_L g12725 ( 
.A(n_10937),
.B(n_11920),
.Y(n_12725)
);

AOI22xp33_ASAP7_75t_L g12726 ( 
.A1(n_11874),
.A2(n_7045),
.B1(n_7046),
.B2(n_7040),
.Y(n_12726)
);

AND2x2_ASAP7_75t_L g12727 ( 
.A(n_11874),
.B(n_9450),
.Y(n_12727)
);

AO31x2_ASAP7_75t_L g12728 ( 
.A1(n_11223),
.A2(n_10541),
.A3(n_10563),
.B(n_10534),
.Y(n_12728)
);

AOI22xp33_ASAP7_75t_L g12729 ( 
.A1(n_10972),
.A2(n_7045),
.B1(n_7046),
.B2(n_7040),
.Y(n_12729)
);

INVx11_ASAP7_75t_L g12730 ( 
.A(n_10734),
.Y(n_12730)
);

INVx2_ASAP7_75t_SL g12731 ( 
.A(n_10754),
.Y(n_12731)
);

AND2x2_ASAP7_75t_L g12732 ( 
.A(n_10991),
.B(n_9450),
.Y(n_12732)
);

CKINVDCx5p33_ASAP7_75t_R g12733 ( 
.A(n_10757),
.Y(n_12733)
);

AND2x4_ASAP7_75t_L g12734 ( 
.A(n_10991),
.B(n_10849),
.Y(n_12734)
);

AND2x4_ASAP7_75t_L g12735 ( 
.A(n_10849),
.B(n_9345),
.Y(n_12735)
);

INVx1_ASAP7_75t_L g12736 ( 
.A(n_10766),
.Y(n_12736)
);

AND2x2_ASAP7_75t_L g12737 ( 
.A(n_11628),
.B(n_9521),
.Y(n_12737)
);

OR2x6_ASAP7_75t_L g12738 ( 
.A(n_10757),
.B(n_8813),
.Y(n_12738)
);

AOI222xp33_ASAP7_75t_L g12739 ( 
.A1(n_10727),
.A2(n_8272),
.B1(n_8117),
.B2(n_8099),
.C1(n_8127),
.C2(n_8118),
.Y(n_12739)
);

AND2x2_ASAP7_75t_L g12740 ( 
.A(n_11631),
.B(n_9521),
.Y(n_12740)
);

AND2x2_ASAP7_75t_L g12741 ( 
.A(n_11645),
.B(n_9525),
.Y(n_12741)
);

AOI22xp33_ASAP7_75t_L g12742 ( 
.A1(n_10923),
.A2(n_7045),
.B1(n_7046),
.B2(n_7040),
.Y(n_12742)
);

AND2x2_ASAP7_75t_L g12743 ( 
.A(n_10736),
.B(n_9525),
.Y(n_12743)
);

AND2x2_ASAP7_75t_L g12744 ( 
.A(n_10736),
.B(n_9540),
.Y(n_12744)
);

OAI22xp5_ASAP7_75t_L g12745 ( 
.A1(n_10923),
.A2(n_8693),
.B1(n_8661),
.B2(n_8296),
.Y(n_12745)
);

AO221x2_ASAP7_75t_L g12746 ( 
.A1(n_10937),
.A2(n_9332),
.B1(n_9348),
.B2(n_9338),
.C(n_9326),
.Y(n_12746)
);

OAI211xp5_ASAP7_75t_L g12747 ( 
.A1(n_11194),
.A2(n_10265),
.B(n_8408),
.C(n_10439),
.Y(n_12747)
);

AOI221xp5_ASAP7_75t_L g12748 ( 
.A1(n_11710),
.A2(n_9363),
.B1(n_9381),
.B2(n_9376),
.C(n_9352),
.Y(n_12748)
);

A2O1A1Ixp33_ASAP7_75t_L g12749 ( 
.A1(n_11135),
.A2(n_8099),
.B(n_8117),
.C(n_8109),
.Y(n_12749)
);

AO21x2_ASAP7_75t_L g12750 ( 
.A1(n_10923),
.A2(n_10563),
.B(n_10541),
.Y(n_12750)
);

OR2x2_ASAP7_75t_L g12751 ( 
.A(n_11927),
.B(n_9135),
.Y(n_12751)
);

AOI22xp33_ASAP7_75t_L g12752 ( 
.A1(n_11194),
.A2(n_7046),
.B1(n_7045),
.B2(n_8846),
.Y(n_12752)
);

HB1xp67_ASAP7_75t_L g12753 ( 
.A(n_10937),
.Y(n_12753)
);

OAI22xp5_ASAP7_75t_L g12754 ( 
.A1(n_11530),
.A2(n_8661),
.B1(n_8296),
.B2(n_8325),
.Y(n_12754)
);

OAI221xp5_ASAP7_75t_L g12755 ( 
.A1(n_11335),
.A2(n_8119),
.B1(n_10265),
.B2(n_8698),
.C(n_8735),
.Y(n_12755)
);

NOR3xp33_ASAP7_75t_L g12756 ( 
.A(n_10757),
.B(n_10517),
.C(n_10463),
.Y(n_12756)
);

AOI221xp5_ASAP7_75t_L g12757 ( 
.A1(n_10768),
.A2(n_9363),
.B1(n_9381),
.B2(n_9376),
.C(n_9352),
.Y(n_12757)
);

AOI22xp5_ASAP7_75t_L g12758 ( 
.A1(n_11732),
.A2(n_7046),
.B1(n_7216),
.B2(n_7109),
.Y(n_12758)
);

OR2x2_ASAP7_75t_L g12759 ( 
.A(n_11572),
.B(n_9152),
.Y(n_12759)
);

HB1xp67_ASAP7_75t_L g12760 ( 
.A(n_10937),
.Y(n_12760)
);

AOI22xp33_ASAP7_75t_SL g12761 ( 
.A1(n_11468),
.A2(n_8360),
.B1(n_9114),
.B2(n_9092),
.Y(n_12761)
);

INVx2_ASAP7_75t_L g12762 ( 
.A(n_11530),
.Y(n_12762)
);

AOI22xp33_ASAP7_75t_L g12763 ( 
.A1(n_11530),
.A2(n_7046),
.B1(n_8846),
.B2(n_8408),
.Y(n_12763)
);

INVx1_ASAP7_75t_L g12764 ( 
.A(n_10780),
.Y(n_12764)
);

INVx1_ASAP7_75t_L g12765 ( 
.A(n_10781),
.Y(n_12765)
);

AND2x4_ASAP7_75t_L g12766 ( 
.A(n_11544),
.B(n_9345),
.Y(n_12766)
);

AOI22xp5_ASAP7_75t_L g12767 ( 
.A1(n_11746),
.A2(n_7216),
.B1(n_7331),
.B2(n_7109),
.Y(n_12767)
);

AOI22xp33_ASAP7_75t_L g12768 ( 
.A1(n_11544),
.A2(n_8846),
.B1(n_8408),
.B2(n_9241),
.Y(n_12768)
);

NOR2xp33_ASAP7_75t_L g12769 ( 
.A(n_11916),
.B(n_7728),
.Y(n_12769)
);

INVx2_ASAP7_75t_L g12770 ( 
.A(n_11544),
.Y(n_12770)
);

A2O1A1Ixp33_ASAP7_75t_L g12771 ( 
.A1(n_11623),
.A2(n_8109),
.B(n_8118),
.C(n_8117),
.Y(n_12771)
);

OAI221xp5_ASAP7_75t_L g12772 ( 
.A1(n_11174),
.A2(n_11190),
.B1(n_11209),
.B2(n_11203),
.C(n_11188),
.Y(n_12772)
);

INVx2_ASAP7_75t_L g12773 ( 
.A(n_11577),
.Y(n_12773)
);

AOI22xp33_ASAP7_75t_L g12774 ( 
.A1(n_11577),
.A2(n_8846),
.B1(n_8408),
.B2(n_9241),
.Y(n_12774)
);

BUFx2_ASAP7_75t_L g12775 ( 
.A(n_11577),
.Y(n_12775)
);

OAI211xp5_ASAP7_75t_L g12776 ( 
.A1(n_11264),
.A2(n_10439),
.B(n_8358),
.C(n_9747),
.Y(n_12776)
);

AOI22xp33_ASAP7_75t_SL g12777 ( 
.A1(n_11468),
.A2(n_8360),
.B1(n_9114),
.B2(n_9092),
.Y(n_12777)
);

INVx2_ASAP7_75t_L g12778 ( 
.A(n_10777),
.Y(n_12778)
);

AOI22xp33_ASAP7_75t_L g12779 ( 
.A1(n_11760),
.A2(n_8846),
.B1(n_9272),
.B2(n_9241),
.Y(n_12779)
);

INVx1_ASAP7_75t_L g12780 ( 
.A(n_10782),
.Y(n_12780)
);

INVx2_ASAP7_75t_L g12781 ( 
.A(n_10777),
.Y(n_12781)
);

BUFx2_ASAP7_75t_L g12782 ( 
.A(n_11541),
.Y(n_12782)
);

OAI221xp5_ASAP7_75t_L g12783 ( 
.A1(n_11174),
.A2(n_8119),
.B1(n_8698),
.B2(n_8735),
.C(n_8676),
.Y(n_12783)
);

INVx1_ASAP7_75t_L g12784 ( 
.A(n_10787),
.Y(n_12784)
);

INVx1_ASAP7_75t_L g12785 ( 
.A(n_10791),
.Y(n_12785)
);

CKINVDCx20_ASAP7_75t_R g12786 ( 
.A(n_11831),
.Y(n_12786)
);

AOI22xp33_ASAP7_75t_SL g12787 ( 
.A1(n_11477),
.A2(n_9114),
.B1(n_9179),
.B2(n_9092),
.Y(n_12787)
);

AOI221x1_ASAP7_75t_SL g12788 ( 
.A1(n_11921),
.A2(n_10306),
.B1(n_9376),
.B2(n_9381),
.C(n_9363),
.Y(n_12788)
);

OAI21x1_ASAP7_75t_L g12789 ( 
.A1(n_11623),
.A2(n_10517),
.B(n_10463),
.Y(n_12789)
);

AOI22xp33_ASAP7_75t_L g12790 ( 
.A1(n_11833),
.A2(n_8846),
.B1(n_9272),
.B2(n_9241),
.Y(n_12790)
);

AND2x2_ASAP7_75t_L g12791 ( 
.A(n_11844),
.B(n_9540),
.Y(n_12791)
);

AOI322xp5_ASAP7_75t_L g12792 ( 
.A1(n_11223),
.A2(n_9396),
.A3(n_9393),
.B1(n_9401),
.B2(n_9409),
.C1(n_9394),
.C2(n_9352),
.Y(n_12792)
);

OA21x2_ASAP7_75t_L g12793 ( 
.A1(n_11227),
.A2(n_10565),
.B(n_10563),
.Y(n_12793)
);

AOI22xp33_ASAP7_75t_L g12794 ( 
.A1(n_11854),
.A2(n_9241),
.B1(n_9272),
.B2(n_8119),
.Y(n_12794)
);

INVx3_ASAP7_75t_L g12795 ( 
.A(n_10777),
.Y(n_12795)
);

OAI21x1_ASAP7_75t_L g12796 ( 
.A1(n_11255),
.A2(n_10530),
.B(n_10517),
.Y(n_12796)
);

NAND2xp5_ASAP7_75t_L g12797 ( 
.A(n_11881),
.B(n_8258),
.Y(n_12797)
);

NAND2x1p5_ASAP7_75t_L g12798 ( 
.A(n_10830),
.B(n_8813),
.Y(n_12798)
);

AND2x4_ASAP7_75t_L g12799 ( 
.A(n_11693),
.B(n_9347),
.Y(n_12799)
);

AOI22xp33_ASAP7_75t_L g12800 ( 
.A1(n_11892),
.A2(n_9241),
.B1(n_9272),
.B2(n_8119),
.Y(n_12800)
);

NAND3xp33_ASAP7_75t_L g12801 ( 
.A(n_11264),
.B(n_8358),
.C(n_8374),
.Y(n_12801)
);

OAI22xp5_ASAP7_75t_L g12802 ( 
.A1(n_11174),
.A2(n_8661),
.B1(n_8296),
.B2(n_8325),
.Y(n_12802)
);

OR2x2_ASAP7_75t_L g12803 ( 
.A(n_10796),
.B(n_9152),
.Y(n_12803)
);

AOI22xp33_ASAP7_75t_L g12804 ( 
.A1(n_11895),
.A2(n_9272),
.B1(n_9241),
.B2(n_7216),
.Y(n_12804)
);

AOI22xp5_ASAP7_75t_L g12805 ( 
.A1(n_11907),
.A2(n_7216),
.B1(n_7331),
.B2(n_7109),
.Y(n_12805)
);

OR2x2_ASAP7_75t_L g12806 ( 
.A(n_10808),
.B(n_9157),
.Y(n_12806)
);

AOI221xp5_ASAP7_75t_L g12807 ( 
.A1(n_10810),
.A2(n_10820),
.B1(n_10823),
.B2(n_10817),
.C(n_10816),
.Y(n_12807)
);

NOR2xp33_ASAP7_75t_L g12808 ( 
.A(n_11918),
.B(n_7728),
.Y(n_12808)
);

AOI22xp33_ASAP7_75t_SL g12809 ( 
.A1(n_11477),
.A2(n_9114),
.B1(n_9179),
.B2(n_9092),
.Y(n_12809)
);

OAI22xp5_ASAP7_75t_L g12810 ( 
.A1(n_11188),
.A2(n_8661),
.B1(n_8296),
.B2(n_8325),
.Y(n_12810)
);

AOI22xp33_ASAP7_75t_L g12811 ( 
.A1(n_11923),
.A2(n_9272),
.B1(n_7331),
.B2(n_7373),
.Y(n_12811)
);

NAND3xp33_ASAP7_75t_L g12812 ( 
.A(n_11264),
.B(n_8358),
.C(n_8374),
.Y(n_12812)
);

NAND2xp5_ASAP7_75t_L g12813 ( 
.A(n_11929),
.B(n_8258),
.Y(n_12813)
);

OAI21x1_ASAP7_75t_L g12814 ( 
.A1(n_11887),
.A2(n_10546),
.B(n_10530),
.Y(n_12814)
);

AOI22xp33_ASAP7_75t_L g12815 ( 
.A1(n_11188),
.A2(n_9272),
.B1(n_7331),
.B2(n_7373),
.Y(n_12815)
);

NAND2xp5_ASAP7_75t_L g12816 ( 
.A(n_11769),
.B(n_8302),
.Y(n_12816)
);

AOI22xp33_ASAP7_75t_L g12817 ( 
.A1(n_11190),
.A2(n_7331),
.B1(n_7373),
.B2(n_7216),
.Y(n_12817)
);

AOI22xp33_ASAP7_75t_L g12818 ( 
.A1(n_11190),
.A2(n_7331),
.B1(n_7373),
.B2(n_7216),
.Y(n_12818)
);

NAND2xp5_ASAP7_75t_L g12819 ( 
.A(n_10827),
.B(n_8302),
.Y(n_12819)
);

INVx2_ASAP7_75t_L g12820 ( 
.A(n_10830),
.Y(n_12820)
);

BUFx12f_ASAP7_75t_L g12821 ( 
.A(n_10830),
.Y(n_12821)
);

AOI22xp33_ASAP7_75t_L g12822 ( 
.A1(n_11203),
.A2(n_7331),
.B1(n_7373),
.B2(n_7216),
.Y(n_12822)
);

INVx1_ASAP7_75t_L g12823 ( 
.A(n_10831),
.Y(n_12823)
);

BUFx2_ASAP7_75t_L g12824 ( 
.A(n_11541),
.Y(n_12824)
);

AOI221xp5_ASAP7_75t_L g12825 ( 
.A1(n_10835),
.A2(n_9394),
.B1(n_9401),
.B2(n_9396),
.C(n_9393),
.Y(n_12825)
);

AOI21xp5_ASAP7_75t_L g12826 ( 
.A1(n_11502),
.A2(n_8514),
.B(n_7733),
.Y(n_12826)
);

OAI22xp33_ASAP7_75t_SL g12827 ( 
.A1(n_10898),
.A2(n_10530),
.B1(n_10553),
.B2(n_10546),
.Y(n_12827)
);

OR2x2_ASAP7_75t_L g12828 ( 
.A(n_10836),
.B(n_9157),
.Y(n_12828)
);

NOR2xp33_ASAP7_75t_L g12829 ( 
.A(n_11203),
.B(n_7733),
.Y(n_12829)
);

AOI21xp33_ASAP7_75t_L g12830 ( 
.A1(n_11502),
.A2(n_8514),
.B(n_7996),
.Y(n_12830)
);

CKINVDCx5p33_ASAP7_75t_R g12831 ( 
.A(n_10898),
.Y(n_12831)
);

INVx2_ASAP7_75t_L g12832 ( 
.A(n_10898),
.Y(n_12832)
);

AND2x2_ASAP7_75t_L g12833 ( 
.A(n_11209),
.B(n_9544),
.Y(n_12833)
);

OR2x2_ASAP7_75t_L g12834 ( 
.A(n_10838),
.B(n_9167),
.Y(n_12834)
);

BUFx5_ASAP7_75t_L g12835 ( 
.A(n_10839),
.Y(n_12835)
);

OR2x2_ASAP7_75t_L g12836 ( 
.A(n_10854),
.B(n_9167),
.Y(n_12836)
);

AOI22xp33_ASAP7_75t_L g12837 ( 
.A1(n_11209),
.A2(n_7373),
.B1(n_7331),
.B2(n_7019),
.Y(n_12837)
);

AOI22xp33_ASAP7_75t_SL g12838 ( 
.A1(n_11229),
.A2(n_9114),
.B1(n_9179),
.B2(n_9092),
.Y(n_12838)
);

OAI22xp5_ASAP7_75t_L g12839 ( 
.A1(n_11229),
.A2(n_8661),
.B1(n_8087),
.B2(n_8325),
.Y(n_12839)
);

NAND2xp5_ASAP7_75t_L g12840 ( 
.A(n_10855),
.B(n_8316),
.Y(n_12840)
);

OAI22xp5_ASAP7_75t_L g12841 ( 
.A1(n_11229),
.A2(n_8661),
.B1(n_8087),
.B2(n_8325),
.Y(n_12841)
);

OAI22xp5_ASAP7_75t_L g12842 ( 
.A1(n_10899),
.A2(n_8087),
.B1(n_8325),
.B2(n_8296),
.Y(n_12842)
);

AOI21xp5_ASAP7_75t_L g12843 ( 
.A1(n_11502),
.A2(n_8514),
.B(n_10049),
.Y(n_12843)
);

AOI222xp33_ASAP7_75t_L g12844 ( 
.A1(n_11227),
.A2(n_8127),
.B1(n_8109),
.B2(n_8134),
.C1(n_8118),
.C2(n_9255),
.Y(n_12844)
);

INVx2_ASAP7_75t_L g12845 ( 
.A(n_10899),
.Y(n_12845)
);

BUFx2_ASAP7_75t_L g12846 ( 
.A(n_11541),
.Y(n_12846)
);

BUFx5_ASAP7_75t_L g12847 ( 
.A(n_10856),
.Y(n_12847)
);

INVx2_ASAP7_75t_L g12848 ( 
.A(n_10899),
.Y(n_12848)
);

AND2x2_ASAP7_75t_L g12849 ( 
.A(n_11541),
.B(n_9544),
.Y(n_12849)
);

AND2x4_ASAP7_75t_L g12850 ( 
.A(n_10913),
.B(n_9347),
.Y(n_12850)
);

OAI22xp5_ASAP7_75t_L g12851 ( 
.A1(n_10913),
.A2(n_8087),
.B1(n_8325),
.B2(n_8296),
.Y(n_12851)
);

AOI21xp5_ASAP7_75t_L g12852 ( 
.A1(n_11514),
.A2(n_8514),
.B(n_10049),
.Y(n_12852)
);

NAND2xp5_ASAP7_75t_L g12853 ( 
.A(n_10857),
.B(n_8316),
.Y(n_12853)
);

INVx2_ASAP7_75t_L g12854 ( 
.A(n_10913),
.Y(n_12854)
);

OR2x6_ASAP7_75t_L g12855 ( 
.A(n_10929),
.B(n_8813),
.Y(n_12855)
);

AND2x2_ASAP7_75t_L g12856 ( 
.A(n_11599),
.B(n_9552),
.Y(n_12856)
);

NAND2xp5_ASAP7_75t_L g12857 ( 
.A(n_10859),
.B(n_8557),
.Y(n_12857)
);

AOI22xp33_ASAP7_75t_L g12858 ( 
.A1(n_11514),
.A2(n_7373),
.B1(n_7019),
.B2(n_7063),
.Y(n_12858)
);

BUFx3_ASAP7_75t_L g12859 ( 
.A(n_10929),
.Y(n_12859)
);

AOI22xp33_ASAP7_75t_SL g12860 ( 
.A1(n_10929),
.A2(n_9179),
.B1(n_8127),
.B2(n_8134),
.Y(n_12860)
);

INVx2_ASAP7_75t_L g12861 ( 
.A(n_10950),
.Y(n_12861)
);

AOI22xp5_ASAP7_75t_L g12862 ( 
.A1(n_11514),
.A2(n_7373),
.B1(n_8379),
.B2(n_8253),
.Y(n_12862)
);

OAI22xp5_ASAP7_75t_L g12863 ( 
.A1(n_10950),
.A2(n_8469),
.B1(n_8651),
.B2(n_8087),
.Y(n_12863)
);

AOI33xp33_ASAP7_75t_L g12864 ( 
.A1(n_10865),
.A2(n_9133),
.A3(n_9393),
.B1(n_9401),
.B2(n_9396),
.B3(n_9394),
.Y(n_12864)
);

NOR2xp33_ASAP7_75t_L g12865 ( 
.A(n_10950),
.B(n_7550),
.Y(n_12865)
);

AOI22xp33_ASAP7_75t_L g12866 ( 
.A1(n_10959),
.A2(n_7019),
.B1(n_7063),
.B2(n_6946),
.Y(n_12866)
);

OAI22xp5_ASAP7_75t_L g12867 ( 
.A1(n_10959),
.A2(n_8651),
.B1(n_9234),
.B2(n_8469),
.Y(n_12867)
);

NAND3xp33_ASAP7_75t_L g12868 ( 
.A(n_11783),
.B(n_8358),
.C(n_8374),
.Y(n_12868)
);

INVx2_ASAP7_75t_L g12869 ( 
.A(n_10959),
.Y(n_12869)
);

OAI22xp5_ASAP7_75t_L g12870 ( 
.A1(n_11003),
.A2(n_8651),
.B1(n_9234),
.B2(n_8469),
.Y(n_12870)
);

AOI22xp33_ASAP7_75t_L g12871 ( 
.A1(n_11003),
.A2(n_7019),
.B1(n_7063),
.B2(n_6946),
.Y(n_12871)
);

AND2x2_ASAP7_75t_L g12872 ( 
.A(n_11599),
.B(n_9552),
.Y(n_12872)
);

AOI21xp33_ASAP7_75t_L g12873 ( 
.A1(n_11003),
.A2(n_8514),
.B(n_11005),
.Y(n_12873)
);

OAI211xp5_ASAP7_75t_L g12874 ( 
.A1(n_11661),
.A2(n_10439),
.B(n_8358),
.C(n_9747),
.Y(n_12874)
);

OAI21xp5_ASAP7_75t_L g12875 ( 
.A1(n_10988),
.A2(n_8330),
.B(n_7994),
.Y(n_12875)
);

NOR2xp33_ASAP7_75t_L g12876 ( 
.A(n_11005),
.B(n_7550),
.Y(n_12876)
);

AOI21x1_ASAP7_75t_L g12877 ( 
.A1(n_11245),
.A2(n_10329),
.B(n_10325),
.Y(n_12877)
);

AOI31xp33_ASAP7_75t_L g12878 ( 
.A1(n_10742),
.A2(n_7543),
.A3(n_7541),
.B(n_9209),
.Y(n_12878)
);

OAI22xp5_ASAP7_75t_L g12879 ( 
.A1(n_11005),
.A2(n_8651),
.B1(n_9234),
.B2(n_8469),
.Y(n_12879)
);

AOI222xp33_ASAP7_75t_L g12880 ( 
.A1(n_11245),
.A2(n_8134),
.B1(n_9255),
.B2(n_8163),
.C1(n_8330),
.C2(n_7095),
.Y(n_12880)
);

AOI22xp33_ASAP7_75t_L g12881 ( 
.A1(n_11023),
.A2(n_7019),
.B1(n_7063),
.B2(n_6946),
.Y(n_12881)
);

AO21x2_ASAP7_75t_L g12882 ( 
.A1(n_11251),
.A2(n_11254),
.B(n_11253),
.Y(n_12882)
);

AOI22xp33_ASAP7_75t_L g12883 ( 
.A1(n_11023),
.A2(n_7019),
.B1(n_7063),
.B2(n_6946),
.Y(n_12883)
);

AND2x2_ASAP7_75t_L g12884 ( 
.A(n_11599),
.B(n_9562),
.Y(n_12884)
);

AOI22xp33_ASAP7_75t_L g12885 ( 
.A1(n_11023),
.A2(n_7019),
.B1(n_7063),
.B2(n_6946),
.Y(n_12885)
);

OAI21xp5_ASAP7_75t_L g12886 ( 
.A1(n_10988),
.A2(n_8330),
.B(n_8163),
.Y(n_12886)
);

AND2x2_ASAP7_75t_L g12887 ( 
.A(n_11599),
.B(n_9562),
.Y(n_12887)
);

INVx1_ASAP7_75t_L g12888 ( 
.A(n_10866),
.Y(n_12888)
);

AOI221xp5_ASAP7_75t_L g12889 ( 
.A1(n_10868),
.A2(n_9409),
.B1(n_9425),
.B2(n_9415),
.C(n_9410),
.Y(n_12889)
);

OAI21x1_ASAP7_75t_L g12890 ( 
.A1(n_11887),
.A2(n_10546),
.B(n_10530),
.Y(n_12890)
);

INVx2_ASAP7_75t_L g12891 ( 
.A(n_11086),
.Y(n_12891)
);

NAND2xp5_ASAP7_75t_L g12892 ( 
.A(n_10873),
.B(n_8557),
.Y(n_12892)
);

AOI221x1_ASAP7_75t_L g12893 ( 
.A1(n_11086),
.A2(n_10579),
.B1(n_10602),
.B2(n_10553),
.C(n_10546),
.Y(n_12893)
);

AND2x2_ASAP7_75t_L g12894 ( 
.A(n_11404),
.B(n_9598),
.Y(n_12894)
);

OR2x2_ASAP7_75t_L g12895 ( 
.A(n_10880),
.B(n_9218),
.Y(n_12895)
);

NAND3xp33_ASAP7_75t_L g12896 ( 
.A(n_11783),
.B(n_8377),
.C(n_8374),
.Y(n_12896)
);

OAI211xp5_ASAP7_75t_SL g12897 ( 
.A1(n_11086),
.A2(n_10579),
.B(n_10602),
.C(n_10553),
.Y(n_12897)
);

INVx1_ASAP7_75t_L g12898 ( 
.A(n_10897),
.Y(n_12898)
);

INVx1_ASAP7_75t_L g12899 ( 
.A(n_10909),
.Y(n_12899)
);

AOI22xp33_ASAP7_75t_L g12900 ( 
.A1(n_11092),
.A2(n_7019),
.B1(n_7063),
.B2(n_6946),
.Y(n_12900)
);

OAI22xp33_ASAP7_75t_L g12901 ( 
.A1(n_11092),
.A2(n_8965),
.B1(n_9074),
.B2(n_8813),
.Y(n_12901)
);

AND2x2_ASAP7_75t_L g12902 ( 
.A(n_11404),
.B(n_9598),
.Y(n_12902)
);

OAI221xp5_ASAP7_75t_L g12903 ( 
.A1(n_11092),
.A2(n_8528),
.B1(n_8556),
.B2(n_8447),
.C(n_8443),
.Y(n_12903)
);

INVx1_ASAP7_75t_L g12904 ( 
.A(n_10910),
.Y(n_12904)
);

INVx2_ASAP7_75t_L g12905 ( 
.A(n_11095),
.Y(n_12905)
);

INVx1_ASAP7_75t_L g12906 ( 
.A(n_10914),
.Y(n_12906)
);

AOI22xp33_ASAP7_75t_L g12907 ( 
.A1(n_11095),
.A2(n_7063),
.B1(n_6946),
.B2(n_7996),
.Y(n_12907)
);

AOI221xp5_ASAP7_75t_L g12908 ( 
.A1(n_10915),
.A2(n_9410),
.B1(n_9425),
.B2(n_9415),
.C(n_9409),
.Y(n_12908)
);

OR2x2_ASAP7_75t_L g12909 ( 
.A(n_10916),
.B(n_9218),
.Y(n_12909)
);

OAI22xp5_ASAP7_75t_L g12910 ( 
.A1(n_11095),
.A2(n_8651),
.B1(n_9234),
.B2(n_8469),
.Y(n_12910)
);

OR2x2_ASAP7_75t_L g12911 ( 
.A(n_10921),
.B(n_9229),
.Y(n_12911)
);

OAI22xp5_ASAP7_75t_L g12912 ( 
.A1(n_11133),
.A2(n_8651),
.B1(n_9234),
.B2(n_8469),
.Y(n_12912)
);

INVx1_ASAP7_75t_L g12913 ( 
.A(n_10925),
.Y(n_12913)
);

INVx1_ASAP7_75t_SL g12914 ( 
.A(n_11133),
.Y(n_12914)
);

HB1xp67_ASAP7_75t_SL g12915 ( 
.A(n_10926),
.Y(n_12915)
);

AOI22xp33_ASAP7_75t_L g12916 ( 
.A1(n_11133),
.A2(n_6946),
.B1(n_7996),
.B2(n_9179),
.Y(n_12916)
);

AOI221xp5_ASAP7_75t_L g12917 ( 
.A1(n_10927),
.A2(n_9415),
.B1(n_9443),
.B2(n_9425),
.C(n_9410),
.Y(n_12917)
);

AOI22xp5_ASAP7_75t_L g12918 ( 
.A1(n_11157),
.A2(n_8253),
.B1(n_8379),
.B2(n_10306),
.Y(n_12918)
);

AOI22xp33_ASAP7_75t_L g12919 ( 
.A1(n_11157),
.A2(n_9179),
.B1(n_8845),
.B2(n_9086),
.Y(n_12919)
);

OAI221xp5_ASAP7_75t_L g12920 ( 
.A1(n_11157),
.A2(n_8528),
.B1(n_8556),
.B2(n_8447),
.C(n_8443),
.Y(n_12920)
);

AOI22xp33_ASAP7_75t_L g12921 ( 
.A1(n_11165),
.A2(n_9086),
.B1(n_9060),
.B2(n_8528),
.Y(n_12921)
);

INVx1_ASAP7_75t_L g12922 ( 
.A(n_10936),
.Y(n_12922)
);

AND2x6_ASAP7_75t_L g12923 ( 
.A(n_11165),
.B(n_7757),
.Y(n_12923)
);

OAI221xp5_ASAP7_75t_L g12924 ( 
.A1(n_11165),
.A2(n_11259),
.B1(n_11238),
.B2(n_8653),
.C(n_8681),
.Y(n_12924)
);

AND2x2_ASAP7_75t_L g12925 ( 
.A(n_11404),
.B(n_9617),
.Y(n_12925)
);

INVx1_ASAP7_75t_L g12926 ( 
.A(n_10939),
.Y(n_12926)
);

AOI22xp33_ASAP7_75t_L g12927 ( 
.A1(n_11661),
.A2(n_9086),
.B1(n_9060),
.B2(n_8556),
.Y(n_12927)
);

AOI221xp5_ASAP7_75t_L g12928 ( 
.A1(n_10940),
.A2(n_9445),
.B1(n_9467),
.B2(n_9460),
.C(n_9443),
.Y(n_12928)
);

INVx2_ASAP7_75t_L g12929 ( 
.A(n_11238),
.Y(n_12929)
);

AOI22xp33_ASAP7_75t_L g12930 ( 
.A1(n_11661),
.A2(n_9086),
.B1(n_9060),
.B2(n_8653),
.Y(n_12930)
);

AOI22xp33_ASAP7_75t_L g12931 ( 
.A1(n_10941),
.A2(n_9086),
.B1(n_9060),
.B2(n_8653),
.Y(n_12931)
);

NAND3xp33_ASAP7_75t_L g12932 ( 
.A(n_11783),
.B(n_8377),
.C(n_8374),
.Y(n_12932)
);

INVx1_ASAP7_75t_L g12933 ( 
.A(n_10946),
.Y(n_12933)
);

INVx1_ASAP7_75t_L g12934 ( 
.A(n_10947),
.Y(n_12934)
);

OAI22xp5_ASAP7_75t_L g12935 ( 
.A1(n_11259),
.A2(n_8469),
.B1(n_9234),
.B2(n_8651),
.Y(n_12935)
);

AND2x4_ASAP7_75t_SL g12936 ( 
.A(n_11259),
.B(n_7763),
.Y(n_12936)
);

INVx2_ASAP7_75t_L g12937 ( 
.A(n_11660),
.Y(n_12937)
);

INVx1_ASAP7_75t_L g12938 ( 
.A(n_10948),
.Y(n_12938)
);

OAI21x1_ASAP7_75t_L g12939 ( 
.A1(n_10828),
.A2(n_10579),
.B(n_10553),
.Y(n_12939)
);

AOI22xp33_ASAP7_75t_L g12940 ( 
.A1(n_10952),
.A2(n_9086),
.B1(n_9060),
.B2(n_8681),
.Y(n_12940)
);

AOI21xp33_ASAP7_75t_L g12941 ( 
.A1(n_10962),
.A2(n_8574),
.B(n_8554),
.Y(n_12941)
);

AOI22xp5_ASAP7_75t_L g12942 ( 
.A1(n_10963),
.A2(n_8253),
.B1(n_8379),
.B2(n_7240),
.Y(n_12942)
);

INVx2_ASAP7_75t_L g12943 ( 
.A(n_11660),
.Y(n_12943)
);

AOI22xp33_ASAP7_75t_L g12944 ( 
.A1(n_10967),
.A2(n_9060),
.B1(n_8681),
.B2(n_8763),
.Y(n_12944)
);

INVx1_ASAP7_75t_L g12945 ( 
.A(n_10969),
.Y(n_12945)
);

OAI221xp5_ASAP7_75t_L g12946 ( 
.A1(n_10973),
.A2(n_8792),
.B1(n_8890),
.B2(n_8763),
.C(n_8447),
.Y(n_12946)
);

AND2x2_ASAP7_75t_L g12947 ( 
.A(n_11404),
.B(n_9617),
.Y(n_12947)
);

AND2x2_ASAP7_75t_L g12948 ( 
.A(n_11925),
.B(n_9658),
.Y(n_12948)
);

AOI21xp5_ASAP7_75t_L g12949 ( 
.A1(n_10987),
.A2(n_10049),
.B(n_9747),
.Y(n_12949)
);

INVx1_ASAP7_75t_L g12950 ( 
.A(n_10975),
.Y(n_12950)
);

OAI21x1_ASAP7_75t_L g12951 ( 
.A1(n_10828),
.A2(n_10602),
.B(n_10579),
.Y(n_12951)
);

AOI21xp5_ASAP7_75t_L g12952 ( 
.A1(n_10987),
.A2(n_10049),
.B(n_9747),
.Y(n_12952)
);

CKINVDCx6p67_ASAP7_75t_R g12953 ( 
.A(n_10982),
.Y(n_12953)
);

OAI221xp5_ASAP7_75t_L g12954 ( 
.A1(n_10983),
.A2(n_8890),
.B1(n_9123),
.B2(n_8792),
.C(n_8763),
.Y(n_12954)
);

AOI22xp33_ASAP7_75t_L g12955 ( 
.A1(n_10996),
.A2(n_8890),
.B1(n_9123),
.B2(n_8792),
.Y(n_12955)
);

AOI221xp5_ASAP7_75t_L g12956 ( 
.A1(n_11000),
.A2(n_9445),
.B1(n_9467),
.B2(n_9460),
.C(n_9443),
.Y(n_12956)
);

CKINVDCx5p33_ASAP7_75t_R g12957 ( 
.A(n_11660),
.Y(n_12957)
);

INVx1_ASAP7_75t_L g12958 ( 
.A(n_11007),
.Y(n_12958)
);

NAND3xp33_ASAP7_75t_L g12959 ( 
.A(n_11865),
.B(n_8377),
.C(n_8374),
.Y(n_12959)
);

INVxp67_ASAP7_75t_L g12960 ( 
.A(n_12915),
.Y(n_12960)
);

INVx1_ASAP7_75t_L g12961 ( 
.A(n_11945),
.Y(n_12961)
);

CKINVDCx5p33_ASAP7_75t_R g12962 ( 
.A(n_12028),
.Y(n_12962)
);

NAND2xp5_ASAP7_75t_L g12963 ( 
.A(n_12591),
.B(n_9962),
.Y(n_12963)
);

INVxp67_ASAP7_75t_R g12964 ( 
.A(n_12491),
.Y(n_12964)
);

INVx1_ASAP7_75t_L g12965 ( 
.A(n_12179),
.Y(n_12965)
);

HB1xp67_ASAP7_75t_L g12966 ( 
.A(n_12205),
.Y(n_12966)
);

AND2x2_ASAP7_75t_L g12967 ( 
.A(n_11946),
.B(n_12022),
.Y(n_12967)
);

INVx1_ASAP7_75t_L g12968 ( 
.A(n_12279),
.Y(n_12968)
);

INVx1_ASAP7_75t_SL g12969 ( 
.A(n_12443),
.Y(n_12969)
);

INVxp67_ASAP7_75t_L g12970 ( 
.A(n_12424),
.Y(n_12970)
);

CKINVDCx20_ASAP7_75t_R g12971 ( 
.A(n_12082),
.Y(n_12971)
);

INVx2_ASAP7_75t_L g12972 ( 
.A(n_12075),
.Y(n_12972)
);

NAND2xp5_ASAP7_75t_L g12973 ( 
.A(n_11951),
.B(n_9962),
.Y(n_12973)
);

NAND2xp5_ASAP7_75t_L g12974 ( 
.A(n_11960),
.B(n_9968),
.Y(n_12974)
);

OR2x2_ASAP7_75t_L g12975 ( 
.A(n_11947),
.B(n_11008),
.Y(n_12975)
);

INVx1_ASAP7_75t_L g12976 ( 
.A(n_12295),
.Y(n_12976)
);

INVx1_ASAP7_75t_L g12977 ( 
.A(n_12332),
.Y(n_12977)
);

INVx1_ASAP7_75t_L g12978 ( 
.A(n_12410),
.Y(n_12978)
);

AND2x2_ASAP7_75t_L g12979 ( 
.A(n_11934),
.B(n_9658),
.Y(n_12979)
);

AND2x2_ASAP7_75t_L g12980 ( 
.A(n_11948),
.B(n_9672),
.Y(n_12980)
);

AND2x2_ASAP7_75t_L g12981 ( 
.A(n_12351),
.B(n_12112),
.Y(n_12981)
);

AND2x4_ASAP7_75t_L g12982 ( 
.A(n_12166),
.B(n_9681),
.Y(n_12982)
);

AND2x2_ASAP7_75t_L g12983 ( 
.A(n_11949),
.B(n_9672),
.Y(n_12983)
);

INVx5_ASAP7_75t_SL g12984 ( 
.A(n_12011),
.Y(n_12984)
);

OR2x2_ASAP7_75t_L g12985 ( 
.A(n_11953),
.B(n_11013),
.Y(n_12985)
);

AND2x2_ASAP7_75t_L g12986 ( 
.A(n_12448),
.B(n_9683),
.Y(n_12986)
);

NAND2xp5_ASAP7_75t_L g12987 ( 
.A(n_11982),
.B(n_9968),
.Y(n_12987)
);

OR2x2_ASAP7_75t_L g12988 ( 
.A(n_11983),
.B(n_11015),
.Y(n_12988)
);

INVx2_ASAP7_75t_L g12989 ( 
.A(n_12187),
.Y(n_12989)
);

INVx1_ASAP7_75t_L g12990 ( 
.A(n_12470),
.Y(n_12990)
);

INVx2_ASAP7_75t_L g12991 ( 
.A(n_12259),
.Y(n_12991)
);

AND2x4_ASAP7_75t_L g12992 ( 
.A(n_12166),
.B(n_9681),
.Y(n_12992)
);

AOI22xp33_ASAP7_75t_SL g12993 ( 
.A1(n_12058),
.A2(n_12054),
.B1(n_11941),
.B2(n_11955),
.Y(n_12993)
);

OR2x2_ASAP7_75t_L g12994 ( 
.A(n_11997),
.B(n_11024),
.Y(n_12994)
);

INVx2_ASAP7_75t_L g12995 ( 
.A(n_12423),
.Y(n_12995)
);

BUFx6f_ASAP7_75t_L g12996 ( 
.A(n_12606),
.Y(n_12996)
);

INVx1_ASAP7_75t_SL g12997 ( 
.A(n_12043),
.Y(n_12997)
);

INVx3_ASAP7_75t_L g12998 ( 
.A(n_12337),
.Y(n_12998)
);

NAND2xp5_ASAP7_75t_L g12999 ( 
.A(n_11999),
.B(n_9999),
.Y(n_12999)
);

INVx1_ASAP7_75t_L g13000 ( 
.A(n_12472),
.Y(n_13000)
);

NAND2xp5_ASAP7_75t_L g13001 ( 
.A(n_12004),
.B(n_12041),
.Y(n_13001)
);

AND2x2_ASAP7_75t_L g13002 ( 
.A(n_12108),
.B(n_9683),
.Y(n_13002)
);

INVx1_ASAP7_75t_L g13003 ( 
.A(n_12478),
.Y(n_13003)
);

AND2x2_ASAP7_75t_L g13004 ( 
.A(n_12038),
.B(n_9773),
.Y(n_13004)
);

INVx1_ASAP7_75t_L g13005 ( 
.A(n_12484),
.Y(n_13005)
);

INVx1_ASAP7_75t_L g13006 ( 
.A(n_12553),
.Y(n_13006)
);

INVx3_ASAP7_75t_L g13007 ( 
.A(n_12606),
.Y(n_13007)
);

CKINVDCx20_ASAP7_75t_R g13008 ( 
.A(n_12174),
.Y(n_13008)
);

INVx2_ASAP7_75t_L g13009 ( 
.A(n_12441),
.Y(n_13009)
);

OR2x2_ASAP7_75t_L g13010 ( 
.A(n_11975),
.B(n_11026),
.Y(n_13010)
);

INVx1_ASAP7_75t_L g13011 ( 
.A(n_12655),
.Y(n_13011)
);

NAND2xp5_ASAP7_75t_L g13012 ( 
.A(n_11973),
.B(n_9999),
.Y(n_13012)
);

INVx2_ASAP7_75t_L g13013 ( 
.A(n_12302),
.Y(n_13013)
);

BUFx12f_ASAP7_75t_L g13014 ( 
.A(n_12086),
.Y(n_13014)
);

INVx2_ASAP7_75t_L g13015 ( 
.A(n_12302),
.Y(n_13015)
);

INVx11_ASAP7_75t_L g13016 ( 
.A(n_12086),
.Y(n_13016)
);

CKINVDCx5p33_ASAP7_75t_R g13017 ( 
.A(n_12238),
.Y(n_13017)
);

AND2x2_ASAP7_75t_L g13018 ( 
.A(n_12239),
.B(n_9773),
.Y(n_13018)
);

AND2x2_ASAP7_75t_L g13019 ( 
.A(n_12009),
.B(n_9827),
.Y(n_13019)
);

AND2x2_ASAP7_75t_L g13020 ( 
.A(n_12293),
.B(n_9827),
.Y(n_13020)
);

AND2x2_ASAP7_75t_L g13021 ( 
.A(n_12014),
.B(n_12024),
.Y(n_13021)
);

BUFx6f_ASAP7_75t_L g13022 ( 
.A(n_12606),
.Y(n_13022)
);

INVx1_ASAP7_75t_L g13023 ( 
.A(n_12678),
.Y(n_13023)
);

BUFx2_ASAP7_75t_L g13024 ( 
.A(n_12130),
.Y(n_13024)
);

AND2x2_ASAP7_75t_L g13025 ( 
.A(n_12034),
.B(n_9833),
.Y(n_13025)
);

BUFx2_ASAP7_75t_L g13026 ( 
.A(n_12184),
.Y(n_13026)
);

BUFx2_ASAP7_75t_L g13027 ( 
.A(n_12398),
.Y(n_13027)
);

AND2x2_ASAP7_75t_L g13028 ( 
.A(n_12042),
.B(n_9833),
.Y(n_13028)
);

AND2x2_ASAP7_75t_L g13029 ( 
.A(n_12085),
.B(n_9834),
.Y(n_13029)
);

OR2x2_ASAP7_75t_L g13030 ( 
.A(n_12632),
.B(n_11028),
.Y(n_13030)
);

INVx1_ASAP7_75t_L g13031 ( 
.A(n_12680),
.Y(n_13031)
);

INVxp67_ASAP7_75t_SL g13032 ( 
.A(n_11995),
.Y(n_13032)
);

AOI21xp5_ASAP7_75t_L g13033 ( 
.A1(n_12001),
.A2(n_11968),
.B(n_11980),
.Y(n_13033)
);

INVx1_ASAP7_75t_L g13034 ( 
.A(n_12415),
.Y(n_13034)
);

AND2x2_ASAP7_75t_L g13035 ( 
.A(n_12102),
.B(n_9834),
.Y(n_13035)
);

AND2x2_ASAP7_75t_L g13036 ( 
.A(n_12304),
.B(n_9852),
.Y(n_13036)
);

AND2x4_ASAP7_75t_L g13037 ( 
.A(n_12255),
.B(n_12046),
.Y(n_13037)
);

INVx3_ASAP7_75t_L g13038 ( 
.A(n_12590),
.Y(n_13038)
);

INVx1_ASAP7_75t_L g13039 ( 
.A(n_11984),
.Y(n_13039)
);

AND2x2_ASAP7_75t_L g13040 ( 
.A(n_12319),
.B(n_9852),
.Y(n_13040)
);

CKINVDCx20_ASAP7_75t_R g13041 ( 
.A(n_12127),
.Y(n_13041)
);

CKINVDCx6p67_ASAP7_75t_R g13042 ( 
.A(n_12185),
.Y(n_13042)
);

INVx1_ASAP7_75t_L g13043 ( 
.A(n_11993),
.Y(n_13043)
);

INVx1_ASAP7_75t_L g13044 ( 
.A(n_12015),
.Y(n_13044)
);

OR2x2_ASAP7_75t_L g13045 ( 
.A(n_12641),
.B(n_11032),
.Y(n_13045)
);

BUFx2_ASAP7_75t_L g13046 ( 
.A(n_12821),
.Y(n_13046)
);

AND2x2_ASAP7_75t_L g13047 ( 
.A(n_12123),
.B(n_9702),
.Y(n_13047)
);

INVx1_ASAP7_75t_L g13048 ( 
.A(n_12045),
.Y(n_13048)
);

NAND2xp5_ASAP7_75t_L g13049 ( 
.A(n_12381),
.B(n_10018),
.Y(n_13049)
);

INVx1_ASAP7_75t_L g13050 ( 
.A(n_12057),
.Y(n_13050)
);

INVx1_ASAP7_75t_L g13051 ( 
.A(n_12066),
.Y(n_13051)
);

NAND2xp5_ASAP7_75t_L g13052 ( 
.A(n_11985),
.B(n_10018),
.Y(n_13052)
);

INVx1_ASAP7_75t_L g13053 ( 
.A(n_12091),
.Y(n_13053)
);

AND2x2_ASAP7_75t_L g13054 ( 
.A(n_12139),
.B(n_9702),
.Y(n_13054)
);

BUFx2_ASAP7_75t_L g13055 ( 
.A(n_12011),
.Y(n_13055)
);

INVx2_ASAP7_75t_L g13056 ( 
.A(n_12302),
.Y(n_13056)
);

AND2x2_ASAP7_75t_L g13057 ( 
.A(n_12148),
.B(n_9374),
.Y(n_13057)
);

BUFx2_ASAP7_75t_SL g13058 ( 
.A(n_12614),
.Y(n_13058)
);

INVx2_ASAP7_75t_L g13059 ( 
.A(n_12326),
.Y(n_13059)
);

INVx2_ASAP7_75t_L g13060 ( 
.A(n_12326),
.Y(n_13060)
);

INVx2_ASAP7_75t_L g13061 ( 
.A(n_12326),
.Y(n_13061)
);

AO31x2_ASAP7_75t_L g13062 ( 
.A1(n_12129),
.A2(n_11253),
.A3(n_11254),
.B(n_11251),
.Y(n_13062)
);

OR2x2_ASAP7_75t_L g13063 ( 
.A(n_12518),
.B(n_11033),
.Y(n_13063)
);

INVx1_ASAP7_75t_L g13064 ( 
.A(n_11936),
.Y(n_13064)
);

INVx2_ASAP7_75t_L g13065 ( 
.A(n_12414),
.Y(n_13065)
);

HB1xp67_ASAP7_75t_L g13066 ( 
.A(n_12775),
.Y(n_13066)
);

AND2x2_ASAP7_75t_L g13067 ( 
.A(n_12171),
.B(n_9374),
.Y(n_13067)
);

NAND2xp5_ASAP7_75t_L g13068 ( 
.A(n_12144),
.B(n_10046),
.Y(n_13068)
);

NAND2xp5_ASAP7_75t_L g13069 ( 
.A(n_11963),
.B(n_10046),
.Y(n_13069)
);

AND2x2_ASAP7_75t_L g13070 ( 
.A(n_12191),
.B(n_10114),
.Y(n_13070)
);

OR2x2_ASAP7_75t_L g13071 ( 
.A(n_12050),
.B(n_12037),
.Y(n_13071)
);

HB1xp67_ASAP7_75t_L g13072 ( 
.A(n_11950),
.Y(n_13072)
);

INVx2_ASAP7_75t_L g13073 ( 
.A(n_12414),
.Y(n_13073)
);

INVx2_ASAP7_75t_L g13074 ( 
.A(n_12414),
.Y(n_13074)
);

AND2x2_ASAP7_75t_L g13075 ( 
.A(n_12198),
.B(n_10114),
.Y(n_13075)
);

INVx2_ASAP7_75t_L g13076 ( 
.A(n_12426),
.Y(n_13076)
);

AND2x2_ASAP7_75t_L g13077 ( 
.A(n_12221),
.B(n_10122),
.Y(n_13077)
);

AND2x2_ASAP7_75t_L g13078 ( 
.A(n_12231),
.B(n_12245),
.Y(n_13078)
);

INVx1_ASAP7_75t_L g13079 ( 
.A(n_11976),
.Y(n_13079)
);

INVx1_ASAP7_75t_L g13080 ( 
.A(n_11977),
.Y(n_13080)
);

OR2x2_ASAP7_75t_L g13081 ( 
.A(n_12137),
.B(n_11034),
.Y(n_13081)
);

INVx1_ASAP7_75t_L g13082 ( 
.A(n_12409),
.Y(n_13082)
);

AND2x2_ASAP7_75t_L g13083 ( 
.A(n_12256),
.B(n_10122),
.Y(n_13083)
);

AND2x2_ASAP7_75t_L g13084 ( 
.A(n_12282),
.B(n_10195),
.Y(n_13084)
);

BUFx2_ASAP7_75t_L g13085 ( 
.A(n_12786),
.Y(n_13085)
);

INVx1_ASAP7_75t_L g13086 ( 
.A(n_12413),
.Y(n_13086)
);

INVx1_ASAP7_75t_L g13087 ( 
.A(n_12419),
.Y(n_13087)
);

INVx1_ASAP7_75t_L g13088 ( 
.A(n_12420),
.Y(n_13088)
);

INVx1_ASAP7_75t_L g13089 ( 
.A(n_12432),
.Y(n_13089)
);

INVx1_ASAP7_75t_L g13090 ( 
.A(n_12447),
.Y(n_13090)
);

HB1xp67_ASAP7_75t_L g13091 ( 
.A(n_12452),
.Y(n_13091)
);

INVxp67_ASAP7_75t_L g13092 ( 
.A(n_12227),
.Y(n_13092)
);

HB1xp67_ASAP7_75t_L g13093 ( 
.A(n_12453),
.Y(n_13093)
);

INVx1_ASAP7_75t_L g13094 ( 
.A(n_12473),
.Y(n_13094)
);

INVxp67_ASAP7_75t_SL g13095 ( 
.A(n_11995),
.Y(n_13095)
);

HB1xp67_ASAP7_75t_L g13096 ( 
.A(n_12475),
.Y(n_13096)
);

INVx2_ASAP7_75t_L g13097 ( 
.A(n_12426),
.Y(n_13097)
);

INVx2_ASAP7_75t_L g13098 ( 
.A(n_12426),
.Y(n_13098)
);

NAND2xp5_ASAP7_75t_L g13099 ( 
.A(n_12021),
.B(n_10195),
.Y(n_13099)
);

INVx2_ASAP7_75t_L g13100 ( 
.A(n_12476),
.Y(n_13100)
);

NOR2x1_ASAP7_75t_L g13101 ( 
.A(n_12581),
.B(n_11688),
.Y(n_13101)
);

INVx2_ASAP7_75t_L g13102 ( 
.A(n_12476),
.Y(n_13102)
);

INVx2_ASAP7_75t_L g13103 ( 
.A(n_12476),
.Y(n_13103)
);

HB1xp67_ASAP7_75t_L g13104 ( 
.A(n_12492),
.Y(n_13104)
);

INVx1_ASAP7_75t_L g13105 ( 
.A(n_12493),
.Y(n_13105)
);

AND2x4_ASAP7_75t_L g13106 ( 
.A(n_12255),
.B(n_12046),
.Y(n_13106)
);

INVx2_ASAP7_75t_L g13107 ( 
.A(n_12039),
.Y(n_13107)
);

AND2x2_ASAP7_75t_L g13108 ( 
.A(n_12397),
.B(n_12402),
.Y(n_13108)
);

BUFx2_ASAP7_75t_L g13109 ( 
.A(n_12652),
.Y(n_13109)
);

INVx1_ASAP7_75t_L g13110 ( 
.A(n_12494),
.Y(n_13110)
);

INVx2_ASAP7_75t_L g13111 ( 
.A(n_12068),
.Y(n_13111)
);

INVx1_ASAP7_75t_L g13112 ( 
.A(n_12502),
.Y(n_13112)
);

AND2x2_ASAP7_75t_L g13113 ( 
.A(n_12406),
.B(n_10212),
.Y(n_13113)
);

INVxp67_ASAP7_75t_SL g13114 ( 
.A(n_11969),
.Y(n_13114)
);

INVx1_ASAP7_75t_L g13115 ( 
.A(n_12514),
.Y(n_13115)
);

INVx2_ASAP7_75t_L g13116 ( 
.A(n_12634),
.Y(n_13116)
);

INVx1_ASAP7_75t_L g13117 ( 
.A(n_12541),
.Y(n_13117)
);

BUFx3_ASAP7_75t_L g13118 ( 
.A(n_12216),
.Y(n_13118)
);

INVx2_ASAP7_75t_L g13119 ( 
.A(n_12634),
.Y(n_13119)
);

OR2x2_ASAP7_75t_L g13120 ( 
.A(n_12056),
.B(n_11039),
.Y(n_13120)
);

NOR2x1_ASAP7_75t_L g13121 ( 
.A(n_11942),
.B(n_11688),
.Y(n_13121)
);

HB1xp67_ASAP7_75t_L g13122 ( 
.A(n_12550),
.Y(n_13122)
);

INVx1_ASAP7_75t_L g13123 ( 
.A(n_12552),
.Y(n_13123)
);

INVx1_ASAP7_75t_L g13124 ( 
.A(n_12562),
.Y(n_13124)
);

INVx1_ASAP7_75t_L g13125 ( 
.A(n_12572),
.Y(n_13125)
);

INVx2_ASAP7_75t_L g13126 ( 
.A(n_12645),
.Y(n_13126)
);

INVx1_ASAP7_75t_L g13127 ( 
.A(n_12579),
.Y(n_13127)
);

HB1xp67_ASAP7_75t_L g13128 ( 
.A(n_12582),
.Y(n_13128)
);

NOR2xp33_ASAP7_75t_L g13129 ( 
.A(n_12025),
.B(n_7541),
.Y(n_13129)
);

INVx1_ASAP7_75t_L g13130 ( 
.A(n_12596),
.Y(n_13130)
);

NAND2xp5_ASAP7_75t_L g13131 ( 
.A(n_12211),
.B(n_10212),
.Y(n_13131)
);

AND2x4_ASAP7_75t_L g13132 ( 
.A(n_12069),
.B(n_11688),
.Y(n_13132)
);

INVx2_ASAP7_75t_L g13133 ( 
.A(n_12645),
.Y(n_13133)
);

AND2x2_ASAP7_75t_L g13134 ( 
.A(n_12070),
.B(n_10242),
.Y(n_13134)
);

AND2x2_ASAP7_75t_L g13135 ( 
.A(n_12362),
.B(n_12367),
.Y(n_13135)
);

INVx1_ASAP7_75t_L g13136 ( 
.A(n_12597),
.Y(n_13136)
);

HB1xp67_ASAP7_75t_L g13137 ( 
.A(n_12604),
.Y(n_13137)
);

NAND2xp5_ASAP7_75t_L g13138 ( 
.A(n_12036),
.B(n_10242),
.Y(n_13138)
);

AND2x2_ASAP7_75t_L g13139 ( 
.A(n_12377),
.B(n_10250),
.Y(n_13139)
);

AND2x2_ASAP7_75t_L g13140 ( 
.A(n_12390),
.B(n_10250),
.Y(n_13140)
);

OAI22xp5_ASAP7_75t_L g13141 ( 
.A1(n_11935),
.A2(n_9123),
.B1(n_9158),
.B2(n_9138),
.Y(n_13141)
);

AND2x2_ASAP7_75t_L g13142 ( 
.A(n_12321),
.B(n_10268),
.Y(n_13142)
);

AND2x2_ASAP7_75t_L g13143 ( 
.A(n_12345),
.B(n_10268),
.Y(n_13143)
);

AND2x2_ASAP7_75t_L g13144 ( 
.A(n_12297),
.B(n_10307),
.Y(n_13144)
);

INVx1_ASAP7_75t_L g13145 ( 
.A(n_12612),
.Y(n_13145)
);

AND2x2_ASAP7_75t_L g13146 ( 
.A(n_11966),
.B(n_12103),
.Y(n_13146)
);

AND2x2_ASAP7_75t_L g13147 ( 
.A(n_11978),
.B(n_10307),
.Y(n_13147)
);

INVx1_ASAP7_75t_L g13148 ( 
.A(n_12620),
.Y(n_13148)
);

NAND2xp5_ASAP7_75t_L g13149 ( 
.A(n_12126),
.B(n_12202),
.Y(n_13149)
);

INVx1_ASAP7_75t_L g13150 ( 
.A(n_12637),
.Y(n_13150)
);

INVx1_ASAP7_75t_L g13151 ( 
.A(n_12665),
.Y(n_13151)
);

INVx2_ASAP7_75t_SL g13152 ( 
.A(n_12185),
.Y(n_13152)
);

INVx2_ASAP7_75t_L g13153 ( 
.A(n_12500),
.Y(n_13153)
);

NOR2x1p5_ASAP7_75t_L g13154 ( 
.A(n_12244),
.B(n_7543),
.Y(n_13154)
);

INVx1_ASAP7_75t_L g13155 ( 
.A(n_12672),
.Y(n_13155)
);

INVx2_ASAP7_75t_L g13156 ( 
.A(n_12539),
.Y(n_13156)
);

NAND2xp5_ASAP7_75t_L g13157 ( 
.A(n_12040),
.B(n_10344),
.Y(n_13157)
);

INVx1_ASAP7_75t_L g13158 ( 
.A(n_12707),
.Y(n_13158)
);

AND2x2_ASAP7_75t_L g13159 ( 
.A(n_11992),
.B(n_10344),
.Y(n_13159)
);

INVxp67_ASAP7_75t_SL g13160 ( 
.A(n_12192),
.Y(n_13160)
);

HB1xp67_ASAP7_75t_L g13161 ( 
.A(n_12711),
.Y(n_13161)
);

HB1xp67_ASAP7_75t_L g13162 ( 
.A(n_12721),
.Y(n_13162)
);

BUFx2_ASAP7_75t_L g13163 ( 
.A(n_12712),
.Y(n_13163)
);

INVx1_ASAP7_75t_L g13164 ( 
.A(n_12094),
.Y(n_13164)
);

INVx2_ASAP7_75t_SL g13165 ( 
.A(n_12225),
.Y(n_13165)
);

INVx4_ASAP7_75t_L g13166 ( 
.A(n_11987),
.Y(n_13166)
);

NAND2xp5_ASAP7_75t_L g13167 ( 
.A(n_12136),
.B(n_10366),
.Y(n_13167)
);

INVx1_ASAP7_75t_L g13168 ( 
.A(n_12113),
.Y(n_13168)
);

AND2x2_ASAP7_75t_L g13169 ( 
.A(n_12006),
.B(n_10366),
.Y(n_13169)
);

HB1xp67_ASAP7_75t_L g13170 ( 
.A(n_12914),
.Y(n_13170)
);

AND2x2_ASAP7_75t_L g13171 ( 
.A(n_12535),
.B(n_10401),
.Y(n_13171)
);

AND2x2_ASAP7_75t_L g13172 ( 
.A(n_12354),
.B(n_10401),
.Y(n_13172)
);

INVx2_ASAP7_75t_L g13173 ( 
.A(n_12795),
.Y(n_13173)
);

NAND2xp5_ASAP7_75t_L g13174 ( 
.A(n_11944),
.B(n_10405),
.Y(n_13174)
);

HB1xp67_ASAP7_75t_L g13175 ( 
.A(n_12147),
.Y(n_13175)
);

INVx1_ASAP7_75t_L g13176 ( 
.A(n_12151),
.Y(n_13176)
);

INVx2_ASAP7_75t_L g13177 ( 
.A(n_12795),
.Y(n_13177)
);

AND2x2_ASAP7_75t_L g13178 ( 
.A(n_12629),
.B(n_10405),
.Y(n_13178)
);

NOR2xp33_ASAP7_75t_L g13179 ( 
.A(n_12530),
.B(n_8720),
.Y(n_13179)
);

INVx2_ASAP7_75t_L g13180 ( 
.A(n_12385),
.Y(n_13180)
);

NAND2xp5_ASAP7_75t_L g13181 ( 
.A(n_12509),
.B(n_10497),
.Y(n_13181)
);

BUFx2_ASAP7_75t_L g13182 ( 
.A(n_12069),
.Y(n_13182)
);

INVx2_ASAP7_75t_SL g13183 ( 
.A(n_12225),
.Y(n_13183)
);

INVx1_ASAP7_75t_L g13184 ( 
.A(n_12180),
.Y(n_13184)
);

INVxp67_ASAP7_75t_L g13185 ( 
.A(n_12154),
.Y(n_13185)
);

AND2x2_ASAP7_75t_L g13186 ( 
.A(n_11981),
.B(n_10497),
.Y(n_13186)
);

INVx2_ASAP7_75t_L g13187 ( 
.A(n_12385),
.Y(n_13187)
);

AND2x2_ASAP7_75t_SL g13188 ( 
.A(n_11933),
.B(n_8965),
.Y(n_13188)
);

BUFx2_ASAP7_75t_L g13189 ( 
.A(n_12114),
.Y(n_13189)
);

INVx1_ASAP7_75t_L g13190 ( 
.A(n_12214),
.Y(n_13190)
);

NAND2xp5_ASAP7_75t_L g13191 ( 
.A(n_11996),
.B(n_10518),
.Y(n_13191)
);

AND2x2_ASAP7_75t_L g13192 ( 
.A(n_11981),
.B(n_10518),
.Y(n_13192)
);

INVx1_ASAP7_75t_L g13193 ( 
.A(n_12275),
.Y(n_13193)
);

INVx1_ASAP7_75t_L g13194 ( 
.A(n_12285),
.Y(n_13194)
);

INVx2_ASAP7_75t_L g13195 ( 
.A(n_12405),
.Y(n_13195)
);

AND2x2_ASAP7_75t_L g13196 ( 
.A(n_12369),
.B(n_10555),
.Y(n_13196)
);

INVx3_ASAP7_75t_L g13197 ( 
.A(n_12114),
.Y(n_13197)
);

HB1xp67_ASAP7_75t_L g13198 ( 
.A(n_12286),
.Y(n_13198)
);

INVx2_ASAP7_75t_L g13199 ( 
.A(n_12405),
.Y(n_13199)
);

BUFx2_ASAP7_75t_L g13200 ( 
.A(n_12698),
.Y(n_13200)
);

INVx4_ASAP7_75t_SL g13201 ( 
.A(n_11987),
.Y(n_13201)
);

OR2x2_ASAP7_75t_L g13202 ( 
.A(n_12061),
.B(n_11050),
.Y(n_13202)
);

INVx4_ASAP7_75t_L g13203 ( 
.A(n_11987),
.Y(n_13203)
);

INVx2_ASAP7_75t_L g13204 ( 
.A(n_12416),
.Y(n_13204)
);

INVx2_ASAP7_75t_L g13205 ( 
.A(n_12416),
.Y(n_13205)
);

AND2x2_ASAP7_75t_L g13206 ( 
.A(n_12097),
.B(n_10555),
.Y(n_13206)
);

BUFx2_ASAP7_75t_L g13207 ( 
.A(n_12713),
.Y(n_13207)
);

INVxp67_ASAP7_75t_SL g13208 ( 
.A(n_12175),
.Y(n_13208)
);

HB1xp67_ASAP7_75t_L g13209 ( 
.A(n_12287),
.Y(n_13209)
);

HB1xp67_ASAP7_75t_L g13210 ( 
.A(n_12290),
.Y(n_13210)
);

OR2x2_ASAP7_75t_L g13211 ( 
.A(n_12128),
.B(n_11060),
.Y(n_13211)
);

AND2x4_ASAP7_75t_L g13212 ( 
.A(n_12417),
.B(n_11694),
.Y(n_13212)
);

INVx1_ASAP7_75t_L g13213 ( 
.A(n_12296),
.Y(n_13213)
);

INVx2_ASAP7_75t_L g13214 ( 
.A(n_12664),
.Y(n_13214)
);

OR2x2_ASAP7_75t_L g13215 ( 
.A(n_12200),
.B(n_11062),
.Y(n_13215)
);

INVx2_ASAP7_75t_L g13216 ( 
.A(n_12664),
.Y(n_13216)
);

INVx1_ASAP7_75t_L g13217 ( 
.A(n_12311),
.Y(n_13217)
);

INVx1_ASAP7_75t_L g13218 ( 
.A(n_12314),
.Y(n_13218)
);

INVx1_ASAP7_75t_L g13219 ( 
.A(n_12325),
.Y(n_13219)
);

OR2x2_ASAP7_75t_L g13220 ( 
.A(n_12234),
.B(n_11064),
.Y(n_13220)
);

HB1xp67_ASAP7_75t_L g13221 ( 
.A(n_12335),
.Y(n_13221)
);

INVx2_ASAP7_75t_L g13222 ( 
.A(n_12668),
.Y(n_13222)
);

AND2x2_ASAP7_75t_L g13223 ( 
.A(n_12071),
.B(n_10561),
.Y(n_13223)
);

INVx2_ASAP7_75t_L g13224 ( 
.A(n_12668),
.Y(n_13224)
);

OR2x2_ASAP7_75t_L g13225 ( 
.A(n_12525),
.B(n_11070),
.Y(n_13225)
);

AND2x2_ASAP7_75t_L g13226 ( 
.A(n_12073),
.B(n_10561),
.Y(n_13226)
);

AND2x4_ASAP7_75t_SL g13227 ( 
.A(n_12152),
.B(n_7763),
.Y(n_13227)
);

AND2x2_ASAP7_75t_L g13228 ( 
.A(n_12702),
.B(n_10569),
.Y(n_13228)
);

INVx2_ASAP7_75t_L g13229 ( 
.A(n_12683),
.Y(n_13229)
);

OR2x2_ASAP7_75t_L g13230 ( 
.A(n_12008),
.B(n_11072),
.Y(n_13230)
);

INVx1_ASAP7_75t_L g13231 ( 
.A(n_12338),
.Y(n_13231)
);

INVx1_ASAP7_75t_L g13232 ( 
.A(n_12341),
.Y(n_13232)
);

AND2x2_ASAP7_75t_L g13233 ( 
.A(n_12706),
.B(n_10569),
.Y(n_13233)
);

INVx3_ASAP7_75t_L g13234 ( 
.A(n_12766),
.Y(n_13234)
);

OR2x2_ASAP7_75t_L g13235 ( 
.A(n_12049),
.B(n_11075),
.Y(n_13235)
);

INVx2_ASAP7_75t_L g13236 ( 
.A(n_12683),
.Y(n_13236)
);

OR2x2_ASAP7_75t_L g13237 ( 
.A(n_12196),
.B(n_11082),
.Y(n_13237)
);

OR2x2_ASAP7_75t_L g13238 ( 
.A(n_12240),
.B(n_11083),
.Y(n_13238)
);

AND2x2_ASAP7_75t_L g13239 ( 
.A(n_12727),
.B(n_10618),
.Y(n_13239)
);

AND2x2_ASAP7_75t_L g13240 ( 
.A(n_12865),
.B(n_10618),
.Y(n_13240)
);

INVx2_ASAP7_75t_L g13241 ( 
.A(n_12131),
.Y(n_13241)
);

INVx1_ASAP7_75t_L g13242 ( 
.A(n_12347),
.Y(n_13242)
);

AND2x2_ASAP7_75t_L g13243 ( 
.A(n_12876),
.B(n_10672),
.Y(n_13243)
);

INVx2_ASAP7_75t_L g13244 ( 
.A(n_12131),
.Y(n_13244)
);

HB1xp67_ASAP7_75t_L g13245 ( 
.A(n_12360),
.Y(n_13245)
);

INVx2_ASAP7_75t_L g13246 ( 
.A(n_12131),
.Y(n_13246)
);

AND2x2_ASAP7_75t_L g13247 ( 
.A(n_12585),
.B(n_10672),
.Y(n_13247)
);

AND2x2_ASAP7_75t_L g13248 ( 
.A(n_12723),
.B(n_12257),
.Y(n_13248)
);

INVx2_ASAP7_75t_L g13249 ( 
.A(n_12850),
.Y(n_13249)
);

NAND2xp5_ASAP7_75t_L g13250 ( 
.A(n_12169),
.B(n_10702),
.Y(n_13250)
);

INVx2_ASAP7_75t_SL g13251 ( 
.A(n_12730),
.Y(n_13251)
);

INVxp67_ASAP7_75t_L g13252 ( 
.A(n_12160),
.Y(n_13252)
);

AND2x4_ASAP7_75t_L g13253 ( 
.A(n_12417),
.B(n_11694),
.Y(n_13253)
);

AND2x2_ASAP7_75t_L g13254 ( 
.A(n_12723),
.B(n_10702),
.Y(n_13254)
);

AND2x4_ASAP7_75t_L g13255 ( 
.A(n_12713),
.B(n_11694),
.Y(n_13255)
);

AND2x4_ASAP7_75t_L g13256 ( 
.A(n_12734),
.B(n_11727),
.Y(n_13256)
);

HB1xp67_ASAP7_75t_L g13257 ( 
.A(n_12370),
.Y(n_13257)
);

BUFx2_ASAP7_75t_L g13258 ( 
.A(n_12734),
.Y(n_13258)
);

INVx1_ASAP7_75t_L g13259 ( 
.A(n_12720),
.Y(n_13259)
);

AND2x2_ASAP7_75t_L g13260 ( 
.A(n_12262),
.B(n_10712),
.Y(n_13260)
);

AND2x2_ASAP7_75t_L g13261 ( 
.A(n_12732),
.B(n_10712),
.Y(n_13261)
);

INVx4_ASAP7_75t_L g13262 ( 
.A(n_12407),
.Y(n_13262)
);

AND2x2_ASAP7_75t_L g13263 ( 
.A(n_12644),
.B(n_9960),
.Y(n_13263)
);

BUFx6f_ASAP7_75t_L g13264 ( 
.A(n_12244),
.Y(n_13264)
);

INVx1_ASAP7_75t_L g13265 ( 
.A(n_12736),
.Y(n_13265)
);

NAND2xp5_ASAP7_75t_SL g13266 ( 
.A(n_11940),
.B(n_8881),
.Y(n_13266)
);

OR2x2_ASAP7_75t_L g13267 ( 
.A(n_12241),
.B(n_11085),
.Y(n_13267)
);

OR2x2_ASAP7_75t_L g13268 ( 
.A(n_12294),
.B(n_11093),
.Y(n_13268)
);

INVx1_ASAP7_75t_L g13269 ( 
.A(n_12764),
.Y(n_13269)
);

HB1xp67_ASAP7_75t_L g13270 ( 
.A(n_12753),
.Y(n_13270)
);

HB1xp67_ASAP7_75t_L g13271 ( 
.A(n_12760),
.Y(n_13271)
);

INVx1_ASAP7_75t_L g13272 ( 
.A(n_12765),
.Y(n_13272)
);

INVx2_ASAP7_75t_L g13273 ( 
.A(n_12850),
.Y(n_13273)
);

AO21x2_ASAP7_75t_L g13274 ( 
.A1(n_12646),
.A2(n_11100),
.B(n_11098),
.Y(n_13274)
);

AND2x4_ASAP7_75t_L g13275 ( 
.A(n_12648),
.B(n_11727),
.Y(n_13275)
);

AND2x2_ASAP7_75t_L g13276 ( 
.A(n_12651),
.B(n_9960),
.Y(n_13276)
);

INVx2_ASAP7_75t_L g13277 ( 
.A(n_12859),
.Y(n_13277)
);

HB1xp67_ASAP7_75t_L g13278 ( 
.A(n_12778),
.Y(n_13278)
);

INVx2_ASAP7_75t_L g13279 ( 
.A(n_12766),
.Y(n_13279)
);

INVx3_ASAP7_75t_L g13280 ( 
.A(n_12674),
.Y(n_13280)
);

INVx2_ASAP7_75t_L g13281 ( 
.A(n_12407),
.Y(n_13281)
);

OR2x2_ASAP7_75t_L g13282 ( 
.A(n_12310),
.B(n_11104),
.Y(n_13282)
);

AND2x2_ASAP7_75t_L g13283 ( 
.A(n_12663),
.B(n_9138),
.Y(n_13283)
);

BUFx3_ASAP7_75t_L g13284 ( 
.A(n_12315),
.Y(n_13284)
);

INVx1_ASAP7_75t_L g13285 ( 
.A(n_12780),
.Y(n_13285)
);

BUFx6f_ASAP7_75t_L g13286 ( 
.A(n_12283),
.Y(n_13286)
);

HB1xp67_ASAP7_75t_L g13287 ( 
.A(n_12781),
.Y(n_13287)
);

INVx1_ASAP7_75t_L g13288 ( 
.A(n_12784),
.Y(n_13288)
);

INVx2_ASAP7_75t_L g13289 ( 
.A(n_12134),
.Y(n_13289)
);

INVx2_ASAP7_75t_SL g13290 ( 
.A(n_12059),
.Y(n_13290)
);

AND2x2_ASAP7_75t_L g13291 ( 
.A(n_12673),
.B(n_9138),
.Y(n_13291)
);

AND2x2_ASAP7_75t_L g13292 ( 
.A(n_12808),
.B(n_9158),
.Y(n_13292)
);

AND2x4_ASAP7_75t_L g13293 ( 
.A(n_12650),
.B(n_11727),
.Y(n_13293)
);

INVx1_ASAP7_75t_L g13294 ( 
.A(n_12785),
.Y(n_13294)
);

INVx2_ASAP7_75t_L g13295 ( 
.A(n_12134),
.Y(n_13295)
);

INVxp67_ASAP7_75t_L g13296 ( 
.A(n_12769),
.Y(n_13296)
);

INVx1_ASAP7_75t_L g13297 ( 
.A(n_12823),
.Y(n_13297)
);

AOI22xp33_ASAP7_75t_L g13298 ( 
.A1(n_12027),
.A2(n_8699),
.B1(n_8665),
.B2(n_8554),
.Y(n_13298)
);

INVx2_ASAP7_75t_L g13299 ( 
.A(n_12135),
.Y(n_13299)
);

AND2x2_ASAP7_75t_L g13300 ( 
.A(n_12829),
.B(n_9158),
.Y(n_13300)
);

INVx1_ASAP7_75t_L g13301 ( 
.A(n_12888),
.Y(n_13301)
);

BUFx3_ASAP7_75t_L g13302 ( 
.A(n_12434),
.Y(n_13302)
);

AND2x2_ASAP7_75t_L g13303 ( 
.A(n_12350),
.B(n_12064),
.Y(n_13303)
);

INVx1_ASAP7_75t_L g13304 ( 
.A(n_12898),
.Y(n_13304)
);

OR2x2_ASAP7_75t_L g13305 ( 
.A(n_12053),
.B(n_11106),
.Y(n_13305)
);

INVx2_ASAP7_75t_L g13306 ( 
.A(n_12135),
.Y(n_13306)
);

BUFx6f_ASAP7_75t_L g13307 ( 
.A(n_12095),
.Y(n_13307)
);

INVx1_ASAP7_75t_L g13308 ( 
.A(n_12899),
.Y(n_13308)
);

INVx1_ASAP7_75t_L g13309 ( 
.A(n_12904),
.Y(n_13309)
);

AND2x2_ASAP7_75t_L g13310 ( 
.A(n_12186),
.B(n_12333),
.Y(n_13310)
);

AND2x2_ASAP7_75t_L g13311 ( 
.A(n_12340),
.B(n_12122),
.Y(n_13311)
);

INVx1_ASAP7_75t_L g13312 ( 
.A(n_12906),
.Y(n_13312)
);

AND2x2_ASAP7_75t_L g13313 ( 
.A(n_12316),
.B(n_9174),
.Y(n_13313)
);

OR2x2_ASAP7_75t_L g13314 ( 
.A(n_12055),
.B(n_11109),
.Y(n_13314)
);

INVx1_ASAP7_75t_L g13315 ( 
.A(n_12913),
.Y(n_13315)
);

INVx1_ASAP7_75t_L g13316 ( 
.A(n_12922),
.Y(n_13316)
);

AND2x2_ASAP7_75t_L g13317 ( 
.A(n_12538),
.B(n_9174),
.Y(n_13317)
);

AOI22xp33_ASAP7_75t_L g13318 ( 
.A1(n_11971),
.A2(n_8699),
.B1(n_8665),
.B2(n_8554),
.Y(n_13318)
);

OR2x2_ASAP7_75t_L g13319 ( 
.A(n_12560),
.B(n_11112),
.Y(n_13319)
);

INVx2_ASAP7_75t_L g13320 ( 
.A(n_12161),
.Y(n_13320)
);

AND2x2_ASAP7_75t_L g13321 ( 
.A(n_12352),
.B(n_9174),
.Y(n_13321)
);

NAND2xp5_ASAP7_75t_L g13322 ( 
.A(n_11954),
.B(n_11113),
.Y(n_13322)
);

INVx5_ASAP7_75t_L g13323 ( 
.A(n_12280),
.Y(n_13323)
);

AND2x4_ASAP7_75t_L g13324 ( 
.A(n_12694),
.B(n_11779),
.Y(n_13324)
);

OR2x2_ASAP7_75t_L g13325 ( 
.A(n_12173),
.B(n_11115),
.Y(n_13325)
);

AND2x4_ASAP7_75t_SL g13326 ( 
.A(n_12547),
.B(n_7763),
.Y(n_13326)
);

OAI22xp5_ASAP7_75t_SL g13327 ( 
.A1(n_11932),
.A2(n_8965),
.B1(n_9074),
.B2(n_8881),
.Y(n_13327)
);

NOR2x1_ASAP7_75t_L g13328 ( 
.A(n_12016),
.B(n_11779),
.Y(n_13328)
);

AND2x2_ASAP7_75t_L g13329 ( 
.A(n_12357),
.B(n_9186),
.Y(n_13329)
);

INVx1_ASAP7_75t_SL g13330 ( 
.A(n_12224),
.Y(n_13330)
);

BUFx6f_ASAP7_75t_L g13331 ( 
.A(n_11974),
.Y(n_13331)
);

INVx3_ASAP7_75t_L g13332 ( 
.A(n_12674),
.Y(n_13332)
);

AND2x2_ASAP7_75t_L g13333 ( 
.A(n_12359),
.B(n_9186),
.Y(n_13333)
);

OR2x2_ASAP7_75t_L g13334 ( 
.A(n_12018),
.B(n_11116),
.Y(n_13334)
);

NAND2xp5_ASAP7_75t_L g13335 ( 
.A(n_12155),
.B(n_11118),
.Y(n_13335)
);

NAND2xp5_ASAP7_75t_L g13336 ( 
.A(n_12342),
.B(n_11120),
.Y(n_13336)
);

AND2x2_ASAP7_75t_L g13337 ( 
.A(n_12361),
.B(n_9186),
.Y(n_13337)
);

INVx1_ASAP7_75t_L g13338 ( 
.A(n_12926),
.Y(n_13338)
);

INVx1_ASAP7_75t_L g13339 ( 
.A(n_12933),
.Y(n_13339)
);

AND2x2_ASAP7_75t_L g13340 ( 
.A(n_12368),
.B(n_9196),
.Y(n_13340)
);

AND2x2_ASAP7_75t_L g13341 ( 
.A(n_12373),
.B(n_9196),
.Y(n_13341)
);

INVx1_ASAP7_75t_SL g13342 ( 
.A(n_12635),
.Y(n_13342)
);

INVx1_ASAP7_75t_L g13343 ( 
.A(n_12934),
.Y(n_13343)
);

AND2x2_ASAP7_75t_L g13344 ( 
.A(n_12376),
.B(n_12383),
.Y(n_13344)
);

AND2x4_ASAP7_75t_SL g13345 ( 
.A(n_12280),
.B(n_7763),
.Y(n_13345)
);

OR2x2_ASAP7_75t_L g13346 ( 
.A(n_11959),
.B(n_11125),
.Y(n_13346)
);

INVx1_ASAP7_75t_L g13347 ( 
.A(n_12938),
.Y(n_13347)
);

INVx1_ASAP7_75t_L g13348 ( 
.A(n_12945),
.Y(n_13348)
);

INVx2_ASAP7_75t_R g13349 ( 
.A(n_12016),
.Y(n_13349)
);

AND2x2_ASAP7_75t_L g13350 ( 
.A(n_12386),
.B(n_9196),
.Y(n_13350)
);

INVx1_ASAP7_75t_L g13351 ( 
.A(n_12950),
.Y(n_13351)
);

BUFx2_ASAP7_75t_L g13352 ( 
.A(n_11994),
.Y(n_13352)
);

NAND2xp5_ASAP7_75t_L g13353 ( 
.A(n_12455),
.B(n_11129),
.Y(n_13353)
);

INVx1_ASAP7_75t_L g13354 ( 
.A(n_12958),
.Y(n_13354)
);

AND2x2_ASAP7_75t_L g13355 ( 
.A(n_12307),
.B(n_9220),
.Y(n_13355)
);

NOR2x1_ASAP7_75t_L g13356 ( 
.A(n_12063),
.B(n_11779),
.Y(n_13356)
);

INVx2_ASAP7_75t_L g13357 ( 
.A(n_12161),
.Y(n_13357)
);

INVx1_ASAP7_75t_L g13358 ( 
.A(n_12882),
.Y(n_13358)
);

AND2x2_ASAP7_75t_L g13359 ( 
.A(n_12456),
.B(n_9220),
.Y(n_13359)
);

INVx1_ASAP7_75t_SL g13360 ( 
.A(n_12630),
.Y(n_13360)
);

BUFx3_ASAP7_75t_L g13361 ( 
.A(n_12639),
.Y(n_13361)
);

INVx2_ASAP7_75t_L g13362 ( 
.A(n_12735),
.Y(n_13362)
);

AND2x2_ASAP7_75t_L g13363 ( 
.A(n_12457),
.B(n_12479),
.Y(n_13363)
);

INVx2_ASAP7_75t_L g13364 ( 
.A(n_12735),
.Y(n_13364)
);

AND2x4_ASAP7_75t_L g13365 ( 
.A(n_12428),
.B(n_11784),
.Y(n_13365)
);

INVx1_ASAP7_75t_L g13366 ( 
.A(n_12882),
.Y(n_13366)
);

INVx1_ASAP7_75t_L g13367 ( 
.A(n_12408),
.Y(n_13367)
);

AO31x2_ASAP7_75t_L g13368 ( 
.A1(n_11989),
.A2(n_11339),
.A3(n_11340),
.B(n_11337),
.Y(n_13368)
);

INVx2_ASAP7_75t_L g13369 ( 
.A(n_12835),
.Y(n_13369)
);

AND2x2_ASAP7_75t_L g13370 ( 
.A(n_12488),
.B(n_12489),
.Y(n_13370)
);

INVx3_ASAP7_75t_L g13371 ( 
.A(n_12438),
.Y(n_13371)
);

AND2x4_ASAP7_75t_L g13372 ( 
.A(n_12428),
.B(n_11784),
.Y(n_13372)
);

INVx2_ASAP7_75t_L g13373 ( 
.A(n_12835),
.Y(n_13373)
);

AOI21xp33_ASAP7_75t_L g13374 ( 
.A1(n_11957),
.A2(n_11889),
.B(n_11865),
.Y(n_13374)
);

INVx1_ASAP7_75t_L g13375 ( 
.A(n_12953),
.Y(n_13375)
);

NAND2xp5_ASAP7_75t_L g13376 ( 
.A(n_12005),
.B(n_12430),
.Y(n_13376)
);

INVx2_ASAP7_75t_SL g13377 ( 
.A(n_12699),
.Y(n_13377)
);

INVx2_ASAP7_75t_SL g13378 ( 
.A(n_12699),
.Y(n_13378)
);

INVx2_ASAP7_75t_L g13379 ( 
.A(n_12835),
.Y(n_13379)
);

INVx1_ASAP7_75t_L g13380 ( 
.A(n_12613),
.Y(n_13380)
);

AND2x2_ASAP7_75t_L g13381 ( 
.A(n_12495),
.B(n_12506),
.Y(n_13381)
);

INVx2_ASAP7_75t_L g13382 ( 
.A(n_12835),
.Y(n_13382)
);

NAND2xp5_ASAP7_75t_L g13383 ( 
.A(n_11956),
.B(n_11136),
.Y(n_13383)
);

INVx1_ASAP7_75t_L g13384 ( 
.A(n_12803),
.Y(n_13384)
);

NOR3xp33_ASAP7_75t_SL g13385 ( 
.A(n_12157),
.B(n_12172),
.C(n_12733),
.Y(n_13385)
);

AND2x4_ASAP7_75t_L g13386 ( 
.A(n_11994),
.B(n_11784),
.Y(n_13386)
);

INVx1_ASAP7_75t_L g13387 ( 
.A(n_12806),
.Y(n_13387)
);

BUFx2_ASAP7_75t_L g13388 ( 
.A(n_12007),
.Y(n_13388)
);

INVx4_ASAP7_75t_L g13389 ( 
.A(n_12098),
.Y(n_13389)
);

INVxp67_ASAP7_75t_L g13390 ( 
.A(n_12497),
.Y(n_13390)
);

NAND2xp5_ASAP7_75t_L g13391 ( 
.A(n_11952),
.B(n_11137),
.Y(n_13391)
);

AND2x2_ASAP7_75t_L g13392 ( 
.A(n_12507),
.B(n_9220),
.Y(n_13392)
);

INVx2_ASAP7_75t_L g13393 ( 
.A(n_12835),
.Y(n_13393)
);

INVx2_ASAP7_75t_L g13394 ( 
.A(n_12847),
.Y(n_13394)
);

AND2x2_ASAP7_75t_L g13395 ( 
.A(n_12543),
.B(n_8898),
.Y(n_13395)
);

OR2x2_ASAP7_75t_L g13396 ( 
.A(n_11938),
.B(n_11142),
.Y(n_13396)
);

AND2x2_ASAP7_75t_L g13397 ( 
.A(n_12615),
.B(n_12580),
.Y(n_13397)
);

INVx1_ASAP7_75t_L g13398 ( 
.A(n_12828),
.Y(n_13398)
);

AND2x2_ASAP7_75t_L g13399 ( 
.A(n_12936),
.B(n_8898),
.Y(n_13399)
);

INVx1_ASAP7_75t_L g13400 ( 
.A(n_12836),
.Y(n_13400)
);

INVx2_ASAP7_75t_L g13401 ( 
.A(n_12847),
.Y(n_13401)
);

AND2x4_ASAP7_75t_L g13402 ( 
.A(n_12007),
.B(n_11849),
.Y(n_13402)
);

INVx1_ASAP7_75t_L g13403 ( 
.A(n_12834),
.Y(n_13403)
);

AND2x2_ASAP7_75t_L g13404 ( 
.A(n_12305),
.B(n_8898),
.Y(n_13404)
);

INVx1_ASAP7_75t_SL g13405 ( 
.A(n_12715),
.Y(n_13405)
);

INVx1_ASAP7_75t_L g13406 ( 
.A(n_12895),
.Y(n_13406)
);

AND2x4_ASAP7_75t_SL g13407 ( 
.A(n_12697),
.B(n_8965),
.Y(n_13407)
);

INVx1_ASAP7_75t_L g13408 ( 
.A(n_12909),
.Y(n_13408)
);

INVxp67_ASAP7_75t_L g13409 ( 
.A(n_12268),
.Y(n_13409)
);

BUFx2_ASAP7_75t_SL g13410 ( 
.A(n_12471),
.Y(n_13410)
);

AND2x2_ASAP7_75t_L g13411 ( 
.A(n_12125),
.B(n_8931),
.Y(n_13411)
);

INVx2_ASAP7_75t_L g13412 ( 
.A(n_12847),
.Y(n_13412)
);

INVx1_ASAP7_75t_L g13413 ( 
.A(n_12911),
.Y(n_13413)
);

HB1xp67_ASAP7_75t_L g13414 ( 
.A(n_12820),
.Y(n_13414)
);

AND2x4_ASAP7_75t_L g13415 ( 
.A(n_12117),
.B(n_11849),
.Y(n_13415)
);

INVx1_ASAP7_75t_L g13416 ( 
.A(n_12561),
.Y(n_13416)
);

INVx2_ASAP7_75t_L g13417 ( 
.A(n_12847),
.Y(n_13417)
);

AOI22xp33_ASAP7_75t_L g13418 ( 
.A1(n_12356),
.A2(n_8699),
.B1(n_8665),
.B2(n_8554),
.Y(n_13418)
);

OR2x2_ASAP7_75t_L g13419 ( 
.A(n_12065),
.B(n_11146),
.Y(n_13419)
);

INVx1_ASAP7_75t_SL g13420 ( 
.A(n_12098),
.Y(n_13420)
);

AND2x2_ASAP7_75t_L g13421 ( 
.A(n_12132),
.B(n_8931),
.Y(n_13421)
);

AND2x2_ASAP7_75t_L g13422 ( 
.A(n_12078),
.B(n_8931),
.Y(n_13422)
);

BUFx2_ASAP7_75t_L g13423 ( 
.A(n_12438),
.Y(n_13423)
);

INVx3_ASAP7_75t_L g13424 ( 
.A(n_12439),
.Y(n_13424)
);

INVx1_ASAP7_75t_L g13425 ( 
.A(n_12587),
.Y(n_13425)
);

AND2x2_ASAP7_75t_L g13426 ( 
.A(n_12312),
.B(n_8935),
.Y(n_13426)
);

AND2x2_ASAP7_75t_L g13427 ( 
.A(n_12312),
.B(n_8935),
.Y(n_13427)
);

INVx2_ASAP7_75t_L g13428 ( 
.A(n_12847),
.Y(n_13428)
);

INVx1_ASAP7_75t_L g13429 ( 
.A(n_12877),
.Y(n_13429)
);

INVx2_ASAP7_75t_L g13430 ( 
.A(n_12799),
.Y(n_13430)
);

INVx2_ASAP7_75t_L g13431 ( 
.A(n_12799),
.Y(n_13431)
);

INVx2_ASAP7_75t_L g13432 ( 
.A(n_12251),
.Y(n_13432)
);

AND2x2_ASAP7_75t_L g13433 ( 
.A(n_12704),
.B(n_8935),
.Y(n_13433)
);

INVx4_ASAP7_75t_L g13434 ( 
.A(n_12355),
.Y(n_13434)
);

INVx1_ASAP7_75t_L g13435 ( 
.A(n_12857),
.Y(n_13435)
);

AND2x4_ASAP7_75t_L g13436 ( 
.A(n_12117),
.B(n_11849),
.Y(n_13436)
);

AND2x2_ASAP7_75t_L g13437 ( 
.A(n_12449),
.B(n_8960),
.Y(n_13437)
);

AND2x2_ASAP7_75t_L g13438 ( 
.A(n_12099),
.B(n_8960),
.Y(n_13438)
);

INVx2_ASAP7_75t_L g13439 ( 
.A(n_12145),
.Y(n_13439)
);

BUFx2_ASAP7_75t_L g13440 ( 
.A(n_12439),
.Y(n_13440)
);

INVx2_ASAP7_75t_L g13441 ( 
.A(n_12167),
.Y(n_13441)
);

NAND2xp5_ASAP7_75t_L g13442 ( 
.A(n_11961),
.B(n_11148),
.Y(n_13442)
);

INVx4_ASAP7_75t_SL g13443 ( 
.A(n_12584),
.Y(n_13443)
);

NAND2xp5_ASAP7_75t_L g13444 ( 
.A(n_12486),
.B(n_11150),
.Y(n_13444)
);

INVx2_ASAP7_75t_L g13445 ( 
.A(n_12206),
.Y(n_13445)
);

BUFx2_ASAP7_75t_L g13446 ( 
.A(n_12831),
.Y(n_13446)
);

INVx3_ASAP7_75t_SL g13447 ( 
.A(n_12355),
.Y(n_13447)
);

INVx2_ASAP7_75t_L g13448 ( 
.A(n_12229),
.Y(n_13448)
);

INVx1_ASAP7_75t_L g13449 ( 
.A(n_12892),
.Y(n_13449)
);

AND2x2_ASAP7_75t_L g13450 ( 
.A(n_12141),
.B(n_8960),
.Y(n_13450)
);

BUFx2_ASAP7_75t_L g13451 ( 
.A(n_12923),
.Y(n_13451)
);

INVx2_ASAP7_75t_L g13452 ( 
.A(n_12248),
.Y(n_13452)
);

INVx2_ASAP7_75t_L g13453 ( 
.A(n_12266),
.Y(n_13453)
);

INVx1_ASAP7_75t_L g13454 ( 
.A(n_12832),
.Y(n_13454)
);

NAND2xp5_ASAP7_75t_L g13455 ( 
.A(n_12498),
.B(n_11154),
.Y(n_13455)
);

BUFx6f_ASAP7_75t_L g13456 ( 
.A(n_12517),
.Y(n_13456)
);

AND2x2_ASAP7_75t_L g13457 ( 
.A(n_12149),
.B(n_9012),
.Y(n_13457)
);

BUFx2_ASAP7_75t_L g13458 ( 
.A(n_12923),
.Y(n_13458)
);

INVx1_ASAP7_75t_L g13459 ( 
.A(n_12845),
.Y(n_13459)
);

INVx2_ASAP7_75t_L g13460 ( 
.A(n_12269),
.Y(n_13460)
);

AND2x2_ASAP7_75t_L g13461 ( 
.A(n_12555),
.B(n_9012),
.Y(n_13461)
);

INVx2_ASAP7_75t_L g13462 ( 
.A(n_12292),
.Y(n_13462)
);

INVx1_ASAP7_75t_L g13463 ( 
.A(n_12848),
.Y(n_13463)
);

OR2x2_ASAP7_75t_L g13464 ( 
.A(n_12556),
.B(n_11155),
.Y(n_13464)
);

INVx1_ASAP7_75t_L g13465 ( 
.A(n_12854),
.Y(n_13465)
);

AND2x2_ASAP7_75t_L g13466 ( 
.A(n_12153),
.B(n_9012),
.Y(n_13466)
);

INVx2_ASAP7_75t_L g13467 ( 
.A(n_12298),
.Y(n_13467)
);

OR2x2_ASAP7_75t_L g13468 ( 
.A(n_12684),
.B(n_11156),
.Y(n_13468)
);

AND2x2_ASAP7_75t_L g13469 ( 
.A(n_12480),
.B(n_9015),
.Y(n_13469)
);

HB1xp67_ASAP7_75t_L g13470 ( 
.A(n_12861),
.Y(n_13470)
);

OR2x2_ASAP7_75t_L g13471 ( 
.A(n_12701),
.B(n_12523),
.Y(n_13471)
);

HB1xp67_ASAP7_75t_L g13472 ( 
.A(n_12869),
.Y(n_13472)
);

INVx2_ASAP7_75t_L g13473 ( 
.A(n_12348),
.Y(n_13473)
);

AND2x2_ASAP7_75t_L g13474 ( 
.A(n_12499),
.B(n_9015),
.Y(n_13474)
);

INVx1_ASAP7_75t_L g13475 ( 
.A(n_12891),
.Y(n_13475)
);

INVx1_ASAP7_75t_L g13476 ( 
.A(n_12905),
.Y(n_13476)
);

BUFx3_ASAP7_75t_L g13477 ( 
.A(n_12653),
.Y(n_13477)
);

INVx4_ASAP7_75t_L g13478 ( 
.A(n_12923),
.Y(n_13478)
);

OR2x2_ASAP7_75t_L g13479 ( 
.A(n_12751),
.B(n_11159),
.Y(n_13479)
);

HB1xp67_ASAP7_75t_L g13480 ( 
.A(n_12396),
.Y(n_13480)
);

INVx2_ASAP7_75t_L g13481 ( 
.A(n_12440),
.Y(n_13481)
);

NAND2xp5_ASAP7_75t_L g13482 ( 
.A(n_12667),
.B(n_11163),
.Y(n_13482)
);

INVx3_ASAP7_75t_L g13483 ( 
.A(n_12517),
.Y(n_13483)
);

INVx1_ASAP7_75t_L g13484 ( 
.A(n_12819),
.Y(n_13484)
);

AND2x2_ASAP7_75t_L g13485 ( 
.A(n_12505),
.B(n_9015),
.Y(n_13485)
);

INVx2_ASAP7_75t_L g13486 ( 
.A(n_12446),
.Y(n_13486)
);

INVx1_ASAP7_75t_L g13487 ( 
.A(n_12840),
.Y(n_13487)
);

INVx2_ASAP7_75t_L g13488 ( 
.A(n_12468),
.Y(n_13488)
);

INVx1_ASAP7_75t_L g13489 ( 
.A(n_12853),
.Y(n_13489)
);

BUFx3_ASAP7_75t_L g13490 ( 
.A(n_12460),
.Y(n_13490)
);

INVx1_ASAP7_75t_L g13491 ( 
.A(n_11990),
.Y(n_13491)
);

AND2x2_ASAP7_75t_L g13492 ( 
.A(n_12508),
.B(n_9050),
.Y(n_13492)
);

AND2x2_ASAP7_75t_L g13493 ( 
.A(n_12511),
.B(n_9050),
.Y(n_13493)
);

INVx1_ASAP7_75t_L g13494 ( 
.A(n_11990),
.Y(n_13494)
);

AND2x2_ASAP7_75t_L g13495 ( 
.A(n_12513),
.B(n_9050),
.Y(n_13495)
);

AND2x4_ASAP7_75t_L g13496 ( 
.A(n_12731),
.B(n_11856),
.Y(n_13496)
);

INVx1_ASAP7_75t_L g13497 ( 
.A(n_12642),
.Y(n_13497)
);

BUFx2_ASAP7_75t_L g13498 ( 
.A(n_12923),
.Y(n_13498)
);

INVx1_ASAP7_75t_L g13499 ( 
.A(n_12666),
.Y(n_13499)
);

HB1xp67_ASAP7_75t_L g13500 ( 
.A(n_12483),
.Y(n_13500)
);

BUFx3_ASAP7_75t_L g13501 ( 
.A(n_12460),
.Y(n_13501)
);

NAND2xp5_ASAP7_75t_L g13502 ( 
.A(n_12689),
.B(n_11164),
.Y(n_13502)
);

NOR2xp33_ASAP7_75t_L g13503 ( 
.A(n_12189),
.B(n_8720),
.Y(n_13503)
);

INVx2_ASAP7_75t_L g13504 ( 
.A(n_12510),
.Y(n_13504)
);

INVx2_ASAP7_75t_L g13505 ( 
.A(n_12564),
.Y(n_13505)
);

BUFx2_ASAP7_75t_L g13506 ( 
.A(n_12957),
.Y(n_13506)
);

INVxp67_ASAP7_75t_L g13507 ( 
.A(n_12272),
.Y(n_13507)
);

INVxp67_ASAP7_75t_L g13508 ( 
.A(n_12382),
.Y(n_13508)
);

INVx2_ASAP7_75t_L g13509 ( 
.A(n_12568),
.Y(n_13509)
);

INVx1_ASAP7_75t_L g13510 ( 
.A(n_12793),
.Y(n_13510)
);

INVx1_ASAP7_75t_L g13511 ( 
.A(n_12793),
.Y(n_13511)
);

AND2x2_ASAP7_75t_L g13512 ( 
.A(n_12521),
.B(n_9061),
.Y(n_13512)
);

INVx3_ASAP7_75t_L g13513 ( 
.A(n_12194),
.Y(n_13513)
);

AND2x2_ASAP7_75t_L g13514 ( 
.A(n_12322),
.B(n_9061),
.Y(n_13514)
);

INVx2_ASAP7_75t_SL g13515 ( 
.A(n_12738),
.Y(n_13515)
);

INVx2_ASAP7_75t_L g13516 ( 
.A(n_12576),
.Y(n_13516)
);

INVx1_ASAP7_75t_L g13517 ( 
.A(n_12728),
.Y(n_13517)
);

INVx2_ASAP7_75t_L g13518 ( 
.A(n_12602),
.Y(n_13518)
);

INVx2_ASAP7_75t_SL g13519 ( 
.A(n_12738),
.Y(n_13519)
);

AND2x4_ASAP7_75t_L g13520 ( 
.A(n_12267),
.B(n_11856),
.Y(n_13520)
);

BUFx2_ASAP7_75t_L g13521 ( 
.A(n_12855),
.Y(n_13521)
);

AND2x2_ASAP7_75t_L g13522 ( 
.A(n_12308),
.B(n_9061),
.Y(n_13522)
);

INVxp67_ASAP7_75t_L g13523 ( 
.A(n_12062),
.Y(n_13523)
);

BUFx6f_ASAP7_75t_L g13524 ( 
.A(n_12855),
.Y(n_13524)
);

INVx1_ASAP7_75t_L g13525 ( 
.A(n_12728),
.Y(n_13525)
);

INVx2_ASAP7_75t_L g13526 ( 
.A(n_12607),
.Y(n_13526)
);

INVx2_ASAP7_75t_L g13527 ( 
.A(n_12622),
.Y(n_13527)
);

NAND2xp5_ASAP7_75t_L g13528 ( 
.A(n_11970),
.B(n_11166),
.Y(n_13528)
);

INVx3_ASAP7_75t_L g13529 ( 
.A(n_12194),
.Y(n_13529)
);

AND2x2_ASAP7_75t_L g13530 ( 
.A(n_12100),
.B(n_9095),
.Y(n_13530)
);

INVx1_ASAP7_75t_L g13531 ( 
.A(n_12728),
.Y(n_13531)
);

INVx1_ASAP7_75t_L g13532 ( 
.A(n_12115),
.Y(n_13532)
);

AND2x2_ASAP7_75t_L g13533 ( 
.A(n_12299),
.B(n_9095),
.Y(n_13533)
);

INVx1_ASAP7_75t_L g13534 ( 
.A(n_12115),
.Y(n_13534)
);

INVx2_ASAP7_75t_L g13535 ( 
.A(n_12638),
.Y(n_13535)
);

AND2x2_ASAP7_75t_L g13536 ( 
.A(n_12301),
.B(n_9095),
.Y(n_13536)
);

INVx1_ASAP7_75t_L g13537 ( 
.A(n_12247),
.Y(n_13537)
);

BUFx3_ASAP7_75t_L g13538 ( 
.A(n_12363),
.Y(n_13538)
);

AND2x2_ASAP7_75t_L g13539 ( 
.A(n_12692),
.B(n_12208),
.Y(n_13539)
);

INVx2_ASAP7_75t_L g13540 ( 
.A(n_12677),
.Y(n_13540)
);

AND2x2_ASAP7_75t_L g13541 ( 
.A(n_12210),
.B(n_9100),
.Y(n_13541)
);

INVx1_ASAP7_75t_L g13542 ( 
.A(n_12247),
.Y(n_13542)
);

INVx1_ASAP7_75t_L g13543 ( 
.A(n_12343),
.Y(n_13543)
);

AND2x2_ASAP7_75t_L g13544 ( 
.A(n_12228),
.B(n_9100),
.Y(n_13544)
);

INVx3_ASAP7_75t_L g13545 ( 
.A(n_12278),
.Y(n_13545)
);

INVx3_ASAP7_75t_L g13546 ( 
.A(n_12278),
.Y(n_13546)
);

INVxp67_ASAP7_75t_SL g13547 ( 
.A(n_12594),
.Y(n_13547)
);

BUFx3_ASAP7_75t_L g13548 ( 
.A(n_12193),
.Y(n_13548)
);

BUFx2_ASAP7_75t_L g13549 ( 
.A(n_12798),
.Y(n_13549)
);

INVx2_ASAP7_75t_L g13550 ( 
.A(n_12688),
.Y(n_13550)
);

INVx2_ASAP7_75t_L g13551 ( 
.A(n_12693),
.Y(n_13551)
);

AND2x2_ASAP7_75t_L g13552 ( 
.A(n_12230),
.B(n_9100),
.Y(n_13552)
);

HB1xp67_ASAP7_75t_L g13553 ( 
.A(n_12695),
.Y(n_13553)
);

INVx3_ASAP7_75t_L g13554 ( 
.A(n_12318),
.Y(n_13554)
);

INVx1_ASAP7_75t_L g13555 ( 
.A(n_12343),
.Y(n_13555)
);

INVx2_ASAP7_75t_L g13556 ( 
.A(n_12762),
.Y(n_13556)
);

INVx2_ASAP7_75t_L g13557 ( 
.A(n_12770),
.Y(n_13557)
);

AND2x2_ASAP7_75t_L g13558 ( 
.A(n_12537),
.B(n_9161),
.Y(n_13558)
);

INVx2_ASAP7_75t_L g13559 ( 
.A(n_12773),
.Y(n_13559)
);

AND2x2_ASAP7_75t_L g13560 ( 
.A(n_12323),
.B(n_9161),
.Y(n_13560)
);

INVx2_ASAP7_75t_L g13561 ( 
.A(n_12929),
.Y(n_13561)
);

AND2x4_ASAP7_75t_L g13562 ( 
.A(n_12183),
.B(n_12199),
.Y(n_13562)
);

INVx2_ASAP7_75t_L g13563 ( 
.A(n_12318),
.Y(n_13563)
);

INVx3_ASAP7_75t_L g13564 ( 
.A(n_12384),
.Y(n_13564)
);

NAND2xp5_ASAP7_75t_L g13565 ( 
.A(n_11972),
.B(n_11167),
.Y(n_13565)
);

HB1xp67_ASAP7_75t_L g13566 ( 
.A(n_12782),
.Y(n_13566)
);

INVx1_ASAP7_75t_L g13567 ( 
.A(n_12346),
.Y(n_13567)
);

INVx1_ASAP7_75t_L g13568 ( 
.A(n_12346),
.Y(n_13568)
);

AND2x2_ASAP7_75t_L g13569 ( 
.A(n_12329),
.B(n_9161),
.Y(n_13569)
);

INVx1_ASAP7_75t_L g13570 ( 
.A(n_12392),
.Y(n_13570)
);

OR2x2_ASAP7_75t_L g13571 ( 
.A(n_12797),
.B(n_11170),
.Y(n_13571)
);

AND2x2_ASAP7_75t_L g13572 ( 
.A(n_12019),
.B(n_9162),
.Y(n_13572)
);

BUFx2_ASAP7_75t_L g13573 ( 
.A(n_12527),
.Y(n_13573)
);

NAND2xp5_ASAP7_75t_L g13574 ( 
.A(n_12520),
.B(n_11176),
.Y(n_13574)
);

INVx2_ASAP7_75t_L g13575 ( 
.A(n_12611),
.Y(n_13575)
);

INVx1_ASAP7_75t_L g13576 ( 
.A(n_12392),
.Y(n_13576)
);

INVx1_ASAP7_75t_L g13577 ( 
.A(n_12393),
.Y(n_13577)
);

NOR2x1_ASAP7_75t_SL g13578 ( 
.A(n_12165),
.B(n_12219),
.Y(n_13578)
);

INVx1_ASAP7_75t_L g13579 ( 
.A(n_12393),
.Y(n_13579)
);

OA21x2_ASAP7_75t_L g13580 ( 
.A1(n_12893),
.A2(n_11079),
.B(n_11076),
.Y(n_13580)
);

AND2x2_ASAP7_75t_L g13581 ( 
.A(n_12074),
.B(n_9162),
.Y(n_13581)
);

INVx2_ASAP7_75t_L g13582 ( 
.A(n_12618),
.Y(n_13582)
);

AND2x2_ASAP7_75t_L g13583 ( 
.A(n_12074),
.B(n_9162),
.Y(n_13583)
);

INVx1_ASAP7_75t_L g13584 ( 
.A(n_12395),
.Y(n_13584)
);

AND2x2_ASAP7_75t_L g13585 ( 
.A(n_12545),
.B(n_9166),
.Y(n_13585)
);

INVx2_ASAP7_75t_L g13586 ( 
.A(n_12937),
.Y(n_13586)
);

AND2x2_ASAP7_75t_L g13587 ( 
.A(n_12076),
.B(n_9166),
.Y(n_13587)
);

AND2x2_ASAP7_75t_L g13588 ( 
.A(n_12422),
.B(n_9166),
.Y(n_13588)
);

AND2x2_ASAP7_75t_L g13589 ( 
.A(n_12170),
.B(n_9206),
.Y(n_13589)
);

AND2x2_ASAP7_75t_L g13590 ( 
.A(n_12176),
.B(n_9206),
.Y(n_13590)
);

NAND2xp5_ASAP7_75t_L g13591 ( 
.A(n_12000),
.B(n_11179),
.Y(n_13591)
);

BUFx6f_ASAP7_75t_L g13592 ( 
.A(n_12943),
.Y(n_13592)
);

BUFx3_ASAP7_75t_L g13593 ( 
.A(n_12254),
.Y(n_13593)
);

INVx2_ASAP7_75t_L g13594 ( 
.A(n_12833),
.Y(n_13594)
);

AND2x2_ASAP7_75t_L g13595 ( 
.A(n_12195),
.B(n_9206),
.Y(n_13595)
);

AND2x4_ASAP7_75t_L g13596 ( 
.A(n_12496),
.B(n_11856),
.Y(n_13596)
);

AND2x2_ASAP7_75t_L g13597 ( 
.A(n_12201),
.B(n_9140),
.Y(n_13597)
);

INVx1_ASAP7_75t_L g13598 ( 
.A(n_12395),
.Y(n_13598)
);

OR2x2_ASAP7_75t_L g13599 ( 
.A(n_12813),
.B(n_11185),
.Y(n_13599)
);

INVx1_ASAP7_75t_L g13600 ( 
.A(n_12178),
.Y(n_13600)
);

INVx2_ASAP7_75t_L g13601 ( 
.A(n_12791),
.Y(n_13601)
);

INVx2_ASAP7_75t_L g13602 ( 
.A(n_12737),
.Y(n_13602)
);

INVx2_ASAP7_75t_L g13603 ( 
.A(n_12740),
.Y(n_13603)
);

BUFx3_ASAP7_75t_L g13604 ( 
.A(n_12331),
.Y(n_13604)
);

AND2x2_ASAP7_75t_L g13605 ( 
.A(n_12207),
.B(n_9140),
.Y(n_13605)
);

HB1xp67_ASAP7_75t_L g13606 ( 
.A(n_12824),
.Y(n_13606)
);

HB1xp67_ASAP7_75t_L g13607 ( 
.A(n_12846),
.Y(n_13607)
);

BUFx2_ASAP7_75t_SL g13608 ( 
.A(n_12412),
.Y(n_13608)
);

INVx1_ASAP7_75t_L g13609 ( 
.A(n_12178),
.Y(n_13609)
);

AND2x2_ASAP7_75t_L g13610 ( 
.A(n_12536),
.B(n_9140),
.Y(n_13610)
);

AND2x2_ASAP7_75t_L g13611 ( 
.A(n_12162),
.B(n_12291),
.Y(n_13611)
);

INVx2_ASAP7_75t_L g13612 ( 
.A(n_12741),
.Y(n_13612)
);

OR2x2_ASAP7_75t_L g13613 ( 
.A(n_12685),
.B(n_11186),
.Y(n_13613)
);

OR2x2_ASAP7_75t_L g13614 ( 
.A(n_12759),
.B(n_11193),
.Y(n_13614)
);

INVx1_ASAP7_75t_SL g13615 ( 
.A(n_12250),
.Y(n_13615)
);

INVx2_ASAP7_75t_L g13616 ( 
.A(n_12743),
.Y(n_13616)
);

INVx1_ASAP7_75t_L g13617 ( 
.A(n_12309),
.Y(n_13617)
);

HB1xp67_ASAP7_75t_L g13618 ( 
.A(n_12084),
.Y(n_13618)
);

OR2x6_ASAP7_75t_L g13619 ( 
.A(n_12158),
.B(n_9074),
.Y(n_13619)
);

INVx1_ASAP7_75t_L g13620 ( 
.A(n_12309),
.Y(n_13620)
);

INVx1_ASAP7_75t_L g13621 ( 
.A(n_12807),
.Y(n_13621)
);

OR2x2_ASAP7_75t_L g13622 ( 
.A(n_12563),
.B(n_11196),
.Y(n_13622)
);

NAND2xp5_ASAP7_75t_L g13623 ( 
.A(n_12371),
.B(n_11198),
.Y(n_13623)
);

BUFx2_ASAP7_75t_L g13624 ( 
.A(n_12619),
.Y(n_13624)
);

OR2x2_ASAP7_75t_L g13625 ( 
.A(n_12628),
.B(n_11200),
.Y(n_13625)
);

HB1xp67_ASAP7_75t_L g13626 ( 
.A(n_12084),
.Y(n_13626)
);

BUFx3_ASAP7_75t_L g13627 ( 
.A(n_12249),
.Y(n_13627)
);

AND2x2_ASAP7_75t_L g13628 ( 
.A(n_12598),
.B(n_8652),
.Y(n_13628)
);

INVx2_ASAP7_75t_L g13629 ( 
.A(n_12744),
.Y(n_13629)
);

INVx1_ASAP7_75t_L g13630 ( 
.A(n_12501),
.Y(n_13630)
);

INVx1_ASAP7_75t_L g13631 ( 
.A(n_12501),
.Y(n_13631)
);

HB1xp67_ASAP7_75t_L g13632 ( 
.A(n_12788),
.Y(n_13632)
);

INVx1_ASAP7_75t_L g13633 ( 
.A(n_12501),
.Y(n_13633)
);

AND2x2_ASAP7_75t_L g13634 ( 
.A(n_12948),
.B(n_8652),
.Y(n_13634)
);

INVx2_ASAP7_75t_L g13635 ( 
.A(n_12849),
.Y(n_13635)
);

NAND2xp5_ASAP7_75t_L g13636 ( 
.A(n_11965),
.B(n_11201),
.Y(n_13636)
);

AND2x2_ASAP7_75t_L g13637 ( 
.A(n_12636),
.B(n_8652),
.Y(n_13637)
);

OR2x2_ASAP7_75t_L g13638 ( 
.A(n_12661),
.B(n_11207),
.Y(n_13638)
);

OR2x2_ASAP7_75t_L g13639 ( 
.A(n_12681),
.B(n_11210),
.Y(n_13639)
);

AND2x4_ASAP7_75t_L g13640 ( 
.A(n_12512),
.B(n_12624),
.Y(n_13640)
);

AND2x2_ASAP7_75t_L g13641 ( 
.A(n_12544),
.B(n_8721),
.Y(n_13641)
);

AOI22xp33_ASAP7_75t_L g13642 ( 
.A1(n_12017),
.A2(n_8699),
.B1(n_8665),
.B2(n_8554),
.Y(n_13642)
);

AND2x2_ASAP7_75t_L g13643 ( 
.A(n_12411),
.B(n_8721),
.Y(n_13643)
);

INVx2_ASAP7_75t_L g13644 ( 
.A(n_12856),
.Y(n_13644)
);

INVx2_ASAP7_75t_L g13645 ( 
.A(n_12872),
.Y(n_13645)
);

INVx1_ASAP7_75t_L g13646 ( 
.A(n_12313),
.Y(n_13646)
);

INVx1_ASAP7_75t_L g13647 ( 
.A(n_12418),
.Y(n_13647)
);

INVx2_ASAP7_75t_L g13648 ( 
.A(n_12884),
.Y(n_13648)
);

INVx2_ASAP7_75t_L g13649 ( 
.A(n_12887),
.Y(n_13649)
);

INVx1_ASAP7_75t_L g13650 ( 
.A(n_12217),
.Y(n_13650)
);

INVx1_ASAP7_75t_L g13651 ( 
.A(n_12454),
.Y(n_13651)
);

AND2x2_ASAP7_75t_L g13652 ( 
.A(n_12026),
.B(n_8721),
.Y(n_13652)
);

AND2x2_ASAP7_75t_L g13653 ( 
.A(n_12232),
.B(n_8079),
.Y(n_13653)
);

HB1xp67_ASAP7_75t_L g13654 ( 
.A(n_12401),
.Y(n_13654)
);

AND2x2_ASAP7_75t_L g13655 ( 
.A(n_12023),
.B(n_12242),
.Y(n_13655)
);

INVx2_ASAP7_75t_L g13656 ( 
.A(n_12796),
.Y(n_13656)
);

AND2x2_ASAP7_75t_L g13657 ( 
.A(n_12031),
.B(n_8079),
.Y(n_13657)
);

INVx1_ASAP7_75t_L g13658 ( 
.A(n_12750),
.Y(n_13658)
);

AND2x2_ASAP7_75t_L g13659 ( 
.A(n_12469),
.B(n_12577),
.Y(n_13659)
);

INVx2_ASAP7_75t_L g13660 ( 
.A(n_12750),
.Y(n_13660)
);

INVx1_ASAP7_75t_L g13661 ( 
.A(n_12816),
.Y(n_13661)
);

INVx1_ASAP7_75t_L g13662 ( 
.A(n_12725),
.Y(n_13662)
);

INVx3_ASAP7_75t_L g13663 ( 
.A(n_12570),
.Y(n_13663)
);

AND2x2_ASAP7_75t_L g13664 ( 
.A(n_12588),
.B(n_8079),
.Y(n_13664)
);

INVx2_ASAP7_75t_L g13665 ( 
.A(n_12939),
.Y(n_13665)
);

CKINVDCx14_ASAP7_75t_R g13666 ( 
.A(n_12142),
.Y(n_13666)
);

AND2x2_ASAP7_75t_L g13667 ( 
.A(n_12589),
.B(n_8079),
.Y(n_13667)
);

AND2x2_ASAP7_75t_L g13668 ( 
.A(n_12519),
.B(n_8079),
.Y(n_13668)
);

AND2x2_ASAP7_75t_L g13669 ( 
.A(n_12163),
.B(n_8079),
.Y(n_13669)
);

OAI22xp5_ASAP7_75t_SL g13670 ( 
.A1(n_11939),
.A2(n_12002),
.B1(n_12003),
.B2(n_11998),
.Y(n_13670)
);

AND2x2_ASAP7_75t_L g13671 ( 
.A(n_12252),
.B(n_11964),
.Y(n_13671)
);

INVx1_ASAP7_75t_L g13672 ( 
.A(n_12288),
.Y(n_13672)
);

INVx2_ASAP7_75t_L g13673 ( 
.A(n_12951),
.Y(n_13673)
);

HB1xp67_ASAP7_75t_L g13674 ( 
.A(n_12746),
.Y(n_13674)
);

AND2x2_ASAP7_75t_L g13675 ( 
.A(n_12258),
.B(n_8082),
.Y(n_13675)
);

INVx2_ASAP7_75t_L g13676 ( 
.A(n_12894),
.Y(n_13676)
);

INVx1_ASAP7_75t_L g13677 ( 
.A(n_12529),
.Y(n_13677)
);

NOR2x1p5_ASAP7_75t_L g13678 ( 
.A(n_11986),
.B(n_9074),
.Y(n_13678)
);

AND2x2_ASAP7_75t_L g13679 ( 
.A(n_12261),
.B(n_8082),
.Y(n_13679)
);

INVx1_ASAP7_75t_L g13680 ( 
.A(n_12531),
.Y(n_13680)
);

OR2x2_ASAP7_75t_L g13681 ( 
.A(n_12030),
.B(n_11211),
.Y(n_13681)
);

INVx1_ASAP7_75t_L g13682 ( 
.A(n_12546),
.Y(n_13682)
);

INVx1_ASAP7_75t_L g13683 ( 
.A(n_12557),
.Y(n_13683)
);

AND2x4_ASAP7_75t_L g13684 ( 
.A(n_12756),
.B(n_11860),
.Y(n_13684)
);

AND2x2_ASAP7_75t_L g13685 ( 
.A(n_11967),
.B(n_8082),
.Y(n_13685)
);

BUFx3_ASAP7_75t_L g13686 ( 
.A(n_12253),
.Y(n_13686)
);

AND2x2_ASAP7_75t_L g13687 ( 
.A(n_12273),
.B(n_8082),
.Y(n_13687)
);

NAND2xp5_ASAP7_75t_L g13688 ( 
.A(n_12020),
.B(n_11213),
.Y(n_13688)
);

AND2x2_ASAP7_75t_L g13689 ( 
.A(n_12276),
.B(n_8082),
.Y(n_13689)
);

AND2x2_ASAP7_75t_L g13690 ( 
.A(n_12277),
.B(n_8082),
.Y(n_13690)
);

AND2x2_ASAP7_75t_L g13691 ( 
.A(n_12281),
.B(n_8244),
.Y(n_13691)
);

INVx2_ASAP7_75t_L g13692 ( 
.A(n_12902),
.Y(n_13692)
);

AO31x2_ASAP7_75t_L g13693 ( 
.A1(n_12403),
.A2(n_11339),
.A3(n_11340),
.B(n_11337),
.Y(n_13693)
);

AND2x4_ASAP7_75t_L g13694 ( 
.A(n_12542),
.B(n_11860),
.Y(n_13694)
);

HB1xp67_ASAP7_75t_L g13695 ( 
.A(n_12746),
.Y(n_13695)
);

HB1xp67_ASAP7_75t_L g13696 ( 
.A(n_12925),
.Y(n_13696)
);

INVx1_ASAP7_75t_L g13697 ( 
.A(n_12461),
.Y(n_13697)
);

HB1xp67_ASAP7_75t_L g13698 ( 
.A(n_12947),
.Y(n_13698)
);

HB1xp67_ASAP7_75t_L g13699 ( 
.A(n_12088),
.Y(n_13699)
);

INVx2_ASAP7_75t_L g13700 ( 
.A(n_12609),
.Y(n_13700)
);

INVx1_ASAP7_75t_L g13701 ( 
.A(n_12461),
.Y(n_13701)
);

INVx1_ASAP7_75t_L g13702 ( 
.A(n_12601),
.Y(n_13702)
);

AND2x2_ASAP7_75t_L g13703 ( 
.A(n_12425),
.B(n_8244),
.Y(n_13703)
);

AND2x4_ASAP7_75t_L g13704 ( 
.A(n_12264),
.B(n_11860),
.Y(n_13704)
);

AND2x2_ASAP7_75t_L g13705 ( 
.A(n_12271),
.B(n_12654),
.Y(n_13705)
);

INVx2_ASAP7_75t_L g13706 ( 
.A(n_12789),
.Y(n_13706)
);

INVx1_ASAP7_75t_L g13707 ( 
.A(n_12601),
.Y(n_13707)
);

INVx2_ASAP7_75t_L g13708 ( 
.A(n_12814),
.Y(n_13708)
);

NAND2xp5_ASAP7_75t_SL g13709 ( 
.A(n_12366),
.B(n_8095),
.Y(n_13709)
);

INVx2_ASAP7_75t_L g13710 ( 
.A(n_12890),
.Y(n_13710)
);

AOI22xp5_ASAP7_75t_L g13711 ( 
.A1(n_12110),
.A2(n_12081),
.B1(n_12093),
.B2(n_12067),
.Y(n_13711)
);

INVx2_ASAP7_75t_L g13712 ( 
.A(n_12265),
.Y(n_13712)
);

AND2x2_ASAP7_75t_L g13713 ( 
.A(n_12662),
.B(n_8244),
.Y(n_13713)
);

BUFx2_ASAP7_75t_L g13714 ( 
.A(n_12274),
.Y(n_13714)
);

INVx2_ASAP7_75t_L g13715 ( 
.A(n_12349),
.Y(n_13715)
);

HB1xp67_ASAP7_75t_L g13716 ( 
.A(n_12522),
.Y(n_13716)
);

INVx2_ASAP7_75t_L g13717 ( 
.A(n_12772),
.Y(n_13717)
);

AND2x2_ASAP7_75t_L g13718 ( 
.A(n_12532),
.B(n_8244),
.Y(n_13718)
);

AND2x2_ASAP7_75t_L g13719 ( 
.A(n_12533),
.B(n_8244),
.Y(n_13719)
);

AND2x2_ASAP7_75t_L g13720 ( 
.A(n_11958),
.B(n_8244),
.Y(n_13720)
);

INVx2_ASAP7_75t_L g13721 ( 
.A(n_12344),
.Y(n_13721)
);

NAND2xp5_ASAP7_75t_L g13722 ( 
.A(n_12107),
.B(n_11218),
.Y(n_13722)
);

AND2x2_ASAP7_75t_L g13723 ( 
.A(n_12605),
.B(n_8349),
.Y(n_13723)
);

INVx2_ASAP7_75t_L g13724 ( 
.A(n_12603),
.Y(n_13724)
);

INVx2_ASAP7_75t_L g13725 ( 
.A(n_12603),
.Y(n_13725)
);

INVx1_ASAP7_75t_L g13726 ( 
.A(n_12353),
.Y(n_13726)
);

INVx2_ASAP7_75t_L g13727 ( 
.A(n_12060),
.Y(n_13727)
);

INVx2_ASAP7_75t_L g13728 ( 
.A(n_12551),
.Y(n_13728)
);

INVx1_ASAP7_75t_L g13729 ( 
.A(n_12111),
.Y(n_13729)
);

AND2x4_ASAP7_75t_L g13730 ( 
.A(n_12220),
.B(n_11861),
.Y(n_13730)
);

BUFx6f_ASAP7_75t_L g13731 ( 
.A(n_12111),
.Y(n_13731)
);

INVx4_ASAP7_75t_R g13732 ( 
.A(n_12188),
.Y(n_13732)
);

BUFx2_ASAP7_75t_L g13733 ( 
.A(n_12284),
.Y(n_13733)
);

INVx1_ASAP7_75t_L g13734 ( 
.A(n_12101),
.Y(n_13734)
);

AND2x2_ASAP7_75t_L g13735 ( 
.A(n_12616),
.B(n_8349),
.Y(n_13735)
);

INVx1_ASAP7_75t_L g13736 ( 
.A(n_12105),
.Y(n_13736)
);

INVx1_ASAP7_75t_L g13737 ( 
.A(n_12051),
.Y(n_13737)
);

OR2x2_ASAP7_75t_L g13738 ( 
.A(n_12047),
.B(n_11221),
.Y(n_13738)
);

INVx2_ASAP7_75t_L g13739 ( 
.A(n_12924),
.Y(n_13739)
);

NAND2xp5_ASAP7_75t_L g13740 ( 
.A(n_12182),
.B(n_11222),
.Y(n_13740)
);

INVx1_ASAP7_75t_L g13741 ( 
.A(n_12458),
.Y(n_13741)
);

AND2x2_ASAP7_75t_L g13742 ( 
.A(n_12421),
.B(n_8349),
.Y(n_13742)
);

INVx2_ASAP7_75t_L g13743 ( 
.A(n_12458),
.Y(n_13743)
);

HB1xp67_ASAP7_75t_L g13744 ( 
.A(n_12389),
.Y(n_13744)
);

INVx2_ASAP7_75t_L g13745 ( 
.A(n_12540),
.Y(n_13745)
);

AND2x2_ASAP7_75t_L g13746 ( 
.A(n_12842),
.B(n_8349),
.Y(n_13746)
);

OR2x2_ASAP7_75t_L g13747 ( 
.A(n_12090),
.B(n_11230),
.Y(n_13747)
);

AND2x2_ASAP7_75t_L g13748 ( 
.A(n_12851),
.B(n_8349),
.Y(n_13748)
);

OAI21xp5_ASAP7_75t_SL g13749 ( 
.A1(n_11937),
.A2(n_9209),
.B(n_8862),
.Y(n_13749)
);

AND2x2_ASAP7_75t_L g13750 ( 
.A(n_12863),
.B(n_8349),
.Y(n_13750)
);

INVx1_ASAP7_75t_L g13751 ( 
.A(n_12540),
.Y(n_13751)
);

AND2x2_ASAP7_75t_L g13752 ( 
.A(n_12867),
.B(n_8412),
.Y(n_13752)
);

INVx2_ASAP7_75t_L g13753 ( 
.A(n_12918),
.Y(n_13753)
);

INVx2_ASAP7_75t_L g13754 ( 
.A(n_12610),
.Y(n_13754)
);

INVx1_ASAP7_75t_L g13755 ( 
.A(n_12896),
.Y(n_13755)
);

INVx1_ASAP7_75t_L g13756 ( 
.A(n_12932),
.Y(n_13756)
);

AND2x2_ASAP7_75t_L g13757 ( 
.A(n_12870),
.B(n_8412),
.Y(n_13757)
);

AND2x2_ASAP7_75t_L g13758 ( 
.A(n_12879),
.B(n_12910),
.Y(n_13758)
);

INVx1_ASAP7_75t_L g13759 ( 
.A(n_12289),
.Y(n_13759)
);

OR2x2_ASAP7_75t_L g13760 ( 
.A(n_12029),
.B(n_11234),
.Y(n_13760)
);

OR2x2_ASAP7_75t_L g13761 ( 
.A(n_12083),
.B(n_11235),
.Y(n_13761)
);

INVx3_ASAP7_75t_L g13762 ( 
.A(n_12827),
.Y(n_13762)
);

AOI22xp33_ASAP7_75t_L g13763 ( 
.A1(n_11979),
.A2(n_8699),
.B1(n_8665),
.B2(n_8574),
.Y(n_13763)
);

AND2x2_ASAP7_75t_L g13764 ( 
.A(n_12912),
.B(n_8412),
.Y(n_13764)
);

INVx1_ASAP7_75t_L g13765 ( 
.A(n_12235),
.Y(n_13765)
);

AND2x2_ASAP7_75t_SL g13766 ( 
.A(n_12012),
.B(n_7991),
.Y(n_13766)
);

INVx2_ASAP7_75t_L g13767 ( 
.A(n_12625),
.Y(n_13767)
);

NAND2xp5_ASAP7_75t_L g13768 ( 
.A(n_12118),
.B(n_11242),
.Y(n_13768)
);

BUFx2_ASAP7_75t_L g13769 ( 
.A(n_12119),
.Y(n_13769)
);

INVx2_ASAP7_75t_L g13770 ( 
.A(n_12640),
.Y(n_13770)
);

INVx1_ASAP7_75t_L g13771 ( 
.A(n_12270),
.Y(n_13771)
);

INVx1_ASAP7_75t_L g13772 ( 
.A(n_12372),
.Y(n_13772)
);

INVx1_ASAP7_75t_L g13773 ( 
.A(n_12380),
.Y(n_13773)
);

AND2x2_ASAP7_75t_L g13774 ( 
.A(n_12623),
.B(n_8412),
.Y(n_13774)
);

NAND2xp5_ASAP7_75t_L g13775 ( 
.A(n_12087),
.B(n_11243),
.Y(n_13775)
);

INVx1_ASAP7_75t_L g13776 ( 
.A(n_12864),
.Y(n_13776)
);

AND2x2_ASAP7_75t_L g13777 ( 
.A(n_12626),
.B(n_8412),
.Y(n_13777)
);

AND2x2_ASAP7_75t_L g13778 ( 
.A(n_12631),
.B(n_12676),
.Y(n_13778)
);

AND2x2_ASAP7_75t_L g13779 ( 
.A(n_12682),
.B(n_8412),
.Y(n_13779)
);

HB1xp67_ASAP7_75t_L g13780 ( 
.A(n_12400),
.Y(n_13780)
);

INVx2_ASAP7_75t_L g13781 ( 
.A(n_12657),
.Y(n_13781)
);

AND2x4_ASAP7_75t_SL g13782 ( 
.A(n_12451),
.B(n_8210),
.Y(n_13782)
);

AND2x2_ASAP7_75t_L g13783 ( 
.A(n_12691),
.B(n_8424),
.Y(n_13783)
);

OR2x2_ASAP7_75t_L g13784 ( 
.A(n_12246),
.B(n_11244),
.Y(n_13784)
);

BUFx6f_ASAP7_75t_L g13785 ( 
.A(n_12092),
.Y(n_13785)
);

OR2x2_ASAP7_75t_L g13786 ( 
.A(n_12010),
.B(n_11246),
.Y(n_13786)
);

BUFx3_ASAP7_75t_L g13787 ( 
.A(n_12394),
.Y(n_13787)
);

INVx3_ASAP7_75t_L g13788 ( 
.A(n_12643),
.Y(n_13788)
);

INVx3_ASAP7_75t_L g13789 ( 
.A(n_12687),
.Y(n_13789)
);

INVx2_ASAP7_75t_L g13790 ( 
.A(n_12600),
.Y(n_13790)
);

INVx1_ASAP7_75t_L g13791 ( 
.A(n_12659),
.Y(n_13791)
);

INVx2_ASAP7_75t_L g13792 ( 
.A(n_12660),
.Y(n_13792)
);

OR2x2_ASAP7_75t_L g13793 ( 
.A(n_12374),
.B(n_11249),
.Y(n_13793)
);

AND2x4_ASAP7_75t_L g13794 ( 
.A(n_12558),
.B(n_11861),
.Y(n_13794)
);

NOR2x1_ASAP7_75t_L g13795 ( 
.A(n_12237),
.B(n_11861),
.Y(n_13795)
);

INVx1_ASAP7_75t_L g13796 ( 
.A(n_12089),
.Y(n_13796)
);

INVxp67_ASAP7_75t_L g13797 ( 
.A(n_12072),
.Y(n_13797)
);

AO21x2_ASAP7_75t_L g13798 ( 
.A1(n_12077),
.A2(n_11252),
.B(n_11250),
.Y(n_13798)
);

INVx1_ASAP7_75t_L g13799 ( 
.A(n_12104),
.Y(n_13799)
);

INVx1_ASAP7_75t_L g13800 ( 
.A(n_12080),
.Y(n_13800)
);

AND2x2_ASAP7_75t_L g13801 ( 
.A(n_12696),
.B(n_8424),
.Y(n_13801)
);

NAND2xp5_ASAP7_75t_L g13802 ( 
.A(n_12358),
.B(n_11261),
.Y(n_13802)
);

AND2x4_ASAP7_75t_L g13803 ( 
.A(n_12675),
.B(n_11914),
.Y(n_13803)
);

AND2x2_ASAP7_75t_L g13804 ( 
.A(n_11988),
.B(n_8424),
.Y(n_13804)
);

AND2x2_ASAP7_75t_L g13805 ( 
.A(n_12935),
.B(n_8424),
.Y(n_13805)
);

INVx1_ASAP7_75t_SL g13806 ( 
.A(n_12013),
.Y(n_13806)
);

AND2x2_ASAP7_75t_L g13807 ( 
.A(n_12794),
.B(n_8424),
.Y(n_13807)
);

AND2x2_ASAP7_75t_L g13808 ( 
.A(n_12800),
.B(n_12463),
.Y(n_13808)
);

INVx1_ASAP7_75t_L g13809 ( 
.A(n_12391),
.Y(n_13809)
);

INVx1_ASAP7_75t_L g13810 ( 
.A(n_11943),
.Y(n_13810)
);

BUFx3_ASAP7_75t_L g13811 ( 
.A(n_12116),
.Y(n_13811)
);

INVx1_ASAP7_75t_L g13812 ( 
.A(n_12757),
.Y(n_13812)
);

INVx3_ASAP7_75t_L g13813 ( 
.A(n_12573),
.Y(n_13813)
);

INVx2_ASAP7_75t_L g13814 ( 
.A(n_12300),
.Y(n_13814)
);

INVx1_ASAP7_75t_L g13815 ( 
.A(n_12825),
.Y(n_13815)
);

INVx2_ASAP7_75t_L g13816 ( 
.A(n_12459),
.Y(n_13816)
);

AND2x2_ASAP7_75t_L g13817 ( 
.A(n_12467),
.B(n_8424),
.Y(n_13817)
);

AND2x2_ASAP7_75t_L g13818 ( 
.A(n_12528),
.B(n_8500),
.Y(n_13818)
);

BUFx3_ASAP7_75t_L g13819 ( 
.A(n_12236),
.Y(n_13819)
);

AND2x2_ASAP7_75t_L g13820 ( 
.A(n_12703),
.B(n_8500),
.Y(n_13820)
);

OR2x2_ASAP7_75t_L g13821 ( 
.A(n_12378),
.B(n_11262),
.Y(n_13821)
);

INVx3_ASAP7_75t_L g13822 ( 
.A(n_12427),
.Y(n_13822)
);

AND2x2_ASAP7_75t_L g13823 ( 
.A(n_12722),
.B(n_8500),
.Y(n_13823)
);

INVx2_ASAP7_75t_L g13824 ( 
.A(n_12466),
.Y(n_13824)
);

INVx1_ASAP7_75t_L g13825 ( 
.A(n_12889),
.Y(n_13825)
);

AO31x2_ASAP7_75t_L g13826 ( 
.A1(n_12204),
.A2(n_11347),
.A3(n_11349),
.B(n_11342),
.Y(n_13826)
);

AO31x2_ASAP7_75t_L g13827 ( 
.A1(n_12303),
.A2(n_11347),
.A3(n_11349),
.B(n_11342),
.Y(n_13827)
);

INVx2_ASAP7_75t_L g13828 ( 
.A(n_12783),
.Y(n_13828)
);

BUFx2_ASAP7_75t_L g13829 ( 
.A(n_12197),
.Y(n_13829)
);

INVx1_ASAP7_75t_L g13830 ( 
.A(n_12908),
.Y(n_13830)
);

INVx1_ASAP7_75t_L g13831 ( 
.A(n_12917),
.Y(n_13831)
);

AND2x2_ASAP7_75t_L g13832 ( 
.A(n_11962),
.B(n_8500),
.Y(n_13832)
);

AND2x2_ASAP7_75t_L g13833 ( 
.A(n_12779),
.B(n_8500),
.Y(n_13833)
);

INVx2_ASAP7_75t_SL g13834 ( 
.A(n_12745),
.Y(n_13834)
);

BUFx2_ASAP7_75t_L g13835 ( 
.A(n_12218),
.Y(n_13835)
);

INVx2_ASAP7_75t_SL g13836 ( 
.A(n_12334),
.Y(n_13836)
);

NAND2xp5_ASAP7_75t_L g13837 ( 
.A(n_12052),
.B(n_11263),
.Y(n_13837)
);

NAND2xp5_ASAP7_75t_L g13838 ( 
.A(n_12327),
.B(n_11266),
.Y(n_13838)
);

AND2x2_ASAP7_75t_L g13839 ( 
.A(n_12790),
.B(n_8500),
.Y(n_13839)
);

INVx2_ASAP7_75t_L g13840 ( 
.A(n_12903),
.Y(n_13840)
);

INVxp67_ASAP7_75t_L g13841 ( 
.A(n_12534),
.Y(n_13841)
);

BUFx3_ASAP7_75t_L g13842 ( 
.A(n_12140),
.Y(n_13842)
);

AND2x2_ASAP7_75t_L g13843 ( 
.A(n_12742),
.B(n_8508),
.Y(n_13843)
);

INVx1_ASAP7_75t_L g13844 ( 
.A(n_12928),
.Y(n_13844)
);

INVx1_ASAP7_75t_L g13845 ( 
.A(n_12956),
.Y(n_13845)
);

INVx2_ASAP7_75t_L g13846 ( 
.A(n_12920),
.Y(n_13846)
);

BUFx2_ASAP7_75t_SL g13847 ( 
.A(n_12336),
.Y(n_13847)
);

INVx1_ASAP7_75t_L g13848 ( 
.A(n_12260),
.Y(n_13848)
);

INVx2_ASAP7_75t_L g13849 ( 
.A(n_12159),
.Y(n_13849)
);

AND2x2_ASAP7_75t_L g13850 ( 
.A(n_12726),
.B(n_8508),
.Y(n_13850)
);

AND2x4_ASAP7_75t_L g13851 ( 
.A(n_12942),
.B(n_11914),
.Y(n_13851)
);

AND2x4_ASAP7_75t_L g13852 ( 
.A(n_12758),
.B(n_11914),
.Y(n_13852)
);

INVx1_ASAP7_75t_L g13853 ( 
.A(n_12243),
.Y(n_13853)
);

INVx1_ASAP7_75t_L g13854 ( 
.A(n_12959),
.Y(n_13854)
);

BUFx2_ASAP7_75t_L g13855 ( 
.A(n_12146),
.Y(n_13855)
);

NAND2xp5_ASAP7_75t_L g13856 ( 
.A(n_12317),
.B(n_12133),
.Y(n_13856)
);

INVx1_ASAP7_75t_L g13857 ( 
.A(n_12868),
.Y(n_13857)
);

AND2x2_ASAP7_75t_L g13858 ( 
.A(n_12729),
.B(n_8508),
.Y(n_13858)
);

BUFx2_ASAP7_75t_L g13859 ( 
.A(n_12901),
.Y(n_13859)
);

INVx2_ASAP7_75t_L g13860 ( 
.A(n_12177),
.Y(n_13860)
);

HB1xp67_ASAP7_75t_L g13861 ( 
.A(n_12339),
.Y(n_13861)
);

INVx1_ASAP7_75t_L g13862 ( 
.A(n_12096),
.Y(n_13862)
);

INVx1_ASAP7_75t_L g13863 ( 
.A(n_12801),
.Y(n_13863)
);

OR2x2_ASAP7_75t_L g13864 ( 
.A(n_12431),
.B(n_11272),
.Y(n_13864)
);

AND2x2_ASAP7_75t_L g13865 ( 
.A(n_12330),
.B(n_8508),
.Y(n_13865)
);

INVx1_ASAP7_75t_L g13866 ( 
.A(n_12812),
.Y(n_13866)
);

INVx1_ASAP7_75t_L g13867 ( 
.A(n_12669),
.Y(n_13867)
);

INVx2_ASAP7_75t_L g13868 ( 
.A(n_12946),
.Y(n_13868)
);

BUFx3_ASAP7_75t_L g13869 ( 
.A(n_12032),
.Y(n_13869)
);

INVx1_ASAP7_75t_L g13870 ( 
.A(n_12716),
.Y(n_13870)
);

NAND2xp5_ASAP7_75t_L g13871 ( 
.A(n_12079),
.B(n_11273),
.Y(n_13871)
);

INVx1_ASAP7_75t_L g13872 ( 
.A(n_12574),
.Y(n_13872)
);

INVx2_ASAP7_75t_L g13873 ( 
.A(n_12954),
.Y(n_13873)
);

BUFx3_ASAP7_75t_L g13874 ( 
.A(n_12033),
.Y(n_13874)
);

NAND2xp5_ASAP7_75t_L g13875 ( 
.A(n_12106),
.B(n_11275),
.Y(n_13875)
);

INVx2_ASAP7_75t_L g13876 ( 
.A(n_12754),
.Y(n_13876)
);

BUFx2_ASAP7_75t_L g13877 ( 
.A(n_12150),
.Y(n_13877)
);

AND2x2_ASAP7_75t_L g13878 ( 
.A(n_12804),
.B(n_8508),
.Y(n_13878)
);

INVx1_ASAP7_75t_L g13879 ( 
.A(n_12718),
.Y(n_13879)
);

INVx1_ASAP7_75t_L g13880 ( 
.A(n_12747),
.Y(n_13880)
);

HB1xp67_ASAP7_75t_L g13881 ( 
.A(n_12445),
.Y(n_13881)
);

BUFx3_ASAP7_75t_L g13882 ( 
.A(n_12433),
.Y(n_13882)
);

AND2x2_ASAP7_75t_L g13883 ( 
.A(n_12399),
.B(n_8508),
.Y(n_13883)
);

INVx2_ASAP7_75t_L g13884 ( 
.A(n_12802),
.Y(n_13884)
);

AND2x2_ASAP7_75t_L g13885 ( 
.A(n_12404),
.B(n_12811),
.Y(n_13885)
);

AND2x2_ASAP7_75t_L g13886 ( 
.A(n_12815),
.B(n_8579),
.Y(n_13886)
);

NAND2xp5_ASAP7_75t_L g13887 ( 
.A(n_12364),
.B(n_11279),
.Y(n_13887)
);

NAND3xp33_ASAP7_75t_L g13888 ( 
.A(n_12554),
.B(n_11889),
.C(n_11865),
.Y(n_13888)
);

BUFx6f_ASAP7_75t_L g13889 ( 
.A(n_12481),
.Y(n_13889)
);

AND2x2_ASAP7_75t_L g13890 ( 
.A(n_12817),
.B(n_8579),
.Y(n_13890)
);

NAND2xp5_ASAP7_75t_L g13891 ( 
.A(n_12223),
.B(n_11283),
.Y(n_13891)
);

INVx2_ASAP7_75t_L g13892 ( 
.A(n_12810),
.Y(n_13892)
);

INVx2_ASAP7_75t_L g13893 ( 
.A(n_12839),
.Y(n_13893)
);

AND2x2_ASAP7_75t_L g13894 ( 
.A(n_12818),
.B(n_8579),
.Y(n_13894)
);

BUFx2_ASAP7_75t_SL g13895 ( 
.A(n_12365),
.Y(n_13895)
);

BUFx3_ASAP7_75t_L g13896 ( 
.A(n_12755),
.Y(n_13896)
);

INVx2_ASAP7_75t_L g13897 ( 
.A(n_12841),
.Y(n_13897)
);

INVx2_ASAP7_75t_L g13898 ( 
.A(n_12767),
.Y(n_13898)
);

INVx1_ASAP7_75t_L g13899 ( 
.A(n_12578),
.Y(n_13899)
);

INVx2_ASAP7_75t_L g13900 ( 
.A(n_12805),
.Y(n_13900)
);

AND2x4_ASAP7_75t_L g13901 ( 
.A(n_12575),
.B(n_11924),
.Y(n_13901)
);

OR2x2_ASAP7_75t_L g13902 ( 
.A(n_12621),
.B(n_11286),
.Y(n_13902)
);

AND2x2_ASAP7_75t_L g13903 ( 
.A(n_12822),
.B(n_8579),
.Y(n_13903)
);

INVx1_ASAP7_75t_L g13904 ( 
.A(n_12787),
.Y(n_13904)
);

BUFx2_ASAP7_75t_L g13905 ( 
.A(n_12109),
.Y(n_13905)
);

INVx1_ASAP7_75t_L g13906 ( 
.A(n_12809),
.Y(n_13906)
);

BUFx2_ASAP7_75t_L g13907 ( 
.A(n_12679),
.Y(n_13907)
);

INVx2_ASAP7_75t_SL g13908 ( 
.A(n_12724),
.Y(n_13908)
);

AND2x2_ASAP7_75t_L g13909 ( 
.A(n_12837),
.B(n_8579),
.Y(n_13909)
);

OR2x2_ASAP7_75t_L g13910 ( 
.A(n_12569),
.B(n_12437),
.Y(n_13910)
);

INVxp67_ASAP7_75t_SL g13911 ( 
.A(n_12048),
.Y(n_13911)
);

AND2x2_ASAP7_75t_L g13912 ( 
.A(n_12044),
.B(n_8579),
.Y(n_13912)
);

AND2x2_ASAP7_75t_L g13913 ( 
.A(n_12670),
.B(n_8615),
.Y(n_13913)
);

INVx1_ASAP7_75t_L g13914 ( 
.A(n_12709),
.Y(n_13914)
);

INVx5_ASAP7_75t_L g13915 ( 
.A(n_12388),
.Y(n_13915)
);

INVx2_ASAP7_75t_L g13916 ( 
.A(n_12862),
.Y(n_13916)
);

INVx2_ASAP7_75t_L g13917 ( 
.A(n_12700),
.Y(n_13917)
);

BUFx2_ASAP7_75t_L g13918 ( 
.A(n_12485),
.Y(n_13918)
);

NAND2xp5_ASAP7_75t_L g13919 ( 
.A(n_12168),
.B(n_11290),
.Y(n_13919)
);

AND2x2_ASAP7_75t_L g13920 ( 
.A(n_12671),
.B(n_8615),
.Y(n_13920)
);

INVx1_ASAP7_75t_L g13921 ( 
.A(n_12966),
.Y(n_13921)
);

NAND2xp5_ASAP7_75t_L g13922 ( 
.A(n_13024),
.B(n_12233),
.Y(n_13922)
);

NAND2xp5_ASAP7_75t_L g13923 ( 
.A(n_13026),
.B(n_12549),
.Y(n_13923)
);

AND2x2_ASAP7_75t_L g13924 ( 
.A(n_12969),
.B(n_12955),
.Y(n_13924)
);

INVx2_ASAP7_75t_L g13925 ( 
.A(n_13118),
.Y(n_13925)
);

AND2x2_ASAP7_75t_L g13926 ( 
.A(n_12981),
.B(n_12907),
.Y(n_13926)
);

INVxp67_ASAP7_75t_SL g13927 ( 
.A(n_12960),
.Y(n_13927)
);

AOI22xp33_ASAP7_75t_L g13928 ( 
.A1(n_13847),
.A2(n_13670),
.B1(n_13869),
.B2(n_12993),
.Y(n_13928)
);

INVx1_ASAP7_75t_L g13929 ( 
.A(n_13162),
.Y(n_13929)
);

AND2x2_ASAP7_75t_L g13930 ( 
.A(n_12967),
.B(n_12566),
.Y(n_13930)
);

HB1xp67_ASAP7_75t_L g13931 ( 
.A(n_13066),
.Y(n_13931)
);

INVx1_ASAP7_75t_L g13932 ( 
.A(n_13072),
.Y(n_13932)
);

AND2x2_ASAP7_75t_L g13933 ( 
.A(n_13027),
.B(n_12866),
.Y(n_13933)
);

AND2x2_ASAP7_75t_L g13934 ( 
.A(n_13200),
.B(n_12871),
.Y(n_13934)
);

NAND2xp5_ASAP7_75t_L g13935 ( 
.A(n_12970),
.B(n_12586),
.Y(n_13935)
);

INVx1_ASAP7_75t_L g13936 ( 
.A(n_13091),
.Y(n_13936)
);

AND2x2_ASAP7_75t_L g13937 ( 
.A(n_13085),
.B(n_12881),
.Y(n_13937)
);

AND2x2_ASAP7_75t_L g13938 ( 
.A(n_13405),
.B(n_12883),
.Y(n_13938)
);

INVxp67_ASAP7_75t_SL g13939 ( 
.A(n_12996),
.Y(n_13939)
);

NAND2xp5_ASAP7_75t_L g13940 ( 
.A(n_13342),
.B(n_12464),
.Y(n_13940)
);

INVx1_ASAP7_75t_L g13941 ( 
.A(n_13093),
.Y(n_13941)
);

OAI22xp33_ASAP7_75t_L g13942 ( 
.A1(n_13915),
.A2(n_12212),
.B1(n_12263),
.B2(n_12035),
.Y(n_13942)
);

AND2x2_ASAP7_75t_L g13943 ( 
.A(n_13186),
.B(n_12885),
.Y(n_13943)
);

AND2x2_ASAP7_75t_L g13944 ( 
.A(n_13192),
.B(n_12900),
.Y(n_13944)
);

AND2x2_ASAP7_75t_L g13945 ( 
.A(n_12964),
.B(n_12768),
.Y(n_13945)
);

AND2x4_ASAP7_75t_L g13946 ( 
.A(n_13037),
.B(n_11924),
.Y(n_13946)
);

BUFx2_ASAP7_75t_L g13947 ( 
.A(n_13037),
.Y(n_13947)
);

INVx2_ASAP7_75t_L g13948 ( 
.A(n_13284),
.Y(n_13948)
);

AND2x2_ASAP7_75t_L g13949 ( 
.A(n_12984),
.B(n_12774),
.Y(n_13949)
);

INVx2_ASAP7_75t_L g13950 ( 
.A(n_13302),
.Y(n_13950)
);

INVx2_ASAP7_75t_L g13951 ( 
.A(n_13041),
.Y(n_13951)
);

INVx1_ASAP7_75t_L g13952 ( 
.A(n_13096),
.Y(n_13952)
);

AND2x2_ASAP7_75t_L g13953 ( 
.A(n_12984),
.B(n_12328),
.Y(n_13953)
);

NAND2xp5_ASAP7_75t_L g13954 ( 
.A(n_12972),
.B(n_12880),
.Y(n_13954)
);

NAND2xp33_ASAP7_75t_L g13955 ( 
.A(n_13915),
.B(n_12504),
.Y(n_13955)
);

AND2x4_ASAP7_75t_L g13956 ( 
.A(n_13106),
.B(n_11924),
.Y(n_13956)
);

AOI22xp33_ASAP7_75t_L g13957 ( 
.A1(n_13847),
.A2(n_12320),
.B1(n_12215),
.B2(n_12124),
.Y(n_13957)
);

INVx1_ASAP7_75t_L g13958 ( 
.A(n_13104),
.Y(n_13958)
);

INVx1_ASAP7_75t_L g13959 ( 
.A(n_13122),
.Y(n_13959)
);

AOI22xp33_ASAP7_75t_L g13960 ( 
.A1(n_13874),
.A2(n_12450),
.B1(n_11991),
.B2(n_12444),
.Y(n_13960)
);

INVx1_ASAP7_75t_L g13961 ( 
.A(n_13128),
.Y(n_13961)
);

INVx1_ASAP7_75t_SL g13962 ( 
.A(n_13058),
.Y(n_13962)
);

AOI22xp33_ASAP7_75t_L g13963 ( 
.A1(n_13811),
.A2(n_12181),
.B1(n_12222),
.B2(n_12203),
.Y(n_13963)
);

AND2x4_ASAP7_75t_L g13964 ( 
.A(n_13106),
.B(n_10602),
.Y(n_13964)
);

HB1xp67_ASAP7_75t_L g13965 ( 
.A(n_13352),
.Y(n_13965)
);

AND2x2_ASAP7_75t_L g13966 ( 
.A(n_12997),
.B(n_12567),
.Y(n_13966)
);

INVx1_ASAP7_75t_L g13967 ( 
.A(n_13137),
.Y(n_13967)
);

INVx1_ASAP7_75t_L g13968 ( 
.A(n_13161),
.Y(n_13968)
);

INVx1_ASAP7_75t_L g13969 ( 
.A(n_13034),
.Y(n_13969)
);

NOR2xp33_ASAP7_75t_L g13970 ( 
.A(n_13014),
.B(n_12878),
.Y(n_13970)
);

NOR2x1_ASAP7_75t_L g13971 ( 
.A(n_13491),
.B(n_12897),
.Y(n_13971)
);

NAND2xp5_ASAP7_75t_L g13972 ( 
.A(n_13388),
.B(n_12477),
.Y(n_13972)
);

INVx1_ASAP7_75t_L g13973 ( 
.A(n_13034),
.Y(n_13973)
);

INVx1_ASAP7_75t_L g13974 ( 
.A(n_12961),
.Y(n_13974)
);

INVx1_ASAP7_75t_L g13975 ( 
.A(n_12961),
.Y(n_13975)
);

INVx2_ASAP7_75t_L g13976 ( 
.A(n_13262),
.Y(n_13976)
);

INVx1_ASAP7_75t_L g13977 ( 
.A(n_12990),
.Y(n_13977)
);

AOI22xp33_ASAP7_75t_L g13978 ( 
.A1(n_13915),
.A2(n_12226),
.B1(n_12462),
.B2(n_12306),
.Y(n_13978)
);

INVx3_ASAP7_75t_L g13979 ( 
.A(n_13016),
.Y(n_13979)
);

INVx2_ASAP7_75t_L g13980 ( 
.A(n_13262),
.Y(n_13980)
);

OR2x2_ASAP7_75t_L g13981 ( 
.A(n_13761),
.B(n_12120),
.Y(n_13981)
);

AOI22xp33_ASAP7_75t_SL g13982 ( 
.A1(n_13895),
.A2(n_13789),
.B1(n_13578),
.B2(n_13877),
.Y(n_13982)
);

INVx1_ASAP7_75t_L g13983 ( 
.A(n_12990),
.Y(n_13983)
);

AND2x2_ASAP7_75t_L g13984 ( 
.A(n_13046),
.B(n_12571),
.Y(n_13984)
);

AOI22xp33_ASAP7_75t_L g13985 ( 
.A1(n_13810),
.A2(n_12324),
.B1(n_12599),
.B2(n_12595),
.Y(n_13985)
);

INVx2_ASAP7_75t_SL g13986 ( 
.A(n_12996),
.Y(n_13986)
);

OAI21xp5_ASAP7_75t_L g13987 ( 
.A1(n_13711),
.A2(n_12826),
.B(n_12164),
.Y(n_13987)
);

NAND2xp5_ASAP7_75t_L g13988 ( 
.A(n_13107),
.B(n_12526),
.Y(n_13988)
);

OR2x2_ASAP7_75t_L g13989 ( 
.A(n_13747),
.B(n_12121),
.Y(n_13989)
);

AND2x2_ASAP7_75t_L g13990 ( 
.A(n_13021),
.B(n_12752),
.Y(n_13990)
);

NAND2x1_ASAP7_75t_L g13991 ( 
.A(n_13038),
.B(n_12658),
.Y(n_13991)
);

INVx1_ASAP7_75t_L g13992 ( 
.A(n_13000),
.Y(n_13992)
);

INVx2_ASAP7_75t_L g13993 ( 
.A(n_12996),
.Y(n_13993)
);

OR2x2_ASAP7_75t_L g13994 ( 
.A(n_13170),
.B(n_12465),
.Y(n_13994)
);

INVx2_ASAP7_75t_L g13995 ( 
.A(n_13022),
.Y(n_13995)
);

INVx1_ASAP7_75t_L g13996 ( 
.A(n_13000),
.Y(n_13996)
);

AOI222xp33_ASAP7_75t_L g13997 ( 
.A1(n_13856),
.A2(n_12156),
.B1(n_12617),
.B2(n_12592),
.C1(n_12647),
.C2(n_12627),
.Y(n_13997)
);

NOR2xp33_ASAP7_75t_SL g13998 ( 
.A(n_13058),
.B(n_12516),
.Y(n_13998)
);

AND2x4_ASAP7_75t_L g13999 ( 
.A(n_13201),
.B(n_10625),
.Y(n_13999)
);

NAND2xp5_ASAP7_75t_L g14000 ( 
.A(n_13111),
.B(n_12474),
.Y(n_14000)
);

INVx2_ASAP7_75t_L g14001 ( 
.A(n_13022),
.Y(n_14001)
);

INVx2_ASAP7_75t_L g14002 ( 
.A(n_13022),
.Y(n_14002)
);

NAND2xp5_ASAP7_75t_L g14003 ( 
.A(n_13013),
.B(n_12838),
.Y(n_14003)
);

INVx2_ASAP7_75t_L g14004 ( 
.A(n_13331),
.Y(n_14004)
);

INVx1_ASAP7_75t_L g14005 ( 
.A(n_13003),
.Y(n_14005)
);

OR2x2_ASAP7_75t_L g14006 ( 
.A(n_13796),
.B(n_12442),
.Y(n_14006)
);

AND2x2_ASAP7_75t_L g14007 ( 
.A(n_13078),
.B(n_12429),
.Y(n_14007)
);

AOI22xp33_ASAP7_75t_L g14008 ( 
.A1(n_13769),
.A2(n_12482),
.B1(n_12714),
.B2(n_12705),
.Y(n_14008)
);

INVx2_ASAP7_75t_L g14009 ( 
.A(n_13331),
.Y(n_14009)
);

AOI22xp33_ASAP7_75t_L g14010 ( 
.A1(n_13789),
.A2(n_12583),
.B1(n_12593),
.B2(n_12503),
.Y(n_14010)
);

NAND2xp5_ASAP7_75t_L g14011 ( 
.A(n_13015),
.B(n_12931),
.Y(n_14011)
);

NOR2xp33_ASAP7_75t_L g14012 ( 
.A(n_12998),
.B(n_12559),
.Y(n_14012)
);

BUFx2_ASAP7_75t_L g14013 ( 
.A(n_13674),
.Y(n_14013)
);

INVx4_ASAP7_75t_L g14014 ( 
.A(n_13331),
.Y(n_14014)
);

INVx2_ASAP7_75t_L g14015 ( 
.A(n_13456),
.Y(n_14015)
);

INVxp67_ASAP7_75t_SL g14016 ( 
.A(n_13695),
.Y(n_14016)
);

NOR2xp33_ASAP7_75t_L g14017 ( 
.A(n_12998),
.B(n_13389),
.Y(n_14017)
);

AOI22xp33_ASAP7_75t_L g14018 ( 
.A1(n_13799),
.A2(n_12387),
.B1(n_12436),
.B2(n_12435),
.Y(n_14018)
);

AND2x2_ASAP7_75t_L g14019 ( 
.A(n_13248),
.B(n_12858),
.Y(n_14019)
);

INVx2_ASAP7_75t_L g14020 ( 
.A(n_13456),
.Y(n_14020)
);

NAND2xp5_ASAP7_75t_SL g14021 ( 
.A(n_13813),
.B(n_13323),
.Y(n_14021)
);

INVx1_ASAP7_75t_L g14022 ( 
.A(n_13003),
.Y(n_14022)
);

INVx1_ASAP7_75t_L g14023 ( 
.A(n_13005),
.Y(n_14023)
);

AND2x4_ASAP7_75t_L g14024 ( 
.A(n_13201),
.B(n_10625),
.Y(n_14024)
);

INVx1_ASAP7_75t_L g14025 ( 
.A(n_13005),
.Y(n_14025)
);

INVx1_ASAP7_75t_L g14026 ( 
.A(n_13006),
.Y(n_14026)
);

OR2x2_ASAP7_75t_L g14027 ( 
.A(n_13591),
.B(n_12763),
.Y(n_14027)
);

AND2x2_ASAP7_75t_L g14028 ( 
.A(n_13135),
.B(n_12916),
.Y(n_14028)
);

INVx1_ASAP7_75t_L g14029 ( 
.A(n_13006),
.Y(n_14029)
);

INVx1_ASAP7_75t_L g14030 ( 
.A(n_13011),
.Y(n_14030)
);

INVx2_ASAP7_75t_L g14031 ( 
.A(n_13456),
.Y(n_14031)
);

AOI22xp5_ASAP7_75t_L g14032 ( 
.A1(n_13862),
.A2(n_12379),
.B1(n_12490),
.B2(n_12487),
.Y(n_14032)
);

HB1xp67_ASAP7_75t_L g14033 ( 
.A(n_13423),
.Y(n_14033)
);

INVx2_ASAP7_75t_L g14034 ( 
.A(n_13038),
.Y(n_14034)
);

OR2x2_ASAP7_75t_L g14035 ( 
.A(n_13012),
.B(n_11297),
.Y(n_14035)
);

AOI22xp33_ASAP7_75t_L g14036 ( 
.A1(n_13666),
.A2(n_12515),
.B1(n_12844),
.B2(n_12686),
.Y(n_14036)
);

INVx1_ASAP7_75t_L g14037 ( 
.A(n_13011),
.Y(n_14037)
);

NOR2xp33_ASAP7_75t_L g14038 ( 
.A(n_13389),
.B(n_12633),
.Y(n_14038)
);

OAI22xp5_ASAP7_75t_L g14039 ( 
.A1(n_13298),
.A2(n_12940),
.B1(n_12921),
.B2(n_12944),
.Y(n_14039)
);

INVx2_ASAP7_75t_L g14040 ( 
.A(n_13234),
.Y(n_14040)
);

AND2x4_ASAP7_75t_L g14041 ( 
.A(n_13258),
.B(n_10625),
.Y(n_14041)
);

INVx1_ASAP7_75t_L g14042 ( 
.A(n_13023),
.Y(n_14042)
);

INVxp67_ASAP7_75t_SL g14043 ( 
.A(n_13286),
.Y(n_14043)
);

INVx1_ASAP7_75t_L g14044 ( 
.A(n_13023),
.Y(n_14044)
);

INVx2_ASAP7_75t_L g14045 ( 
.A(n_13234),
.Y(n_14045)
);

AND2x2_ASAP7_75t_L g14046 ( 
.A(n_13108),
.B(n_12708),
.Y(n_14046)
);

INVx1_ASAP7_75t_L g14047 ( 
.A(n_13031),
.Y(n_14047)
);

NOR2x1_ASAP7_75t_SL g14048 ( 
.A(n_13619),
.B(n_12138),
.Y(n_14048)
);

NAND2x1p5_ASAP7_75t_L g14049 ( 
.A(n_13323),
.B(n_7757),
.Y(n_14049)
);

NAND2x1p5_ASAP7_75t_L g14050 ( 
.A(n_13323),
.B(n_7757),
.Y(n_14050)
);

AND2x4_ASAP7_75t_L g14051 ( 
.A(n_13207),
.B(n_10625),
.Y(n_14051)
);

OR2x2_ASAP7_75t_L g14052 ( 
.A(n_13784),
.B(n_11298),
.Y(n_14052)
);

INVx2_ASAP7_75t_L g14053 ( 
.A(n_13280),
.Y(n_14053)
);

BUFx2_ASAP7_75t_L g14054 ( 
.A(n_13440),
.Y(n_14054)
);

INVx1_ASAP7_75t_L g14055 ( 
.A(n_13031),
.Y(n_14055)
);

AND2x2_ASAP7_75t_L g14056 ( 
.A(n_13153),
.B(n_12565),
.Y(n_14056)
);

INVx1_ASAP7_75t_L g14057 ( 
.A(n_13175),
.Y(n_14057)
);

INVx2_ASAP7_75t_L g14058 ( 
.A(n_13280),
.Y(n_14058)
);

NAND2xp5_ASAP7_75t_L g14059 ( 
.A(n_13056),
.B(n_11306),
.Y(n_14059)
);

INVx2_ASAP7_75t_L g14060 ( 
.A(n_13332),
.Y(n_14060)
);

INVx3_ASAP7_75t_L g14061 ( 
.A(n_13307),
.Y(n_14061)
);

INVx1_ASAP7_75t_L g14062 ( 
.A(n_13198),
.Y(n_14062)
);

INVx1_ASAP7_75t_L g14063 ( 
.A(n_13209),
.Y(n_14063)
);

INVx1_ASAP7_75t_L g14064 ( 
.A(n_13210),
.Y(n_14064)
);

INVx1_ASAP7_75t_L g14065 ( 
.A(n_13221),
.Y(n_14065)
);

NAND2xp5_ASAP7_75t_L g14066 ( 
.A(n_13059),
.B(n_11307),
.Y(n_14066)
);

AND2x2_ASAP7_75t_L g14067 ( 
.A(n_13156),
.B(n_10629),
.Y(n_14067)
);

INVx2_ASAP7_75t_L g14068 ( 
.A(n_13332),
.Y(n_14068)
);

AND2x2_ASAP7_75t_L g14069 ( 
.A(n_13109),
.B(n_13447),
.Y(n_14069)
);

INVx4_ASAP7_75t_L g14070 ( 
.A(n_13307),
.Y(n_14070)
);

INVx1_ASAP7_75t_L g14071 ( 
.A(n_13245),
.Y(n_14071)
);

INVx3_ASAP7_75t_L g14072 ( 
.A(n_13307),
.Y(n_14072)
);

AND3x1_ASAP7_75t_L g14073 ( 
.A(n_13385),
.B(n_12656),
.C(n_12649),
.Y(n_14073)
);

NAND2xp5_ASAP7_75t_L g14074 ( 
.A(n_13060),
.B(n_11311),
.Y(n_14074)
);

CKINVDCx5p33_ASAP7_75t_R g14075 ( 
.A(n_12962),
.Y(n_14075)
);

OR2x2_ASAP7_75t_L g14076 ( 
.A(n_13071),
.B(n_11316),
.Y(n_14076)
);

NOR2xp33_ASAP7_75t_L g14077 ( 
.A(n_13185),
.B(n_12719),
.Y(n_14077)
);

HB1xp67_ASAP7_75t_L g14078 ( 
.A(n_13566),
.Y(n_14078)
);

INVx1_ASAP7_75t_SL g14079 ( 
.A(n_12971),
.Y(n_14079)
);

INVx2_ASAP7_75t_L g14080 ( 
.A(n_13371),
.Y(n_14080)
);

NAND2xp5_ASAP7_75t_L g14081 ( 
.A(n_13061),
.B(n_11324),
.Y(n_14081)
);

INVx2_ASAP7_75t_L g14082 ( 
.A(n_13371),
.Y(n_14082)
);

NAND2xp5_ASAP7_75t_L g14083 ( 
.A(n_13065),
.B(n_11327),
.Y(n_14083)
);

NAND2xp5_ASAP7_75t_L g14084 ( 
.A(n_13073),
.B(n_11328),
.Y(n_14084)
);

OR2x2_ASAP7_75t_L g14085 ( 
.A(n_13335),
.B(n_11330),
.Y(n_14085)
);

AND2x4_ASAP7_75t_L g14086 ( 
.A(n_13197),
.B(n_10629),
.Y(n_14086)
);

AOI221xp5_ASAP7_75t_L g14087 ( 
.A1(n_13862),
.A2(n_13033),
.B1(n_13841),
.B2(n_13632),
.C(n_13734),
.Y(n_14087)
);

AND2x2_ASAP7_75t_L g14088 ( 
.A(n_13116),
.B(n_13119),
.Y(n_14088)
);

BUFx3_ASAP7_75t_L g14089 ( 
.A(n_13008),
.Y(n_14089)
);

INVx2_ASAP7_75t_L g14090 ( 
.A(n_13424),
.Y(n_14090)
);

INVx1_ASAP7_75t_L g14091 ( 
.A(n_13257),
.Y(n_14091)
);

INVx1_ASAP7_75t_L g14092 ( 
.A(n_13270),
.Y(n_14092)
);

INVx1_ASAP7_75t_L g14093 ( 
.A(n_13271),
.Y(n_14093)
);

AND2x2_ASAP7_75t_L g14094 ( 
.A(n_13126),
.B(n_10629),
.Y(n_14094)
);

AND2x2_ASAP7_75t_L g14095 ( 
.A(n_13133),
.B(n_10629),
.Y(n_14095)
);

NAND2xp5_ASAP7_75t_L g14096 ( 
.A(n_13074),
.B(n_11332),
.Y(n_14096)
);

AND2x2_ASAP7_75t_L g14097 ( 
.A(n_12986),
.B(n_10665),
.Y(n_14097)
);

AND2x2_ASAP7_75t_L g14098 ( 
.A(n_13007),
.B(n_10665),
.Y(n_14098)
);

AOI22xp33_ASAP7_75t_L g14099 ( 
.A1(n_13882),
.A2(n_12608),
.B1(n_12860),
.B2(n_12717),
.Y(n_14099)
);

AND2x2_ASAP7_75t_L g14100 ( 
.A(n_13007),
.B(n_10665),
.Y(n_14100)
);

INVx1_ASAP7_75t_L g14101 ( 
.A(n_13358),
.Y(n_14101)
);

INVx1_ASAP7_75t_L g14102 ( 
.A(n_13366),
.Y(n_14102)
);

HB1xp67_ASAP7_75t_L g14103 ( 
.A(n_13606),
.Y(n_14103)
);

INVx1_ASAP7_75t_L g14104 ( 
.A(n_13607),
.Y(n_14104)
);

NOR2xp67_ASAP7_75t_L g14105 ( 
.A(n_13813),
.B(n_12776),
.Y(n_14105)
);

INVx1_ASAP7_75t_L g14106 ( 
.A(n_12965),
.Y(n_14106)
);

INVx1_ASAP7_75t_L g14107 ( 
.A(n_12968),
.Y(n_14107)
);

AND2x4_ASAP7_75t_L g14108 ( 
.A(n_13197),
.B(n_13281),
.Y(n_14108)
);

AND2x4_ASAP7_75t_SL g14109 ( 
.A(n_13042),
.B(n_8210),
.Y(n_14109)
);

AND2x2_ASAP7_75t_L g14110 ( 
.A(n_12989),
.B(n_10665),
.Y(n_14110)
);

AND2x2_ASAP7_75t_L g14111 ( 
.A(n_12991),
.B(n_11336),
.Y(n_14111)
);

INVx1_ASAP7_75t_L g14112 ( 
.A(n_12976),
.Y(n_14112)
);

AND2x2_ASAP7_75t_L g14113 ( 
.A(n_12995),
.B(n_11344),
.Y(n_14113)
);

INVx1_ASAP7_75t_L g14114 ( 
.A(n_12977),
.Y(n_14114)
);

OR2x2_ASAP7_75t_L g14115 ( 
.A(n_13052),
.B(n_11352),
.Y(n_14115)
);

INVx2_ASAP7_75t_L g14116 ( 
.A(n_13424),
.Y(n_14116)
);

AND2x2_ASAP7_75t_L g14117 ( 
.A(n_13009),
.B(n_11356),
.Y(n_14117)
);

OR2x2_ASAP7_75t_L g14118 ( 
.A(n_13902),
.B(n_11358),
.Y(n_14118)
);

AND2x2_ASAP7_75t_L g14119 ( 
.A(n_13182),
.B(n_11366),
.Y(n_14119)
);

AND2x2_ASAP7_75t_L g14120 ( 
.A(n_13189),
.B(n_11369),
.Y(n_14120)
);

INVx1_ASAP7_75t_L g14121 ( 
.A(n_12978),
.Y(n_14121)
);

AND2x2_ASAP7_75t_L g14122 ( 
.A(n_13134),
.B(n_11372),
.Y(n_14122)
);

INVx1_ASAP7_75t_L g14123 ( 
.A(n_13259),
.Y(n_14123)
);

NAND2xp5_ASAP7_75t_L g14124 ( 
.A(n_13076),
.B(n_11378),
.Y(n_14124)
);

AND2x2_ASAP7_75t_L g14125 ( 
.A(n_13420),
.B(n_11383),
.Y(n_14125)
);

OR2x2_ASAP7_75t_L g14126 ( 
.A(n_13736),
.B(n_11388),
.Y(n_14126)
);

NAND2xp5_ASAP7_75t_L g14127 ( 
.A(n_13097),
.B(n_11390),
.Y(n_14127)
);

INVx1_ASAP7_75t_L g14128 ( 
.A(n_13259),
.Y(n_14128)
);

HB1xp67_ASAP7_75t_L g14129 ( 
.A(n_13483),
.Y(n_14129)
);

INVx1_ASAP7_75t_L g14130 ( 
.A(n_13265),
.Y(n_14130)
);

NOR2xp33_ASAP7_75t_L g14131 ( 
.A(n_13252),
.B(n_12143),
.Y(n_14131)
);

AND2x4_ASAP7_75t_SL g14132 ( 
.A(n_13286),
.B(n_8210),
.Y(n_14132)
);

HB1xp67_ASAP7_75t_L g14133 ( 
.A(n_13483),
.Y(n_14133)
);

INVxp67_ASAP7_75t_L g14134 ( 
.A(n_13578),
.Y(n_14134)
);

OR2x2_ASAP7_75t_L g14135 ( 
.A(n_13736),
.B(n_11391),
.Y(n_14135)
);

NAND2xp5_ASAP7_75t_L g14136 ( 
.A(n_13098),
.B(n_11395),
.Y(n_14136)
);

INVx1_ASAP7_75t_L g14137 ( 
.A(n_13265),
.Y(n_14137)
);

INVx3_ASAP7_75t_L g14138 ( 
.A(n_13286),
.Y(n_14138)
);

AND2x2_ASAP7_75t_L g14139 ( 
.A(n_13055),
.B(n_11397),
.Y(n_14139)
);

INVx4_ASAP7_75t_L g14140 ( 
.A(n_13264),
.Y(n_14140)
);

INVxp67_ASAP7_75t_SL g14141 ( 
.A(n_13356),
.Y(n_14141)
);

AND2x2_ASAP7_75t_L g14142 ( 
.A(n_13163),
.B(n_11399),
.Y(n_14142)
);

INVxp33_ASAP7_75t_L g14143 ( 
.A(n_13129),
.Y(n_14143)
);

NAND2xp5_ASAP7_75t_L g14144 ( 
.A(n_13100),
.B(n_11420),
.Y(n_14144)
);

AND2x4_ASAP7_75t_SL g14145 ( 
.A(n_13264),
.B(n_13434),
.Y(n_14145)
);

HB1xp67_ASAP7_75t_L g14146 ( 
.A(n_13491),
.Y(n_14146)
);

INVx1_ASAP7_75t_L g14147 ( 
.A(n_13269),
.Y(n_14147)
);

AND2x2_ASAP7_75t_L g14148 ( 
.A(n_13330),
.B(n_11422),
.Y(n_14148)
);

AND2x2_ASAP7_75t_L g14149 ( 
.A(n_13290),
.B(n_11426),
.Y(n_14149)
);

AOI221xp5_ASAP7_75t_L g14150 ( 
.A1(n_13734),
.A2(n_12941),
.B1(n_12873),
.B2(n_12919),
.C(n_12213),
.Y(n_14150)
);

OR2x2_ASAP7_75t_L g14151 ( 
.A(n_13864),
.B(n_11428),
.Y(n_14151)
);

INVx1_ASAP7_75t_L g14152 ( 
.A(n_13269),
.Y(n_14152)
);

OR2x2_ASAP7_75t_L g14153 ( 
.A(n_13049),
.B(n_11432),
.Y(n_14153)
);

BUFx4f_ASAP7_75t_L g14154 ( 
.A(n_13264),
.Y(n_14154)
);

OR2x2_ASAP7_75t_L g14155 ( 
.A(n_13776),
.B(n_11435),
.Y(n_14155)
);

AOI22xp33_ASAP7_75t_L g14156 ( 
.A1(n_13855),
.A2(n_12761),
.B1(n_12777),
.B2(n_12739),
.Y(n_14156)
);

AND2x2_ASAP7_75t_L g14157 ( 
.A(n_13443),
.B(n_11436),
.Y(n_14157)
);

OR2x2_ASAP7_75t_L g14158 ( 
.A(n_13001),
.B(n_11438),
.Y(n_14158)
);

INVx2_ASAP7_75t_L g14159 ( 
.A(n_13256),
.Y(n_14159)
);

INVx1_ASAP7_75t_L g14160 ( 
.A(n_13272),
.Y(n_14160)
);

INVx1_ASAP7_75t_L g14161 ( 
.A(n_13272),
.Y(n_14161)
);

INVx1_ASAP7_75t_L g14162 ( 
.A(n_13285),
.Y(n_14162)
);

OAI21xp5_ASAP7_75t_L g14163 ( 
.A1(n_13266),
.A2(n_12209),
.B(n_12190),
.Y(n_14163)
);

OAI22xp5_ASAP7_75t_L g14164 ( 
.A1(n_13523),
.A2(n_12927),
.B1(n_12930),
.B2(n_12749),
.Y(n_14164)
);

INVxp67_ASAP7_75t_SL g14165 ( 
.A(n_13032),
.Y(n_14165)
);

AND2x4_ASAP7_75t_L g14166 ( 
.A(n_13166),
.B(n_13203),
.Y(n_14166)
);

OR2x2_ASAP7_75t_L g14167 ( 
.A(n_13738),
.B(n_11442),
.Y(n_14167)
);

BUFx2_ASAP7_75t_L g14168 ( 
.A(n_13166),
.Y(n_14168)
);

AND2x2_ASAP7_75t_L g14169 ( 
.A(n_13443),
.B(n_11444),
.Y(n_14169)
);

AND2x2_ASAP7_75t_L g14170 ( 
.A(n_13446),
.B(n_11449),
.Y(n_14170)
);

BUFx6f_ASAP7_75t_L g14171 ( 
.A(n_13361),
.Y(n_14171)
);

INVx2_ASAP7_75t_L g14172 ( 
.A(n_13256),
.Y(n_14172)
);

INVx2_ASAP7_75t_L g14173 ( 
.A(n_13255),
.Y(n_14173)
);

AND2x2_ASAP7_75t_L g14174 ( 
.A(n_13360),
.B(n_11454),
.Y(n_14174)
);

AND2x2_ASAP7_75t_L g14175 ( 
.A(n_13260),
.B(n_11458),
.Y(n_14175)
);

INVx1_ASAP7_75t_L g14176 ( 
.A(n_13285),
.Y(n_14176)
);

INVxp67_ASAP7_75t_SL g14177 ( 
.A(n_13095),
.Y(n_14177)
);

INVx2_ASAP7_75t_L g14178 ( 
.A(n_13255),
.Y(n_14178)
);

AND2x2_ASAP7_75t_L g14179 ( 
.A(n_13506),
.B(n_13165),
.Y(n_14179)
);

AND2x2_ASAP7_75t_L g14180 ( 
.A(n_13183),
.B(n_11460),
.Y(n_14180)
);

INVx1_ASAP7_75t_L g14181 ( 
.A(n_13288),
.Y(n_14181)
);

AOI22xp33_ASAP7_75t_SL g14182 ( 
.A1(n_13895),
.A2(n_12375),
.B1(n_12874),
.B2(n_12524),
.Y(n_14182)
);

AND2x2_ASAP7_75t_L g14183 ( 
.A(n_13397),
.B(n_11463),
.Y(n_14183)
);

AND2x2_ASAP7_75t_L g14184 ( 
.A(n_13426),
.B(n_13427),
.Y(n_14184)
);

INVx2_ASAP7_75t_L g14185 ( 
.A(n_13386),
.Y(n_14185)
);

INVx1_ASAP7_75t_L g14186 ( 
.A(n_13288),
.Y(n_14186)
);

NAND2xp5_ASAP7_75t_L g14187 ( 
.A(n_13102),
.B(n_11472),
.Y(n_14187)
);

INVx1_ASAP7_75t_L g14188 ( 
.A(n_13294),
.Y(n_14188)
);

NAND2xp5_ASAP7_75t_L g14189 ( 
.A(n_13103),
.B(n_11474),
.Y(n_14189)
);

AND2x4_ASAP7_75t_L g14190 ( 
.A(n_13203),
.B(n_9223),
.Y(n_14190)
);

INVx2_ASAP7_75t_L g14191 ( 
.A(n_13386),
.Y(n_14191)
);

AND2x2_ASAP7_75t_L g14192 ( 
.A(n_13152),
.B(n_11481),
.Y(n_14192)
);

AND2x2_ASAP7_75t_L g14193 ( 
.A(n_13608),
.B(n_11485),
.Y(n_14193)
);

AND2x2_ASAP7_75t_L g14194 ( 
.A(n_13608),
.B(n_11486),
.Y(n_14194)
);

NAND2xp5_ASAP7_75t_L g14195 ( 
.A(n_13146),
.B(n_11487),
.Y(n_14195)
);

OR2x2_ASAP7_75t_L g14196 ( 
.A(n_13471),
.B(n_11489),
.Y(n_14196)
);

INVx1_ASAP7_75t_L g14197 ( 
.A(n_13294),
.Y(n_14197)
);

INVx1_ASAP7_75t_L g14198 ( 
.A(n_13297),
.Y(n_14198)
);

OAI21xp5_ASAP7_75t_L g14199 ( 
.A1(n_13699),
.A2(n_12875),
.B(n_12852),
.Y(n_14199)
);

NAND2xp5_ASAP7_75t_L g14200 ( 
.A(n_13092),
.B(n_11492),
.Y(n_14200)
);

INVx2_ASAP7_75t_L g14201 ( 
.A(n_13402),
.Y(n_14201)
);

INVx1_ASAP7_75t_L g14202 ( 
.A(n_13297),
.Y(n_14202)
);

HB1xp67_ASAP7_75t_L g14203 ( 
.A(n_13494),
.Y(n_14203)
);

HB1xp67_ASAP7_75t_L g14204 ( 
.A(n_13494),
.Y(n_14204)
);

INVx1_ASAP7_75t_L g14205 ( 
.A(n_13301),
.Y(n_14205)
);

INVx2_ASAP7_75t_L g14206 ( 
.A(n_13402),
.Y(n_14206)
);

INVx2_ASAP7_75t_L g14207 ( 
.A(n_12982),
.Y(n_14207)
);

INVx1_ASAP7_75t_L g14208 ( 
.A(n_13301),
.Y(n_14208)
);

INVx1_ASAP7_75t_L g14209 ( 
.A(n_13618),
.Y(n_14209)
);

INVx1_ASAP7_75t_L g14210 ( 
.A(n_13626),
.Y(n_14210)
);

INVx1_ASAP7_75t_SL g14211 ( 
.A(n_13017),
.Y(n_14211)
);

AND2x2_ASAP7_75t_L g14212 ( 
.A(n_13375),
.B(n_11493),
.Y(n_14212)
);

AND2x2_ASAP7_75t_L g14213 ( 
.A(n_13247),
.B(n_11494),
.Y(n_14213)
);

NOR2x1_ASAP7_75t_SL g14214 ( 
.A(n_13619),
.B(n_10742),
.Y(n_14214)
);

AND2x4_ASAP7_75t_L g14215 ( 
.A(n_13154),
.B(n_9223),
.Y(n_14215)
);

OR2x2_ASAP7_75t_L g14216 ( 
.A(n_13336),
.B(n_13760),
.Y(n_14216)
);

NOR3xp33_ASAP7_75t_L g14217 ( 
.A(n_13149),
.B(n_12710),
.C(n_12690),
.Y(n_14217)
);

AOI22xp33_ASAP7_75t_L g14218 ( 
.A1(n_13737),
.A2(n_12886),
.B1(n_12830),
.B2(n_8574),
.Y(n_14218)
);

HB1xp67_ASAP7_75t_L g14219 ( 
.A(n_13289),
.Y(n_14219)
);

INVx1_ASAP7_75t_L g14220 ( 
.A(n_13039),
.Y(n_14220)
);

INVxp67_ASAP7_75t_SL g14221 ( 
.A(n_13547),
.Y(n_14221)
);

INVx1_ASAP7_75t_L g14222 ( 
.A(n_13039),
.Y(n_14222)
);

AND2x2_ASAP7_75t_L g14223 ( 
.A(n_13490),
.B(n_11498),
.Y(n_14223)
);

AND2x2_ASAP7_75t_L g14224 ( 
.A(n_13501),
.B(n_11503),
.Y(n_14224)
);

INVx2_ASAP7_75t_L g14225 ( 
.A(n_12982),
.Y(n_14225)
);

OAI22xp5_ASAP7_75t_L g14226 ( 
.A1(n_13910),
.A2(n_12548),
.B1(n_12771),
.B2(n_8142),
.Y(n_14226)
);

HB1xp67_ASAP7_75t_L g14227 ( 
.A(n_13295),
.Y(n_14227)
);

INVx1_ASAP7_75t_L g14228 ( 
.A(n_13043),
.Y(n_14228)
);

AOI22xp33_ASAP7_75t_L g14229 ( 
.A1(n_13737),
.A2(n_8574),
.B1(n_8150),
.B2(n_10415),
.Y(n_14229)
);

AOI21xp5_ASAP7_75t_SL g14230 ( 
.A1(n_13160),
.A2(n_12843),
.B(n_12949),
.Y(n_14230)
);

AND2x2_ASAP7_75t_L g14231 ( 
.A(n_13171),
.B(n_11516),
.Y(n_14231)
);

NAND2xp5_ASAP7_75t_L g14232 ( 
.A(n_13241),
.B(n_11518),
.Y(n_14232)
);

INVx2_ASAP7_75t_L g14233 ( 
.A(n_12992),
.Y(n_14233)
);

AND2x4_ASAP7_75t_L g14234 ( 
.A(n_13434),
.B(n_11521),
.Y(n_14234)
);

BUFx3_ASAP7_75t_L g14235 ( 
.A(n_13277),
.Y(n_14235)
);

INVx2_ASAP7_75t_L g14236 ( 
.A(n_12992),
.Y(n_14236)
);

AND2x4_ASAP7_75t_L g14237 ( 
.A(n_13362),
.B(n_13364),
.Y(n_14237)
);

HB1xp67_ASAP7_75t_L g14238 ( 
.A(n_13299),
.Y(n_14238)
);

AND2x4_ASAP7_75t_L g14239 ( 
.A(n_13251),
.B(n_11524),
.Y(n_14239)
);

HB1xp67_ASAP7_75t_L g14240 ( 
.A(n_13306),
.Y(n_14240)
);

NAND2xp5_ASAP7_75t_L g14241 ( 
.A(n_13244),
.B(n_11525),
.Y(n_14241)
);

INVx1_ASAP7_75t_L g14242 ( 
.A(n_13043),
.Y(n_14242)
);

INVx1_ASAP7_75t_L g14243 ( 
.A(n_13044),
.Y(n_14243)
);

NAND2xp67_ASAP7_75t_L g14244 ( 
.A(n_13611),
.B(n_10745),
.Y(n_14244)
);

INVx2_ASAP7_75t_L g14245 ( 
.A(n_13132),
.Y(n_14245)
);

AOI22xp33_ASAP7_75t_SL g14246 ( 
.A1(n_13905),
.A2(n_8377),
.B1(n_8150),
.B2(n_7971),
.Y(n_14246)
);

AND2x2_ASAP7_75t_L g14247 ( 
.A(n_13390),
.B(n_11526),
.Y(n_14247)
);

INVx1_ASAP7_75t_L g14248 ( 
.A(n_13044),
.Y(n_14248)
);

INVx2_ASAP7_75t_L g14249 ( 
.A(n_13132),
.Y(n_14249)
);

BUFx2_ASAP7_75t_L g14250 ( 
.A(n_13208),
.Y(n_14250)
);

HB1xp67_ASAP7_75t_L g14251 ( 
.A(n_13320),
.Y(n_14251)
);

OR2x2_ASAP7_75t_L g14252 ( 
.A(n_13174),
.B(n_11532),
.Y(n_14252)
);

OR2x2_ASAP7_75t_L g14253 ( 
.A(n_13616),
.B(n_11533),
.Y(n_14253)
);

AND2x2_ASAP7_75t_L g14254 ( 
.A(n_13581),
.B(n_11535),
.Y(n_14254)
);

AND2x2_ASAP7_75t_L g14255 ( 
.A(n_13583),
.B(n_11537),
.Y(n_14255)
);

NAND2xp5_ASAP7_75t_L g14256 ( 
.A(n_13246),
.B(n_11538),
.Y(n_14256)
);

AND2x2_ASAP7_75t_L g14257 ( 
.A(n_13249),
.B(n_11539),
.Y(n_14257)
);

INVx4_ASAP7_75t_L g14258 ( 
.A(n_13524),
.Y(n_14258)
);

INVx1_ASAP7_75t_L g14259 ( 
.A(n_13048),
.Y(n_14259)
);

NOR2xp67_ASAP7_75t_L g14260 ( 
.A(n_13788),
.B(n_12952),
.Y(n_14260)
);

AND2x2_ASAP7_75t_L g14261 ( 
.A(n_13273),
.B(n_11543),
.Y(n_14261)
);

INVx1_ASAP7_75t_L g14262 ( 
.A(n_13048),
.Y(n_14262)
);

NAND2xp5_ASAP7_75t_L g14263 ( 
.A(n_13861),
.B(n_11545),
.Y(n_14263)
);

INVx1_ASAP7_75t_L g14264 ( 
.A(n_13050),
.Y(n_14264)
);

BUFx2_ASAP7_75t_L g14265 ( 
.A(n_13114),
.Y(n_14265)
);

INVx1_ASAP7_75t_L g14266 ( 
.A(n_13050),
.Y(n_14266)
);

INVxp67_ASAP7_75t_SL g14267 ( 
.A(n_13795),
.Y(n_14267)
);

HB1xp67_ASAP7_75t_L g14268 ( 
.A(n_13357),
.Y(n_14268)
);

INVx2_ASAP7_75t_L g14269 ( 
.A(n_13212),
.Y(n_14269)
);

AND2x2_ASAP7_75t_L g14270 ( 
.A(n_13196),
.B(n_11549),
.Y(n_14270)
);

NAND3xp33_ASAP7_75t_L g14271 ( 
.A(n_13870),
.B(n_12748),
.C(n_11889),
.Y(n_14271)
);

INVx1_ASAP7_75t_L g14272 ( 
.A(n_13051),
.Y(n_14272)
);

OAI22xp5_ASAP7_75t_L g14273 ( 
.A1(n_13318),
.A2(n_8142),
.B1(n_8295),
.B2(n_8095),
.Y(n_14273)
);

NAND2xp5_ASAP7_75t_L g14274 ( 
.A(n_13797),
.B(n_11551),
.Y(n_14274)
);

HB1xp67_ASAP7_75t_L g14275 ( 
.A(n_13693),
.Y(n_14275)
);

CKINVDCx5p33_ASAP7_75t_R g14276 ( 
.A(n_13477),
.Y(n_14276)
);

OR2x2_ASAP7_75t_L g14277 ( 
.A(n_13629),
.B(n_11553),
.Y(n_14277)
);

AND2x4_ASAP7_75t_L g14278 ( 
.A(n_13180),
.B(n_11557),
.Y(n_14278)
);

INVx4_ASAP7_75t_L g14279 ( 
.A(n_13524),
.Y(n_14279)
);

HB1xp67_ASAP7_75t_L g14280 ( 
.A(n_13693),
.Y(n_14280)
);

AND2x2_ASAP7_75t_L g14281 ( 
.A(n_13279),
.B(n_11559),
.Y(n_14281)
);

AND2x2_ASAP7_75t_L g14282 ( 
.A(n_13640),
.B(n_11570),
.Y(n_14282)
);

INVx1_ASAP7_75t_L g14283 ( 
.A(n_13051),
.Y(n_14283)
);

NAND2xp5_ASAP7_75t_L g14284 ( 
.A(n_13507),
.B(n_11576),
.Y(n_14284)
);

INVx1_ASAP7_75t_L g14285 ( 
.A(n_13053),
.Y(n_14285)
);

INVx1_ASAP7_75t_L g14286 ( 
.A(n_13053),
.Y(n_14286)
);

INVxp67_ASAP7_75t_L g14287 ( 
.A(n_13714),
.Y(n_14287)
);

INVx1_ASAP7_75t_L g14288 ( 
.A(n_13063),
.Y(n_14288)
);

INVxp67_ASAP7_75t_SL g14289 ( 
.A(n_13788),
.Y(n_14289)
);

INVx1_ASAP7_75t_L g14290 ( 
.A(n_13064),
.Y(n_14290)
);

AND2x2_ASAP7_75t_L g14291 ( 
.A(n_13640),
.B(n_13363),
.Y(n_14291)
);

AND2x2_ASAP7_75t_L g14292 ( 
.A(n_13370),
.B(n_11583),
.Y(n_14292)
);

INVx2_ASAP7_75t_L g14293 ( 
.A(n_13212),
.Y(n_14293)
);

INVx1_ASAP7_75t_L g14294 ( 
.A(n_13079),
.Y(n_14294)
);

INVx1_ASAP7_75t_L g14295 ( 
.A(n_13080),
.Y(n_14295)
);

OR2x2_ASAP7_75t_L g14296 ( 
.A(n_13069),
.B(n_11587),
.Y(n_14296)
);

INVx1_ASAP7_75t_L g14297 ( 
.A(n_13082),
.Y(n_14297)
);

AND2x2_ASAP7_75t_L g14298 ( 
.A(n_13381),
.B(n_11589),
.Y(n_14298)
);

AND2x2_ASAP7_75t_L g14299 ( 
.A(n_13627),
.B(n_11594),
.Y(n_14299)
);

AND2x2_ASAP7_75t_L g14300 ( 
.A(n_13686),
.B(n_11595),
.Y(n_14300)
);

INVx2_ASAP7_75t_L g14301 ( 
.A(n_13253),
.Y(n_14301)
);

INVx2_ASAP7_75t_L g14302 ( 
.A(n_13253),
.Y(n_14302)
);

OR2x2_ASAP7_75t_L g14303 ( 
.A(n_13775),
.B(n_11602),
.Y(n_14303)
);

NAND2xp5_ASAP7_75t_L g14304 ( 
.A(n_13508),
.B(n_11603),
.Y(n_14304)
);

AND2x2_ASAP7_75t_L g14305 ( 
.A(n_13344),
.B(n_11606),
.Y(n_14305)
);

AND2x4_ASAP7_75t_L g14306 ( 
.A(n_13187),
.B(n_11610),
.Y(n_14306)
);

NAND2xp5_ASAP7_75t_L g14307 ( 
.A(n_13836),
.B(n_11612),
.Y(n_14307)
);

BUFx6f_ASAP7_75t_SL g14308 ( 
.A(n_13562),
.Y(n_14308)
);

AND2x2_ASAP7_75t_L g14309 ( 
.A(n_13430),
.B(n_11614),
.Y(n_14309)
);

INVx1_ASAP7_75t_L g14310 ( 
.A(n_13086),
.Y(n_14310)
);

INVx1_ASAP7_75t_L g14311 ( 
.A(n_13087),
.Y(n_14311)
);

INVx2_ASAP7_75t_L g14312 ( 
.A(n_13365),
.Y(n_14312)
);

INVx1_ASAP7_75t_L g14313 ( 
.A(n_13088),
.Y(n_14313)
);

OR2x2_ASAP7_75t_L g14314 ( 
.A(n_13181),
.B(n_11617),
.Y(n_14314)
);

AND2x2_ASAP7_75t_L g14315 ( 
.A(n_13431),
.B(n_11622),
.Y(n_14315)
);

AOI22xp33_ASAP7_75t_L g14316 ( 
.A1(n_13787),
.A2(n_8574),
.B1(n_8150),
.B2(n_10415),
.Y(n_14316)
);

AND2x2_ASAP7_75t_L g14317 ( 
.A(n_13615),
.B(n_11624),
.Y(n_14317)
);

INVx2_ASAP7_75t_L g14318 ( 
.A(n_13365),
.Y(n_14318)
);

BUFx2_ASAP7_75t_L g14319 ( 
.A(n_13704),
.Y(n_14319)
);

AND2x2_ASAP7_75t_L g14320 ( 
.A(n_13705),
.B(n_11625),
.Y(n_14320)
);

BUFx3_ASAP7_75t_L g14321 ( 
.A(n_13377),
.Y(n_14321)
);

INVx1_ASAP7_75t_L g14322 ( 
.A(n_13089),
.Y(n_14322)
);

INVx1_ASAP7_75t_L g14323 ( 
.A(n_13090),
.Y(n_14323)
);

AOI22xp5_ASAP7_75t_L g14324 ( 
.A1(n_13800),
.A2(n_8150),
.B1(n_8641),
.B2(n_8626),
.Y(n_14324)
);

INVx1_ASAP7_75t_SL g14325 ( 
.A(n_13733),
.Y(n_14325)
);

AND2x2_ASAP7_75t_L g14326 ( 
.A(n_13404),
.B(n_11627),
.Y(n_14326)
);

INVx1_ASAP7_75t_L g14327 ( 
.A(n_13094),
.Y(n_14327)
);

INVxp67_ASAP7_75t_SL g14328 ( 
.A(n_13101),
.Y(n_14328)
);

INVx2_ASAP7_75t_L g14329 ( 
.A(n_13372),
.Y(n_14329)
);

AND2x2_ASAP7_75t_L g14330 ( 
.A(n_13378),
.B(n_11634),
.Y(n_14330)
);

NAND2xp5_ASAP7_75t_L g14331 ( 
.A(n_13780),
.B(n_11639),
.Y(n_14331)
);

NOR2xp33_ASAP7_75t_L g14332 ( 
.A(n_13296),
.B(n_9229),
.Y(n_14332)
);

INVx2_ASAP7_75t_L g14333 ( 
.A(n_13372),
.Y(n_14333)
);

NAND2xp5_ASAP7_75t_L g14334 ( 
.A(n_13744),
.B(n_11640),
.Y(n_14334)
);

NAND2xp5_ASAP7_75t_L g14335 ( 
.A(n_13409),
.B(n_11641),
.Y(n_14335)
);

AND2x2_ASAP7_75t_L g14336 ( 
.A(n_13573),
.B(n_11644),
.Y(n_14336)
);

OR2x2_ASAP7_75t_L g14337 ( 
.A(n_12975),
.B(n_11649),
.Y(n_14337)
);

AND2x2_ASAP7_75t_L g14338 ( 
.A(n_13653),
.B(n_11651),
.Y(n_14338)
);

INVx1_ASAP7_75t_L g14339 ( 
.A(n_13105),
.Y(n_14339)
);

AND2x4_ASAP7_75t_L g14340 ( 
.A(n_13195),
.B(n_11653),
.Y(n_14340)
);

INVx1_ASAP7_75t_SL g14341 ( 
.A(n_13704),
.Y(n_14341)
);

AND2x2_ASAP7_75t_L g14342 ( 
.A(n_13223),
.B(n_13226),
.Y(n_14342)
);

INVx2_ASAP7_75t_L g14343 ( 
.A(n_13496),
.Y(n_14343)
);

INVx1_ASAP7_75t_L g14344 ( 
.A(n_13110),
.Y(n_14344)
);

AND2x2_ASAP7_75t_L g14345 ( 
.A(n_13227),
.B(n_11655),
.Y(n_14345)
);

INVx4_ASAP7_75t_L g14346 ( 
.A(n_13524),
.Y(n_14346)
);

AND2x4_ASAP7_75t_L g14347 ( 
.A(n_13199),
.B(n_11659),
.Y(n_14347)
);

INVx1_ASAP7_75t_L g14348 ( 
.A(n_13112),
.Y(n_14348)
);

INVx1_ASAP7_75t_L g14349 ( 
.A(n_13115),
.Y(n_14349)
);

INVx1_ASAP7_75t_L g14350 ( 
.A(n_13117),
.Y(n_14350)
);

BUFx6f_ASAP7_75t_L g14351 ( 
.A(n_13592),
.Y(n_14351)
);

INVx1_ASAP7_75t_L g14352 ( 
.A(n_13123),
.Y(n_14352)
);

INVx2_ASAP7_75t_L g14353 ( 
.A(n_13496),
.Y(n_14353)
);

HB1xp67_ASAP7_75t_L g14354 ( 
.A(n_13693),
.Y(n_14354)
);

NAND2xp5_ASAP7_75t_L g14355 ( 
.A(n_13881),
.B(n_11665),
.Y(n_14355)
);

AND2x2_ASAP7_75t_L g14356 ( 
.A(n_13326),
.B(n_11671),
.Y(n_14356)
);

INVx2_ASAP7_75t_L g14357 ( 
.A(n_13415),
.Y(n_14357)
);

INVx1_ASAP7_75t_L g14358 ( 
.A(n_13124),
.Y(n_14358)
);

INVx2_ASAP7_75t_L g14359 ( 
.A(n_13415),
.Y(n_14359)
);

AOI22xp5_ASAP7_75t_L g14360 ( 
.A1(n_13904),
.A2(n_8150),
.B1(n_8641),
.B2(n_8626),
.Y(n_14360)
);

INVx1_ASAP7_75t_L g14361 ( 
.A(n_13125),
.Y(n_14361)
);

OR2x2_ASAP7_75t_L g14362 ( 
.A(n_12985),
.B(n_11674),
.Y(n_14362)
);

NAND2xp5_ASAP7_75t_L g14363 ( 
.A(n_13672),
.B(n_11675),
.Y(n_14363)
);

OR2x2_ASAP7_75t_L g14364 ( 
.A(n_13391),
.B(n_11676),
.Y(n_14364)
);

INVx1_ASAP7_75t_L g14365 ( 
.A(n_13127),
.Y(n_14365)
);

NAND2xp5_ASAP7_75t_L g14366 ( 
.A(n_13677),
.B(n_11697),
.Y(n_14366)
);

NAND2xp5_ASAP7_75t_L g14367 ( 
.A(n_13680),
.B(n_11699),
.Y(n_14367)
);

INVx2_ASAP7_75t_L g14368 ( 
.A(n_13436),
.Y(n_14368)
);

INVx1_ASAP7_75t_L g14369 ( 
.A(n_13130),
.Y(n_14369)
);

AOI22xp33_ASAP7_75t_L g14370 ( 
.A1(n_13671),
.A2(n_10415),
.B1(n_8626),
.B2(n_8655),
.Y(n_14370)
);

BUFx2_ASAP7_75t_L g14371 ( 
.A(n_13368),
.Y(n_14371)
);

AOI22xp33_ASAP7_75t_L g14372 ( 
.A1(n_13621),
.A2(n_10415),
.B1(n_8626),
.B2(n_8655),
.Y(n_14372)
);

AND2x2_ASAP7_75t_L g14373 ( 
.A(n_13865),
.B(n_11700),
.Y(n_14373)
);

AND2x4_ASAP7_75t_L g14374 ( 
.A(n_13204),
.B(n_13205),
.Y(n_14374)
);

AND2x2_ASAP7_75t_L g14375 ( 
.A(n_13575),
.B(n_11701),
.Y(n_14375)
);

INVx1_ASAP7_75t_L g14376 ( 
.A(n_13136),
.Y(n_14376)
);

AND2x2_ASAP7_75t_L g14377 ( 
.A(n_13582),
.B(n_11709),
.Y(n_14377)
);

AND2x2_ASAP7_75t_L g14378 ( 
.A(n_13594),
.B(n_11714),
.Y(n_14378)
);

INVx2_ASAP7_75t_L g14379 ( 
.A(n_13436),
.Y(n_14379)
);

NAND2xp5_ASAP7_75t_L g14380 ( 
.A(n_13682),
.B(n_11715),
.Y(n_14380)
);

AND2x2_ASAP7_75t_L g14381 ( 
.A(n_13758),
.B(n_13593),
.Y(n_14381)
);

INVx2_ASAP7_75t_L g14382 ( 
.A(n_13592),
.Y(n_14382)
);

INVx1_ASAP7_75t_L g14383 ( 
.A(n_13145),
.Y(n_14383)
);

INVx1_ASAP7_75t_L g14384 ( 
.A(n_13148),
.Y(n_14384)
);

INVx2_ASAP7_75t_L g14385 ( 
.A(n_13592),
.Y(n_14385)
);

AND2x2_ASAP7_75t_L g14386 ( 
.A(n_13539),
.B(n_13604),
.Y(n_14386)
);

AND2x2_ASAP7_75t_L g14387 ( 
.A(n_13601),
.B(n_11718),
.Y(n_14387)
);

NAND2xp5_ASAP7_75t_L g14388 ( 
.A(n_13683),
.B(n_11723),
.Y(n_14388)
);

INVx1_ASAP7_75t_L g14389 ( 
.A(n_13150),
.Y(n_14389)
);

INVx2_ASAP7_75t_L g14390 ( 
.A(n_13275),
.Y(n_14390)
);

NAND2xp5_ASAP7_75t_L g14391 ( 
.A(n_13726),
.B(n_11733),
.Y(n_14391)
);

INVx1_ASAP7_75t_L g14392 ( 
.A(n_13151),
.Y(n_14392)
);

AND2x4_ASAP7_75t_L g14393 ( 
.A(n_13214),
.B(n_11736),
.Y(n_14393)
);

INVx1_ASAP7_75t_SL g14394 ( 
.A(n_13730),
.Y(n_14394)
);

INVx2_ASAP7_75t_L g14395 ( 
.A(n_13275),
.Y(n_14395)
);

AND2x2_ASAP7_75t_L g14396 ( 
.A(n_13311),
.B(n_11741),
.Y(n_14396)
);

INVx2_ASAP7_75t_L g14397 ( 
.A(n_13293),
.Y(n_14397)
);

INVxp67_ASAP7_75t_SL g14398 ( 
.A(n_13121),
.Y(n_14398)
);

INVx1_ASAP7_75t_L g14399 ( 
.A(n_13155),
.Y(n_14399)
);

AOI22xp33_ASAP7_75t_L g14400 ( 
.A1(n_13655),
.A2(n_8626),
.B1(n_8655),
.B2(n_8641),
.Y(n_14400)
);

AND2x4_ASAP7_75t_SL g14401 ( 
.A(n_13562),
.B(n_8210),
.Y(n_14401)
);

INVx3_ASAP7_75t_L g14402 ( 
.A(n_13293),
.Y(n_14402)
);

AOI22xp33_ASAP7_75t_L g14403 ( 
.A1(n_13904),
.A2(n_8641),
.B1(n_8657),
.B2(n_8655),
.Y(n_14403)
);

INVx1_ASAP7_75t_L g14404 ( 
.A(n_13158),
.Y(n_14404)
);

AND2x2_ASAP7_75t_L g14405 ( 
.A(n_13002),
.B(n_11742),
.Y(n_14405)
);

INVx1_ASAP7_75t_L g14406 ( 
.A(n_13278),
.Y(n_14406)
);

INVx1_ASAP7_75t_L g14407 ( 
.A(n_13287),
.Y(n_14407)
);

AND2x2_ASAP7_75t_L g14408 ( 
.A(n_13602),
.B(n_11744),
.Y(n_14408)
);

AND2x4_ASAP7_75t_L g14409 ( 
.A(n_13216),
.B(n_11747),
.Y(n_14409)
);

INVx2_ASAP7_75t_L g14410 ( 
.A(n_13324),
.Y(n_14410)
);

AND2x2_ASAP7_75t_L g14411 ( 
.A(n_13603),
.B(n_11752),
.Y(n_14411)
);

INVxp67_ASAP7_75t_SL g14412 ( 
.A(n_13654),
.Y(n_14412)
);

OAI22xp5_ASAP7_75t_L g14413 ( 
.A1(n_13749),
.A2(n_8142),
.B1(n_8295),
.B2(n_8095),
.Y(n_14413)
);

INVx2_ASAP7_75t_L g14414 ( 
.A(n_13324),
.Y(n_14414)
);

INVx1_ASAP7_75t_L g14415 ( 
.A(n_13414),
.Y(n_14415)
);

INVx2_ASAP7_75t_L g14416 ( 
.A(n_13222),
.Y(n_14416)
);

BUFx3_ASAP7_75t_L g14417 ( 
.A(n_13521),
.Y(n_14417)
);

NAND2xp5_ASAP7_75t_L g14418 ( 
.A(n_13911),
.B(n_13806),
.Y(n_14418)
);

BUFx2_ASAP7_75t_L g14419 ( 
.A(n_13368),
.Y(n_14419)
);

OR2x2_ASAP7_75t_L g14420 ( 
.A(n_12963),
.B(n_11754),
.Y(n_14420)
);

INVx2_ASAP7_75t_L g14421 ( 
.A(n_13224),
.Y(n_14421)
);

INVx3_ASAP7_75t_L g14422 ( 
.A(n_13478),
.Y(n_14422)
);

OR2x2_ASAP7_75t_L g14423 ( 
.A(n_13793),
.B(n_13821),
.Y(n_14423)
);

AND2x2_ASAP7_75t_L g14424 ( 
.A(n_13612),
.B(n_11756),
.Y(n_14424)
);

AOI211x1_ASAP7_75t_SL g14425 ( 
.A1(n_13919),
.A2(n_10747),
.B(n_10751),
.C(n_10745),
.Y(n_14425)
);

AND2x2_ASAP7_75t_L g14426 ( 
.A(n_13310),
.B(n_13019),
.Y(n_14426)
);

INVx2_ASAP7_75t_L g14427 ( 
.A(n_13229),
.Y(n_14427)
);

AND2x2_ASAP7_75t_L g14428 ( 
.A(n_13147),
.B(n_13159),
.Y(n_14428)
);

NOR2x1_ASAP7_75t_R g14429 ( 
.A(n_13548),
.B(n_7757),
.Y(n_14429)
);

CKINVDCx5p33_ASAP7_75t_R g14430 ( 
.A(n_13345),
.Y(n_14430)
);

INVx2_ASAP7_75t_L g14431 ( 
.A(n_13236),
.Y(n_14431)
);

AND2x4_ASAP7_75t_L g14432 ( 
.A(n_13520),
.B(n_13173),
.Y(n_14432)
);

OR2x2_ASAP7_75t_L g14433 ( 
.A(n_13906),
.B(n_11757),
.Y(n_14433)
);

INVx2_ASAP7_75t_L g14434 ( 
.A(n_13513),
.Y(n_14434)
);

NOR2xp33_ASAP7_75t_SL g14435 ( 
.A(n_13327),
.B(n_7582),
.Y(n_14435)
);

HB1xp67_ASAP7_75t_L g14436 ( 
.A(n_13470),
.Y(n_14436)
);

INVx1_ASAP7_75t_L g14437 ( 
.A(n_13472),
.Y(n_14437)
);

AND2x4_ASAP7_75t_L g14438 ( 
.A(n_13520),
.B(n_11759),
.Y(n_14438)
);

AND2x2_ASAP7_75t_L g14439 ( 
.A(n_13169),
.B(n_11762),
.Y(n_14439)
);

OR2x2_ASAP7_75t_L g14440 ( 
.A(n_13906),
.B(n_11766),
.Y(n_14440)
);

AND2x2_ASAP7_75t_L g14441 ( 
.A(n_13303),
.B(n_13560),
.Y(n_14441)
);

INVx1_ASAP7_75t_L g14442 ( 
.A(n_13304),
.Y(n_14442)
);

INVx1_ASAP7_75t_L g14443 ( 
.A(n_13308),
.Y(n_14443)
);

AND2x2_ASAP7_75t_L g14444 ( 
.A(n_13569),
.B(n_13254),
.Y(n_14444)
);

INVx2_ASAP7_75t_L g14445 ( 
.A(n_13513),
.Y(n_14445)
);

OR2x2_ASAP7_75t_L g14446 ( 
.A(n_13768),
.B(n_13871),
.Y(n_14446)
);

AND2x2_ASAP7_75t_L g14447 ( 
.A(n_13047),
.B(n_11767),
.Y(n_14447)
);

INVx2_ASAP7_75t_L g14448 ( 
.A(n_13529),
.Y(n_14448)
);

INVx1_ASAP7_75t_L g14449 ( 
.A(n_13309),
.Y(n_14449)
);

AND2x2_ASAP7_75t_L g14450 ( 
.A(n_13054),
.B(n_11776),
.Y(n_14450)
);

INVx2_ASAP7_75t_L g14451 ( 
.A(n_13529),
.Y(n_14451)
);

INVx2_ASAP7_75t_L g14452 ( 
.A(n_13545),
.Y(n_14452)
);

INVx1_ASAP7_75t_L g14453 ( 
.A(n_13312),
.Y(n_14453)
);

NAND2xp5_ASAP7_75t_L g14454 ( 
.A(n_13179),
.B(n_11777),
.Y(n_14454)
);

AND2x4_ASAP7_75t_L g14455 ( 
.A(n_13177),
.B(n_11778),
.Y(n_14455)
);

INVxp67_ASAP7_75t_SL g14456 ( 
.A(n_13762),
.Y(n_14456)
);

BUFx3_ASAP7_75t_L g14457 ( 
.A(n_13407),
.Y(n_14457)
);

INVx1_ASAP7_75t_L g14458 ( 
.A(n_13315),
.Y(n_14458)
);

OR2x2_ASAP7_75t_L g14459 ( 
.A(n_13250),
.B(n_11780),
.Y(n_14459)
);

INVx1_ASAP7_75t_L g14460 ( 
.A(n_13316),
.Y(n_14460)
);

AOI22xp33_ASAP7_75t_SL g14461 ( 
.A1(n_13624),
.A2(n_8377),
.B1(n_8432),
.B2(n_8392),
.Y(n_14461)
);

AND2x2_ASAP7_75t_L g14462 ( 
.A(n_13791),
.B(n_11781),
.Y(n_14462)
);

INVxp67_ASAP7_75t_L g14463 ( 
.A(n_13829),
.Y(n_14463)
);

INVx1_ASAP7_75t_L g14464 ( 
.A(n_13338),
.Y(n_14464)
);

INVx1_ASAP7_75t_L g14465 ( 
.A(n_13339),
.Y(n_14465)
);

HB1xp67_ASAP7_75t_L g14466 ( 
.A(n_13480),
.Y(n_14466)
);

OR2x6_ASAP7_75t_L g14467 ( 
.A(n_13432),
.B(n_7790),
.Y(n_14467)
);

BUFx2_ASAP7_75t_L g14468 ( 
.A(n_13730),
.Y(n_14468)
);

INVx2_ASAP7_75t_L g14469 ( 
.A(n_13545),
.Y(n_14469)
);

AND2x4_ASAP7_75t_L g14470 ( 
.A(n_13515),
.B(n_11785),
.Y(n_14470)
);

INVx1_ASAP7_75t_L g14471 ( 
.A(n_13343),
.Y(n_14471)
);

AND2x2_ASAP7_75t_L g14472 ( 
.A(n_13240),
.B(n_11788),
.Y(n_14472)
);

HB1xp67_ASAP7_75t_L g14473 ( 
.A(n_13500),
.Y(n_14473)
);

INVx2_ASAP7_75t_L g14474 ( 
.A(n_13546),
.Y(n_14474)
);

AND2x4_ASAP7_75t_L g14475 ( 
.A(n_13519),
.B(n_11789),
.Y(n_14475)
);

INVx1_ASAP7_75t_L g14476 ( 
.A(n_13347),
.Y(n_14476)
);

INVx1_ASAP7_75t_L g14477 ( 
.A(n_13348),
.Y(n_14477)
);

INVx2_ASAP7_75t_L g14478 ( 
.A(n_13546),
.Y(n_14478)
);

INVxp67_ASAP7_75t_L g14479 ( 
.A(n_13835),
.Y(n_14479)
);

AND2x4_ASAP7_75t_L g14480 ( 
.A(n_13478),
.B(n_11792),
.Y(n_14480)
);

AND2x2_ASAP7_75t_L g14481 ( 
.A(n_13243),
.B(n_11796),
.Y(n_14481)
);

INVx1_ASAP7_75t_L g14482 ( 
.A(n_13351),
.Y(n_14482)
);

INVx4_ASAP7_75t_L g14483 ( 
.A(n_13451),
.Y(n_14483)
);

AND2x2_ASAP7_75t_L g14484 ( 
.A(n_13057),
.B(n_11798),
.Y(n_14484)
);

NAND2xp5_ASAP7_75t_L g14485 ( 
.A(n_13759),
.B(n_11803),
.Y(n_14485)
);

INVx1_ASAP7_75t_L g14486 ( 
.A(n_13354),
.Y(n_14486)
);

BUFx6f_ASAP7_75t_L g14487 ( 
.A(n_13458),
.Y(n_14487)
);

OR2x2_ASAP7_75t_L g14488 ( 
.A(n_13837),
.B(n_11804),
.Y(n_14488)
);

HB1xp67_ASAP7_75t_L g14489 ( 
.A(n_13553),
.Y(n_14489)
);

INVx1_ASAP7_75t_L g14490 ( 
.A(n_13396),
.Y(n_14490)
);

AND2x4_ASAP7_75t_L g14491 ( 
.A(n_13498),
.B(n_11807),
.Y(n_14491)
);

INVxp67_ASAP7_75t_SL g14492 ( 
.A(n_13762),
.Y(n_14492)
);

INVx1_ASAP7_75t_L g14493 ( 
.A(n_13334),
.Y(n_14493)
);

AND2x2_ASAP7_75t_L g14494 ( 
.A(n_13067),
.B(n_11811),
.Y(n_14494)
);

INVx1_ASAP7_75t_L g14495 ( 
.A(n_13346),
.Y(n_14495)
);

OAI21xp5_ASAP7_75t_SL g14496 ( 
.A1(n_13763),
.A2(n_8862),
.B(n_8183),
.Y(n_14496)
);

HB1xp67_ASAP7_75t_L g14497 ( 
.A(n_13696),
.Y(n_14497)
);

OR2x2_ASAP7_75t_L g14498 ( 
.A(n_13191),
.B(n_11812),
.Y(n_14498)
);

BUFx12f_ASAP7_75t_L g14499 ( 
.A(n_13678),
.Y(n_14499)
);

AOI22xp33_ASAP7_75t_L g14500 ( 
.A1(n_13896),
.A2(n_8641),
.B1(n_8657),
.B2(n_8655),
.Y(n_14500)
);

AND2x2_ASAP7_75t_L g14501 ( 
.A(n_12983),
.B(n_11814),
.Y(n_14501)
);

AND2x4_ASAP7_75t_L g14502 ( 
.A(n_13554),
.B(n_11815),
.Y(n_14502)
);

INVx1_ASAP7_75t_L g14503 ( 
.A(n_12988),
.Y(n_14503)
);

INVxp67_ASAP7_75t_L g14504 ( 
.A(n_13907),
.Y(n_14504)
);

NAND2xp5_ASAP7_75t_L g14505 ( 
.A(n_13765),
.B(n_11817),
.Y(n_14505)
);

INVx2_ASAP7_75t_L g14506 ( 
.A(n_13554),
.Y(n_14506)
);

INVx2_ASAP7_75t_L g14507 ( 
.A(n_12979),
.Y(n_14507)
);

NAND2xp5_ASAP7_75t_L g14508 ( 
.A(n_13367),
.B(n_11818),
.Y(n_14508)
);

INVx1_ASAP7_75t_L g14509 ( 
.A(n_12994),
.Y(n_14509)
);

AND2x2_ASAP7_75t_L g14510 ( 
.A(n_13538),
.B(n_11821),
.Y(n_14510)
);

BUFx2_ASAP7_75t_L g14511 ( 
.A(n_13368),
.Y(n_14511)
);

INVxp67_ASAP7_75t_L g14512 ( 
.A(n_13859),
.Y(n_14512)
);

HB1xp67_ASAP7_75t_L g14513 ( 
.A(n_13698),
.Y(n_14513)
);

INVxp67_ASAP7_75t_L g14514 ( 
.A(n_13716),
.Y(n_14514)
);

INVxp67_ASAP7_75t_SL g14515 ( 
.A(n_13819),
.Y(n_14515)
);

BUFx2_ASAP7_75t_L g14516 ( 
.A(n_13274),
.Y(n_14516)
);

NAND2xp5_ASAP7_75t_L g14517 ( 
.A(n_13380),
.B(n_11823),
.Y(n_14517)
);

INVx1_ASAP7_75t_L g14518 ( 
.A(n_13164),
.Y(n_14518)
);

INVx2_ASAP7_75t_SL g14519 ( 
.A(n_13596),
.Y(n_14519)
);

AND2x2_ASAP7_75t_L g14520 ( 
.A(n_13025),
.B(n_11824),
.Y(n_14520)
);

OR2x2_ASAP7_75t_L g14521 ( 
.A(n_13528),
.B(n_11829),
.Y(n_14521)
);

HB1xp67_ASAP7_75t_L g14522 ( 
.A(n_13062),
.Y(n_14522)
);

OR2x2_ASAP7_75t_L g14523 ( 
.A(n_13157),
.B(n_11830),
.Y(n_14523)
);

INVx2_ASAP7_75t_L g14524 ( 
.A(n_12980),
.Y(n_14524)
);

HB1xp67_ASAP7_75t_L g14525 ( 
.A(n_13062),
.Y(n_14525)
);

INVx1_ASAP7_75t_L g14526 ( 
.A(n_13168),
.Y(n_14526)
);

NAND2x1p5_ASAP7_75t_SL g14527 ( 
.A(n_13717),
.B(n_7916),
.Y(n_14527)
);

INVx1_ASAP7_75t_L g14528 ( 
.A(n_13176),
.Y(n_14528)
);

INVx1_ASAP7_75t_L g14529 ( 
.A(n_13184),
.Y(n_14529)
);

INVx1_ASAP7_75t_L g14530 ( 
.A(n_13190),
.Y(n_14530)
);

INVx2_ASAP7_75t_L g14531 ( 
.A(n_13036),
.Y(n_14531)
);

NOR2x1_ASAP7_75t_SL g14532 ( 
.A(n_13410),
.B(n_10747),
.Y(n_14532)
);

AND2x4_ASAP7_75t_L g14533 ( 
.A(n_13561),
.B(n_11832),
.Y(n_14533)
);

INVx1_ASAP7_75t_L g14534 ( 
.A(n_13193),
.Y(n_14534)
);

INVx2_ASAP7_75t_L g14535 ( 
.A(n_13040),
.Y(n_14535)
);

AND2x2_ASAP7_75t_L g14536 ( 
.A(n_13028),
.B(n_11836),
.Y(n_14536)
);

NAND2xp5_ASAP7_75t_L g14537 ( 
.A(n_13772),
.B(n_13773),
.Y(n_14537)
);

OR2x2_ASAP7_75t_L g14538 ( 
.A(n_13623),
.B(n_11839),
.Y(n_14538)
);

INVx1_ASAP7_75t_L g14539 ( 
.A(n_13194),
.Y(n_14539)
);

INVx2_ASAP7_75t_L g14540 ( 
.A(n_13029),
.Y(n_14540)
);

OR2x2_ASAP7_75t_L g14541 ( 
.A(n_13068),
.B(n_11840),
.Y(n_14541)
);

AND2x2_ASAP7_75t_L g14542 ( 
.A(n_13035),
.B(n_11852),
.Y(n_14542)
);

INVx1_ASAP7_75t_L g14543 ( 
.A(n_13213),
.Y(n_14543)
);

HB1xp67_ASAP7_75t_L g14544 ( 
.A(n_13062),
.Y(n_14544)
);

AND2x2_ASAP7_75t_L g14545 ( 
.A(n_13514),
.B(n_13178),
.Y(n_14545)
);

AND2x2_ASAP7_75t_L g14546 ( 
.A(n_13771),
.B(n_11855),
.Y(n_14546)
);

INVx1_ASAP7_75t_L g14547 ( 
.A(n_13217),
.Y(n_14547)
);

BUFx6f_ASAP7_75t_L g14548 ( 
.A(n_13596),
.Y(n_14548)
);

NAND2xp5_ASAP7_75t_L g14549 ( 
.A(n_13870),
.B(n_13376),
.Y(n_14549)
);

HB1xp67_ASAP7_75t_L g14550 ( 
.A(n_13429),
.Y(n_14550)
);

INVx2_ASAP7_75t_L g14551 ( 
.A(n_13020),
.Y(n_14551)
);

AND2x2_ASAP7_75t_L g14552 ( 
.A(n_13641),
.B(n_11859),
.Y(n_14552)
);

AND2x4_ASAP7_75t_L g14553 ( 
.A(n_13563),
.B(n_11863),
.Y(n_14553)
);

OR2x2_ASAP7_75t_SL g14554 ( 
.A(n_13721),
.B(n_9369),
.Y(n_14554)
);

OR2x2_ASAP7_75t_L g14555 ( 
.A(n_13225),
.B(n_11867),
.Y(n_14555)
);

INVx2_ASAP7_75t_L g14556 ( 
.A(n_13004),
.Y(n_14556)
);

HB1xp67_ASAP7_75t_L g14557 ( 
.A(n_13635),
.Y(n_14557)
);

AND2x2_ASAP7_75t_L g14558 ( 
.A(n_13144),
.B(n_13522),
.Y(n_14558)
);

INVx1_ASAP7_75t_L g14559 ( 
.A(n_13218),
.Y(n_14559)
);

INVx2_ASAP7_75t_L g14560 ( 
.A(n_13018),
.Y(n_14560)
);

NOR2xp33_ASAP7_75t_L g14561 ( 
.A(n_13322),
.B(n_13383),
.Y(n_14561)
);

INVxp33_ASAP7_75t_L g14562 ( 
.A(n_13503),
.Y(n_14562)
);

INVx1_ASAP7_75t_L g14563 ( 
.A(n_13219),
.Y(n_14563)
);

INVx1_ASAP7_75t_L g14564 ( 
.A(n_13231),
.Y(n_14564)
);

BUFx2_ASAP7_75t_L g14565 ( 
.A(n_13826),
.Y(n_14565)
);

NAND2xp5_ASAP7_75t_L g14566 ( 
.A(n_13872),
.B(n_11870),
.Y(n_14566)
);

AND2x2_ASAP7_75t_L g14567 ( 
.A(n_13070),
.B(n_11873),
.Y(n_14567)
);

OR2x2_ASAP7_75t_L g14568 ( 
.A(n_13636),
.B(n_11879),
.Y(n_14568)
);

AND2x4_ASAP7_75t_SL g14569 ( 
.A(n_13650),
.B(n_8210),
.Y(n_14569)
);

NAND2xp5_ASAP7_75t_L g14570 ( 
.A(n_13872),
.B(n_11886),
.Y(n_14570)
);

NAND2xp5_ASAP7_75t_L g14571 ( 
.A(n_13646),
.B(n_11891),
.Y(n_14571)
);

NAND2xp5_ASAP7_75t_L g14572 ( 
.A(n_13647),
.B(n_11897),
.Y(n_14572)
);

INVx1_ASAP7_75t_L g14573 ( 
.A(n_13232),
.Y(n_14573)
);

INVx3_ASAP7_75t_L g14574 ( 
.A(n_13684),
.Y(n_14574)
);

INVx1_ASAP7_75t_L g14575 ( 
.A(n_13242),
.Y(n_14575)
);

NAND2xp5_ASAP7_75t_L g14576 ( 
.A(n_13651),
.B(n_11898),
.Y(n_14576)
);

INVx2_ASAP7_75t_L g14577 ( 
.A(n_13075),
.Y(n_14577)
);

INVxp67_ASAP7_75t_SL g14578 ( 
.A(n_13889),
.Y(n_14578)
);

AND2x2_ASAP7_75t_L g14579 ( 
.A(n_13077),
.B(n_11905),
.Y(n_14579)
);

OR2x2_ASAP7_75t_L g14580 ( 
.A(n_13565),
.B(n_11909),
.Y(n_14580)
);

OR2x2_ASAP7_75t_L g14581 ( 
.A(n_13010),
.B(n_11911),
.Y(n_14581)
);

AND2x2_ASAP7_75t_L g14582 ( 
.A(n_13083),
.B(n_11913),
.Y(n_14582)
);

AND2x2_ASAP7_75t_L g14583 ( 
.A(n_13084),
.B(n_11915),
.Y(n_14583)
);

INVx1_ASAP7_75t_SL g14584 ( 
.A(n_13549),
.Y(n_14584)
);

NAND2xp5_ASAP7_75t_L g14585 ( 
.A(n_13879),
.B(n_11917),
.Y(n_14585)
);

INVx2_ASAP7_75t_L g14586 ( 
.A(n_13901),
.Y(n_14586)
);

HB1xp67_ASAP7_75t_L g14587 ( 
.A(n_13644),
.Y(n_14587)
);

INVxp67_ASAP7_75t_L g14588 ( 
.A(n_13659),
.Y(n_14588)
);

INVx2_ASAP7_75t_L g14589 ( 
.A(n_13901),
.Y(n_14589)
);

INVx2_ASAP7_75t_L g14590 ( 
.A(n_13663),
.Y(n_14590)
);

INVx1_ASAP7_75t_L g14591 ( 
.A(n_13081),
.Y(n_14591)
);

INVx2_ASAP7_75t_L g14592 ( 
.A(n_13663),
.Y(n_14592)
);

INVx1_ASAP7_75t_L g14593 ( 
.A(n_13419),
.Y(n_14593)
);

NAND2xp5_ASAP7_75t_L g14594 ( 
.A(n_13879),
.B(n_11928),
.Y(n_14594)
);

INVx1_ASAP7_75t_L g14595 ( 
.A(n_13622),
.Y(n_14595)
);

AND2x2_ASAP7_75t_L g14596 ( 
.A(n_13637),
.B(n_8590),
.Y(n_14596)
);

NAND2xp5_ASAP7_75t_SL g14597 ( 
.A(n_13188),
.B(n_8095),
.Y(n_14597)
);

INVx1_ASAP7_75t_L g14598 ( 
.A(n_13625),
.Y(n_14598)
);

AND2x4_ASAP7_75t_SL g14599 ( 
.A(n_13754),
.B(n_8210),
.Y(n_14599)
);

NAND2xp5_ASAP7_75t_L g14600 ( 
.A(n_13880),
.B(n_11353),
.Y(n_14600)
);

INVx3_ASAP7_75t_L g14601 ( 
.A(n_13684),
.Y(n_14601)
);

INVx2_ASAP7_75t_L g14602 ( 
.A(n_13142),
.Y(n_14602)
);

AND2x2_ASAP7_75t_L g14603 ( 
.A(n_13804),
.B(n_8590),
.Y(n_14603)
);

INVx2_ASAP7_75t_L g14604 ( 
.A(n_13143),
.Y(n_14604)
);

INVxp67_ASAP7_75t_L g14605 ( 
.A(n_13410),
.Y(n_14605)
);

INVx1_ASAP7_75t_L g14606 ( 
.A(n_13638),
.Y(n_14606)
);

INVx1_ASAP7_75t_L g14607 ( 
.A(n_13639),
.Y(n_14607)
);

AND2x2_ASAP7_75t_L g14608 ( 
.A(n_13433),
.B(n_8590),
.Y(n_14608)
);

NAND2xp5_ASAP7_75t_L g14609 ( 
.A(n_13880),
.B(n_11353),
.Y(n_14609)
);

BUFx3_ASAP7_75t_L g14610 ( 
.A(n_13767),
.Y(n_14610)
);

INVx2_ASAP7_75t_L g14611 ( 
.A(n_13139),
.Y(n_14611)
);

AND2x2_ASAP7_75t_L g14612 ( 
.A(n_13782),
.B(n_8645),
.Y(n_14612)
);

AND2x4_ASAP7_75t_L g14613 ( 
.A(n_13439),
.B(n_11355),
.Y(n_14613)
);

NAND2xp5_ASAP7_75t_L g14614 ( 
.A(n_13899),
.B(n_11355),
.Y(n_14614)
);

INVx2_ASAP7_75t_L g14615 ( 
.A(n_13140),
.Y(n_14615)
);

INVx2_ASAP7_75t_L g14616 ( 
.A(n_13113),
.Y(n_14616)
);

AND2x2_ASAP7_75t_L g14617 ( 
.A(n_13770),
.B(n_8645),
.Y(n_14617)
);

INVxp67_ASAP7_75t_SL g14618 ( 
.A(n_13889),
.Y(n_14618)
);

INVx2_ASAP7_75t_L g14619 ( 
.A(n_13694),
.Y(n_14619)
);

OR2x2_ASAP7_75t_L g14620 ( 
.A(n_13681),
.B(n_8238),
.Y(n_14620)
);

NOR2xp67_ASAP7_75t_L g14621 ( 
.A(n_13822),
.B(n_10751),
.Y(n_14621)
);

INVx1_ASAP7_75t_L g14622 ( 
.A(n_13319),
.Y(n_14622)
);

AND2x2_ASAP7_75t_L g14623 ( 
.A(n_13781),
.B(n_8645),
.Y(n_14623)
);

OAI22xp5_ASAP7_75t_L g14624 ( 
.A1(n_13899),
.A2(n_13812),
.B1(n_13825),
.B2(n_13815),
.Y(n_14624)
);

INVx2_ASAP7_75t_L g14625 ( 
.A(n_13694),
.Y(n_14625)
);

AOI22xp33_ASAP7_75t_L g14626 ( 
.A1(n_13830),
.A2(n_8657),
.B1(n_8096),
.B2(n_7265),
.Y(n_14626)
);

INVx1_ASAP7_75t_L g14627 ( 
.A(n_13120),
.Y(n_14627)
);

INVx2_ASAP7_75t_L g14628 ( 
.A(n_13228),
.Y(n_14628)
);

BUFx2_ASAP7_75t_L g14629 ( 
.A(n_13794),
.Y(n_14629)
);

INVx2_ASAP7_75t_L g14630 ( 
.A(n_13233),
.Y(n_14630)
);

INVx1_ASAP7_75t_L g14631 ( 
.A(n_13482),
.Y(n_14631)
);

INVx2_ASAP7_75t_L g14632 ( 
.A(n_13239),
.Y(n_14632)
);

INVx1_ASAP7_75t_L g14633 ( 
.A(n_13502),
.Y(n_14633)
);

HB1xp67_ASAP7_75t_L g14634 ( 
.A(n_13645),
.Y(n_14634)
);

AND2x2_ASAP7_75t_L g14635 ( 
.A(n_13834),
.B(n_8650),
.Y(n_14635)
);

OR2x2_ASAP7_75t_L g14636 ( 
.A(n_13167),
.B(n_13442),
.Y(n_14636)
);

INVx2_ASAP7_75t_SL g14637 ( 
.A(n_13794),
.Y(n_14637)
);

HB1xp67_ASAP7_75t_L g14638 ( 
.A(n_13648),
.Y(n_14638)
);

INVx1_ASAP7_75t_L g14639 ( 
.A(n_13479),
.Y(n_14639)
);

AND2x4_ASAP7_75t_L g14640 ( 
.A(n_13441),
.B(n_11361),
.Y(n_14640)
);

AND2x2_ASAP7_75t_L g14641 ( 
.A(n_13908),
.B(n_8650),
.Y(n_14641)
);

AND2x2_ASAP7_75t_L g14642 ( 
.A(n_13848),
.B(n_8650),
.Y(n_14642)
);

NOR2xp33_ASAP7_75t_L g14643 ( 
.A(n_13842),
.B(n_8738),
.Y(n_14643)
);

OAI222xp33_ASAP7_75t_L g14644 ( 
.A1(n_13709),
.A2(n_10771),
.B1(n_9470),
.B2(n_9460),
.C1(n_9478),
.C2(n_9467),
.Y(n_14644)
);

NOR2xp33_ASAP7_75t_L g14645 ( 
.A(n_13766),
.B(n_8738),
.Y(n_14645)
);

AND2x2_ASAP7_75t_L g14646 ( 
.A(n_13853),
.B(n_8666),
.Y(n_14646)
);

BUFx6f_ASAP7_75t_L g14647 ( 
.A(n_13445),
.Y(n_14647)
);

INVx1_ASAP7_75t_L g14648 ( 
.A(n_13613),
.Y(n_14648)
);

INVxp67_ASAP7_75t_SL g14649 ( 
.A(n_13889),
.Y(n_14649)
);

INVxp67_ASAP7_75t_L g14650 ( 
.A(n_13138),
.Y(n_14650)
);

OAI21xp5_ASAP7_75t_SL g14651 ( 
.A1(n_13722),
.A2(n_8862),
.B(n_8183),
.Y(n_14651)
);

INVx1_ASAP7_75t_L g14652 ( 
.A(n_13614),
.Y(n_14652)
);

NOR2x1_ASAP7_75t_L g14653 ( 
.A(n_13798),
.B(n_10771),
.Y(n_14653)
);

INVx1_ASAP7_75t_L g14654 ( 
.A(n_13600),
.Y(n_14654)
);

INVxp67_ASAP7_75t_SL g14655 ( 
.A(n_13785),
.Y(n_14655)
);

INVx2_ASAP7_75t_L g14656 ( 
.A(n_13261),
.Y(n_14656)
);

OR2x2_ASAP7_75t_L g14657 ( 
.A(n_13786),
.B(n_8238),
.Y(n_14657)
);

INVx1_ASAP7_75t_L g14658 ( 
.A(n_13600),
.Y(n_14658)
);

INVxp67_ASAP7_75t_SL g14659 ( 
.A(n_13785),
.Y(n_14659)
);

NAND2xp33_ASAP7_75t_SL g14660 ( 
.A(n_13785),
.B(n_8095),
.Y(n_14660)
);

INVx2_ASAP7_75t_L g14661 ( 
.A(n_13172),
.Y(n_14661)
);

AOI21xp33_ASAP7_75t_SL g14662 ( 
.A1(n_13353),
.A2(n_9209),
.B(n_7984),
.Y(n_14662)
);

INVx1_ASAP7_75t_L g14663 ( 
.A(n_13609),
.Y(n_14663)
);

NAND2xp5_ASAP7_75t_L g14664 ( 
.A(n_13435),
.B(n_11361),
.Y(n_14664)
);

INVx1_ASAP7_75t_L g14665 ( 
.A(n_13609),
.Y(n_14665)
);

AND2x2_ASAP7_75t_L g14666 ( 
.A(n_13317),
.B(n_8666),
.Y(n_14666)
);

INVx2_ASAP7_75t_L g14667 ( 
.A(n_13656),
.Y(n_14667)
);

INVx2_ASAP7_75t_L g14668 ( 
.A(n_13263),
.Y(n_14668)
);

AND2x2_ASAP7_75t_L g14669 ( 
.A(n_13558),
.B(n_8666),
.Y(n_14669)
);

NAND2xp5_ASAP7_75t_L g14670 ( 
.A(n_13449),
.B(n_11368),
.Y(n_14670)
);

INVx1_ASAP7_75t_L g14671 ( 
.A(n_13617),
.Y(n_14671)
);

INVx1_ASAP7_75t_L g14672 ( 
.A(n_13617),
.Y(n_14672)
);

BUFx2_ASAP7_75t_L g14673 ( 
.A(n_13827),
.Y(n_14673)
);

INVx2_ASAP7_75t_L g14674 ( 
.A(n_13276),
.Y(n_14674)
);

BUFx2_ASAP7_75t_L g14675 ( 
.A(n_13827),
.Y(n_14675)
);

INVx1_ASAP7_75t_SL g14676 ( 
.A(n_13131),
.Y(n_14676)
);

INVxp67_ASAP7_75t_SL g14677 ( 
.A(n_13822),
.Y(n_14677)
);

NAND2xp5_ASAP7_75t_L g14678 ( 
.A(n_13753),
.B(n_11368),
.Y(n_14678)
);

AND2x2_ASAP7_75t_L g14679 ( 
.A(n_13643),
.B(n_8731),
.Y(n_14679)
);

OR2x2_ASAP7_75t_L g14680 ( 
.A(n_13030),
.B(n_8238),
.Y(n_14680)
);

INVx1_ASAP7_75t_SL g14681 ( 
.A(n_13676),
.Y(n_14681)
);

AND2x2_ASAP7_75t_L g14682 ( 
.A(n_13321),
.B(n_8731),
.Y(n_14682)
);

INVx1_ASAP7_75t_L g14683 ( 
.A(n_13510),
.Y(n_14683)
);

INVx3_ASAP7_75t_L g14684 ( 
.A(n_13803),
.Y(n_14684)
);

INVx1_ASAP7_75t_L g14685 ( 
.A(n_13510),
.Y(n_14685)
);

HB1xp67_ASAP7_75t_L g14686 ( 
.A(n_13649),
.Y(n_14686)
);

OAI22xp5_ASAP7_75t_L g14687 ( 
.A1(n_13831),
.A2(n_8142),
.B1(n_8295),
.B2(n_8095),
.Y(n_14687)
);

NAND2xp5_ASAP7_75t_L g14688 ( 
.A(n_13416),
.B(n_11374),
.Y(n_14688)
);

AOI22xp33_ASAP7_75t_SL g14689 ( 
.A1(n_13918),
.A2(n_8377),
.B1(n_8432),
.B2(n_8392),
.Y(n_14689)
);

AND2x2_ASAP7_75t_L g14690 ( 
.A(n_13329),
.B(n_8731),
.Y(n_14690)
);

OR2x2_ASAP7_75t_L g14691 ( 
.A(n_13045),
.B(n_8238),
.Y(n_14691)
);

AND2x2_ASAP7_75t_L g14692 ( 
.A(n_13333),
.B(n_8736),
.Y(n_14692)
);

NAND2xp5_ASAP7_75t_L g14693 ( 
.A(n_13425),
.B(n_11374),
.Y(n_14693)
);

INVx2_ASAP7_75t_L g14694 ( 
.A(n_13700),
.Y(n_14694)
);

AND2x2_ASAP7_75t_L g14695 ( 
.A(n_13337),
.B(n_8736),
.Y(n_14695)
);

INVx2_ASAP7_75t_SL g14696 ( 
.A(n_13803),
.Y(n_14696)
);

AND2x4_ASAP7_75t_L g14697 ( 
.A(n_13448),
.B(n_11379),
.Y(n_14697)
);

INVx1_ASAP7_75t_L g14698 ( 
.A(n_13511),
.Y(n_14698)
);

OR2x2_ASAP7_75t_L g14699 ( 
.A(n_13099),
.B(n_8238),
.Y(n_14699)
);

AND2x2_ASAP7_75t_L g14700 ( 
.A(n_13340),
.B(n_8736),
.Y(n_14700)
);

NOR2xp33_ASAP7_75t_L g14701 ( 
.A(n_13814),
.B(n_8809),
.Y(n_14701)
);

NOR2xp33_ASAP7_75t_L g14702 ( 
.A(n_13849),
.B(n_8809),
.Y(n_14702)
);

NOR2xp33_ASAP7_75t_L g14703 ( 
.A(n_13860),
.B(n_8818),
.Y(n_14703)
);

AND2x4_ASAP7_75t_L g14704 ( 
.A(n_13452),
.B(n_11379),
.Y(n_14704)
);

AND2x2_ASAP7_75t_L g14705 ( 
.A(n_13341),
.B(n_8743),
.Y(n_14705)
);

INVx2_ASAP7_75t_L g14706 ( 
.A(n_13706),
.Y(n_14706)
);

AND2x2_ASAP7_75t_L g14707 ( 
.A(n_13350),
.B(n_8743),
.Y(n_14707)
);

NAND2xp5_ASAP7_75t_L g14708 ( 
.A(n_13844),
.B(n_13845),
.Y(n_14708)
);

NAND2xp5_ASAP7_75t_L g14709 ( 
.A(n_13497),
.B(n_11380),
.Y(n_14709)
);

AND2x2_ASAP7_75t_L g14710 ( 
.A(n_13313),
.B(n_8743),
.Y(n_14710)
);

OR2x2_ASAP7_75t_L g14711 ( 
.A(n_13444),
.B(n_8238),
.Y(n_14711)
);

NAND2xp5_ASAP7_75t_L g14712 ( 
.A(n_13497),
.B(n_11380),
.Y(n_14712)
);

BUFx2_ASAP7_75t_SL g14713 ( 
.A(n_13453),
.Y(n_14713)
);

INVx1_ASAP7_75t_L g14714 ( 
.A(n_13511),
.Y(n_14714)
);

AND2x4_ASAP7_75t_SL g14715 ( 
.A(n_13206),
.B(n_8338),
.Y(n_14715)
);

INVx1_ASAP7_75t_L g14716 ( 
.A(n_13517),
.Y(n_14716)
);

BUFx2_ASAP7_75t_L g14717 ( 
.A(n_13827),
.Y(n_14717)
);

AND2x2_ASAP7_75t_L g14718 ( 
.A(n_13817),
.B(n_8793),
.Y(n_14718)
);

OR2x2_ASAP7_75t_L g14719 ( 
.A(n_13455),
.B(n_8238),
.Y(n_14719)
);

INVx1_ASAP7_75t_L g14720 ( 
.A(n_13517),
.Y(n_14720)
);

INVx2_ASAP7_75t_L g14721 ( 
.A(n_13369),
.Y(n_14721)
);

INVx1_ASAP7_75t_L g14722 ( 
.A(n_13525),
.Y(n_14722)
);

INVxp67_ASAP7_75t_L g14723 ( 
.A(n_13778),
.Y(n_14723)
);

INVx1_ASAP7_75t_L g14724 ( 
.A(n_13525),
.Y(n_14724)
);

INVx2_ASAP7_75t_L g14725 ( 
.A(n_13373),
.Y(n_14725)
);

INVx1_ASAP7_75t_L g14726 ( 
.A(n_13531),
.Y(n_14726)
);

INVx2_ASAP7_75t_SL g14727 ( 
.A(n_13460),
.Y(n_14727)
);

OR2x2_ASAP7_75t_L g14728 ( 
.A(n_13875),
.B(n_8238),
.Y(n_14728)
);

INVx1_ASAP7_75t_L g14729 ( 
.A(n_13531),
.Y(n_14729)
);

INVx4_ASAP7_75t_L g14730 ( 
.A(n_13462),
.Y(n_14730)
);

AND2x2_ASAP7_75t_L g14731 ( 
.A(n_13572),
.B(n_8793),
.Y(n_14731)
);

INVx2_ASAP7_75t_L g14732 ( 
.A(n_13379),
.Y(n_14732)
);

INVx1_ASAP7_75t_L g14733 ( 
.A(n_13384),
.Y(n_14733)
);

AND2x2_ASAP7_75t_L g14734 ( 
.A(n_13355),
.B(n_8793),
.Y(n_14734)
);

BUFx2_ASAP7_75t_L g14735 ( 
.A(n_13826),
.Y(n_14735)
);

AND2x2_ASAP7_75t_L g14736 ( 
.A(n_13533),
.B(n_8180),
.Y(n_14736)
);

INVxp67_ASAP7_75t_L g14737 ( 
.A(n_13808),
.Y(n_14737)
);

INVx2_ASAP7_75t_L g14738 ( 
.A(n_13382),
.Y(n_14738)
);

AOI22xp33_ASAP7_75t_L g14739 ( 
.A1(n_13688),
.A2(n_8657),
.B1(n_8096),
.B2(n_7265),
.Y(n_14739)
);

AND2x2_ASAP7_75t_L g14740 ( 
.A(n_13536),
.B(n_8180),
.Y(n_14740)
);

INVx2_ASAP7_75t_L g14741 ( 
.A(n_14089),
.Y(n_14741)
);

AND2x2_ASAP7_75t_L g14742 ( 
.A(n_13962),
.B(n_13914),
.Y(n_14742)
);

INVx1_ASAP7_75t_L g14743 ( 
.A(n_13931),
.Y(n_14743)
);

INVx2_ASAP7_75t_L g14744 ( 
.A(n_14532),
.Y(n_14744)
);

INVx1_ASAP7_75t_L g14745 ( 
.A(n_13965),
.Y(n_14745)
);

BUFx6f_ASAP7_75t_L g14746 ( 
.A(n_14154),
.Y(n_14746)
);

OA332x1_ASAP7_75t_L g14747 ( 
.A1(n_14624),
.A2(n_13141),
.A3(n_13732),
.B1(n_13349),
.B2(n_13739),
.B3(n_13917),
.C1(n_13840),
.C2(n_13846),
.Y(n_14747)
);

INVx1_ASAP7_75t_L g14748 ( 
.A(n_14436),
.Y(n_14748)
);

OR2x2_ASAP7_75t_L g14749 ( 
.A(n_13927),
.B(n_13740),
.Y(n_14749)
);

AOI22xp5_ASAP7_75t_L g14750 ( 
.A1(n_14217),
.A2(n_13867),
.B1(n_13838),
.B2(n_13809),
.Y(n_14750)
);

OR2x2_ASAP7_75t_L g14751 ( 
.A(n_14325),
.B(n_13574),
.Y(n_14751)
);

BUFx6f_ASAP7_75t_L g14752 ( 
.A(n_14171),
.Y(n_14752)
);

INVx1_ASAP7_75t_L g14753 ( 
.A(n_14466),
.Y(n_14753)
);

INVx2_ASAP7_75t_L g14754 ( 
.A(n_14014),
.Y(n_14754)
);

NAND2xp5_ASAP7_75t_L g14755 ( 
.A(n_14054),
.B(n_13454),
.Y(n_14755)
);

NAND2x1_ASAP7_75t_L g14756 ( 
.A(n_14230),
.B(n_13580),
.Y(n_14756)
);

AND2x4_ASAP7_75t_L g14757 ( 
.A(n_14043),
.B(n_13467),
.Y(n_14757)
);

INVx2_ASAP7_75t_L g14758 ( 
.A(n_14319),
.Y(n_14758)
);

NOR3xp33_ASAP7_75t_L g14759 ( 
.A(n_14087),
.B(n_13828),
.C(n_13891),
.Y(n_14759)
);

HB1xp67_ASAP7_75t_L g14760 ( 
.A(n_13947),
.Y(n_14760)
);

AND2x2_ASAP7_75t_L g14761 ( 
.A(n_14069),
.B(n_13790),
.Y(n_14761)
);

AOI22xp5_ASAP7_75t_L g14762 ( 
.A1(n_13942),
.A2(n_13867),
.B1(n_13802),
.B2(n_13884),
.Y(n_14762)
);

INVx1_ASAP7_75t_L g14763 ( 
.A(n_14473),
.Y(n_14763)
);

AND2x2_ASAP7_75t_L g14764 ( 
.A(n_14291),
.B(n_13792),
.Y(n_14764)
);

HB1xp67_ASAP7_75t_L g14765 ( 
.A(n_14033),
.Y(n_14765)
);

HB1xp67_ASAP7_75t_L g14766 ( 
.A(n_14129),
.Y(n_14766)
);

INVx1_ASAP7_75t_L g14767 ( 
.A(n_14489),
.Y(n_14767)
);

INVxp67_ASAP7_75t_SL g14768 ( 
.A(n_14134),
.Y(n_14768)
);

INVx1_ASAP7_75t_L g14769 ( 
.A(n_14146),
.Y(n_14769)
);

AND2x2_ASAP7_75t_L g14770 ( 
.A(n_14079),
.B(n_13876),
.Y(n_14770)
);

HB1xp67_ASAP7_75t_L g14771 ( 
.A(n_14133),
.Y(n_14771)
);

AND2x2_ASAP7_75t_L g14772 ( 
.A(n_13951),
.B(n_13661),
.Y(n_14772)
);

BUFx3_ASAP7_75t_L g14773 ( 
.A(n_13979),
.Y(n_14773)
);

INVx1_ASAP7_75t_L g14774 ( 
.A(n_14203),
.Y(n_14774)
);

OR2x2_ASAP7_75t_L g14775 ( 
.A(n_14423),
.B(n_13202),
.Y(n_14775)
);

INVx1_ASAP7_75t_L g14776 ( 
.A(n_14204),
.Y(n_14776)
);

NAND2xp5_ASAP7_75t_SL g14777 ( 
.A(n_13998),
.B(n_13852),
.Y(n_14777)
);

INVx2_ASAP7_75t_L g14778 ( 
.A(n_14629),
.Y(n_14778)
);

INVx1_ASAP7_75t_L g14779 ( 
.A(n_14078),
.Y(n_14779)
);

INVx1_ASAP7_75t_L g14780 ( 
.A(n_14103),
.Y(n_14780)
);

AND2x2_ASAP7_75t_L g14781 ( 
.A(n_14211),
.B(n_13892),
.Y(n_14781)
);

NAND2xp5_ASAP7_75t_L g14782 ( 
.A(n_14515),
.B(n_13459),
.Y(n_14782)
);

AND2x2_ASAP7_75t_L g14783 ( 
.A(n_14179),
.B(n_13893),
.Y(n_14783)
);

AND2x2_ASAP7_75t_L g14784 ( 
.A(n_14004),
.B(n_13897),
.Y(n_14784)
);

AND2x2_ASAP7_75t_L g14785 ( 
.A(n_14009),
.B(n_13816),
.Y(n_14785)
);

OAI21xp5_ASAP7_75t_L g14786 ( 
.A1(n_13982),
.A2(n_13887),
.B(n_13866),
.Y(n_14786)
);

NOR2xp33_ASAP7_75t_L g14787 ( 
.A(n_14070),
.B(n_13387),
.Y(n_14787)
);

INVx2_ASAP7_75t_L g14788 ( 
.A(n_14548),
.Y(n_14788)
);

BUFx2_ASAP7_75t_L g14789 ( 
.A(n_14516),
.Y(n_14789)
);

HB1xp67_ASAP7_75t_L g14790 ( 
.A(n_14468),
.Y(n_14790)
);

AND2x2_ASAP7_75t_L g14791 ( 
.A(n_14138),
.B(n_13925),
.Y(n_14791)
);

INVx2_ASAP7_75t_L g14792 ( 
.A(n_14548),
.Y(n_14792)
);

INVx5_ASAP7_75t_L g14793 ( 
.A(n_14140),
.Y(n_14793)
);

AOI22xp33_ASAP7_75t_L g14794 ( 
.A1(n_14561),
.A2(n_13824),
.B1(n_13916),
.B2(n_13900),
.Y(n_14794)
);

NAND2xp5_ASAP7_75t_L g14795 ( 
.A(n_13939),
.B(n_13463),
.Y(n_14795)
);

BUFx6f_ASAP7_75t_L g14796 ( 
.A(n_14171),
.Y(n_14796)
);

NAND2xp5_ASAP7_75t_L g14797 ( 
.A(n_14412),
.B(n_13465),
.Y(n_14797)
);

INVx2_ASAP7_75t_L g14798 ( 
.A(n_14351),
.Y(n_14798)
);

INVx1_ASAP7_75t_L g14799 ( 
.A(n_14497),
.Y(n_14799)
);

AND2x2_ASAP7_75t_L g14800 ( 
.A(n_13948),
.B(n_13588),
.Y(n_14800)
);

AND2x2_ASAP7_75t_L g14801 ( 
.A(n_13950),
.B(n_13675),
.Y(n_14801)
);

INVx2_ASAP7_75t_L g14802 ( 
.A(n_14351),
.Y(n_14802)
);

INVx1_ASAP7_75t_L g14803 ( 
.A(n_14513),
.Y(n_14803)
);

AND2x2_ASAP7_75t_L g14804 ( 
.A(n_14061),
.B(n_13679),
.Y(n_14804)
);

NAND2xp5_ASAP7_75t_L g14805 ( 
.A(n_14221),
.B(n_13475),
.Y(n_14805)
);

INVx1_ASAP7_75t_L g14806 ( 
.A(n_14683),
.Y(n_14806)
);

AND2x2_ASAP7_75t_L g14807 ( 
.A(n_14072),
.B(n_13685),
.Y(n_14807)
);

AND2x2_ASAP7_75t_L g14808 ( 
.A(n_14444),
.B(n_13398),
.Y(n_14808)
);

INVx2_ASAP7_75t_SL g14809 ( 
.A(n_14145),
.Y(n_14809)
);

NAND2xp5_ASAP7_75t_L g14810 ( 
.A(n_14463),
.B(n_13476),
.Y(n_14810)
);

NAND2xp5_ASAP7_75t_L g14811 ( 
.A(n_14479),
.B(n_13499),
.Y(n_14811)
);

INVx1_ASAP7_75t_L g14812 ( 
.A(n_14685),
.Y(n_14812)
);

INVx3_ASAP7_75t_L g14813 ( 
.A(n_14166),
.Y(n_14813)
);

OR2x2_ASAP7_75t_L g14814 ( 
.A(n_14418),
.B(n_13211),
.Y(n_14814)
);

AND2x4_ASAP7_75t_L g14815 ( 
.A(n_14108),
.B(n_13473),
.Y(n_14815)
);

INVx1_ASAP7_75t_L g14816 ( 
.A(n_14698),
.Y(n_14816)
);

AND2x2_ASAP7_75t_L g14817 ( 
.A(n_14321),
.B(n_13400),
.Y(n_14817)
);

AND2x2_ASAP7_75t_L g14818 ( 
.A(n_14017),
.B(n_13403),
.Y(n_14818)
);

BUFx2_ASAP7_75t_L g14819 ( 
.A(n_14516),
.Y(n_14819)
);

AND2x2_ASAP7_75t_L g14820 ( 
.A(n_14088),
.B(n_13406),
.Y(n_14820)
);

NAND2xp5_ASAP7_75t_L g14821 ( 
.A(n_14456),
.B(n_14492),
.Y(n_14821)
);

INVx3_ASAP7_75t_L g14822 ( 
.A(n_14166),
.Y(n_14822)
);

INVx1_ASAP7_75t_L g14823 ( 
.A(n_14714),
.Y(n_14823)
);

INVx1_ASAP7_75t_L g14824 ( 
.A(n_14522),
.Y(n_14824)
);

AND2x2_ASAP7_75t_L g14825 ( 
.A(n_14402),
.B(n_13408),
.Y(n_14825)
);

INVx2_ASAP7_75t_L g14826 ( 
.A(n_13946),
.Y(n_14826)
);

INVx2_ASAP7_75t_L g14827 ( 
.A(n_13946),
.Y(n_14827)
);

AND2x2_ASAP7_75t_L g14828 ( 
.A(n_14428),
.B(n_13413),
.Y(n_14828)
);

BUFx3_ASAP7_75t_L g14829 ( 
.A(n_14108),
.Y(n_14829)
);

AND2x4_ASAP7_75t_L g14830 ( 
.A(n_14417),
.B(n_13481),
.Y(n_14830)
);

AO21x2_ASAP7_75t_L g14831 ( 
.A1(n_14525),
.A2(n_13701),
.B(n_13697),
.Y(n_14831)
);

INVx2_ASAP7_75t_L g14832 ( 
.A(n_13956),
.Y(n_14832)
);

INVx2_ASAP7_75t_L g14833 ( 
.A(n_13956),
.Y(n_14833)
);

INVx2_ASAP7_75t_L g14834 ( 
.A(n_14049),
.Y(n_14834)
);

AND2x2_ASAP7_75t_L g14835 ( 
.A(n_14558),
.B(n_13669),
.Y(n_14835)
);

INVx2_ASAP7_75t_L g14836 ( 
.A(n_14050),
.Y(n_14836)
);

INVx1_ASAP7_75t_L g14837 ( 
.A(n_14544),
.Y(n_14837)
);

AND2x2_ASAP7_75t_L g14838 ( 
.A(n_14545),
.B(n_13585),
.Y(n_14838)
);

BUFx6f_ASAP7_75t_L g14839 ( 
.A(n_14168),
.Y(n_14839)
);

INVx1_ASAP7_75t_L g14840 ( 
.A(n_14557),
.Y(n_14840)
);

INVx2_ASAP7_75t_L g14841 ( 
.A(n_14637),
.Y(n_14841)
);

NAND2xp5_ASAP7_75t_L g14842 ( 
.A(n_14287),
.B(n_13499),
.Y(n_14842)
);

AO21x2_ASAP7_75t_L g14843 ( 
.A1(n_14275),
.A2(n_13707),
.B(n_13702),
.Y(n_14843)
);

NAND2xp5_ASAP7_75t_L g14844 ( 
.A(n_14677),
.B(n_13484),
.Y(n_14844)
);

BUFx3_ASAP7_75t_L g14845 ( 
.A(n_14075),
.Y(n_14845)
);

AND2x2_ASAP7_75t_L g14846 ( 
.A(n_14426),
.B(n_14184),
.Y(n_14846)
);

NOR2x1_ASAP7_75t_L g14847 ( 
.A(n_14565),
.B(n_14735),
.Y(n_14847)
);

INVx2_ASAP7_75t_L g14848 ( 
.A(n_14343),
.Y(n_14848)
);

OR2x2_ASAP7_75t_L g14849 ( 
.A(n_13929),
.B(n_13994),
.Y(n_14849)
);

AND2x2_ASAP7_75t_L g14850 ( 
.A(n_14159),
.B(n_13668),
.Y(n_14850)
);

AND2x2_ASAP7_75t_L g14851 ( 
.A(n_14172),
.B(n_13541),
.Y(n_14851)
);

AND2x2_ASAP7_75t_L g14852 ( 
.A(n_14173),
.B(n_13544),
.Y(n_14852)
);

INVx2_ASAP7_75t_L g14853 ( 
.A(n_14353),
.Y(n_14853)
);

INVx1_ASAP7_75t_L g14854 ( 
.A(n_14587),
.Y(n_14854)
);

AND2x4_ASAP7_75t_L g14855 ( 
.A(n_14040),
.B(n_13486),
.Y(n_14855)
);

INVx1_ASAP7_75t_L g14856 ( 
.A(n_14634),
.Y(n_14856)
);

INVx1_ASAP7_75t_L g14857 ( 
.A(n_14638),
.Y(n_14857)
);

HB1xp67_ASAP7_75t_L g14858 ( 
.A(n_14250),
.Y(n_14858)
);

NOR2xp67_ASAP7_75t_L g14859 ( 
.A(n_14684),
.B(n_13564),
.Y(n_14859)
);

INVx1_ASAP7_75t_L g14860 ( 
.A(n_14686),
.Y(n_14860)
);

INVx2_ASAP7_75t_L g14861 ( 
.A(n_14207),
.Y(n_14861)
);

NAND2xp5_ASAP7_75t_L g14862 ( 
.A(n_14265),
.B(n_13484),
.Y(n_14862)
);

AND2x2_ASAP7_75t_L g14863 ( 
.A(n_14178),
.B(n_13552),
.Y(n_14863)
);

INVx1_ASAP7_75t_L g14864 ( 
.A(n_14716),
.Y(n_14864)
);

INVx3_ASAP7_75t_L g14865 ( 
.A(n_14432),
.Y(n_14865)
);

AND2x2_ASAP7_75t_L g14866 ( 
.A(n_14185),
.B(n_13868),
.Y(n_14866)
);

AND2x2_ASAP7_75t_L g14867 ( 
.A(n_14191),
.B(n_13873),
.Y(n_14867)
);

INVx2_ASAP7_75t_L g14868 ( 
.A(n_14225),
.Y(n_14868)
);

INVx1_ASAP7_75t_L g14869 ( 
.A(n_14720),
.Y(n_14869)
);

NAND2xp5_ASAP7_75t_L g14870 ( 
.A(n_14578),
.B(n_13487),
.Y(n_14870)
);

AO21x2_ASAP7_75t_L g14871 ( 
.A1(n_14280),
.A2(n_13658),
.B(n_13660),
.Y(n_14871)
);

INVx2_ASAP7_75t_L g14872 ( 
.A(n_14233),
.Y(n_14872)
);

INVx5_ASAP7_75t_SL g14873 ( 
.A(n_14467),
.Y(n_14873)
);

INVx2_ASAP7_75t_L g14874 ( 
.A(n_14236),
.Y(n_14874)
);

AND2x4_ASAP7_75t_L g14875 ( 
.A(n_14045),
.B(n_13488),
.Y(n_14875)
);

HB1xp67_ASAP7_75t_L g14876 ( 
.A(n_14621),
.Y(n_14876)
);

OR2x2_ASAP7_75t_L g14877 ( 
.A(n_14537),
.B(n_14504),
.Y(n_14877)
);

NAND2xp5_ASAP7_75t_L g14878 ( 
.A(n_14618),
.B(n_13487),
.Y(n_14878)
);

INVxp67_ASAP7_75t_SL g14879 ( 
.A(n_14429),
.Y(n_14879)
);

BUFx6f_ASAP7_75t_L g14880 ( 
.A(n_13986),
.Y(n_14880)
);

INVx1_ASAP7_75t_L g14881 ( 
.A(n_14722),
.Y(n_14881)
);

INVx1_ASAP7_75t_L g14882 ( 
.A(n_14724),
.Y(n_14882)
);

INVx1_ASAP7_75t_L g14883 ( 
.A(n_14726),
.Y(n_14883)
);

INVx2_ASAP7_75t_L g14884 ( 
.A(n_13976),
.Y(n_14884)
);

INVx2_ASAP7_75t_SL g14885 ( 
.A(n_14432),
.Y(n_14885)
);

INVx2_ASAP7_75t_L g14886 ( 
.A(n_13980),
.Y(n_14886)
);

NAND2xp5_ASAP7_75t_L g14887 ( 
.A(n_14649),
.B(n_13489),
.Y(n_14887)
);

INVx3_ASAP7_75t_L g14888 ( 
.A(n_14258),
.Y(n_14888)
);

AND2x2_ASAP7_75t_L g14889 ( 
.A(n_14201),
.B(n_13466),
.Y(n_14889)
);

INVx5_ASAP7_75t_L g14890 ( 
.A(n_14279),
.Y(n_14890)
);

INVx2_ASAP7_75t_L g14891 ( 
.A(n_14487),
.Y(n_14891)
);

AND2x2_ASAP7_75t_L g14892 ( 
.A(n_14206),
.B(n_13469),
.Y(n_14892)
);

AOI22xp33_ASAP7_75t_L g14893 ( 
.A1(n_13955),
.A2(n_13898),
.B1(n_13642),
.B2(n_13885),
.Y(n_14893)
);

INVx2_ASAP7_75t_SL g14894 ( 
.A(n_14401),
.Y(n_14894)
);

INVx2_ASAP7_75t_L g14895 ( 
.A(n_14487),
.Y(n_14895)
);

INVxp67_ASAP7_75t_L g14896 ( 
.A(n_14308),
.Y(n_14896)
);

INVx3_ASAP7_75t_L g14897 ( 
.A(n_14346),
.Y(n_14897)
);

INVx2_ASAP7_75t_L g14898 ( 
.A(n_14519),
.Y(n_14898)
);

AND2x2_ASAP7_75t_L g14899 ( 
.A(n_13953),
.B(n_13474),
.Y(n_14899)
);

AND2x2_ASAP7_75t_L g14900 ( 
.A(n_14381),
.B(n_13485),
.Y(n_14900)
);

NAND2xp5_ASAP7_75t_L g14901 ( 
.A(n_14386),
.B(n_13489),
.Y(n_14901)
);

INVx2_ASAP7_75t_L g14902 ( 
.A(n_14053),
.Y(n_14902)
);

BUFx2_ASAP7_75t_L g14903 ( 
.A(n_14565),
.Y(n_14903)
);

AND2x2_ASAP7_75t_L g14904 ( 
.A(n_14235),
.B(n_13492),
.Y(n_14904)
);

INVx4_ASAP7_75t_L g14905 ( 
.A(n_13993),
.Y(n_14905)
);

INVx2_ASAP7_75t_L g14906 ( 
.A(n_14058),
.Y(n_14906)
);

BUFx3_ASAP7_75t_L g14907 ( 
.A(n_14015),
.Y(n_14907)
);

AND2x2_ASAP7_75t_L g14908 ( 
.A(n_14357),
.B(n_13493),
.Y(n_14908)
);

INVx1_ASAP7_75t_L g14909 ( 
.A(n_14729),
.Y(n_14909)
);

INVx1_ASAP7_75t_L g14910 ( 
.A(n_14654),
.Y(n_14910)
);

INVx1_ASAP7_75t_L g14911 ( 
.A(n_14658),
.Y(n_14911)
);

INVx1_ASAP7_75t_L g14912 ( 
.A(n_14663),
.Y(n_14912)
);

INVx2_ASAP7_75t_L g14913 ( 
.A(n_14060),
.Y(n_14913)
);

OR2x2_ASAP7_75t_L g14914 ( 
.A(n_14118),
.B(n_13215),
.Y(n_14914)
);

AND2x2_ASAP7_75t_L g14915 ( 
.A(n_14359),
.B(n_13495),
.Y(n_14915)
);

INVx1_ASAP7_75t_L g14916 ( 
.A(n_14665),
.Y(n_14916)
);

NAND2xp5_ASAP7_75t_L g14917 ( 
.A(n_14165),
.B(n_13504),
.Y(n_14917)
);

INVx5_ASAP7_75t_L g14918 ( 
.A(n_14735),
.Y(n_14918)
);

INVx2_ASAP7_75t_L g14919 ( 
.A(n_14068),
.Y(n_14919)
);

INVx4_ASAP7_75t_L g14920 ( 
.A(n_13995),
.Y(n_14920)
);

BUFx2_ASAP7_75t_L g14921 ( 
.A(n_14141),
.Y(n_14921)
);

INVx2_ASAP7_75t_L g14922 ( 
.A(n_14574),
.Y(n_14922)
);

OR2x2_ASAP7_75t_L g14923 ( 
.A(n_14216),
.B(n_13220),
.Y(n_14923)
);

INVx1_ASAP7_75t_L g14924 ( 
.A(n_14671),
.Y(n_14924)
);

HB1xp67_ASAP7_75t_L g14925 ( 
.A(n_14696),
.Y(n_14925)
);

HB1xp67_ASAP7_75t_L g14926 ( 
.A(n_14394),
.Y(n_14926)
);

INVx2_ASAP7_75t_L g14927 ( 
.A(n_14601),
.Y(n_14927)
);

AND2x2_ASAP7_75t_L g14928 ( 
.A(n_14368),
.B(n_13512),
.Y(n_14928)
);

INVx1_ASAP7_75t_L g14929 ( 
.A(n_14672),
.Y(n_14929)
);

BUFx2_ASAP7_75t_L g14930 ( 
.A(n_14177),
.Y(n_14930)
);

INVx2_ASAP7_75t_L g14931 ( 
.A(n_14586),
.Y(n_14931)
);

INVx1_ASAP7_75t_L g14932 ( 
.A(n_13921),
.Y(n_14932)
);

NAND2xp5_ASAP7_75t_L g14933 ( 
.A(n_14512),
.B(n_13505),
.Y(n_14933)
);

BUFx3_ASAP7_75t_L g14934 ( 
.A(n_14020),
.Y(n_14934)
);

AND2x2_ASAP7_75t_L g14935 ( 
.A(n_14379),
.B(n_13818),
.Y(n_14935)
);

HB1xp67_ASAP7_75t_L g14936 ( 
.A(n_14193),
.Y(n_14936)
);

INVxp67_ASAP7_75t_L g14937 ( 
.A(n_14267),
.Y(n_14937)
);

INVx2_ASAP7_75t_L g14938 ( 
.A(n_14589),
.Y(n_14938)
);

INVx2_ASAP7_75t_L g14939 ( 
.A(n_14034),
.Y(n_14939)
);

AND2x2_ASAP7_75t_L g14940 ( 
.A(n_14245),
.B(n_13719),
.Y(n_14940)
);

INVx1_ASAP7_75t_L g14941 ( 
.A(n_14101),
.Y(n_14941)
);

INVx1_ASAP7_75t_L g14942 ( 
.A(n_14102),
.Y(n_14942)
);

INVx1_ASAP7_75t_L g14943 ( 
.A(n_14013),
.Y(n_14943)
);

BUFx2_ASAP7_75t_L g14944 ( 
.A(n_14398),
.Y(n_14944)
);

INVx2_ASAP7_75t_L g14945 ( 
.A(n_14249),
.Y(n_14945)
);

AND2x2_ASAP7_75t_L g14946 ( 
.A(n_14390),
.B(n_13411),
.Y(n_14946)
);

INVx2_ASAP7_75t_L g14947 ( 
.A(n_14080),
.Y(n_14947)
);

INVxp67_ASAP7_75t_SL g14948 ( 
.A(n_14328),
.Y(n_14948)
);

AO21x2_ASAP7_75t_L g14949 ( 
.A1(n_14354),
.A2(n_13729),
.B(n_13863),
.Y(n_14949)
);

AOI22xp5_ASAP7_75t_L g14950 ( 
.A1(n_14073),
.A2(n_13863),
.B1(n_13866),
.B2(n_13854),
.Y(n_14950)
);

BUFx3_ASAP7_75t_L g14951 ( 
.A(n_14031),
.Y(n_14951)
);

OR2x2_ASAP7_75t_L g14952 ( 
.A(n_14541),
.B(n_13230),
.Y(n_14952)
);

INVx2_ASAP7_75t_L g14953 ( 
.A(n_14082),
.Y(n_14953)
);

INVx2_ASAP7_75t_L g14954 ( 
.A(n_14090),
.Y(n_14954)
);

NAND2xp5_ASAP7_75t_L g14955 ( 
.A(n_14016),
.B(n_13509),
.Y(n_14955)
);

NAND2xp5_ASAP7_75t_L g14956 ( 
.A(n_14289),
.B(n_13516),
.Y(n_14956)
);

INVx3_ASAP7_75t_L g14957 ( 
.A(n_14041),
.Y(n_14957)
);

INVx1_ASAP7_75t_L g14958 ( 
.A(n_14013),
.Y(n_14958)
);

NAND2xp5_ASAP7_75t_L g14959 ( 
.A(n_14655),
.B(n_13518),
.Y(n_14959)
);

INVxp67_ASAP7_75t_SL g14960 ( 
.A(n_14021),
.Y(n_14960)
);

HB1xp67_ASAP7_75t_L g14961 ( 
.A(n_14194),
.Y(n_14961)
);

NAND2x1p5_ASAP7_75t_L g14962 ( 
.A(n_14422),
.B(n_14584),
.Y(n_14962)
);

AND2x2_ASAP7_75t_L g14963 ( 
.A(n_14395),
.B(n_13718),
.Y(n_14963)
);

BUFx6f_ASAP7_75t_L g14964 ( 
.A(n_14001),
.Y(n_14964)
);

AND2x2_ASAP7_75t_L g14965 ( 
.A(n_14397),
.B(n_13652),
.Y(n_14965)
);

HB1xp67_ASAP7_75t_L g14966 ( 
.A(n_14341),
.Y(n_14966)
);

INVx1_ASAP7_75t_L g14967 ( 
.A(n_14209),
.Y(n_14967)
);

HB1xp67_ASAP7_75t_L g14968 ( 
.A(n_14210),
.Y(n_14968)
);

NOR2xp33_ASAP7_75t_L g14969 ( 
.A(n_14276),
.B(n_13235),
.Y(n_14969)
);

OR2x2_ASAP7_75t_L g14970 ( 
.A(n_14459),
.B(n_13237),
.Y(n_14970)
);

INVx2_ASAP7_75t_L g14971 ( 
.A(n_14116),
.Y(n_14971)
);

INVx1_ASAP7_75t_L g14972 ( 
.A(n_13932),
.Y(n_14972)
);

INVx1_ASAP7_75t_L g14973 ( 
.A(n_13936),
.Y(n_14973)
);

INVx1_ASAP7_75t_L g14974 ( 
.A(n_13941),
.Y(n_14974)
);

INVx1_ASAP7_75t_L g14975 ( 
.A(n_13952),
.Y(n_14975)
);

AND2x2_ASAP7_75t_L g14976 ( 
.A(n_14410),
.B(n_13587),
.Y(n_14976)
);

AND2x2_ASAP7_75t_L g14977 ( 
.A(n_14414),
.B(n_13292),
.Y(n_14977)
);

INVx2_ASAP7_75t_L g14978 ( 
.A(n_14269),
.Y(n_14978)
);

INVx4_ASAP7_75t_L g14979 ( 
.A(n_14002),
.Y(n_14979)
);

INVxp67_ASAP7_75t_SL g14980 ( 
.A(n_14214),
.Y(n_14980)
);

BUFx2_ASAP7_75t_L g14981 ( 
.A(n_14371),
.Y(n_14981)
);

INVx2_ASAP7_75t_L g14982 ( 
.A(n_14293),
.Y(n_14982)
);

INVx1_ASAP7_75t_L g14983 ( 
.A(n_13958),
.Y(n_14983)
);

INVx2_ASAP7_75t_SL g14984 ( 
.A(n_14132),
.Y(n_14984)
);

NAND2xp5_ASAP7_75t_L g14985 ( 
.A(n_14659),
.B(n_13526),
.Y(n_14985)
);

INVx1_ASAP7_75t_L g14986 ( 
.A(n_13959),
.Y(n_14986)
);

AND2x4_ASAP7_75t_L g14987 ( 
.A(n_14301),
.B(n_14302),
.Y(n_14987)
);

INVx1_ASAP7_75t_L g14988 ( 
.A(n_13961),
.Y(n_14988)
);

INVx2_ASAP7_75t_L g14989 ( 
.A(n_14312),
.Y(n_14989)
);

AND2x2_ASAP7_75t_L g14990 ( 
.A(n_14318),
.B(n_13421),
.Y(n_14990)
);

OR2x2_ASAP7_75t_L g14991 ( 
.A(n_14195),
.B(n_13238),
.Y(n_14991)
);

AND2x2_ASAP7_75t_L g14992 ( 
.A(n_14329),
.B(n_13438),
.Y(n_14992)
);

AND2x2_ASAP7_75t_L g14993 ( 
.A(n_14333),
.B(n_13530),
.Y(n_14993)
);

NAND2xp5_ASAP7_75t_L g14994 ( 
.A(n_14441),
.B(n_13527),
.Y(n_14994)
);

INVx1_ASAP7_75t_L g14995 ( 
.A(n_13967),
.Y(n_14995)
);

INVx2_ASAP7_75t_SL g14996 ( 
.A(n_13964),
.Y(n_14996)
);

AND2x4_ASAP7_75t_L g14997 ( 
.A(n_14237),
.B(n_13535),
.Y(n_14997)
);

INVx1_ASAP7_75t_L g14998 ( 
.A(n_13968),
.Y(n_14998)
);

INVx2_ASAP7_75t_L g14999 ( 
.A(n_14619),
.Y(n_14999)
);

NAND2xp5_ASAP7_75t_L g15000 ( 
.A(n_14588),
.B(n_14374),
.Y(n_15000)
);

INVx1_ASAP7_75t_L g15001 ( 
.A(n_14057),
.Y(n_15001)
);

AND2x2_ASAP7_75t_L g15002 ( 
.A(n_13938),
.B(n_13450),
.Y(n_15002)
);

INVx2_ASAP7_75t_L g15003 ( 
.A(n_14625),
.Y(n_15003)
);

INVx1_ASAP7_75t_L g15004 ( 
.A(n_14062),
.Y(n_15004)
);

INVx4_ASAP7_75t_R g15005 ( 
.A(n_14610),
.Y(n_15005)
);

AND2x2_ASAP7_75t_L g15006 ( 
.A(n_13949),
.B(n_13457),
.Y(n_15006)
);

INVx2_ASAP7_75t_L g15007 ( 
.A(n_14483),
.Y(n_15007)
);

INVx2_ASAP7_75t_L g15008 ( 
.A(n_13999),
.Y(n_15008)
);

INVx8_ASAP7_75t_L g15009 ( 
.A(n_14430),
.Y(n_15009)
);

HB1xp67_ASAP7_75t_L g15010 ( 
.A(n_14244),
.Y(n_15010)
);

OR2x2_ASAP7_75t_L g15011 ( 
.A(n_14514),
.B(n_13267),
.Y(n_15011)
);

HB1xp67_ASAP7_75t_L g15012 ( 
.A(n_14219),
.Y(n_15012)
);

OR2x2_ASAP7_75t_L g15013 ( 
.A(n_14661),
.B(n_13268),
.Y(n_15013)
);

NAND2xp5_ASAP7_75t_L g15014 ( 
.A(n_14374),
.B(n_13540),
.Y(n_15014)
);

NAND2xp5_ASAP7_75t_L g15015 ( 
.A(n_14237),
.B(n_13550),
.Y(n_15015)
);

AND2x2_ASAP7_75t_L g15016 ( 
.A(n_13966),
.B(n_13422),
.Y(n_15016)
);

INVx2_ASAP7_75t_L g15017 ( 
.A(n_13999),
.Y(n_15017)
);

AO21x2_ASAP7_75t_L g15018 ( 
.A1(n_14260),
.A2(n_13729),
.B(n_13755),
.Y(n_15018)
);

INVx2_ASAP7_75t_L g15019 ( 
.A(n_14024),
.Y(n_15019)
);

AND2x2_ASAP7_75t_L g15020 ( 
.A(n_13924),
.B(n_13551),
.Y(n_15020)
);

AND2x2_ASAP7_75t_L g15021 ( 
.A(n_13934),
.B(n_13556),
.Y(n_15021)
);

INVx2_ASAP7_75t_L g15022 ( 
.A(n_14024),
.Y(n_15022)
);

BUFx2_ASAP7_75t_L g15023 ( 
.A(n_14605),
.Y(n_15023)
);

AND2x2_ASAP7_75t_L g15024 ( 
.A(n_13937),
.B(n_14056),
.Y(n_15024)
);

OR2x6_ASAP7_75t_L g15025 ( 
.A(n_14499),
.B(n_14713),
.Y(n_15025)
);

OR2x6_ASAP7_75t_L g15026 ( 
.A(n_14382),
.B(n_13557),
.Y(n_15026)
);

INVx2_ASAP7_75t_L g15027 ( 
.A(n_13964),
.Y(n_15027)
);

INVx2_ASAP7_75t_L g15028 ( 
.A(n_14434),
.Y(n_15028)
);

INVx3_ASAP7_75t_L g15029 ( 
.A(n_14041),
.Y(n_15029)
);

INVx1_ASAP7_75t_SL g15030 ( 
.A(n_14282),
.Y(n_15030)
);

INVx1_ASAP7_75t_L g15031 ( 
.A(n_14063),
.Y(n_15031)
);

INVx2_ASAP7_75t_L g15032 ( 
.A(n_14445),
.Y(n_15032)
);

INVx2_ASAP7_75t_L g15033 ( 
.A(n_14448),
.Y(n_15033)
);

AND2x4_ASAP7_75t_L g15034 ( 
.A(n_14239),
.B(n_13559),
.Y(n_15034)
);

HB1xp67_ASAP7_75t_L g15035 ( 
.A(n_14227),
.Y(n_15035)
);

AND3x1_ASAP7_75t_L g15036 ( 
.A(n_13928),
.B(n_13970),
.C(n_14038),
.Y(n_15036)
);

INVx2_ASAP7_75t_L g15037 ( 
.A(n_14451),
.Y(n_15037)
);

INVxp67_ASAP7_75t_SL g15038 ( 
.A(n_14105),
.Y(n_15038)
);

NAND3xp33_ASAP7_75t_L g15039 ( 
.A(n_13978),
.B(n_13756),
.C(n_13755),
.Y(n_15039)
);

INVx2_ASAP7_75t_L g15040 ( 
.A(n_14452),
.Y(n_15040)
);

BUFx3_ASAP7_75t_L g15041 ( 
.A(n_14239),
.Y(n_15041)
);

INVx2_ASAP7_75t_SL g15042 ( 
.A(n_14051),
.Y(n_15042)
);

AND2x2_ASAP7_75t_L g15043 ( 
.A(n_13984),
.B(n_13657),
.Y(n_15043)
);

INVx1_ASAP7_75t_L g15044 ( 
.A(n_14064),
.Y(n_15044)
);

HB1xp67_ASAP7_75t_L g15045 ( 
.A(n_14238),
.Y(n_15045)
);

INVx2_ASAP7_75t_L g15046 ( 
.A(n_14469),
.Y(n_15046)
);

BUFx3_ASAP7_75t_L g15047 ( 
.A(n_14457),
.Y(n_15047)
);

AND2x2_ASAP7_75t_L g15048 ( 
.A(n_13933),
.B(n_13742),
.Y(n_15048)
);

AND2x2_ASAP7_75t_L g15049 ( 
.A(n_14342),
.B(n_13589),
.Y(n_15049)
);

AND2x2_ASAP7_75t_L g15050 ( 
.A(n_14531),
.B(n_13590),
.Y(n_15050)
);

INVx2_ASAP7_75t_L g15051 ( 
.A(n_14474),
.Y(n_15051)
);

HB1xp67_ASAP7_75t_L g15052 ( 
.A(n_14240),
.Y(n_15052)
);

AND2x2_ASAP7_75t_L g15053 ( 
.A(n_14535),
.B(n_13595),
.Y(n_15053)
);

INVx2_ASAP7_75t_L g15054 ( 
.A(n_14478),
.Y(n_15054)
);

HB1xp67_ASAP7_75t_L g15055 ( 
.A(n_14251),
.Y(n_15055)
);

HB1xp67_ASAP7_75t_L g15056 ( 
.A(n_14268),
.Y(n_15056)
);

AND2x2_ASAP7_75t_L g15057 ( 
.A(n_14507),
.B(n_13687),
.Y(n_15057)
);

BUFx2_ASAP7_75t_L g15058 ( 
.A(n_14371),
.Y(n_15058)
);

INVx1_ASAP7_75t_SL g15059 ( 
.A(n_14157),
.Y(n_15059)
);

HB1xp67_ASAP7_75t_L g15060 ( 
.A(n_13971),
.Y(n_15060)
);

INVx1_ASAP7_75t_L g15061 ( 
.A(n_14065),
.Y(n_15061)
);

HB1xp67_ASAP7_75t_L g15062 ( 
.A(n_14419),
.Y(n_15062)
);

AND2x2_ASAP7_75t_L g15063 ( 
.A(n_14524),
.B(n_13689),
.Y(n_15063)
);

INVx1_ASAP7_75t_L g15064 ( 
.A(n_14071),
.Y(n_15064)
);

INVx1_ASAP7_75t_L g15065 ( 
.A(n_14091),
.Y(n_15065)
);

INVx1_ASAP7_75t_L g15066 ( 
.A(n_14104),
.Y(n_15066)
);

OR2x6_ASAP7_75t_L g15067 ( 
.A(n_14385),
.B(n_14730),
.Y(n_15067)
);

INVx1_ASAP7_75t_L g15068 ( 
.A(n_14550),
.Y(n_15068)
);

INVx2_ASAP7_75t_L g15069 ( 
.A(n_14506),
.Y(n_15069)
);

INVx1_ASAP7_75t_L g15070 ( 
.A(n_13974),
.Y(n_15070)
);

AND2x4_ASAP7_75t_L g15071 ( 
.A(n_14170),
.B(n_13586),
.Y(n_15071)
);

INVx1_ASAP7_75t_L g15072 ( 
.A(n_13975),
.Y(n_15072)
);

INVx2_ASAP7_75t_L g15073 ( 
.A(n_14086),
.Y(n_15073)
);

AND2x2_ASAP7_75t_L g15074 ( 
.A(n_14143),
.B(n_13690),
.Y(n_15074)
);

OR2x2_ASAP7_75t_L g15075 ( 
.A(n_14681),
.B(n_13282),
.Y(n_15075)
);

NOR2x1_ASAP7_75t_L g15076 ( 
.A(n_14419),
.B(n_13328),
.Y(n_15076)
);

INVx1_ASAP7_75t_L g15077 ( 
.A(n_13977),
.Y(n_15077)
);

INVx1_ASAP7_75t_L g15078 ( 
.A(n_13983),
.Y(n_15078)
);

AND2x2_ASAP7_75t_L g15079 ( 
.A(n_14540),
.B(n_13691),
.Y(n_15079)
);

INVx2_ASAP7_75t_L g15080 ( 
.A(n_14086),
.Y(n_15080)
);

AND2x2_ASAP7_75t_L g15081 ( 
.A(n_14551),
.B(n_13720),
.Y(n_15081)
);

AND2x2_ASAP7_75t_L g15082 ( 
.A(n_14556),
.B(n_13300),
.Y(n_15082)
);

AND2x2_ASAP7_75t_L g15083 ( 
.A(n_14560),
.B(n_13703),
.Y(n_15083)
);

INVx3_ASAP7_75t_L g15084 ( 
.A(n_14051),
.Y(n_15084)
);

AOI21xp5_ASAP7_75t_L g15085 ( 
.A1(n_13987),
.A2(n_13957),
.B(n_13922),
.Y(n_15085)
);

AO21x2_ASAP7_75t_L g15086 ( 
.A1(n_14199),
.A2(n_13857),
.B(n_13756),
.Y(n_15086)
);

INVx1_ASAP7_75t_L g15087 ( 
.A(n_13992),
.Y(n_15087)
);

OR2x2_ASAP7_75t_L g15088 ( 
.A(n_14406),
.B(n_13305),
.Y(n_15088)
);

AND2x2_ASAP7_75t_L g15089 ( 
.A(n_14602),
.B(n_13692),
.Y(n_15089)
);

INVx1_ASAP7_75t_L g15090 ( 
.A(n_13996),
.Y(n_15090)
);

INVx1_ASAP7_75t_L g15091 ( 
.A(n_14005),
.Y(n_15091)
);

INVx1_ASAP7_75t_L g15092 ( 
.A(n_14022),
.Y(n_15092)
);

INVx5_ASAP7_75t_L g15093 ( 
.A(n_14511),
.Y(n_15093)
);

INVx1_ASAP7_75t_L g15094 ( 
.A(n_14023),
.Y(n_15094)
);

NAND2x1p5_ASAP7_75t_L g15095 ( 
.A(n_14148),
.B(n_13564),
.Y(n_15095)
);

INVx1_ASAP7_75t_L g15096 ( 
.A(n_14025),
.Y(n_15096)
);

AND2x4_ASAP7_75t_L g15097 ( 
.A(n_14125),
.B(n_13399),
.Y(n_15097)
);

INVx1_ASAP7_75t_L g15098 ( 
.A(n_14026),
.Y(n_15098)
);

BUFx3_ASAP7_75t_L g15099 ( 
.A(n_14647),
.Y(n_15099)
);

AND2x4_ASAP7_75t_L g15100 ( 
.A(n_14416),
.B(n_13852),
.Y(n_15100)
);

INVx1_ASAP7_75t_L g15101 ( 
.A(n_14029),
.Y(n_15101)
);

OR2x2_ASAP7_75t_L g15102 ( 
.A(n_14407),
.B(n_13314),
.Y(n_15102)
);

INVx4_ASAP7_75t_L g15103 ( 
.A(n_14647),
.Y(n_15103)
);

INVx2_ASAP7_75t_L g15104 ( 
.A(n_14590),
.Y(n_15104)
);

AND2x2_ASAP7_75t_L g15105 ( 
.A(n_14604),
.B(n_13628),
.Y(n_15105)
);

NAND2xp5_ASAP7_75t_L g15106 ( 
.A(n_14723),
.B(n_13662),
.Y(n_15106)
);

BUFx3_ASAP7_75t_L g15107 ( 
.A(n_14067),
.Y(n_15107)
);

INVx2_ASAP7_75t_L g15108 ( 
.A(n_14592),
.Y(n_15108)
);

OR2x2_ASAP7_75t_L g15109 ( 
.A(n_14415),
.B(n_13325),
.Y(n_15109)
);

INVx2_ASAP7_75t_L g15110 ( 
.A(n_14467),
.Y(n_15110)
);

AND2x2_ASAP7_75t_L g15111 ( 
.A(n_14611),
.B(n_13912),
.Y(n_15111)
);

AND2x2_ASAP7_75t_L g15112 ( 
.A(n_14615),
.B(n_13664),
.Y(n_15112)
);

NAND2xp5_ASAP7_75t_L g15113 ( 
.A(n_14737),
.B(n_13826),
.Y(n_15113)
);

INVx3_ASAP7_75t_L g15114 ( 
.A(n_14234),
.Y(n_15114)
);

AND2x2_ASAP7_75t_L g15115 ( 
.A(n_14616),
.B(n_13667),
.Y(n_15115)
);

AND2x2_ASAP7_75t_L g15116 ( 
.A(n_14320),
.B(n_13774),
.Y(n_15116)
);

AND2x2_ASAP7_75t_L g15117 ( 
.A(n_14577),
.B(n_13777),
.Y(n_15117)
);

BUFx2_ASAP7_75t_L g15118 ( 
.A(n_14511),
.Y(n_15118)
);

INVx1_ASAP7_75t_L g15119 ( 
.A(n_14030),
.Y(n_15119)
);

INVx1_ASAP7_75t_L g15120 ( 
.A(n_14037),
.Y(n_15120)
);

OAI22xp33_ASAP7_75t_L g15121 ( 
.A1(n_14032),
.A2(n_13991),
.B1(n_14562),
.B2(n_14446),
.Y(n_15121)
);

INVxp67_ASAP7_75t_SL g15122 ( 
.A(n_14048),
.Y(n_15122)
);

INVx1_ASAP7_75t_L g15123 ( 
.A(n_14042),
.Y(n_15123)
);

AND2x2_ASAP7_75t_L g15124 ( 
.A(n_13926),
.B(n_13779),
.Y(n_15124)
);

INVx1_ASAP7_75t_L g15125 ( 
.A(n_14044),
.Y(n_15125)
);

INVx3_ASAP7_75t_L g15126 ( 
.A(n_14234),
.Y(n_15126)
);

INVxp67_ASAP7_75t_L g15127 ( 
.A(n_14012),
.Y(n_15127)
);

AND2x2_ASAP7_75t_L g15128 ( 
.A(n_14628),
.B(n_13783),
.Y(n_15128)
);

AND2x2_ASAP7_75t_L g15129 ( 
.A(n_14630),
.B(n_13801),
.Y(n_15129)
);

NOR2x1_ASAP7_75t_L g15130 ( 
.A(n_14673),
.B(n_13857),
.Y(n_15130)
);

BUFx6f_ASAP7_75t_L g15131 ( 
.A(n_14727),
.Y(n_15131)
);

OR2x2_ASAP7_75t_L g15132 ( 
.A(n_14437),
.B(n_13464),
.Y(n_15132)
);

INVx2_ASAP7_75t_SL g15133 ( 
.A(n_14109),
.Y(n_15133)
);

AND2x4_ASAP7_75t_L g15134 ( 
.A(n_14421),
.B(n_12973),
.Y(n_15134)
);

AND2x2_ASAP7_75t_L g15135 ( 
.A(n_14632),
.B(n_13723),
.Y(n_15135)
);

AND2x2_ASAP7_75t_SL g15136 ( 
.A(n_14636),
.B(n_13580),
.Y(n_15136)
);

AND2x2_ASAP7_75t_L g15137 ( 
.A(n_14656),
.B(n_13735),
.Y(n_15137)
);

AND2x2_ASAP7_75t_L g15138 ( 
.A(n_13990),
.B(n_13610),
.Y(n_15138)
);

INVx2_ASAP7_75t_L g15139 ( 
.A(n_14438),
.Y(n_15139)
);

INVxp67_ASAP7_75t_L g15140 ( 
.A(n_14169),
.Y(n_15140)
);

OR2x2_ASAP7_75t_L g15141 ( 
.A(n_14288),
.B(n_13571),
.Y(n_15141)
);

BUFx3_ASAP7_75t_L g15142 ( 
.A(n_14212),
.Y(n_15142)
);

OR2x2_ASAP7_75t_L g15143 ( 
.A(n_14427),
.B(n_13599),
.Y(n_15143)
);

AO21x2_ASAP7_75t_L g15144 ( 
.A1(n_14549),
.A2(n_13620),
.B(n_13630),
.Y(n_15144)
);

INVx2_ASAP7_75t_L g15145 ( 
.A(n_14438),
.Y(n_15145)
);

INVx2_ASAP7_75t_L g15146 ( 
.A(n_14502),
.Y(n_15146)
);

OR2x2_ASAP7_75t_L g15147 ( 
.A(n_14431),
.B(n_13468),
.Y(n_15147)
);

AND2x4_ASAP7_75t_L g15148 ( 
.A(n_14174),
.B(n_12974),
.Y(n_15148)
);

AND2x2_ASAP7_75t_L g15149 ( 
.A(n_14019),
.B(n_13832),
.Y(n_15149)
);

AND2x2_ASAP7_75t_L g15150 ( 
.A(n_14668),
.B(n_13597),
.Y(n_15150)
);

AND2x2_ASAP7_75t_L g15151 ( 
.A(n_14674),
.B(n_13605),
.Y(n_15151)
);

INVx2_ASAP7_75t_L g15152 ( 
.A(n_14502),
.Y(n_15152)
);

INVx1_ASAP7_75t_L g15153 ( 
.A(n_14047),
.Y(n_15153)
);

HB1xp67_ASAP7_75t_L g15154 ( 
.A(n_14119),
.Y(n_15154)
);

INVx2_ASAP7_75t_L g15155 ( 
.A(n_14190),
.Y(n_15155)
);

AND2x2_ASAP7_75t_L g15156 ( 
.A(n_13943),
.B(n_13883),
.Y(n_15156)
);

AND2x2_ASAP7_75t_L g15157 ( 
.A(n_13944),
.B(n_13833),
.Y(n_15157)
);

AO21x2_ASAP7_75t_L g15158 ( 
.A1(n_14271),
.A2(n_13633),
.B(n_13631),
.Y(n_15158)
);

AND2x2_ASAP7_75t_L g15159 ( 
.A(n_14299),
.B(n_13839),
.Y(n_15159)
);

INVx2_ASAP7_75t_L g15160 ( 
.A(n_14190),
.Y(n_15160)
);

NAND2xp5_ASAP7_75t_L g15161 ( 
.A(n_14142),
.B(n_12987),
.Y(n_15161)
);

INVx2_ASAP7_75t_L g15162 ( 
.A(n_14470),
.Y(n_15162)
);

NAND2xp5_ASAP7_75t_L g15163 ( 
.A(n_14676),
.B(n_12999),
.Y(n_15163)
);

INVx2_ASAP7_75t_L g15164 ( 
.A(n_14470),
.Y(n_15164)
);

AND2x4_ASAP7_75t_L g15165 ( 
.A(n_14149),
.B(n_13851),
.Y(n_15165)
);

BUFx2_ASAP7_75t_L g15166 ( 
.A(n_14675),
.Y(n_15166)
);

INVx1_ASAP7_75t_L g15167 ( 
.A(n_14055),
.Y(n_15167)
);

INVx1_ASAP7_75t_L g15168 ( 
.A(n_13969),
.Y(n_15168)
);

INVx1_ASAP7_75t_SL g15169 ( 
.A(n_14336),
.Y(n_15169)
);

AO21x2_ASAP7_75t_L g15170 ( 
.A1(n_13923),
.A2(n_13374),
.B(n_13532),
.Y(n_15170)
);

AND2x2_ASAP7_75t_L g15171 ( 
.A(n_14300),
.B(n_13713),
.Y(n_15171)
);

AND2x2_ASAP7_75t_L g15172 ( 
.A(n_14183),
.B(n_13746),
.Y(n_15172)
);

INVx1_ASAP7_75t_L g15173 ( 
.A(n_13973),
.Y(n_15173)
);

OR2x2_ASAP7_75t_L g15174 ( 
.A(n_14490),
.B(n_13727),
.Y(n_15174)
);

INVx2_ASAP7_75t_L g15175 ( 
.A(n_14475),
.Y(n_15175)
);

AND2x2_ASAP7_75t_L g15176 ( 
.A(n_13930),
.B(n_13748),
.Y(n_15176)
);

BUFx3_ASAP7_75t_L g15177 ( 
.A(n_14192),
.Y(n_15177)
);

INVx1_ASAP7_75t_L g15178 ( 
.A(n_14092),
.Y(n_15178)
);

INVx1_ASAP7_75t_L g15179 ( 
.A(n_14093),
.Y(n_15179)
);

NAND2x1_ASAP7_75t_L g15180 ( 
.A(n_14475),
.B(n_14215),
.Y(n_15180)
);

AND2x2_ASAP7_75t_L g15181 ( 
.A(n_14231),
.B(n_13750),
.Y(n_15181)
);

NAND2xp5_ASAP7_75t_L g15182 ( 
.A(n_14650),
.B(n_14139),
.Y(n_15182)
);

INVx1_ASAP7_75t_L g15183 ( 
.A(n_14220),
.Y(n_15183)
);

NAND2xp5_ASAP7_75t_L g15184 ( 
.A(n_14396),
.B(n_13634),
.Y(n_15184)
);

BUFx2_ASAP7_75t_L g15185 ( 
.A(n_14717),
.Y(n_15185)
);

AND2x2_ASAP7_75t_L g15186 ( 
.A(n_14635),
.B(n_13752),
.Y(n_15186)
);

HB1xp67_ASAP7_75t_L g15187 ( 
.A(n_14120),
.Y(n_15187)
);

AND2x4_ASAP7_75t_SL g15188 ( 
.A(n_14247),
.B(n_13757),
.Y(n_15188)
);

AND2x2_ASAP7_75t_L g15189 ( 
.A(n_14305),
.B(n_13764),
.Y(n_15189)
);

NAND2xp5_ASAP7_75t_L g15190 ( 
.A(n_14510),
.B(n_13461),
.Y(n_15190)
);

INVx1_ASAP7_75t_SL g15191 ( 
.A(n_13981),
.Y(n_15191)
);

OR2x2_ASAP7_75t_L g15192 ( 
.A(n_14493),
.B(n_13712),
.Y(n_15192)
);

AND2x2_ASAP7_75t_L g15193 ( 
.A(n_14642),
.B(n_13807),
.Y(n_15193)
);

INVx1_ASAP7_75t_L g15194 ( 
.A(n_14222),
.Y(n_15194)
);

OAI33xp33_ASAP7_75t_L g15195 ( 
.A1(n_13940),
.A2(n_13888),
.A3(n_13751),
.B1(n_13741),
.B2(n_13576),
.B3(n_13568),
.Y(n_15195)
);

AND2x2_ASAP7_75t_L g15196 ( 
.A(n_14646),
.B(n_14641),
.Y(n_15196)
);

INVx1_ASAP7_75t_L g15197 ( 
.A(n_14228),
.Y(n_15197)
);

AND2x2_ASAP7_75t_L g15198 ( 
.A(n_14599),
.B(n_13805),
.Y(n_15198)
);

OR2x2_ASAP7_75t_L g15199 ( 
.A(n_14495),
.B(n_13715),
.Y(n_15199)
);

AND2x2_ASAP7_75t_L g15200 ( 
.A(n_14617),
.B(n_13820),
.Y(n_15200)
);

INVx1_ASAP7_75t_L g15201 ( 
.A(n_14242),
.Y(n_15201)
);

AND2x2_ASAP7_75t_L g15202 ( 
.A(n_14623),
.B(n_13823),
.Y(n_15202)
);

INVxp67_ASAP7_75t_L g15203 ( 
.A(n_13945),
.Y(n_15203)
);

AND2x2_ASAP7_75t_L g15204 ( 
.A(n_14317),
.B(n_13878),
.Y(n_15204)
);

AND2x4_ASAP7_75t_L g15205 ( 
.A(n_14595),
.B(n_13851),
.Y(n_15205)
);

AND2x4_ASAP7_75t_L g15206 ( 
.A(n_14598),
.B(n_13850),
.Y(n_15206)
);

AND2x2_ASAP7_75t_L g15207 ( 
.A(n_14110),
.B(n_13283),
.Y(n_15207)
);

HB1xp67_ASAP7_75t_L g15208 ( 
.A(n_14491),
.Y(n_15208)
);

INVx4_ASAP7_75t_L g15209 ( 
.A(n_14480),
.Y(n_15209)
);

INVx1_ASAP7_75t_L g15210 ( 
.A(n_14243),
.Y(n_15210)
);

AND2x2_ASAP7_75t_L g15211 ( 
.A(n_14175),
.B(n_13291),
.Y(n_15211)
);

INVx2_ASAP7_75t_L g15212 ( 
.A(n_14491),
.Y(n_15212)
);

INVx1_ASAP7_75t_L g15213 ( 
.A(n_14248),
.Y(n_15213)
);

AND2x2_ASAP7_75t_L g15214 ( 
.A(n_14462),
.B(n_13913),
.Y(n_15214)
);

AND2x2_ASAP7_75t_L g15215 ( 
.A(n_14292),
.B(n_13920),
.Y(n_15215)
);

HB1xp67_ASAP7_75t_L g15216 ( 
.A(n_14480),
.Y(n_15216)
);

INVx2_ASAP7_75t_L g15217 ( 
.A(n_14097),
.Y(n_15217)
);

INVxp67_ASAP7_75t_L g15218 ( 
.A(n_13989),
.Y(n_15218)
);

INVx2_ASAP7_75t_L g15219 ( 
.A(n_14098),
.Y(n_15219)
);

INVxp67_ASAP7_75t_L g15220 ( 
.A(n_14131),
.Y(n_15220)
);

BUFx3_ASAP7_75t_L g15221 ( 
.A(n_14330),
.Y(n_15221)
);

AND2x4_ASAP7_75t_L g15222 ( 
.A(n_14606),
.B(n_13858),
.Y(n_15222)
);

INVx1_ASAP7_75t_L g15223 ( 
.A(n_14259),
.Y(n_15223)
);

INVx1_ASAP7_75t_SL g15224 ( 
.A(n_14167),
.Y(n_15224)
);

INVx2_ASAP7_75t_L g15225 ( 
.A(n_14100),
.Y(n_15225)
);

AND2x2_ASAP7_75t_L g15226 ( 
.A(n_14298),
.B(n_13395),
.Y(n_15226)
);

AND2x2_ASAP7_75t_L g15227 ( 
.A(n_14213),
.B(n_13437),
.Y(n_15227)
);

BUFx2_ASAP7_75t_L g15228 ( 
.A(n_14527),
.Y(n_15228)
);

OAI31xp33_ASAP7_75t_L g15229 ( 
.A1(n_14008),
.A2(n_14164),
.A3(n_14039),
.B(n_13960),
.Y(n_15229)
);

INVx1_ASAP7_75t_L g15230 ( 
.A(n_14262),
.Y(n_15230)
);

AND2x2_ASAP7_75t_L g15231 ( 
.A(n_14472),
.B(n_13843),
.Y(n_15231)
);

BUFx3_ASAP7_75t_L g15232 ( 
.A(n_14180),
.Y(n_15232)
);

INVx1_ASAP7_75t_L g15233 ( 
.A(n_14264),
.Y(n_15233)
);

HB1xp67_ASAP7_75t_L g15234 ( 
.A(n_14503),
.Y(n_15234)
);

AND2x2_ASAP7_75t_L g15235 ( 
.A(n_14481),
.B(n_13886),
.Y(n_15235)
);

INVx1_ASAP7_75t_L g15236 ( 
.A(n_14266),
.Y(n_15236)
);

INVx2_ASAP7_75t_L g15237 ( 
.A(n_14613),
.Y(n_15237)
);

INVx1_ASAP7_75t_SL g15238 ( 
.A(n_14151),
.Y(n_15238)
);

INVx1_ASAP7_75t_L g15239 ( 
.A(n_14272),
.Y(n_15239)
);

INVx1_ASAP7_75t_SL g15240 ( 
.A(n_14052),
.Y(n_15240)
);

AND2x2_ASAP7_75t_L g15241 ( 
.A(n_14546),
.B(n_13890),
.Y(n_15241)
);

OR2x2_ASAP7_75t_L g15242 ( 
.A(n_13935),
.B(n_13418),
.Y(n_15242)
);

INVx1_ASAP7_75t_L g15243 ( 
.A(n_14283),
.Y(n_15243)
);

BUFx2_ASAP7_75t_L g15244 ( 
.A(n_14509),
.Y(n_15244)
);

AND2x2_ASAP7_75t_L g15245 ( 
.A(n_14007),
.B(n_13894),
.Y(n_15245)
);

INVx1_ASAP7_75t_L g15246 ( 
.A(n_14285),
.Y(n_15246)
);

NAND3xp33_ASAP7_75t_L g15247 ( 
.A(n_13997),
.B(n_13731),
.C(n_13741),
.Y(n_15247)
);

OR2x2_ASAP7_75t_L g15248 ( 
.A(n_14538),
.B(n_13728),
.Y(n_15248)
);

INVxp67_ASAP7_75t_SL g15249 ( 
.A(n_14653),
.Y(n_15249)
);

INVx2_ASAP7_75t_L g15250 ( 
.A(n_14613),
.Y(n_15250)
);

OR2x2_ASAP7_75t_L g15251 ( 
.A(n_14607),
.B(n_13708),
.Y(n_15251)
);

INVxp67_ASAP7_75t_SL g15252 ( 
.A(n_13972),
.Y(n_15252)
);

AND2x2_ASAP7_75t_L g15253 ( 
.A(n_14122),
.B(n_13903),
.Y(n_15253)
);

BUFx2_ASAP7_75t_L g15254 ( 
.A(n_14278),
.Y(n_15254)
);

INVx2_ASAP7_75t_L g15255 ( 
.A(n_14640),
.Y(n_15255)
);

AND2x2_ASAP7_75t_L g15256 ( 
.A(n_14270),
.B(n_13909),
.Y(n_15256)
);

INVx1_ASAP7_75t_L g15257 ( 
.A(n_14286),
.Y(n_15257)
);

AND2x4_ASAP7_75t_L g15258 ( 
.A(n_14639),
.B(n_13359),
.Y(n_15258)
);

INVx1_ASAP7_75t_L g15259 ( 
.A(n_14123),
.Y(n_15259)
);

AND2x2_ASAP7_75t_L g15260 ( 
.A(n_14345),
.B(n_13392),
.Y(n_15260)
);

AND2x2_ASAP7_75t_L g15261 ( 
.A(n_14356),
.B(n_13710),
.Y(n_15261)
);

AND2x4_ASAP7_75t_L g15262 ( 
.A(n_14648),
.B(n_13665),
.Y(n_15262)
);

AND2x4_ASAP7_75t_L g15263 ( 
.A(n_14652),
.B(n_13673),
.Y(n_15263)
);

INVx1_ASAP7_75t_L g15264 ( 
.A(n_14128),
.Y(n_15264)
);

BUFx3_ASAP7_75t_L g15265 ( 
.A(n_14111),
.Y(n_15265)
);

AND2x4_ASAP7_75t_L g15266 ( 
.A(n_14591),
.B(n_13393),
.Y(n_15266)
);

OAI211xp5_ASAP7_75t_L g15267 ( 
.A1(n_13963),
.A2(n_13751),
.B(n_13570),
.C(n_13577),
.Y(n_15267)
);

INVxp67_ASAP7_75t_L g15268 ( 
.A(n_14077),
.Y(n_15268)
);

OR2x2_ASAP7_75t_L g15269 ( 
.A(n_14331),
.B(n_13724),
.Y(n_15269)
);

INVx1_ASAP7_75t_L g15270 ( 
.A(n_14130),
.Y(n_15270)
);

INVx2_ASAP7_75t_L g15271 ( 
.A(n_14640),
.Y(n_15271)
);

NOR2x1p5_ASAP7_75t_L g15272 ( 
.A(n_13988),
.B(n_13394),
.Y(n_15272)
);

INVx3_ASAP7_75t_L g15273 ( 
.A(n_14215),
.Y(n_15273)
);

INVx2_ASAP7_75t_L g15274 ( 
.A(n_14697),
.Y(n_15274)
);

AND2x2_ASAP7_75t_L g15275 ( 
.A(n_14373),
.B(n_13401),
.Y(n_15275)
);

BUFx2_ASAP7_75t_L g15276 ( 
.A(n_14278),
.Y(n_15276)
);

BUFx3_ASAP7_75t_L g15277 ( 
.A(n_14113),
.Y(n_15277)
);

OR2x6_ASAP7_75t_L g15278 ( 
.A(n_14627),
.B(n_13731),
.Y(n_15278)
);

AND2x2_ASAP7_75t_L g15279 ( 
.A(n_14552),
.B(n_13412),
.Y(n_15279)
);

AND2x2_ASAP7_75t_L g15280 ( 
.A(n_14484),
.B(n_13417),
.Y(n_15280)
);

NAND2xp5_ASAP7_75t_L g15281 ( 
.A(n_14223),
.B(n_14224),
.Y(n_15281)
);

OR2x2_ASAP7_75t_L g15282 ( 
.A(n_14252),
.B(n_13725),
.Y(n_15282)
);

INVx2_ASAP7_75t_L g15283 ( 
.A(n_14697),
.Y(n_15283)
);

OAI21xp5_ASAP7_75t_L g15284 ( 
.A1(n_14182),
.A2(n_13579),
.B(n_13567),
.Y(n_15284)
);

INVx2_ASAP7_75t_L g15285 ( 
.A(n_14704),
.Y(n_15285)
);

INVx2_ASAP7_75t_L g15286 ( 
.A(n_14704),
.Y(n_15286)
);

INVx1_ASAP7_75t_L g15287 ( 
.A(n_14137),
.Y(n_15287)
);

INVx1_ASAP7_75t_L g15288 ( 
.A(n_14147),
.Y(n_15288)
);

INVx3_ASAP7_75t_L g15289 ( 
.A(n_14715),
.Y(n_15289)
);

INVx1_ASAP7_75t_L g15290 ( 
.A(n_14152),
.Y(n_15290)
);

AND2x2_ASAP7_75t_L g15291 ( 
.A(n_14494),
.B(n_13428),
.Y(n_15291)
);

NAND2xp5_ASAP7_75t_L g15292 ( 
.A(n_14593),
.B(n_13743),
.Y(n_15292)
);

INVx1_ASAP7_75t_L g15293 ( 
.A(n_14160),
.Y(n_15293)
);

INVx2_ASAP7_75t_L g15294 ( 
.A(n_14608),
.Y(n_15294)
);

INVx1_ASAP7_75t_L g15295 ( 
.A(n_14161),
.Y(n_15295)
);

INVx1_ASAP7_75t_L g15296 ( 
.A(n_14162),
.Y(n_15296)
);

INVx1_ASAP7_75t_L g15297 ( 
.A(n_14176),
.Y(n_15297)
);

AND2x2_ASAP7_75t_L g15298 ( 
.A(n_14405),
.B(n_13745),
.Y(n_15298)
);

INVx1_ASAP7_75t_L g15299 ( 
.A(n_14181),
.Y(n_15299)
);

INVx1_ASAP7_75t_L g15300 ( 
.A(n_14186),
.Y(n_15300)
);

INVx1_ASAP7_75t_L g15301 ( 
.A(n_14188),
.Y(n_15301)
);

INVx1_ASAP7_75t_L g15302 ( 
.A(n_14197),
.Y(n_15302)
);

HB1xp67_ASAP7_75t_L g15303 ( 
.A(n_14306),
.Y(n_15303)
);

BUFx3_ASAP7_75t_L g15304 ( 
.A(n_14117),
.Y(n_15304)
);

BUFx2_ASAP7_75t_L g15305 ( 
.A(n_14306),
.Y(n_15305)
);

INVx2_ASAP7_75t_L g15306 ( 
.A(n_14094),
.Y(n_15306)
);

OA21x2_ASAP7_75t_L g15307 ( 
.A1(n_14156),
.A2(n_13534),
.B(n_13532),
.Y(n_15307)
);

OR2x2_ASAP7_75t_L g15308 ( 
.A(n_14296),
.B(n_13534),
.Y(n_15308)
);

NAND2xp5_ASAP7_75t_L g15309 ( 
.A(n_14106),
.B(n_14107),
.Y(n_15309)
);

INVx2_ASAP7_75t_L g15310 ( 
.A(n_14095),
.Y(n_15310)
);

INVx1_ASAP7_75t_L g15311 ( 
.A(n_14198),
.Y(n_15311)
);

HB1xp67_ASAP7_75t_L g15312 ( 
.A(n_14340),
.Y(n_15312)
);

AND2x2_ASAP7_75t_L g15313 ( 
.A(n_14520),
.B(n_13537),
.Y(n_15313)
);

HB1xp67_ASAP7_75t_L g15314 ( 
.A(n_14340),
.Y(n_15314)
);

NAND2xp5_ASAP7_75t_L g15315 ( 
.A(n_14112),
.B(n_13537),
.Y(n_15315)
);

INVx2_ASAP7_75t_L g15316 ( 
.A(n_14347),
.Y(n_15316)
);

AND2x2_ASAP7_75t_L g15317 ( 
.A(n_14536),
.B(n_13542),
.Y(n_15317)
);

AND2x2_ASAP7_75t_L g15318 ( 
.A(n_14542),
.B(n_13542),
.Y(n_15318)
);

INVx1_ASAP7_75t_L g15319 ( 
.A(n_14202),
.Y(n_15319)
);

AND2x2_ASAP7_75t_L g15320 ( 
.A(n_14326),
.B(n_13543),
.Y(n_15320)
);

OR2x2_ASAP7_75t_L g15321 ( 
.A(n_14035),
.B(n_13543),
.Y(n_15321)
);

AND2x2_ASAP7_75t_L g15322 ( 
.A(n_14439),
.B(n_13555),
.Y(n_15322)
);

INVxp67_ASAP7_75t_L g15323 ( 
.A(n_14000),
.Y(n_15323)
);

AND2x2_ASAP7_75t_L g15324 ( 
.A(n_14501),
.B(n_13555),
.Y(n_15324)
);

OR2x2_ASAP7_75t_L g15325 ( 
.A(n_14498),
.B(n_13584),
.Y(n_15325)
);

AND2x2_ASAP7_75t_L g15326 ( 
.A(n_14447),
.B(n_13584),
.Y(n_15326)
);

AND2x2_ASAP7_75t_L g15327 ( 
.A(n_14450),
.B(n_13598),
.Y(n_15327)
);

AND2x2_ASAP7_75t_L g15328 ( 
.A(n_14338),
.B(n_13598),
.Y(n_15328)
);

NOR2x1_ASAP7_75t_R g15329 ( 
.A(n_14708),
.B(n_14200),
.Y(n_15329)
);

INVx2_ASAP7_75t_L g15330 ( 
.A(n_14347),
.Y(n_15330)
);

INVx5_ASAP7_75t_SL g15331 ( 
.A(n_14553),
.Y(n_15331)
);

INVx1_ASAP7_75t_L g15332 ( 
.A(n_14205),
.Y(n_15332)
);

INVx1_ASAP7_75t_L g15333 ( 
.A(n_14208),
.Y(n_15333)
);

AND2x2_ASAP7_75t_L g15334 ( 
.A(n_14567),
.B(n_11382),
.Y(n_15334)
);

AND2x2_ASAP7_75t_L g15335 ( 
.A(n_14579),
.B(n_11382),
.Y(n_15335)
);

INVx5_ASAP7_75t_L g15336 ( 
.A(n_14393),
.Y(n_15336)
);

AND2x2_ASAP7_75t_L g15337 ( 
.A(n_14582),
.B(n_11385),
.Y(n_15337)
);

AND2x4_ASAP7_75t_L g15338 ( 
.A(n_14733),
.B(n_8615),
.Y(n_15338)
);

INVx3_ASAP7_75t_L g15339 ( 
.A(n_14569),
.Y(n_15339)
);

INVx2_ASAP7_75t_L g15340 ( 
.A(n_14393),
.Y(n_15340)
);

INVx2_ASAP7_75t_SL g15341 ( 
.A(n_14409),
.Y(n_15341)
);

NAND2x1_ASAP7_75t_L g15342 ( 
.A(n_14409),
.B(n_14455),
.Y(n_15342)
);

AND2x2_ASAP7_75t_L g15343 ( 
.A(n_14583),
.B(n_14028),
.Y(n_15343)
);

AND2x2_ASAP7_75t_L g15344 ( 
.A(n_14046),
.B(n_14631),
.Y(n_15344)
);

INVxp67_ASAP7_75t_L g15345 ( 
.A(n_14643),
.Y(n_15345)
);

INVxp67_ASAP7_75t_L g15346 ( 
.A(n_14126),
.Y(n_15346)
);

INVx4_ASAP7_75t_L g15347 ( 
.A(n_14114),
.Y(n_15347)
);

AND2x2_ASAP7_75t_L g15348 ( 
.A(n_14633),
.B(n_11385),
.Y(n_15348)
);

INVx2_ASAP7_75t_L g15349 ( 
.A(n_14666),
.Y(n_15349)
);

AND2x2_ASAP7_75t_L g15350 ( 
.A(n_14254),
.B(n_11386),
.Y(n_15350)
);

AND2x2_ASAP7_75t_L g15351 ( 
.A(n_14255),
.B(n_11386),
.Y(n_15351)
);

INVx2_ASAP7_75t_L g15352 ( 
.A(n_14455),
.Y(n_15352)
);

INVx2_ASAP7_75t_L g15353 ( 
.A(n_14734),
.Y(n_15353)
);

OR2x2_ASAP7_75t_L g15354 ( 
.A(n_14334),
.B(n_13731),
.Y(n_15354)
);

INVx2_ASAP7_75t_L g15355 ( 
.A(n_14553),
.Y(n_15355)
);

AND2x4_ASAP7_75t_L g15356 ( 
.A(n_14121),
.B(n_8615),
.Y(n_15356)
);

AND2x2_ASAP7_75t_L g15357 ( 
.A(n_14603),
.B(n_14622),
.Y(n_15357)
);

BUFx2_ASAP7_75t_L g15358 ( 
.A(n_14660),
.Y(n_15358)
);

AND2x2_ASAP7_75t_L g15359 ( 
.A(n_14612),
.B(n_11417),
.Y(n_15359)
);

INVx2_ASAP7_75t_L g15360 ( 
.A(n_14710),
.Y(n_15360)
);

AOI22xp33_ASAP7_75t_SL g15361 ( 
.A1(n_14435),
.A2(n_8432),
.B1(n_8392),
.B2(n_8095),
.Y(n_15361)
);

INVx1_ASAP7_75t_L g15362 ( 
.A(n_14135),
.Y(n_15362)
);

OR2x2_ASAP7_75t_L g15363 ( 
.A(n_14314),
.B(n_11417),
.Y(n_15363)
);

AND2x2_ASAP7_75t_L g15364 ( 
.A(n_14309),
.B(n_11425),
.Y(n_15364)
);

OAI211xp5_ASAP7_75t_L g15365 ( 
.A1(n_13985),
.A2(n_12792),
.B(n_11065),
.C(n_11066),
.Y(n_15365)
);

NOR2x1_ASAP7_75t_L g15366 ( 
.A(n_14667),
.B(n_14694),
.Y(n_15366)
);

AND2x2_ASAP7_75t_L g15367 ( 
.A(n_14315),
.B(n_14332),
.Y(n_15367)
);

INVx2_ASAP7_75t_L g15368 ( 
.A(n_14682),
.Y(n_15368)
);

BUFx6f_ASAP7_75t_L g15369 ( 
.A(n_14721),
.Y(n_15369)
);

INVx1_ASAP7_75t_L g15370 ( 
.A(n_14196),
.Y(n_15370)
);

NAND2xp5_ASAP7_75t_L g15371 ( 
.A(n_14701),
.B(n_11425),
.Y(n_15371)
);

NAND3xp33_ASAP7_75t_L g15372 ( 
.A(n_14036),
.B(n_11065),
.C(n_11059),
.Y(n_15372)
);

INVx2_ASAP7_75t_L g15373 ( 
.A(n_14690),
.Y(n_15373)
);

OR2x2_ASAP7_75t_L g15374 ( 
.A(n_14115),
.B(n_11427),
.Y(n_15374)
);

HB1xp67_ASAP7_75t_L g15375 ( 
.A(n_14533),
.Y(n_15375)
);

HB1xp67_ASAP7_75t_L g15376 ( 
.A(n_14533),
.Y(n_15376)
);

INVx2_ASAP7_75t_L g15377 ( 
.A(n_14692),
.Y(n_15377)
);

INVx3_ASAP7_75t_L g15378 ( 
.A(n_14257),
.Y(n_15378)
);

OR2x6_ASAP7_75t_L g15379 ( 
.A(n_14307),
.B(n_14274),
.Y(n_15379)
);

HB1xp67_ASAP7_75t_L g15380 ( 
.A(n_14433),
.Y(n_15380)
);

AND2x2_ASAP7_75t_L g15381 ( 
.A(n_14731),
.B(n_11427),
.Y(n_15381)
);

AND2x2_ASAP7_75t_L g15382 ( 
.A(n_14261),
.B(n_11429),
.Y(n_15382)
);

AOI22xp33_ASAP7_75t_SL g15383 ( 
.A1(n_14163),
.A2(n_8095),
.B1(n_8295),
.B2(n_8142),
.Y(n_15383)
);

AND2x2_ASAP7_75t_L g15384 ( 
.A(n_14281),
.B(n_11429),
.Y(n_15384)
);

AND2x2_ASAP7_75t_L g15385 ( 
.A(n_14669),
.B(n_14695),
.Y(n_15385)
);

INVx3_ASAP7_75t_L g15386 ( 
.A(n_14253),
.Y(n_15386)
);

INVx1_ASAP7_75t_L g15387 ( 
.A(n_14076),
.Y(n_15387)
);

INVx2_ASAP7_75t_L g15388 ( 
.A(n_14700),
.Y(n_15388)
);

INVx2_ASAP7_75t_L g15389 ( 
.A(n_14705),
.Y(n_15389)
);

INVx1_ASAP7_75t_L g15390 ( 
.A(n_14337),
.Y(n_15390)
);

INVx2_ASAP7_75t_L g15391 ( 
.A(n_14707),
.Y(n_15391)
);

HB1xp67_ASAP7_75t_L g15392 ( 
.A(n_14440),
.Y(n_15392)
);

AND2x2_ASAP7_75t_L g15393 ( 
.A(n_14387),
.B(n_11434),
.Y(n_15393)
);

INVx2_ASAP7_75t_L g15394 ( 
.A(n_14596),
.Y(n_15394)
);

INVx1_ASAP7_75t_L g15395 ( 
.A(n_14362),
.Y(n_15395)
);

INVx1_ASAP7_75t_L g15396 ( 
.A(n_14375),
.Y(n_15396)
);

CKINVDCx6p67_ASAP7_75t_R g15397 ( 
.A(n_14391),
.Y(n_15397)
);

INVx1_ASAP7_75t_L g15398 ( 
.A(n_14377),
.Y(n_15398)
);

INVx4_ASAP7_75t_L g15399 ( 
.A(n_14155),
.Y(n_15399)
);

OAI33xp33_ASAP7_75t_L g15400 ( 
.A1(n_14006),
.A2(n_11066),
.A3(n_11059),
.B1(n_11295),
.B2(n_11300),
.B3(n_11289),
.Y(n_15400)
);

AND2x2_ASAP7_75t_L g15401 ( 
.A(n_14408),
.B(n_11434),
.Y(n_15401)
);

INVx1_ASAP7_75t_L g15402 ( 
.A(n_14555),
.Y(n_15402)
);

INVx1_ASAP7_75t_L g15403 ( 
.A(n_14378),
.Y(n_15403)
);

AND2x2_ASAP7_75t_L g15404 ( 
.A(n_14411),
.B(n_11439),
.Y(n_15404)
);

OR2x2_ASAP7_75t_L g15405 ( 
.A(n_14580),
.B(n_11439),
.Y(n_15405)
);

AOI221xp5_ASAP7_75t_L g15406 ( 
.A1(n_14018),
.A2(n_11300),
.B1(n_11301),
.B2(n_11295),
.C(n_11289),
.Y(n_15406)
);

INVx2_ASAP7_75t_L g15407 ( 
.A(n_14706),
.Y(n_15407)
);

OAI22xp33_ASAP7_75t_L g15408 ( 
.A1(n_14657),
.A2(n_8295),
.B1(n_8430),
.B2(n_8142),
.Y(n_15408)
);

AND2x2_ASAP7_75t_L g15409 ( 
.A(n_14424),
.B(n_14003),
.Y(n_15409)
);

INVx1_ASAP7_75t_L g15410 ( 
.A(n_14581),
.Y(n_15410)
);

AND2x2_ASAP7_75t_L g15411 ( 
.A(n_14718),
.B(n_11448),
.Y(n_15411)
);

INVx1_ASAP7_75t_L g15412 ( 
.A(n_14678),
.Y(n_15412)
);

HB1xp67_ASAP7_75t_L g15413 ( 
.A(n_14263),
.Y(n_15413)
);

NOR2xp67_ASAP7_75t_L g15414 ( 
.A(n_14597),
.B(n_11448),
.Y(n_15414)
);

INVx5_ASAP7_75t_L g15415 ( 
.A(n_14725),
.Y(n_15415)
);

INVx1_ASAP7_75t_L g15416 ( 
.A(n_14277),
.Y(n_15416)
);

AND2x2_ASAP7_75t_L g15417 ( 
.A(n_14679),
.B(n_11450),
.Y(n_15417)
);

HB1xp67_ASAP7_75t_L g15418 ( 
.A(n_14355),
.Y(n_15418)
);

INVx2_ASAP7_75t_L g15419 ( 
.A(n_14732),
.Y(n_15419)
);

INVx2_ASAP7_75t_L g15420 ( 
.A(n_14738),
.Y(n_15420)
);

INVx1_ASAP7_75t_L g15421 ( 
.A(n_14232),
.Y(n_15421)
);

HB1xp67_ASAP7_75t_L g15422 ( 
.A(n_14614),
.Y(n_15422)
);

NAND2x1p5_ASAP7_75t_L g15423 ( 
.A(n_14290),
.B(n_7790),
.Y(n_15423)
);

AND2x2_ASAP7_75t_L g15424 ( 
.A(n_14645),
.B(n_11450),
.Y(n_15424)
);

AND2x2_ASAP7_75t_L g15425 ( 
.A(n_14702),
.B(n_11452),
.Y(n_15425)
);

AOI22xp33_ASAP7_75t_SL g15426 ( 
.A1(n_14027),
.A2(n_8142),
.B1(n_8430),
.B2(n_8295),
.Y(n_15426)
);

INVx2_ASAP7_75t_L g15427 ( 
.A(n_14158),
.Y(n_15427)
);

AND2x2_ASAP7_75t_L g15428 ( 
.A(n_14703),
.B(n_11452),
.Y(n_15428)
);

BUFx2_ASAP7_75t_L g15429 ( 
.A(n_14600),
.Y(n_15429)
);

BUFx2_ASAP7_75t_L g15430 ( 
.A(n_14609),
.Y(n_15430)
);

BUFx2_ASAP7_75t_L g15431 ( 
.A(n_14554),
.Y(n_15431)
);

NOR3xp33_ASAP7_75t_L g15432 ( 
.A(n_13954),
.B(n_11302),
.C(n_11301),
.Y(n_15432)
);

AND2x2_ASAP7_75t_L g15433 ( 
.A(n_14011),
.B(n_11455),
.Y(n_15433)
);

CKINVDCx20_ASAP7_75t_R g15434 ( 
.A(n_14284),
.Y(n_15434)
);

INVx1_ASAP7_75t_L g15435 ( 
.A(n_14241),
.Y(n_15435)
);

AND2x4_ASAP7_75t_L g15436 ( 
.A(n_14294),
.B(n_8615),
.Y(n_15436)
);

INVx2_ASAP7_75t_L g15437 ( 
.A(n_14420),
.Y(n_15437)
);

INVx2_ASAP7_75t_L g15438 ( 
.A(n_14153),
.Y(n_15438)
);

INVx2_ASAP7_75t_L g15439 ( 
.A(n_14523),
.Y(n_15439)
);

AND2x2_ASAP7_75t_L g15440 ( 
.A(n_14505),
.B(n_11455),
.Y(n_15440)
);

INVx2_ASAP7_75t_L g15441 ( 
.A(n_14295),
.Y(n_15441)
);

BUFx12f_ASAP7_75t_L g15442 ( 
.A(n_14568),
.Y(n_15442)
);

BUFx6f_ASAP7_75t_L g15443 ( 
.A(n_14059),
.Y(n_15443)
);

INVx3_ASAP7_75t_L g15444 ( 
.A(n_14297),
.Y(n_15444)
);

AND2x2_ASAP7_75t_L g15445 ( 
.A(n_14485),
.B(n_11473),
.Y(n_15445)
);

AND2x2_ASAP7_75t_L g15446 ( 
.A(n_14304),
.B(n_11473),
.Y(n_15446)
);

INVx2_ASAP7_75t_L g15447 ( 
.A(n_14310),
.Y(n_15447)
);

AND2x2_ASAP7_75t_L g15448 ( 
.A(n_14651),
.B(n_11478),
.Y(n_15448)
);

OR2x2_ASAP7_75t_L g15449 ( 
.A(n_14303),
.B(n_11478),
.Y(n_15449)
);

BUFx2_ASAP7_75t_L g15450 ( 
.A(n_14488),
.Y(n_15450)
);

AND2x4_ASAP7_75t_L g15451 ( 
.A(n_14311),
.B(n_8615),
.Y(n_15451)
);

INVx2_ASAP7_75t_L g15452 ( 
.A(n_14313),
.Y(n_15452)
);

INVx2_ASAP7_75t_SL g15453 ( 
.A(n_14066),
.Y(n_15453)
);

INVxp67_ASAP7_75t_L g15454 ( 
.A(n_14566),
.Y(n_15454)
);

AND2x2_ASAP7_75t_L g15455 ( 
.A(n_14366),
.B(n_11483),
.Y(n_15455)
);

INVx2_ASAP7_75t_L g15456 ( 
.A(n_15336),
.Y(n_15456)
);

OR2x2_ASAP7_75t_L g15457 ( 
.A(n_14821),
.B(n_14521),
.Y(n_15457)
);

INVx1_ASAP7_75t_L g15458 ( 
.A(n_14903),
.Y(n_15458)
);

INVx1_ASAP7_75t_L g15459 ( 
.A(n_14903),
.Y(n_15459)
);

OR2x2_ASAP7_75t_L g15460 ( 
.A(n_15191),
.B(n_14335),
.Y(n_15460)
);

OR2x2_ASAP7_75t_L g15461 ( 
.A(n_14760),
.B(n_14364),
.Y(n_15461)
);

OR2x2_ASAP7_75t_L g15462 ( 
.A(n_14790),
.B(n_14085),
.Y(n_15462)
);

AND2x2_ASAP7_75t_L g15463 ( 
.A(n_14846),
.B(n_14367),
.Y(n_15463)
);

INVx1_ASAP7_75t_L g15464 ( 
.A(n_14981),
.Y(n_15464)
);

AND2x2_ASAP7_75t_L g15465 ( 
.A(n_14773),
.B(n_14380),
.Y(n_15465)
);

AND2x2_ASAP7_75t_L g15466 ( 
.A(n_14962),
.B(n_14388),
.Y(n_15466)
);

AND2x2_ASAP7_75t_L g15467 ( 
.A(n_14900),
.B(n_14454),
.Y(n_15467)
);

OR2x2_ASAP7_75t_L g15468 ( 
.A(n_14849),
.B(n_14074),
.Y(n_15468)
);

INVx3_ASAP7_75t_L g15469 ( 
.A(n_15009),
.Y(n_15469)
);

INVx1_ASAP7_75t_L g15470 ( 
.A(n_14981),
.Y(n_15470)
);

AND2x4_ASAP7_75t_L g15471 ( 
.A(n_14829),
.B(n_14322),
.Y(n_15471)
);

INVx1_ASAP7_75t_L g15472 ( 
.A(n_15058),
.Y(n_15472)
);

AND2x4_ASAP7_75t_SL g15473 ( 
.A(n_14746),
.B(n_14323),
.Y(n_15473)
);

NAND2xp5_ASAP7_75t_L g15474 ( 
.A(n_15059),
.B(n_14425),
.Y(n_15474)
);

OR2x2_ASAP7_75t_L g15475 ( 
.A(n_15000),
.B(n_14081),
.Y(n_15475)
);

AND2x2_ASAP7_75t_L g15476 ( 
.A(n_14925),
.B(n_14327),
.Y(n_15476)
);

AND2x4_ASAP7_75t_L g15477 ( 
.A(n_15041),
.B(n_14339),
.Y(n_15477)
);

AND2x2_ASAP7_75t_L g15478 ( 
.A(n_14783),
.B(n_14344),
.Y(n_15478)
);

INVx1_ASAP7_75t_L g15479 ( 
.A(n_15058),
.Y(n_15479)
);

INVx1_ASAP7_75t_L g15480 ( 
.A(n_15118),
.Y(n_15480)
);

HB1xp67_ASAP7_75t_L g15481 ( 
.A(n_15336),
.Y(n_15481)
);

AND2x4_ASAP7_75t_SL g15482 ( 
.A(n_14746),
.B(n_14348),
.Y(n_15482)
);

AND2x2_ASAP7_75t_L g15483 ( 
.A(n_14904),
.B(n_14349),
.Y(n_15483)
);

OR2x2_ASAP7_75t_L g15484 ( 
.A(n_14936),
.B(n_14961),
.Y(n_15484)
);

INVx2_ASAP7_75t_L g15485 ( 
.A(n_15336),
.Y(n_15485)
);

INVx1_ASAP7_75t_L g15486 ( 
.A(n_15118),
.Y(n_15486)
);

AND2x2_ASAP7_75t_L g15487 ( 
.A(n_14764),
.B(n_14350),
.Y(n_15487)
);

INVx1_ASAP7_75t_SL g15488 ( 
.A(n_15009),
.Y(n_15488)
);

INVx2_ASAP7_75t_L g15489 ( 
.A(n_15276),
.Y(n_15489)
);

INVx1_ASAP7_75t_L g15490 ( 
.A(n_14918),
.Y(n_15490)
);

NAND2xp5_ASAP7_75t_L g15491 ( 
.A(n_15038),
.B(n_14885),
.Y(n_15491)
);

AND2x2_ASAP7_75t_L g15492 ( 
.A(n_14761),
.B(n_14352),
.Y(n_15492)
);

INVx1_ASAP7_75t_L g15493 ( 
.A(n_14918),
.Y(n_15493)
);

INVx1_ASAP7_75t_L g15494 ( 
.A(n_14918),
.Y(n_15494)
);

OR2x2_ASAP7_75t_L g15495 ( 
.A(n_15169),
.B(n_14083),
.Y(n_15495)
);

INVx1_ASAP7_75t_L g15496 ( 
.A(n_15093),
.Y(n_15496)
);

AND2x2_ASAP7_75t_L g15497 ( 
.A(n_14813),
.B(n_14822),
.Y(n_15497)
);

INVx2_ASAP7_75t_L g15498 ( 
.A(n_15276),
.Y(n_15498)
);

AND2x2_ASAP7_75t_L g15499 ( 
.A(n_14791),
.B(n_14358),
.Y(n_15499)
);

OR2x2_ASAP7_75t_L g15500 ( 
.A(n_14930),
.B(n_14084),
.Y(n_15500)
);

INVx1_ASAP7_75t_L g15501 ( 
.A(n_15093),
.Y(n_15501)
);

NOR2xp33_ASAP7_75t_SL g15502 ( 
.A(n_15103),
.B(n_14644),
.Y(n_15502)
);

AND2x2_ASAP7_75t_L g15503 ( 
.A(n_14888),
.B(n_14361),
.Y(n_15503)
);

INVx4_ASAP7_75t_L g15504 ( 
.A(n_14890),
.Y(n_15504)
);

NAND2xp5_ASAP7_75t_L g15505 ( 
.A(n_14768),
.B(n_14365),
.Y(n_15505)
);

NAND2xp5_ASAP7_75t_SL g15506 ( 
.A(n_14839),
.B(n_14010),
.Y(n_15506)
);

NAND2xp5_ASAP7_75t_L g15507 ( 
.A(n_14865),
.B(n_14369),
.Y(n_15507)
);

INVx1_ASAP7_75t_L g15508 ( 
.A(n_15093),
.Y(n_15508)
);

INVx1_ASAP7_75t_L g15509 ( 
.A(n_15305),
.Y(n_15509)
);

INVx1_ASAP7_75t_L g15510 ( 
.A(n_15305),
.Y(n_15510)
);

AND2x4_ASAP7_75t_L g15511 ( 
.A(n_14890),
.B(n_14376),
.Y(n_15511)
);

INVx1_ASAP7_75t_L g15512 ( 
.A(n_14847),
.Y(n_15512)
);

AND2x2_ASAP7_75t_L g15513 ( 
.A(n_14897),
.B(n_14383),
.Y(n_15513)
);

OR2x2_ASAP7_75t_L g15514 ( 
.A(n_14758),
.B(n_14778),
.Y(n_15514)
);

AND2x2_ASAP7_75t_L g15515 ( 
.A(n_14838),
.B(n_14384),
.Y(n_15515)
);

AND2x2_ASAP7_75t_L g15516 ( 
.A(n_15049),
.B(n_14389),
.Y(n_15516)
);

AND2x2_ASAP7_75t_L g15517 ( 
.A(n_14809),
.B(n_14392),
.Y(n_15517)
);

HB1xp67_ASAP7_75t_L g15518 ( 
.A(n_15060),
.Y(n_15518)
);

INVx1_ASAP7_75t_L g15519 ( 
.A(n_15375),
.Y(n_15519)
);

INVx1_ASAP7_75t_L g15520 ( 
.A(n_15376),
.Y(n_15520)
);

AND2x4_ASAP7_75t_L g15521 ( 
.A(n_14890),
.B(n_14399),
.Y(n_15521)
);

INVx1_ASAP7_75t_L g15522 ( 
.A(n_15062),
.Y(n_15522)
);

INVx1_ASAP7_75t_L g15523 ( 
.A(n_14766),
.Y(n_15523)
);

AND2x4_ASAP7_75t_L g15524 ( 
.A(n_15142),
.B(n_15177),
.Y(n_15524)
);

INVx2_ASAP7_75t_L g15525 ( 
.A(n_14793),
.Y(n_15525)
);

INVx1_ASAP7_75t_L g15526 ( 
.A(n_14771),
.Y(n_15526)
);

INVx2_ASAP7_75t_L g15527 ( 
.A(n_14793),
.Y(n_15527)
);

INVx1_ASAP7_75t_L g15528 ( 
.A(n_15166),
.Y(n_15528)
);

HB1xp67_ASAP7_75t_L g15529 ( 
.A(n_15208),
.Y(n_15529)
);

NAND2xp5_ASAP7_75t_L g15530 ( 
.A(n_14858),
.B(n_14404),
.Y(n_15530)
);

NAND2xp5_ASAP7_75t_L g15531 ( 
.A(n_15140),
.B(n_14518),
.Y(n_15531)
);

NAND2xp5_ASAP7_75t_L g15532 ( 
.A(n_14765),
.B(n_14526),
.Y(n_15532)
);

OR2x2_ASAP7_75t_L g15533 ( 
.A(n_14751),
.B(n_14096),
.Y(n_15533)
);

OR2x2_ASAP7_75t_L g15534 ( 
.A(n_15154),
.B(n_14124),
.Y(n_15534)
);

INVx1_ASAP7_75t_L g15535 ( 
.A(n_15166),
.Y(n_15535)
);

OR2x2_ASAP7_75t_L g15536 ( 
.A(n_15187),
.B(n_14127),
.Y(n_15536)
);

AND2x4_ASAP7_75t_L g15537 ( 
.A(n_15232),
.B(n_15221),
.Y(n_15537)
);

AND2x2_ASAP7_75t_L g15538 ( 
.A(n_14742),
.B(n_14528),
.Y(n_15538)
);

NAND2xp5_ASAP7_75t_L g15539 ( 
.A(n_14839),
.B(n_14529),
.Y(n_15539)
);

INVx1_ASAP7_75t_L g15540 ( 
.A(n_15185),
.Y(n_15540)
);

NAND2xp5_ASAP7_75t_L g15541 ( 
.A(n_14815),
.B(n_14530),
.Y(n_15541)
);

BUFx2_ASAP7_75t_L g15542 ( 
.A(n_15249),
.Y(n_15542)
);

HB1xp67_ASAP7_75t_L g15543 ( 
.A(n_15342),
.Y(n_15543)
);

HB1xp67_ASAP7_75t_L g15544 ( 
.A(n_15216),
.Y(n_15544)
);

BUFx2_ASAP7_75t_L g15545 ( 
.A(n_14789),
.Y(n_15545)
);

NAND2x1_ASAP7_75t_L g15546 ( 
.A(n_15005),
.B(n_14534),
.Y(n_15546)
);

AND2x2_ASAP7_75t_L g15547 ( 
.A(n_15343),
.B(n_14539),
.Y(n_15547)
);

AND2x2_ASAP7_75t_L g15548 ( 
.A(n_15007),
.B(n_14543),
.Y(n_15548)
);

NOR2xp33_ASAP7_75t_R g15549 ( 
.A(n_15434),
.B(n_14547),
.Y(n_15549)
);

INVx3_ASAP7_75t_L g15550 ( 
.A(n_15209),
.Y(n_15550)
);

AND2x2_ASAP7_75t_L g15551 ( 
.A(n_14770),
.B(n_14559),
.Y(n_15551)
);

INVx1_ASAP7_75t_L g15552 ( 
.A(n_15185),
.Y(n_15552)
);

AND2x2_ASAP7_75t_L g15553 ( 
.A(n_14817),
.B(n_14563),
.Y(n_15553)
);

INVx2_ASAP7_75t_L g15554 ( 
.A(n_14793),
.Y(n_15554)
);

AND2x2_ASAP7_75t_L g15555 ( 
.A(n_15006),
.B(n_14564),
.Y(n_15555)
);

AND2x2_ASAP7_75t_L g15556 ( 
.A(n_14976),
.B(n_14573),
.Y(n_15556)
);

NAND2xp5_ASAP7_75t_L g15557 ( 
.A(n_14948),
.B(n_14575),
.Y(n_15557)
);

NAND2xp5_ASAP7_75t_SL g15558 ( 
.A(n_14752),
.B(n_14099),
.Y(n_15558)
);

AND2x2_ASAP7_75t_L g15559 ( 
.A(n_15196),
.B(n_14442),
.Y(n_15559)
);

OR2x2_ASAP7_75t_L g15560 ( 
.A(n_14745),
.B(n_14136),
.Y(n_15560)
);

NOR2xp67_ASAP7_75t_L g15561 ( 
.A(n_14876),
.B(n_14443),
.Y(n_15561)
);

INVx1_ASAP7_75t_L g15562 ( 
.A(n_14789),
.Y(n_15562)
);

NAND2xp5_ASAP7_75t_L g15563 ( 
.A(n_14943),
.B(n_14144),
.Y(n_15563)
);

NAND2xp5_ASAP7_75t_L g15564 ( 
.A(n_14958),
.B(n_14187),
.Y(n_15564)
);

INVx2_ASAP7_75t_L g15565 ( 
.A(n_15254),
.Y(n_15565)
);

OR2x2_ASAP7_75t_L g15566 ( 
.A(n_14926),
.B(n_14189),
.Y(n_15566)
);

AND2x2_ASAP7_75t_L g15567 ( 
.A(n_14800),
.B(n_14449),
.Y(n_15567)
);

NAND2xp5_ASAP7_75t_L g15568 ( 
.A(n_14966),
.B(n_14570),
.Y(n_15568)
);

NOR2x1_ASAP7_75t_SL g15569 ( 
.A(n_15025),
.B(n_14453),
.Y(n_15569)
);

NOR2xp33_ASAP7_75t_L g15570 ( 
.A(n_14896),
.B(n_14571),
.Y(n_15570)
);

AND2x2_ASAP7_75t_L g15571 ( 
.A(n_15025),
.B(n_14458),
.Y(n_15571)
);

OR2x2_ASAP7_75t_L g15572 ( 
.A(n_14749),
.B(n_14363),
.Y(n_15572)
);

INVx1_ASAP7_75t_L g15573 ( 
.A(n_14819),
.Y(n_15573)
);

AND2x2_ASAP7_75t_L g15574 ( 
.A(n_14899),
.B(n_14460),
.Y(n_15574)
);

INVx2_ASAP7_75t_L g15575 ( 
.A(n_15331),
.Y(n_15575)
);

OR2x2_ASAP7_75t_L g15576 ( 
.A(n_15023),
.B(n_14877),
.Y(n_15576)
);

INVx1_ASAP7_75t_L g15577 ( 
.A(n_14819),
.Y(n_15577)
);

INVx1_ASAP7_75t_L g15578 ( 
.A(n_15303),
.Y(n_15578)
);

INVx1_ASAP7_75t_L g15579 ( 
.A(n_15312),
.Y(n_15579)
);

NAND2xp5_ASAP7_75t_L g15580 ( 
.A(n_15024),
.B(n_14585),
.Y(n_15580)
);

AND2x4_ASAP7_75t_L g15581 ( 
.A(n_15047),
.B(n_14464),
.Y(n_15581)
);

INVx1_ASAP7_75t_L g15582 ( 
.A(n_15314),
.Y(n_15582)
);

OAI21xp33_ASAP7_75t_L g15583 ( 
.A1(n_14762),
.A2(n_14739),
.B(n_14594),
.Y(n_15583)
);

NAND2xp5_ASAP7_75t_L g15584 ( 
.A(n_14921),
.B(n_14256),
.Y(n_15584)
);

NAND2xp5_ASAP7_75t_L g15585 ( 
.A(n_14997),
.B(n_14465),
.Y(n_15585)
);

INVx1_ASAP7_75t_L g15586 ( 
.A(n_15012),
.Y(n_15586)
);

NAND2x1_ASAP7_75t_L g15587 ( 
.A(n_15114),
.B(n_14471),
.Y(n_15587)
);

AND2x2_ASAP7_75t_L g15588 ( 
.A(n_14965),
.B(n_14476),
.Y(n_15588)
);

OR2x2_ASAP7_75t_L g15589 ( 
.A(n_14955),
.B(n_14994),
.Y(n_15589)
);

OAI22xp5_ASAP7_75t_L g15590 ( 
.A1(n_14756),
.A2(n_14728),
.B1(n_14316),
.B2(n_14218),
.Y(n_15590)
);

OR2x2_ASAP7_75t_L g15591 ( 
.A(n_14775),
.B(n_14572),
.Y(n_15591)
);

AND2x4_ASAP7_75t_SL g15592 ( 
.A(n_14752),
.B(n_14477),
.Y(n_15592)
);

INVx2_ASAP7_75t_L g15593 ( 
.A(n_15331),
.Y(n_15593)
);

AND2x2_ASAP7_75t_L g15594 ( 
.A(n_14807),
.B(n_14482),
.Y(n_15594)
);

INVx1_ASAP7_75t_L g15595 ( 
.A(n_15035),
.Y(n_15595)
);

NOR2xp33_ASAP7_75t_L g15596 ( 
.A(n_14796),
.B(n_14576),
.Y(n_15596)
);

NAND2xp5_ASAP7_75t_L g15597 ( 
.A(n_15162),
.B(n_14486),
.Y(n_15597)
);

INVx3_ASAP7_75t_L g15598 ( 
.A(n_14796),
.Y(n_15598)
);

INVx2_ASAP7_75t_L g15599 ( 
.A(n_15126),
.Y(n_15599)
);

INVx2_ASAP7_75t_L g15600 ( 
.A(n_14744),
.Y(n_15600)
);

AND2x2_ASAP7_75t_L g15601 ( 
.A(n_14946),
.B(n_14508),
.Y(n_15601)
);

BUFx3_ASAP7_75t_L g15602 ( 
.A(n_15131),
.Y(n_15602)
);

OR2x2_ASAP7_75t_L g15603 ( 
.A(n_15218),
.B(n_14517),
.Y(n_15603)
);

INVxp67_ASAP7_75t_R g15604 ( 
.A(n_15045),
.Y(n_15604)
);

HB1xp67_ASAP7_75t_L g15605 ( 
.A(n_14859),
.Y(n_15605)
);

NAND2xp5_ASAP7_75t_L g15606 ( 
.A(n_15164),
.B(n_14664),
.Y(n_15606)
);

INVx1_ASAP7_75t_L g15607 ( 
.A(n_15052),
.Y(n_15607)
);

NAND2xp5_ASAP7_75t_L g15608 ( 
.A(n_15175),
.B(n_14670),
.Y(n_15608)
);

NAND2x1p5_ASAP7_75t_L g15609 ( 
.A(n_14845),
.B(n_14688),
.Y(n_15609)
);

INVx1_ASAP7_75t_L g15610 ( 
.A(n_15055),
.Y(n_15610)
);

INVx1_ASAP7_75t_L g15611 ( 
.A(n_15056),
.Y(n_15611)
);

INVxp67_ASAP7_75t_SL g15612 ( 
.A(n_15130),
.Y(n_15612)
);

HB1xp67_ASAP7_75t_L g15613 ( 
.A(n_15380),
.Y(n_15613)
);

NAND2xp5_ASAP7_75t_L g15614 ( 
.A(n_15212),
.B(n_14693),
.Y(n_15614)
);

OR2x2_ASAP7_75t_L g15615 ( 
.A(n_14743),
.B(n_14709),
.Y(n_15615)
);

NAND2xp5_ASAP7_75t_L g15616 ( 
.A(n_14987),
.B(n_14712),
.Y(n_15616)
);

INVx1_ASAP7_75t_L g15617 ( 
.A(n_14968),
.Y(n_15617)
);

INVx2_ASAP7_75t_L g15618 ( 
.A(n_14880),
.Y(n_15618)
);

INVx1_ASAP7_75t_L g15619 ( 
.A(n_15244),
.Y(n_15619)
);

HB1xp67_ASAP7_75t_L g15620 ( 
.A(n_15392),
.Y(n_15620)
);

INVx1_ASAP7_75t_L g15621 ( 
.A(n_15234),
.Y(n_15621)
);

NAND2xp5_ASAP7_75t_L g15622 ( 
.A(n_15002),
.B(n_14150),
.Y(n_15622)
);

AND2x2_ASAP7_75t_L g15623 ( 
.A(n_14781),
.B(n_14736),
.Y(n_15623)
);

NAND2xp5_ASAP7_75t_L g15624 ( 
.A(n_14944),
.B(n_14740),
.Y(n_15624)
);

OR2x2_ASAP7_75t_L g15625 ( 
.A(n_14779),
.B(n_14620),
.Y(n_15625)
);

AND2x2_ASAP7_75t_L g15626 ( 
.A(n_14835),
.B(n_15048),
.Y(n_15626)
);

INVx1_ASAP7_75t_L g15627 ( 
.A(n_14769),
.Y(n_15627)
);

INVx2_ASAP7_75t_L g15628 ( 
.A(n_14880),
.Y(n_15628)
);

AND2x4_ASAP7_75t_L g15629 ( 
.A(n_14907),
.B(n_14680),
.Y(n_15629)
);

INVx2_ASAP7_75t_L g15630 ( 
.A(n_15095),
.Y(n_15630)
);

AND2x4_ASAP7_75t_L g15631 ( 
.A(n_14934),
.B(n_14691),
.Y(n_15631)
);

OR2x2_ASAP7_75t_L g15632 ( 
.A(n_14780),
.B(n_14711),
.Y(n_15632)
);

NOR2xp33_ASAP7_75t_L g15633 ( 
.A(n_15127),
.B(n_14662),
.Y(n_15633)
);

INVx2_ASAP7_75t_L g15634 ( 
.A(n_15131),
.Y(n_15634)
);

NAND2xp5_ASAP7_75t_L g15635 ( 
.A(n_15030),
.B(n_14830),
.Y(n_15635)
);

AND2x2_ASAP7_75t_L g15636 ( 
.A(n_14892),
.B(n_14413),
.Y(n_15636)
);

AND2x2_ASAP7_75t_L g15637 ( 
.A(n_14908),
.B(n_14226),
.Y(n_15637)
);

OR2x2_ASAP7_75t_L g15638 ( 
.A(n_14923),
.B(n_14719),
.Y(n_15638)
);

INVx3_ASAP7_75t_L g15639 ( 
.A(n_15034),
.Y(n_15639)
);

INVxp67_ASAP7_75t_L g15640 ( 
.A(n_15450),
.Y(n_15640)
);

NOR3xp33_ASAP7_75t_L g15641 ( 
.A(n_15121),
.B(n_15039),
.C(n_14786),
.Y(n_15641)
);

INVx1_ASAP7_75t_SL g15642 ( 
.A(n_15450),
.Y(n_15642)
);

AND2x2_ASAP7_75t_L g15643 ( 
.A(n_14915),
.B(n_14699),
.Y(n_15643)
);

INVx1_ASAP7_75t_L g15644 ( 
.A(n_14774),
.Y(n_15644)
);

HB1xp67_ASAP7_75t_L g15645 ( 
.A(n_15026),
.Y(n_15645)
);

HB1xp67_ASAP7_75t_L g15646 ( 
.A(n_15026),
.Y(n_15646)
);

AND2x2_ASAP7_75t_L g15647 ( 
.A(n_14928),
.B(n_14687),
.Y(n_15647)
);

INVx1_ASAP7_75t_L g15648 ( 
.A(n_14776),
.Y(n_15648)
);

INVx1_ASAP7_75t_L g15649 ( 
.A(n_15313),
.Y(n_15649)
);

INVx2_ASAP7_75t_L g15650 ( 
.A(n_14957),
.Y(n_15650)
);

NAND2xp5_ASAP7_75t_L g15651 ( 
.A(n_14922),
.B(n_14496),
.Y(n_15651)
);

NAND2x1p5_ASAP7_75t_L g15652 ( 
.A(n_15099),
.B(n_7790),
.Y(n_15652)
);

INVx2_ASAP7_75t_L g15653 ( 
.A(n_15029),
.Y(n_15653)
);

NAND2x1p5_ASAP7_75t_L g15654 ( 
.A(n_14757),
.B(n_7790),
.Y(n_15654)
);

AND2x4_ASAP7_75t_L g15655 ( 
.A(n_14951),
.B(n_8624),
.Y(n_15655)
);

NAND2xp5_ASAP7_75t_L g15656 ( 
.A(n_14927),
.B(n_14626),
.Y(n_15656)
);

OR2x2_ASAP7_75t_L g15657 ( 
.A(n_14917),
.B(n_14273),
.Y(n_15657)
);

NAND2xp5_ASAP7_75t_L g15658 ( 
.A(n_14905),
.B(n_14324),
.Y(n_15658)
);

INVx1_ASAP7_75t_L g15659 ( 
.A(n_15317),
.Y(n_15659)
);

NAND3x1_ASAP7_75t_SL g15660 ( 
.A(n_15229),
.B(n_14246),
.C(n_14461),
.Y(n_15660)
);

INVx2_ASAP7_75t_L g15661 ( 
.A(n_15084),
.Y(n_15661)
);

AND2x2_ASAP7_75t_L g15662 ( 
.A(n_14889),
.B(n_14689),
.Y(n_15662)
);

AND2x2_ASAP7_75t_L g15663 ( 
.A(n_14992),
.B(n_14229),
.Y(n_15663)
);

AND2x2_ASAP7_75t_L g15664 ( 
.A(n_14993),
.B(n_14370),
.Y(n_15664)
);

NAND2xp5_ASAP7_75t_L g15665 ( 
.A(n_14920),
.B(n_14400),
.Y(n_15665)
);

INVx1_ASAP7_75t_L g15666 ( 
.A(n_15318),
.Y(n_15666)
);

AND2x2_ASAP7_75t_L g15667 ( 
.A(n_14990),
.B(n_14825),
.Y(n_15667)
);

HB1xp67_ASAP7_75t_L g15668 ( 
.A(n_15415),
.Y(n_15668)
);

INVx1_ASAP7_75t_L g15669 ( 
.A(n_15322),
.Y(n_15669)
);

AND2x2_ASAP7_75t_L g15670 ( 
.A(n_14808),
.B(n_11483),
.Y(n_15670)
);

INVx1_ASAP7_75t_L g15671 ( 
.A(n_15324),
.Y(n_15671)
);

NOR3xp33_ASAP7_75t_L g15672 ( 
.A(n_15247),
.B(n_14360),
.C(n_11303),
.Y(n_15672)
);

NAND2xp5_ASAP7_75t_SL g15673 ( 
.A(n_15228),
.B(n_15165),
.Y(n_15673)
);

NOR2xp33_ASAP7_75t_L g15674 ( 
.A(n_14741),
.B(n_11497),
.Y(n_15674)
);

OR2x2_ASAP7_75t_L g15675 ( 
.A(n_14799),
.B(n_14500),
.Y(n_15675)
);

AND2x2_ASAP7_75t_L g15676 ( 
.A(n_14891),
.B(n_14895),
.Y(n_15676)
);

HB1xp67_ASAP7_75t_L g15677 ( 
.A(n_15415),
.Y(n_15677)
);

HB1xp67_ASAP7_75t_L g15678 ( 
.A(n_15415),
.Y(n_15678)
);

AND2x2_ASAP7_75t_L g15679 ( 
.A(n_14804),
.B(n_11497),
.Y(n_15679)
);

BUFx2_ASAP7_75t_L g15680 ( 
.A(n_15076),
.Y(n_15680)
);

HB1xp67_ASAP7_75t_L g15681 ( 
.A(n_15067),
.Y(n_15681)
);

NAND2xp5_ASAP7_75t_L g15682 ( 
.A(n_14979),
.B(n_14372),
.Y(n_15682)
);

AND2x2_ASAP7_75t_L g15683 ( 
.A(n_14851),
.B(n_11500),
.Y(n_15683)
);

INVx1_ASAP7_75t_L g15684 ( 
.A(n_15326),
.Y(n_15684)
);

INVx2_ASAP7_75t_L g15685 ( 
.A(n_15358),
.Y(n_15685)
);

AND2x2_ASAP7_75t_L g15686 ( 
.A(n_14852),
.B(n_14863),
.Y(n_15686)
);

AND2x2_ASAP7_75t_L g15687 ( 
.A(n_15020),
.B(n_11500),
.Y(n_15687)
);

NAND2x1p5_ASAP7_75t_L g15688 ( 
.A(n_14984),
.B(n_7792),
.Y(n_15688)
);

INVx1_ASAP7_75t_L g15689 ( 
.A(n_15327),
.Y(n_15689)
);

INVx1_ASAP7_75t_L g15690 ( 
.A(n_14803),
.Y(n_15690)
);

INVx2_ASAP7_75t_L g15691 ( 
.A(n_15358),
.Y(n_15691)
);

AND2x2_ASAP7_75t_L g15692 ( 
.A(n_14828),
.B(n_11504),
.Y(n_15692)
);

OR2x2_ASAP7_75t_L g15693 ( 
.A(n_14805),
.B(n_14403),
.Y(n_15693)
);

AND2x2_ASAP7_75t_L g15694 ( 
.A(n_14963),
.B(n_11504),
.Y(n_15694)
);

INVx1_ASAP7_75t_L g15695 ( 
.A(n_14871),
.Y(n_15695)
);

INVx1_ASAP7_75t_L g15696 ( 
.A(n_14748),
.Y(n_15696)
);

INVx1_ASAP7_75t_L g15697 ( 
.A(n_14753),
.Y(n_15697)
);

OR2x2_ASAP7_75t_L g15698 ( 
.A(n_14914),
.B(n_11507),
.Y(n_15698)
);

INVx1_ASAP7_75t_L g15699 ( 
.A(n_14763),
.Y(n_15699)
);

AND2x2_ASAP7_75t_L g15700 ( 
.A(n_14801),
.B(n_11507),
.Y(n_15700)
);

OR2x2_ASAP7_75t_L g15701 ( 
.A(n_14755),
.B(n_11509),
.Y(n_15701)
);

OR2x2_ASAP7_75t_L g15702 ( 
.A(n_15224),
.B(n_11509),
.Y(n_15702)
);

AND2x2_ASAP7_75t_L g15703 ( 
.A(n_14820),
.B(n_11513),
.Y(n_15703)
);

OR2x2_ASAP7_75t_L g15704 ( 
.A(n_15238),
.B(n_11513),
.Y(n_15704)
);

INVx1_ASAP7_75t_L g15705 ( 
.A(n_14767),
.Y(n_15705)
);

NOR2xp33_ASAP7_75t_L g15706 ( 
.A(n_14960),
.B(n_11515),
.Y(n_15706)
);

NAND2x1p5_ASAP7_75t_L g15707 ( 
.A(n_15265),
.B(n_7792),
.Y(n_15707)
);

AND2x2_ASAP7_75t_L g15708 ( 
.A(n_14935),
.B(n_11515),
.Y(n_15708)
);

NAND2xp5_ASAP7_75t_L g15709 ( 
.A(n_14841),
.B(n_11527),
.Y(n_15709)
);

HB1xp67_ASAP7_75t_L g15710 ( 
.A(n_15067),
.Y(n_15710)
);

OR2x2_ASAP7_75t_L g15711 ( 
.A(n_15240),
.B(n_11527),
.Y(n_15711)
);

INVx1_ASAP7_75t_L g15712 ( 
.A(n_15320),
.Y(n_15712)
);

INVx1_ASAP7_75t_L g15713 ( 
.A(n_14824),
.Y(n_15713)
);

INVx2_ASAP7_75t_L g15714 ( 
.A(n_15341),
.Y(n_15714)
);

INVxp67_ASAP7_75t_L g15715 ( 
.A(n_14980),
.Y(n_15715)
);

NAND2x1_ASAP7_75t_L g15716 ( 
.A(n_15278),
.B(n_11529),
.Y(n_15716)
);

NOR3xp33_ASAP7_75t_L g15717 ( 
.A(n_15085),
.B(n_15268),
.C(n_15203),
.Y(n_15717)
);

INVx1_ASAP7_75t_L g15718 ( 
.A(n_14837),
.Y(n_15718)
);

INVx1_ASAP7_75t_L g15719 ( 
.A(n_14840),
.Y(n_15719)
);

INVxp67_ASAP7_75t_L g15720 ( 
.A(n_15329),
.Y(n_15720)
);

AND2x2_ASAP7_75t_L g15721 ( 
.A(n_14940),
.B(n_11529),
.Y(n_15721)
);

AND2x4_ASAP7_75t_L g15722 ( 
.A(n_15042),
.B(n_11534),
.Y(n_15722)
);

NAND2xp5_ASAP7_75t_L g15723 ( 
.A(n_14898),
.B(n_11534),
.Y(n_15723)
);

AND2x4_ASAP7_75t_L g15724 ( 
.A(n_15316),
.B(n_11536),
.Y(n_15724)
);

NOR2xp33_ASAP7_75t_L g15725 ( 
.A(n_15345),
.B(n_11536),
.Y(n_15725)
);

AND2x2_ASAP7_75t_L g15726 ( 
.A(n_14977),
.B(n_11548),
.Y(n_15726)
);

BUFx3_ASAP7_75t_L g15727 ( 
.A(n_15277),
.Y(n_15727)
);

NAND2xp5_ASAP7_75t_L g15728 ( 
.A(n_15016),
.B(n_11548),
.Y(n_15728)
);

INVx2_ASAP7_75t_L g15729 ( 
.A(n_14964),
.Y(n_15729)
);

HB1xp67_ASAP7_75t_L g15730 ( 
.A(n_15278),
.Y(n_15730)
);

INVx2_ASAP7_75t_L g15731 ( 
.A(n_14964),
.Y(n_15731)
);

AND2x2_ASAP7_75t_L g15732 ( 
.A(n_14784),
.B(n_11550),
.Y(n_15732)
);

OR2x2_ASAP7_75t_L g15733 ( 
.A(n_14848),
.B(n_11550),
.Y(n_15733)
);

INVx1_ASAP7_75t_L g15734 ( 
.A(n_14854),
.Y(n_15734)
);

OAI22xp33_ASAP7_75t_L g15735 ( 
.A1(n_14950),
.A2(n_14750),
.B1(n_15431),
.B2(n_15122),
.Y(n_15735)
);

OR2x2_ASAP7_75t_L g15736 ( 
.A(n_14853),
.B(n_11564),
.Y(n_15736)
);

INVx1_ASAP7_75t_L g15737 ( 
.A(n_14856),
.Y(n_15737)
);

AND2x4_ASAP7_75t_L g15738 ( 
.A(n_15330),
.B(n_11564),
.Y(n_15738)
);

INVx1_ASAP7_75t_L g15739 ( 
.A(n_14857),
.Y(n_15739)
);

OR2x2_ASAP7_75t_L g15740 ( 
.A(n_14814),
.B(n_11568),
.Y(n_15740)
);

INVx1_ASAP7_75t_L g15741 ( 
.A(n_14860),
.Y(n_15741)
);

INVx2_ASAP7_75t_L g15742 ( 
.A(n_15008),
.Y(n_15742)
);

INVx1_ASAP7_75t_L g15743 ( 
.A(n_14797),
.Y(n_15743)
);

INVx1_ASAP7_75t_L g15744 ( 
.A(n_14843),
.Y(n_15744)
);

INVx2_ASAP7_75t_L g15745 ( 
.A(n_15017),
.Y(n_15745)
);

INVx1_ASAP7_75t_L g15746 ( 
.A(n_14831),
.Y(n_15746)
);

OR2x2_ASAP7_75t_L g15747 ( 
.A(n_15182),
.B(n_14959),
.Y(n_15747)
);

HB1xp67_ASAP7_75t_L g15748 ( 
.A(n_15010),
.Y(n_15748)
);

NAND2xp5_ASAP7_75t_L g15749 ( 
.A(n_15071),
.B(n_11568),
.Y(n_15749)
);

INVx2_ASAP7_75t_L g15750 ( 
.A(n_15019),
.Y(n_15750)
);

INVx1_ASAP7_75t_L g15751 ( 
.A(n_15237),
.Y(n_15751)
);

NOR2x1_ASAP7_75t_L g15752 ( 
.A(n_15086),
.B(n_11569),
.Y(n_15752)
);

INVx1_ASAP7_75t_L g15753 ( 
.A(n_15250),
.Y(n_15753)
);

AND2x2_ASAP7_75t_L g15754 ( 
.A(n_14818),
.B(n_11569),
.Y(n_15754)
);

INVx2_ASAP7_75t_L g15755 ( 
.A(n_15022),
.Y(n_15755)
);

OR2x2_ASAP7_75t_L g15756 ( 
.A(n_14985),
.B(n_11571),
.Y(n_15756)
);

INVx1_ASAP7_75t_L g15757 ( 
.A(n_15255),
.Y(n_15757)
);

NAND2xp5_ASAP7_75t_L g15758 ( 
.A(n_14788),
.B(n_11571),
.Y(n_15758)
);

INVx1_ASAP7_75t_L g15759 ( 
.A(n_15271),
.Y(n_15759)
);

AND2x4_ASAP7_75t_L g15760 ( 
.A(n_15340),
.B(n_11574),
.Y(n_15760)
);

OAI21xp5_ASAP7_75t_SL g15761 ( 
.A1(n_14893),
.A2(n_8862),
.B(n_8183),
.Y(n_15761)
);

INVx2_ASAP7_75t_L g15762 ( 
.A(n_14826),
.Y(n_15762)
);

AND2x2_ASAP7_75t_L g15763 ( 
.A(n_15171),
.B(n_11574),
.Y(n_15763)
);

AND2x2_ASAP7_75t_L g15764 ( 
.A(n_15260),
.B(n_11575),
.Y(n_15764)
);

INVx1_ASAP7_75t_L g15765 ( 
.A(n_15274),
.Y(n_15765)
);

OR2x2_ASAP7_75t_L g15766 ( 
.A(n_14945),
.B(n_11575),
.Y(n_15766)
);

HB1xp67_ASAP7_75t_L g15767 ( 
.A(n_15431),
.Y(n_15767)
);

AND2x2_ASAP7_75t_L g15768 ( 
.A(n_15116),
.B(n_11581),
.Y(n_15768)
);

INVx1_ASAP7_75t_L g15769 ( 
.A(n_15283),
.Y(n_15769)
);

INVx1_ASAP7_75t_L g15770 ( 
.A(n_15285),
.Y(n_15770)
);

AND2x2_ASAP7_75t_L g15771 ( 
.A(n_14792),
.B(n_11581),
.Y(n_15771)
);

INVx2_ASAP7_75t_L g15772 ( 
.A(n_14827),
.Y(n_15772)
);

AND2x2_ASAP7_75t_L g15773 ( 
.A(n_15074),
.B(n_11590),
.Y(n_15773)
);

AND2x2_ASAP7_75t_L g15774 ( 
.A(n_15021),
.B(n_15204),
.Y(n_15774)
);

NAND2xp5_ASAP7_75t_L g15775 ( 
.A(n_15205),
.B(n_11590),
.Y(n_15775)
);

INVx2_ASAP7_75t_L g15776 ( 
.A(n_14832),
.Y(n_15776)
);

AND2x2_ASAP7_75t_L g15777 ( 
.A(n_15159),
.B(n_11592),
.Y(n_15777)
);

INVx1_ASAP7_75t_L g15778 ( 
.A(n_15286),
.Y(n_15778)
);

INVx1_ASAP7_75t_L g15779 ( 
.A(n_15075),
.Y(n_15779)
);

HB1xp67_ASAP7_75t_L g15780 ( 
.A(n_15018),
.Y(n_15780)
);

NOR2x1_ASAP7_75t_SL g15781 ( 
.A(n_15442),
.B(n_11302),
.Y(n_15781)
);

INVx1_ASAP7_75t_L g15782 ( 
.A(n_15357),
.Y(n_15782)
);

INVx1_ASAP7_75t_L g15783 ( 
.A(n_14810),
.Y(n_15783)
);

HB1xp67_ASAP7_75t_L g15784 ( 
.A(n_15304),
.Y(n_15784)
);

HB1xp67_ASAP7_75t_L g15785 ( 
.A(n_15352),
.Y(n_15785)
);

HB1xp67_ASAP7_75t_L g15786 ( 
.A(n_15355),
.Y(n_15786)
);

AND2x4_ASAP7_75t_L g15787 ( 
.A(n_14833),
.B(n_14754),
.Y(n_15787)
);

AND2x2_ASAP7_75t_L g15788 ( 
.A(n_15149),
.B(n_11592),
.Y(n_15788)
);

AND2x2_ASAP7_75t_L g15789 ( 
.A(n_15097),
.B(n_11613),
.Y(n_15789)
);

AND2x2_ASAP7_75t_L g15790 ( 
.A(n_14850),
.B(n_11613),
.Y(n_15790)
);

INVx2_ASAP7_75t_L g15791 ( 
.A(n_14873),
.Y(n_15791)
);

INVx2_ASAP7_75t_L g15792 ( 
.A(n_14873),
.Y(n_15792)
);

AND2x2_ASAP7_75t_L g15793 ( 
.A(n_14866),
.B(n_14867),
.Y(n_15793)
);

HB1xp67_ASAP7_75t_L g15794 ( 
.A(n_15139),
.Y(n_15794)
);

AND2x2_ASAP7_75t_L g15795 ( 
.A(n_14785),
.B(n_11630),
.Y(n_15795)
);

INVx1_ASAP7_75t_L g15796 ( 
.A(n_14933),
.Y(n_15796)
);

INVx2_ASAP7_75t_L g15797 ( 
.A(n_15145),
.Y(n_15797)
);

HB1xp67_ASAP7_75t_L g15798 ( 
.A(n_15146),
.Y(n_15798)
);

OR2x2_ASAP7_75t_L g15799 ( 
.A(n_14978),
.B(n_11630),
.Y(n_15799)
);

INVx2_ASAP7_75t_L g15800 ( 
.A(n_15180),
.Y(n_15800)
);

INVx2_ASAP7_75t_L g15801 ( 
.A(n_15152),
.Y(n_15801)
);

AND2x2_ASAP7_75t_L g15802 ( 
.A(n_15050),
.B(n_11635),
.Y(n_15802)
);

AND2x2_ASAP7_75t_L g15803 ( 
.A(n_15053),
.B(n_11635),
.Y(n_15803)
);

AND2x2_ASAP7_75t_L g15804 ( 
.A(n_15105),
.B(n_11646),
.Y(n_15804)
);

INVx1_ASAP7_75t_L g15805 ( 
.A(n_14844),
.Y(n_15805)
);

AND2x4_ASAP7_75t_L g15806 ( 
.A(n_15107),
.B(n_8624),
.Y(n_15806)
);

INVx1_ASAP7_75t_L g15807 ( 
.A(n_15088),
.Y(n_15807)
);

AOI22xp33_ASAP7_75t_SL g15808 ( 
.A1(n_15136),
.A2(n_8295),
.B1(n_8430),
.B2(n_8142),
.Y(n_15808)
);

NAND2xp5_ASAP7_75t_L g15809 ( 
.A(n_15399),
.B(n_11646),
.Y(n_15809)
);

NAND2xp5_ASAP7_75t_SL g15810 ( 
.A(n_15443),
.B(n_8295),
.Y(n_15810)
);

INVx2_ASAP7_75t_L g15811 ( 
.A(n_14996),
.Y(n_15811)
);

NAND2xp5_ASAP7_75t_L g15812 ( 
.A(n_15100),
.B(n_11652),
.Y(n_15812)
);

INVx1_ASAP7_75t_L g15813 ( 
.A(n_15102),
.Y(n_15813)
);

INVx1_ASAP7_75t_L g15814 ( 
.A(n_15109),
.Y(n_15814)
);

INVx1_ASAP7_75t_L g15815 ( 
.A(n_15132),
.Y(n_15815)
);

INVx3_ASAP7_75t_L g15816 ( 
.A(n_15369),
.Y(n_15816)
);

INVx1_ASAP7_75t_L g15817 ( 
.A(n_15141),
.Y(n_15817)
);

AND2x2_ASAP7_75t_L g15818 ( 
.A(n_15241),
.B(n_11652),
.Y(n_15818)
);

AND2x2_ASAP7_75t_L g15819 ( 
.A(n_15081),
.B(n_11657),
.Y(n_15819)
);

INVxp67_ASAP7_75t_L g15820 ( 
.A(n_14777),
.Y(n_15820)
);

AND2x2_ASAP7_75t_L g15821 ( 
.A(n_15138),
.B(n_11657),
.Y(n_15821)
);

INVx2_ASAP7_75t_L g15822 ( 
.A(n_15073),
.Y(n_15822)
);

NAND2xp5_ASAP7_75t_L g15823 ( 
.A(n_14937),
.B(n_11666),
.Y(n_15823)
);

AND2x2_ASAP7_75t_L g15824 ( 
.A(n_15176),
.B(n_11666),
.Y(n_15824)
);

AND2x2_ASAP7_75t_L g15825 ( 
.A(n_15082),
.B(n_11669),
.Y(n_15825)
);

AND2x2_ASAP7_75t_L g15826 ( 
.A(n_15083),
.B(n_11669),
.Y(n_15826)
);

INVx2_ASAP7_75t_L g15827 ( 
.A(n_15080),
.Y(n_15827)
);

AND2x4_ASAP7_75t_SL g15828 ( 
.A(n_15339),
.B(n_8338),
.Y(n_15828)
);

OR2x2_ASAP7_75t_L g15829 ( 
.A(n_14982),
.B(n_11673),
.Y(n_15829)
);

INVx1_ASAP7_75t_L g15830 ( 
.A(n_15068),
.Y(n_15830)
);

AND2x2_ASAP7_75t_L g15831 ( 
.A(n_15043),
.B(n_15214),
.Y(n_15831)
);

OR2x2_ASAP7_75t_L g15832 ( 
.A(n_14989),
.B(n_11673),
.Y(n_15832)
);

INVx1_ASAP7_75t_L g15833 ( 
.A(n_15328),
.Y(n_15833)
);

AND2x2_ASAP7_75t_L g15834 ( 
.A(n_15057),
.B(n_11683),
.Y(n_15834)
);

AND2x2_ASAP7_75t_L g15835 ( 
.A(n_15063),
.B(n_11683),
.Y(n_15835)
);

NOR2xp33_ASAP7_75t_L g15836 ( 
.A(n_15220),
.B(n_11685),
.Y(n_15836)
);

AND2x2_ASAP7_75t_L g15837 ( 
.A(n_15079),
.B(n_11685),
.Y(n_15837)
);

NOR2xp33_ASAP7_75t_L g15838 ( 
.A(n_15281),
.B(n_11687),
.Y(n_15838)
);

OR2x2_ASAP7_75t_L g15839 ( 
.A(n_14862),
.B(n_11687),
.Y(n_15839)
);

HB1xp67_ASAP7_75t_L g15840 ( 
.A(n_15272),
.Y(n_15840)
);

NAND2xp5_ASAP7_75t_L g15841 ( 
.A(n_15378),
.B(n_11689),
.Y(n_15841)
);

AND2x2_ASAP7_75t_L g15842 ( 
.A(n_15124),
.B(n_11689),
.Y(n_15842)
);

AND2x2_ASAP7_75t_L g15843 ( 
.A(n_15157),
.B(n_11691),
.Y(n_15843)
);

AND2x2_ASAP7_75t_L g15844 ( 
.A(n_15189),
.B(n_11691),
.Y(n_15844)
);

AND2x2_ASAP7_75t_L g15845 ( 
.A(n_15112),
.B(n_11704),
.Y(n_15845)
);

AND2x4_ASAP7_75t_L g15846 ( 
.A(n_14884),
.B(n_8624),
.Y(n_15846)
);

AND2x2_ASAP7_75t_L g15847 ( 
.A(n_15115),
.B(n_11704),
.Y(n_15847)
);

AND2x2_ASAP7_75t_L g15848 ( 
.A(n_15117),
.B(n_11708),
.Y(n_15848)
);

INVx1_ASAP7_75t_L g15849 ( 
.A(n_15362),
.Y(n_15849)
);

INVx1_ASAP7_75t_L g15850 ( 
.A(n_14870),
.Y(n_15850)
);

INVx1_ASAP7_75t_L g15851 ( 
.A(n_14878),
.Y(n_15851)
);

INVx1_ASAP7_75t_L g15852 ( 
.A(n_14887),
.Y(n_15852)
);

INVx1_ASAP7_75t_L g15853 ( 
.A(n_14956),
.Y(n_15853)
);

AND2x2_ASAP7_75t_L g15854 ( 
.A(n_15135),
.B(n_11708),
.Y(n_15854)
);

INVx1_ASAP7_75t_L g15855 ( 
.A(n_14806),
.Y(n_15855)
);

INVx2_ASAP7_75t_L g15856 ( 
.A(n_15027),
.Y(n_15856)
);

OR2x2_ASAP7_75t_L g15857 ( 
.A(n_14931),
.B(n_11726),
.Y(n_15857)
);

AND2x2_ASAP7_75t_L g15858 ( 
.A(n_15137),
.B(n_11726),
.Y(n_15858)
);

OR2x2_ASAP7_75t_L g15859 ( 
.A(n_14938),
.B(n_11728),
.Y(n_15859)
);

NAND2xp5_ASAP7_75t_L g15860 ( 
.A(n_15262),
.B(n_11728),
.Y(n_15860)
);

AND2x2_ASAP7_75t_L g15861 ( 
.A(n_15150),
.B(n_11730),
.Y(n_15861)
);

INVx1_ASAP7_75t_L g15862 ( 
.A(n_14812),
.Y(n_15862)
);

AND2x2_ASAP7_75t_L g15863 ( 
.A(n_15151),
.B(n_11730),
.Y(n_15863)
);

NAND2xp5_ASAP7_75t_L g15864 ( 
.A(n_15263),
.B(n_11731),
.Y(n_15864)
);

OR2x2_ASAP7_75t_L g15865 ( 
.A(n_14999),
.B(n_11731),
.Y(n_15865)
);

INVx1_ASAP7_75t_L g15866 ( 
.A(n_14816),
.Y(n_15866)
);

AND2x2_ASAP7_75t_L g15867 ( 
.A(n_15367),
.B(n_11734),
.Y(n_15867)
);

INVx1_ASAP7_75t_L g15868 ( 
.A(n_14823),
.Y(n_15868)
);

INVx1_ASAP7_75t_L g15869 ( 
.A(n_14861),
.Y(n_15869)
);

HB1xp67_ASAP7_75t_L g15870 ( 
.A(n_15386),
.Y(n_15870)
);

NOR3xp33_ASAP7_75t_L g15871 ( 
.A(n_14969),
.B(n_11305),
.C(n_11303),
.Y(n_15871)
);

NAND2xp5_ASAP7_75t_L g15872 ( 
.A(n_15344),
.B(n_11734),
.Y(n_15872)
);

AND2x2_ASAP7_75t_L g15873 ( 
.A(n_15226),
.B(n_11740),
.Y(n_15873)
);

INVx1_ASAP7_75t_L g15874 ( 
.A(n_14868),
.Y(n_15874)
);

AND2x2_ASAP7_75t_L g15875 ( 
.A(n_15128),
.B(n_11740),
.Y(n_15875)
);

NAND2xp5_ASAP7_75t_L g15876 ( 
.A(n_15409),
.B(n_11748),
.Y(n_15876)
);

AND2x4_ASAP7_75t_SL g15877 ( 
.A(n_15289),
.B(n_8338),
.Y(n_15877)
);

INVx1_ASAP7_75t_L g15878 ( 
.A(n_14872),
.Y(n_15878)
);

INVx1_ASAP7_75t_L g15879 ( 
.A(n_14874),
.Y(n_15879)
);

INVx1_ASAP7_75t_L g15880 ( 
.A(n_15174),
.Y(n_15880)
);

NAND2xp5_ASAP7_75t_L g15881 ( 
.A(n_14855),
.B(n_11748),
.Y(n_15881)
);

NAND2xp5_ASAP7_75t_L g15882 ( 
.A(n_14875),
.B(n_11749),
.Y(n_15882)
);

INVxp67_ASAP7_75t_L g15883 ( 
.A(n_15036),
.Y(n_15883)
);

OR2x2_ASAP7_75t_L g15884 ( 
.A(n_15003),
.B(n_11749),
.Y(n_15884)
);

AND2x2_ASAP7_75t_L g15885 ( 
.A(n_15129),
.B(n_11753),
.Y(n_15885)
);

AND2x2_ASAP7_75t_L g15886 ( 
.A(n_15227),
.B(n_15172),
.Y(n_15886)
);

INVx2_ASAP7_75t_L g15887 ( 
.A(n_15385),
.Y(n_15887)
);

AND2x2_ASAP7_75t_L g15888 ( 
.A(n_14879),
.B(n_11753),
.Y(n_15888)
);

AND2x2_ASAP7_75t_L g15889 ( 
.A(n_15111),
.B(n_11758),
.Y(n_15889)
);

INVx1_ASAP7_75t_L g15890 ( 
.A(n_15199),
.Y(n_15890)
);

AND2x2_ASAP7_75t_L g15891 ( 
.A(n_14798),
.B(n_11758),
.Y(n_15891)
);

INVx2_ASAP7_75t_L g15892 ( 
.A(n_15369),
.Y(n_15892)
);

INVx2_ASAP7_75t_L g15893 ( 
.A(n_15273),
.Y(n_15893)
);

AND2x2_ASAP7_75t_L g15894 ( 
.A(n_14802),
.B(n_11761),
.Y(n_15894)
);

NAND2xp5_ASAP7_75t_L g15895 ( 
.A(n_15258),
.B(n_14886),
.Y(n_15895)
);

NOR2xp33_ASAP7_75t_L g15896 ( 
.A(n_15323),
.B(n_11761),
.Y(n_15896)
);

INVxp67_ASAP7_75t_SL g15897 ( 
.A(n_15346),
.Y(n_15897)
);

INVx1_ASAP7_75t_L g15898 ( 
.A(n_15192),
.Y(n_15898)
);

BUFx2_ASAP7_75t_L g15899 ( 
.A(n_15170),
.Y(n_15899)
);

AND2x4_ASAP7_75t_SL g15900 ( 
.A(n_15110),
.B(n_8338),
.Y(n_15900)
);

INVx1_ASAP7_75t_L g15901 ( 
.A(n_15251),
.Y(n_15901)
);

INVx1_ASAP7_75t_L g15902 ( 
.A(n_15292),
.Y(n_15902)
);

INVx2_ASAP7_75t_L g15903 ( 
.A(n_15211),
.Y(n_15903)
);

NOR3xp33_ASAP7_75t_L g15904 ( 
.A(n_14787),
.B(n_11325),
.C(n_11305),
.Y(n_15904)
);

INVx1_ASAP7_75t_L g15905 ( 
.A(n_15013),
.Y(n_15905)
);

NAND3xp33_ASAP7_75t_L g15906 ( 
.A(n_14759),
.B(n_11325),
.C(n_11682),
.Y(n_15906)
);

AND2x2_ASAP7_75t_L g15907 ( 
.A(n_15181),
.B(n_11763),
.Y(n_15907)
);

INVx2_ASAP7_75t_L g15908 ( 
.A(n_15186),
.Y(n_15908)
);

OR2x2_ASAP7_75t_L g15909 ( 
.A(n_15161),
.B(n_11763),
.Y(n_15909)
);

AND2x2_ASAP7_75t_L g15910 ( 
.A(n_15156),
.B(n_11764),
.Y(n_15910)
);

OR2x2_ASAP7_75t_L g15911 ( 
.A(n_14795),
.B(n_11764),
.Y(n_15911)
);

AND2x2_ASAP7_75t_L g15912 ( 
.A(n_15261),
.B(n_11775),
.Y(n_15912)
);

INVx2_ASAP7_75t_L g15913 ( 
.A(n_15423),
.Y(n_15913)
);

INVx1_ASAP7_75t_L g15914 ( 
.A(n_15298),
.Y(n_15914)
);

INVx2_ASAP7_75t_L g15915 ( 
.A(n_14834),
.Y(n_15915)
);

AND2x2_ASAP7_75t_L g15916 ( 
.A(n_15349),
.B(n_11775),
.Y(n_15916)
);

INVx1_ASAP7_75t_L g15917 ( 
.A(n_14782),
.Y(n_15917)
);

NAND2xp5_ASAP7_75t_SL g15918 ( 
.A(n_15443),
.B(n_8430),
.Y(n_15918)
);

NOR2xp33_ASAP7_75t_L g15919 ( 
.A(n_15397),
.B(n_11791),
.Y(n_15919)
);

OAI21xp33_ASAP7_75t_L g15920 ( 
.A1(n_14794),
.A2(n_10773),
.B(n_10772),
.Y(n_15920)
);

INVx1_ASAP7_75t_L g15921 ( 
.A(n_15011),
.Y(n_15921)
);

NAND2xp5_ASAP7_75t_L g15922 ( 
.A(n_15148),
.B(n_11791),
.Y(n_15922)
);

AND2x2_ASAP7_75t_L g15923 ( 
.A(n_15353),
.B(n_11793),
.Y(n_15923)
);

INVx2_ASAP7_75t_L g15924 ( 
.A(n_14836),
.Y(n_15924)
);

AND2x2_ASAP7_75t_L g15925 ( 
.A(n_15360),
.B(n_11793),
.Y(n_15925)
);

AND2x2_ASAP7_75t_L g15926 ( 
.A(n_15368),
.B(n_11800),
.Y(n_15926)
);

AND2x2_ASAP7_75t_L g15927 ( 
.A(n_15373),
.B(n_11800),
.Y(n_15927)
);

INVxp67_ASAP7_75t_SL g15928 ( 
.A(n_15015),
.Y(n_15928)
);

INVx4_ASAP7_75t_L g15929 ( 
.A(n_15347),
.Y(n_15929)
);

INVx1_ASAP7_75t_L g15930 ( 
.A(n_15147),
.Y(n_15930)
);

INVx2_ASAP7_75t_L g15931 ( 
.A(n_15188),
.Y(n_15931)
);

AND2x2_ASAP7_75t_L g15932 ( 
.A(n_15377),
.B(n_11808),
.Y(n_15932)
);

INVx2_ASAP7_75t_L g15933 ( 
.A(n_15207),
.Y(n_15933)
);

NAND2xp5_ASAP7_75t_L g15934 ( 
.A(n_15206),
.B(n_11808),
.Y(n_15934)
);

NAND2xp5_ASAP7_75t_L g15935 ( 
.A(n_15222),
.B(n_11813),
.Y(n_15935)
);

AND2x4_ASAP7_75t_L g15936 ( 
.A(n_14902),
.B(n_14906),
.Y(n_15936)
);

NAND2x1_ASAP7_75t_L g15937 ( 
.A(n_15366),
.B(n_11813),
.Y(n_15937)
);

HB1xp67_ASAP7_75t_L g15938 ( 
.A(n_15379),
.Y(n_15938)
);

OR2x6_ASAP7_75t_L g15939 ( 
.A(n_14894),
.B(n_7792),
.Y(n_15939)
);

BUFx3_ASAP7_75t_L g15940 ( 
.A(n_14913),
.Y(n_15940)
);

NAND2x1p5_ASAP7_75t_L g15941 ( 
.A(n_15133),
.B(n_7792),
.Y(n_15941)
);

INVx1_ASAP7_75t_L g15942 ( 
.A(n_14967),
.Y(n_15942)
);

INVx1_ASAP7_75t_L g15943 ( 
.A(n_15143),
.Y(n_15943)
);

INVx1_ASAP7_75t_L g15944 ( 
.A(n_14772),
.Y(n_15944)
);

NAND3xp33_ASAP7_75t_L g15945 ( 
.A(n_15284),
.B(n_11743),
.C(n_11682),
.Y(n_15945)
);

INVx2_ASAP7_75t_L g15946 ( 
.A(n_14939),
.Y(n_15946)
);

OR2x2_ASAP7_75t_L g15947 ( 
.A(n_15388),
.B(n_11820),
.Y(n_15947)
);

AND2x2_ASAP7_75t_L g15948 ( 
.A(n_15389),
.B(n_11820),
.Y(n_15948)
);

OR2x2_ASAP7_75t_L g15949 ( 
.A(n_15391),
.B(n_11822),
.Y(n_15949)
);

INVx1_ASAP7_75t_L g15950 ( 
.A(n_15396),
.Y(n_15950)
);

NAND2xp5_ASAP7_75t_L g15951 ( 
.A(n_15252),
.B(n_11822),
.Y(n_15951)
);

INVx1_ASAP7_75t_L g15952 ( 
.A(n_15398),
.Y(n_15952)
);

INVx1_ASAP7_75t_L g15953 ( 
.A(n_15403),
.Y(n_15953)
);

INVx1_ASAP7_75t_L g15954 ( 
.A(n_15387),
.Y(n_15954)
);

AND2x2_ASAP7_75t_L g15955 ( 
.A(n_15193),
.B(n_11837),
.Y(n_15955)
);

AND2x4_ASAP7_75t_L g15956 ( 
.A(n_14919),
.B(n_8624),
.Y(n_15956)
);

AND2x2_ASAP7_75t_L g15957 ( 
.A(n_15089),
.B(n_11837),
.Y(n_15957)
);

INVx1_ASAP7_75t_L g15958 ( 
.A(n_15066),
.Y(n_15958)
);

AOI211xp5_ASAP7_75t_L g15959 ( 
.A1(n_15267),
.A2(n_11046),
.B(n_11067),
.C(n_10755),
.Y(n_15959)
);

INVx1_ASAP7_75t_L g15960 ( 
.A(n_14949),
.Y(n_15960)
);

INVx2_ASAP7_75t_L g15961 ( 
.A(n_14947),
.Y(n_15961)
);

NOR2xp33_ASAP7_75t_L g15962 ( 
.A(n_14901),
.B(n_11841),
.Y(n_15962)
);

OR2x2_ASAP7_75t_L g15963 ( 
.A(n_14953),
.B(n_11841),
.Y(n_15963)
);

NOR2x1_ASAP7_75t_L g15964 ( 
.A(n_15144),
.B(n_11845),
.Y(n_15964)
);

INVx2_ASAP7_75t_L g15965 ( 
.A(n_14954),
.Y(n_15965)
);

AND2x2_ASAP7_75t_L g15966 ( 
.A(n_15198),
.B(n_15231),
.Y(n_15966)
);

NAND2xp5_ASAP7_75t_L g15967 ( 
.A(n_14971),
.B(n_11845),
.Y(n_15967)
);

NOR2xp67_ASAP7_75t_L g15968 ( 
.A(n_15453),
.B(n_11848),
.Y(n_15968)
);

AND2x2_ASAP7_75t_L g15969 ( 
.A(n_15235),
.B(n_15253),
.Y(n_15969)
);

AND2x2_ASAP7_75t_L g15970 ( 
.A(n_15256),
.B(n_11848),
.Y(n_15970)
);

AND2x2_ASAP7_75t_L g15971 ( 
.A(n_15294),
.B(n_11850),
.Y(n_15971)
);

INVx2_ASAP7_75t_L g15972 ( 
.A(n_15155),
.Y(n_15972)
);

INVx1_ASAP7_75t_L g15973 ( 
.A(n_15370),
.Y(n_15973)
);

INVxp67_ASAP7_75t_SL g15974 ( 
.A(n_15014),
.Y(n_15974)
);

INVx2_ASAP7_75t_L g15975 ( 
.A(n_15160),
.Y(n_15975)
);

AND2x2_ASAP7_75t_L g15976 ( 
.A(n_15394),
.B(n_11850),
.Y(n_15976)
);

INVx1_ASAP7_75t_L g15977 ( 
.A(n_14932),
.Y(n_15977)
);

AND2x4_ASAP7_75t_L g15978 ( 
.A(n_15028),
.B(n_8624),
.Y(n_15978)
);

INVx1_ASAP7_75t_L g15979 ( 
.A(n_15178),
.Y(n_15979)
);

OR2x2_ASAP7_75t_L g15980 ( 
.A(n_15184),
.B(n_15032),
.Y(n_15980)
);

AND2x2_ASAP7_75t_L g15981 ( 
.A(n_15217),
.B(n_11866),
.Y(n_15981)
);

AND2x2_ASAP7_75t_L g15982 ( 
.A(n_15245),
.B(n_11866),
.Y(n_15982)
);

INVx1_ASAP7_75t_L g15983 ( 
.A(n_15179),
.Y(n_15983)
);

AND2x2_ASAP7_75t_L g15984 ( 
.A(n_15215),
.B(n_11869),
.Y(n_15984)
);

INVx1_ASAP7_75t_L g15985 ( 
.A(n_14864),
.Y(n_15985)
);

INVx1_ASAP7_75t_L g15986 ( 
.A(n_14869),
.Y(n_15986)
);

INVx1_ASAP7_75t_L g15987 ( 
.A(n_14881),
.Y(n_15987)
);

AND2x4_ASAP7_75t_SL g15988 ( 
.A(n_15134),
.B(n_8338),
.Y(n_15988)
);

AND2x2_ASAP7_75t_L g15989 ( 
.A(n_15200),
.B(n_11869),
.Y(n_15989)
);

INVx2_ASAP7_75t_L g15990 ( 
.A(n_15033),
.Y(n_15990)
);

NAND2xp5_ASAP7_75t_L g15991 ( 
.A(n_15037),
.B(n_11871),
.Y(n_15991)
);

AND2x2_ASAP7_75t_L g15992 ( 
.A(n_15202),
.B(n_11871),
.Y(n_15992)
);

INVx2_ASAP7_75t_L g15993 ( 
.A(n_15040),
.Y(n_15993)
);

INVx1_ASAP7_75t_L g15994 ( 
.A(n_14882),
.Y(n_15994)
);

INVx1_ASAP7_75t_L g15995 ( 
.A(n_14883),
.Y(n_15995)
);

AND2x2_ASAP7_75t_L g15996 ( 
.A(n_15306),
.B(n_11882),
.Y(n_15996)
);

NAND2xp5_ASAP7_75t_L g15997 ( 
.A(n_15046),
.B(n_11882),
.Y(n_15997)
);

OR2x2_ASAP7_75t_L g15998 ( 
.A(n_15051),
.B(n_11884),
.Y(n_15998)
);

INVx1_ASAP7_75t_L g15999 ( 
.A(n_14909),
.Y(n_15999)
);

INVx1_ASAP7_75t_L g16000 ( 
.A(n_15390),
.Y(n_16000)
);

INVx1_ASAP7_75t_L g16001 ( 
.A(n_15395),
.Y(n_16001)
);

AND2x2_ASAP7_75t_L g16002 ( 
.A(n_15310),
.B(n_15219),
.Y(n_16002)
);

OR2x2_ASAP7_75t_L g16003 ( 
.A(n_15054),
.B(n_11884),
.Y(n_16003)
);

NAND2xp5_ASAP7_75t_L g16004 ( 
.A(n_15069),
.B(n_11890),
.Y(n_16004)
);

AND2x2_ASAP7_75t_L g16005 ( 
.A(n_15225),
.B(n_15275),
.Y(n_16005)
);

INVxp67_ASAP7_75t_SL g16006 ( 
.A(n_15113),
.Y(n_16006)
);

INVx1_ASAP7_75t_L g16007 ( 
.A(n_15402),
.Y(n_16007)
);

AND2x6_ASAP7_75t_SL g16008 ( 
.A(n_15106),
.B(n_8818),
.Y(n_16008)
);

NOR2x1_ASAP7_75t_L g16009 ( 
.A(n_15158),
.B(n_11890),
.Y(n_16009)
);

AND2x2_ASAP7_75t_L g16010 ( 
.A(n_15279),
.B(n_11899),
.Y(n_16010)
);

NAND2xp5_ASAP7_75t_L g16011 ( 
.A(n_15266),
.B(n_11899),
.Y(n_16011)
);

AND2x2_ASAP7_75t_L g16012 ( 
.A(n_15280),
.B(n_11900),
.Y(n_16012)
);

INVx2_ASAP7_75t_SL g16013 ( 
.A(n_15364),
.Y(n_16013)
);

AND2x2_ASAP7_75t_L g16014 ( 
.A(n_15291),
.B(n_11900),
.Y(n_16014)
);

OR2x2_ASAP7_75t_L g16015 ( 
.A(n_14952),
.B(n_11901),
.Y(n_16015)
);

NAND2xp5_ASAP7_75t_SL g16016 ( 
.A(n_15383),
.B(n_8430),
.Y(n_16016)
);

INVx2_ASAP7_75t_L g16017 ( 
.A(n_15104),
.Y(n_16017)
);

OR2x2_ASAP7_75t_L g16018 ( 
.A(n_14970),
.B(n_11901),
.Y(n_16018)
);

NAND3xp33_ASAP7_75t_L g16019 ( 
.A(n_15432),
.B(n_11743),
.C(n_11682),
.Y(n_16019)
);

INVx1_ASAP7_75t_SL g16020 ( 
.A(n_15429),
.Y(n_16020)
);

AND2x2_ASAP7_75t_L g16021 ( 
.A(n_15379),
.B(n_11902),
.Y(n_16021)
);

NAND2xp5_ASAP7_75t_L g16022 ( 
.A(n_15108),
.B(n_11902),
.Y(n_16022)
);

INVxp67_ASAP7_75t_L g16023 ( 
.A(n_15430),
.Y(n_16023)
);

INVx1_ASAP7_75t_L g16024 ( 
.A(n_15410),
.Y(n_16024)
);

AND2x2_ASAP7_75t_L g16025 ( 
.A(n_15190),
.B(n_11904),
.Y(n_16025)
);

AND2x2_ASAP7_75t_L g16026 ( 
.A(n_15437),
.B(n_11904),
.Y(n_16026)
);

NAND2xp5_ASAP7_75t_SL g16027 ( 
.A(n_15361),
.B(n_8430),
.Y(n_16027)
);

INVx1_ASAP7_75t_L g16028 ( 
.A(n_15315),
.Y(n_16028)
);

AND2x2_ASAP7_75t_L g16029 ( 
.A(n_15413),
.B(n_11906),
.Y(n_16029)
);

OR2x2_ASAP7_75t_L g16030 ( 
.A(n_14811),
.B(n_11906),
.Y(n_16030)
);

INVx1_ASAP7_75t_L g16031 ( 
.A(n_14910),
.Y(n_16031)
);

NAND2xp5_ASAP7_75t_L g16032 ( 
.A(n_15422),
.B(n_11908),
.Y(n_16032)
);

INVx2_ASAP7_75t_L g16033 ( 
.A(n_15338),
.Y(n_16033)
);

BUFx3_ASAP7_75t_L g16034 ( 
.A(n_15416),
.Y(n_16034)
);

OR2x2_ASAP7_75t_L g16035 ( 
.A(n_14842),
.B(n_11908),
.Y(n_16035)
);

NAND2x1p5_ASAP7_75t_L g16036 ( 
.A(n_15444),
.B(n_14972),
.Y(n_16036)
);

INVx2_ASAP7_75t_L g16037 ( 
.A(n_15356),
.Y(n_16037)
);

OR2x2_ASAP7_75t_L g16038 ( 
.A(n_15163),
.B(n_15248),
.Y(n_16038)
);

AND2x2_ASAP7_75t_L g16039 ( 
.A(n_15418),
.B(n_11910),
.Y(n_16039)
);

AND2x2_ASAP7_75t_L g16040 ( 
.A(n_15438),
.B(n_15439),
.Y(n_16040)
);

OR2x2_ASAP7_75t_L g16041 ( 
.A(n_14991),
.B(n_11910),
.Y(n_16041)
);

INVxp67_ASAP7_75t_SL g16042 ( 
.A(n_15308),
.Y(n_16042)
);

AND2x2_ASAP7_75t_L g16043 ( 
.A(n_15433),
.B(n_11926),
.Y(n_16043)
);

AND2x2_ASAP7_75t_L g16044 ( 
.A(n_15427),
.B(n_11926),
.Y(n_16044)
);

AND2x2_ASAP7_75t_L g16045 ( 
.A(n_15424),
.B(n_8180),
.Y(n_16045)
);

INVx1_ASAP7_75t_L g16046 ( 
.A(n_14911),
.Y(n_16046)
);

OR2x2_ASAP7_75t_L g16047 ( 
.A(n_15282),
.B(n_8973),
.Y(n_16047)
);

AND2x2_ASAP7_75t_L g16048 ( 
.A(n_15425),
.B(n_8180),
.Y(n_16048)
);

INVx1_ASAP7_75t_L g16049 ( 
.A(n_14912),
.Y(n_16049)
);

HB1xp67_ASAP7_75t_L g16050 ( 
.A(n_15321),
.Y(n_16050)
);

AND2x2_ASAP7_75t_L g16051 ( 
.A(n_15428),
.B(n_8180),
.Y(n_16051)
);

AND2x4_ASAP7_75t_SL g16052 ( 
.A(n_15407),
.B(n_8338),
.Y(n_16052)
);

AND2x2_ASAP7_75t_L g16053 ( 
.A(n_14973),
.B(n_8180),
.Y(n_16053)
);

AND2x4_ASAP7_75t_L g16054 ( 
.A(n_14974),
.B(n_8624),
.Y(n_16054)
);

AND2x2_ASAP7_75t_L g16055 ( 
.A(n_14975),
.B(n_14983),
.Y(n_16055)
);

AND2x4_ASAP7_75t_L g16056 ( 
.A(n_15419),
.B(n_11720),
.Y(n_16056)
);

HB1xp67_ASAP7_75t_L g16057 ( 
.A(n_15325),
.Y(n_16057)
);

NOR2xp33_ASAP7_75t_L g16058 ( 
.A(n_15454),
.B(n_8430),
.Y(n_16058)
);

OR2x2_ASAP7_75t_L g16059 ( 
.A(n_15269),
.B(n_8973),
.Y(n_16059)
);

INVx1_ASAP7_75t_L g16060 ( 
.A(n_14916),
.Y(n_16060)
);

INVx1_ASAP7_75t_L g16061 ( 
.A(n_14924),
.Y(n_16061)
);

OR2x2_ASAP7_75t_L g16062 ( 
.A(n_14986),
.B(n_14988),
.Y(n_16062)
);

AND2x2_ASAP7_75t_L g16063 ( 
.A(n_14995),
.B(n_14998),
.Y(n_16063)
);

AOI22xp33_ASAP7_75t_L g16064 ( 
.A1(n_15307),
.A2(n_8096),
.B1(n_8468),
.B2(n_8430),
.Y(n_16064)
);

NAND2xp67_ASAP7_75t_L g16065 ( 
.A(n_15441),
.B(n_10772),
.Y(n_16065)
);

AND2x2_ASAP7_75t_L g16066 ( 
.A(n_15001),
.B(n_8180),
.Y(n_16066)
);

NOR2xp33_ASAP7_75t_L g16067 ( 
.A(n_15412),
.B(n_15421),
.Y(n_16067)
);

AND2x4_ASAP7_75t_L g16068 ( 
.A(n_15004),
.B(n_8686),
.Y(n_16068)
);

NOR2xp33_ASAP7_75t_L g16069 ( 
.A(n_15435),
.B(n_8468),
.Y(n_16069)
);

INVx1_ASAP7_75t_L g16070 ( 
.A(n_14929),
.Y(n_16070)
);

INVx1_ASAP7_75t_L g16071 ( 
.A(n_15309),
.Y(n_16071)
);

OR2x2_ASAP7_75t_L g16072 ( 
.A(n_15031),
.B(n_8989),
.Y(n_16072)
);

INVx1_ASAP7_75t_L g16073 ( 
.A(n_15405),
.Y(n_16073)
);

INVx2_ASAP7_75t_L g16074 ( 
.A(n_15382),
.Y(n_16074)
);

INVx1_ASAP7_75t_L g16075 ( 
.A(n_15449),
.Y(n_16075)
);

INVx2_ASAP7_75t_L g16076 ( 
.A(n_15384),
.Y(n_16076)
);

INVx1_ASAP7_75t_L g16077 ( 
.A(n_15044),
.Y(n_16077)
);

INVx2_ASAP7_75t_L g16078 ( 
.A(n_15436),
.Y(n_16078)
);

NAND2xp5_ASAP7_75t_L g16079 ( 
.A(n_15061),
.B(n_10334),
.Y(n_16079)
);

OR2x2_ASAP7_75t_L g16080 ( 
.A(n_15064),
.B(n_8989),
.Y(n_16080)
);

OR2x2_ASAP7_75t_L g16081 ( 
.A(n_15065),
.B(n_8999),
.Y(n_16081)
);

INVx3_ASAP7_75t_L g16082 ( 
.A(n_15451),
.Y(n_16082)
);

AND2x2_ASAP7_75t_L g16083 ( 
.A(n_15420),
.B(n_8180),
.Y(n_16083)
);

AND2x4_ASAP7_75t_L g16084 ( 
.A(n_15447),
.B(n_11720),
.Y(n_16084)
);

INVx2_ASAP7_75t_L g16085 ( 
.A(n_15411),
.Y(n_16085)
);

INVx2_ASAP7_75t_L g16086 ( 
.A(n_15381),
.Y(n_16086)
);

INVx1_ASAP7_75t_L g16087 ( 
.A(n_15440),
.Y(n_16087)
);

AND2x2_ASAP7_75t_L g16088 ( 
.A(n_15359),
.B(n_8180),
.Y(n_16088)
);

AND2x2_ASAP7_75t_L g16089 ( 
.A(n_15446),
.B(n_8219),
.Y(n_16089)
);

BUFx2_ASAP7_75t_L g16090 ( 
.A(n_15307),
.Y(n_16090)
);

HB1xp67_ASAP7_75t_L g16091 ( 
.A(n_15414),
.Y(n_16091)
);

INVx2_ASAP7_75t_L g16092 ( 
.A(n_15417),
.Y(n_16092)
);

INVx1_ASAP7_75t_L g16093 ( 
.A(n_15445),
.Y(n_16093)
);

INVx1_ASAP7_75t_L g16094 ( 
.A(n_15455),
.Y(n_16094)
);

INVx1_ASAP7_75t_L g16095 ( 
.A(n_15070),
.Y(n_16095)
);

INVx2_ASAP7_75t_L g16096 ( 
.A(n_16090),
.Y(n_16096)
);

AND2x4_ASAP7_75t_L g16097 ( 
.A(n_16090),
.B(n_15452),
.Y(n_16097)
);

AND2x2_ASAP7_75t_L g16098 ( 
.A(n_15469),
.B(n_15348),
.Y(n_16098)
);

INVx1_ASAP7_75t_L g16099 ( 
.A(n_15545),
.Y(n_16099)
);

INVx1_ASAP7_75t_L g16100 ( 
.A(n_15545),
.Y(n_16100)
);

OR2x2_ASAP7_75t_L g16101 ( 
.A(n_15642),
.B(n_15371),
.Y(n_16101)
);

INVx1_ASAP7_75t_L g16102 ( 
.A(n_15780),
.Y(n_16102)
);

OR2x2_ASAP7_75t_L g16103 ( 
.A(n_15484),
.B(n_15529),
.Y(n_16103)
);

AND2x2_ASAP7_75t_L g16104 ( 
.A(n_15488),
.B(n_15072),
.Y(n_16104)
);

INVx1_ASAP7_75t_L g16105 ( 
.A(n_15899),
.Y(n_16105)
);

INVx1_ASAP7_75t_L g16106 ( 
.A(n_15899),
.Y(n_16106)
);

AND2x2_ASAP7_75t_L g16107 ( 
.A(n_15497),
.B(n_15077),
.Y(n_16107)
);

NAND2xp5_ASAP7_75t_L g16108 ( 
.A(n_15544),
.B(n_15078),
.Y(n_16108)
);

INVx2_ASAP7_75t_L g16109 ( 
.A(n_15504),
.Y(n_16109)
);

NAND2xp5_ASAP7_75t_L g16110 ( 
.A(n_15667),
.B(n_15087),
.Y(n_16110)
);

AND2x2_ASAP7_75t_L g16111 ( 
.A(n_15626),
.B(n_15090),
.Y(n_16111)
);

INVx1_ASAP7_75t_SL g16112 ( 
.A(n_15576),
.Y(n_16112)
);

INVx3_ASAP7_75t_L g16113 ( 
.A(n_15929),
.Y(n_16113)
);

INVx1_ASAP7_75t_L g16114 ( 
.A(n_15481),
.Y(n_16114)
);

INVx1_ASAP7_75t_L g16115 ( 
.A(n_15960),
.Y(n_16115)
);

NAND2xp5_ASAP7_75t_L g16116 ( 
.A(n_15639),
.B(n_15091),
.Y(n_16116)
);

AND2x2_ASAP7_75t_L g16117 ( 
.A(n_15831),
.B(n_15774),
.Y(n_16117)
);

NAND2xp5_ASAP7_75t_L g16118 ( 
.A(n_15645),
.B(n_15646),
.Y(n_16118)
);

OR2x2_ASAP7_75t_L g16119 ( 
.A(n_15514),
.B(n_15354),
.Y(n_16119)
);

NAND2xp5_ASAP7_75t_L g16120 ( 
.A(n_15681),
.B(n_15092),
.Y(n_16120)
);

NAND2xp5_ASAP7_75t_L g16121 ( 
.A(n_15710),
.B(n_15094),
.Y(n_16121)
);

AND2x2_ASAP7_75t_L g16122 ( 
.A(n_15686),
.B(n_15096),
.Y(n_16122)
);

AND2x2_ASAP7_75t_L g16123 ( 
.A(n_15886),
.B(n_15098),
.Y(n_16123)
);

INVx1_ASAP7_75t_L g16124 ( 
.A(n_15744),
.Y(n_16124)
);

NAND2xp5_ASAP7_75t_L g16125 ( 
.A(n_15685),
.B(n_15691),
.Y(n_16125)
);

AND2x2_ASAP7_75t_L g16126 ( 
.A(n_15969),
.B(n_15623),
.Y(n_16126)
);

AOI22xp33_ASAP7_75t_L g16127 ( 
.A1(n_15641),
.A2(n_15242),
.B1(n_15195),
.B2(n_15372),
.Y(n_16127)
);

INVx1_ASAP7_75t_L g16128 ( 
.A(n_15746),
.Y(n_16128)
);

INVx1_ASAP7_75t_L g16129 ( 
.A(n_15668),
.Y(n_16129)
);

NAND2x1p5_ASAP7_75t_L g16130 ( 
.A(n_15546),
.B(n_15168),
.Y(n_16130)
);

INVx1_ASAP7_75t_SL g16131 ( 
.A(n_15461),
.Y(n_16131)
);

INVx2_ASAP7_75t_L g16132 ( 
.A(n_15569),
.Y(n_16132)
);

AND2x2_ASAP7_75t_L g16133 ( 
.A(n_15550),
.B(n_15101),
.Y(n_16133)
);

INVx4_ASAP7_75t_L g16134 ( 
.A(n_15598),
.Y(n_16134)
);

INVx1_ASAP7_75t_L g16135 ( 
.A(n_15677),
.Y(n_16135)
);

AND2x2_ASAP7_75t_L g16136 ( 
.A(n_15793),
.B(n_15119),
.Y(n_16136)
);

INVx1_ASAP7_75t_L g16137 ( 
.A(n_15678),
.Y(n_16137)
);

INVx2_ASAP7_75t_L g16138 ( 
.A(n_15781),
.Y(n_16138)
);

INVx1_ASAP7_75t_L g16139 ( 
.A(n_15695),
.Y(n_16139)
);

INVx2_ASAP7_75t_L g16140 ( 
.A(n_15716),
.Y(n_16140)
);

BUFx12f_ASAP7_75t_L g16141 ( 
.A(n_15537),
.Y(n_16141)
);

OR2x2_ASAP7_75t_L g16142 ( 
.A(n_15565),
.B(n_15363),
.Y(n_16142)
);

NAND2xp5_ASAP7_75t_L g16143 ( 
.A(n_15715),
.B(n_15120),
.Y(n_16143)
);

NAND2xp5_ASAP7_75t_L g16144 ( 
.A(n_15640),
.B(n_15123),
.Y(n_16144)
);

INVx3_ASAP7_75t_L g16145 ( 
.A(n_15524),
.Y(n_16145)
);

OR2x2_ASAP7_75t_L g16146 ( 
.A(n_15489),
.B(n_15374),
.Y(n_16146)
);

NAND2xp5_ASAP7_75t_L g16147 ( 
.A(n_15543),
.B(n_15125),
.Y(n_16147)
);

BUFx3_ASAP7_75t_L g16148 ( 
.A(n_15602),
.Y(n_16148)
);

AND2x2_ASAP7_75t_L g16149 ( 
.A(n_15966),
.B(n_15466),
.Y(n_16149)
);

INVx2_ASAP7_75t_L g16150 ( 
.A(n_15498),
.Y(n_16150)
);

OR2x2_ASAP7_75t_L g16151 ( 
.A(n_15624),
.B(n_15153),
.Y(n_16151)
);

AND2x2_ASAP7_75t_L g16152 ( 
.A(n_15893),
.B(n_15167),
.Y(n_16152)
);

INVx1_ASAP7_75t_L g16153 ( 
.A(n_15613),
.Y(n_16153)
);

NAND2xp5_ASAP7_75t_SL g16154 ( 
.A(n_15735),
.B(n_15426),
.Y(n_16154)
);

AND2x2_ASAP7_75t_L g16155 ( 
.A(n_15575),
.B(n_15173),
.Y(n_16155)
);

NAND2xp5_ASAP7_75t_L g16156 ( 
.A(n_15820),
.B(n_16042),
.Y(n_16156)
);

OR2x2_ASAP7_75t_L g16157 ( 
.A(n_15462),
.B(n_15183),
.Y(n_16157)
);

NAND2xp5_ASAP7_75t_L g16158 ( 
.A(n_15883),
.B(n_15393),
.Y(n_16158)
);

INVx1_ASAP7_75t_L g16159 ( 
.A(n_15620),
.Y(n_16159)
);

AND2x2_ASAP7_75t_L g16160 ( 
.A(n_15593),
.B(n_15334),
.Y(n_16160)
);

INVx2_ASAP7_75t_L g16161 ( 
.A(n_15456),
.Y(n_16161)
);

INVx1_ASAP7_75t_SL g16162 ( 
.A(n_15549),
.Y(n_16162)
);

INVx1_ASAP7_75t_L g16163 ( 
.A(n_15509),
.Y(n_16163)
);

AND2x4_ASAP7_75t_L g16164 ( 
.A(n_15510),
.B(n_15194),
.Y(n_16164)
);

INVx2_ASAP7_75t_L g16165 ( 
.A(n_15485),
.Y(n_16165)
);

INVx2_ASAP7_75t_L g16166 ( 
.A(n_15937),
.Y(n_16166)
);

AND2x2_ASAP7_75t_L g16167 ( 
.A(n_15599),
.B(n_15335),
.Y(n_16167)
);

AND2x2_ASAP7_75t_L g16168 ( 
.A(n_15650),
.B(n_15653),
.Y(n_16168)
);

OR2x2_ASAP7_75t_L g16169 ( 
.A(n_15491),
.B(n_15197),
.Y(n_16169)
);

HB1xp67_ASAP7_75t_L g16170 ( 
.A(n_15605),
.Y(n_16170)
);

AND2x2_ASAP7_75t_L g16171 ( 
.A(n_15661),
.B(n_15337),
.Y(n_16171)
);

AND2x2_ASAP7_75t_L g16172 ( 
.A(n_15574),
.B(n_15555),
.Y(n_16172)
);

INVx1_ASAP7_75t_L g16173 ( 
.A(n_15870),
.Y(n_16173)
);

NAND2xp5_ASAP7_75t_L g16174 ( 
.A(n_15840),
.B(n_15401),
.Y(n_16174)
);

AND2x2_ASAP7_75t_L g16175 ( 
.A(n_15487),
.B(n_15404),
.Y(n_16175)
);

INVx1_ASAP7_75t_L g16176 ( 
.A(n_15458),
.Y(n_16176)
);

INVx3_ASAP7_75t_L g16177 ( 
.A(n_15727),
.Y(n_16177)
);

INVx2_ASAP7_75t_L g16178 ( 
.A(n_15587),
.Y(n_16178)
);

AND2x2_ASAP7_75t_L g16179 ( 
.A(n_16005),
.B(n_15448),
.Y(n_16179)
);

OR2x2_ASAP7_75t_L g16180 ( 
.A(n_15649),
.B(n_15201),
.Y(n_16180)
);

AND2x2_ASAP7_75t_L g16181 ( 
.A(n_15811),
.B(n_15350),
.Y(n_16181)
);

INVx2_ASAP7_75t_L g16182 ( 
.A(n_15800),
.Y(n_16182)
);

INVx2_ASAP7_75t_L g16183 ( 
.A(n_16036),
.Y(n_16183)
);

AND2x2_ASAP7_75t_L g16184 ( 
.A(n_15492),
.B(n_15791),
.Y(n_16184)
);

INVx1_ASAP7_75t_L g16185 ( 
.A(n_15459),
.Y(n_16185)
);

AND2x2_ASAP7_75t_L g16186 ( 
.A(n_15792),
.B(n_15351),
.Y(n_16186)
);

NAND2xp5_ASAP7_75t_L g16187 ( 
.A(n_15659),
.B(n_15210),
.Y(n_16187)
);

NAND2xp5_ASAP7_75t_L g16188 ( 
.A(n_15666),
.B(n_15213),
.Y(n_16188)
);

AND2x2_ASAP7_75t_L g16189 ( 
.A(n_15887),
.B(n_15571),
.Y(n_16189)
);

AND2x2_ASAP7_75t_L g16190 ( 
.A(n_15547),
.B(n_15223),
.Y(n_16190)
);

NAND2xp5_ASAP7_75t_L g16191 ( 
.A(n_15669),
.B(n_15230),
.Y(n_16191)
);

INVx2_ASAP7_75t_SL g16192 ( 
.A(n_15592),
.Y(n_16192)
);

INVx1_ASAP7_75t_L g16193 ( 
.A(n_15464),
.Y(n_16193)
);

NAND2xp5_ASAP7_75t_L g16194 ( 
.A(n_15671),
.B(n_15233),
.Y(n_16194)
);

HB1xp67_ASAP7_75t_L g16195 ( 
.A(n_16050),
.Y(n_16195)
);

AND2x2_ASAP7_75t_L g16196 ( 
.A(n_15903),
.B(n_15236),
.Y(n_16196)
);

AND2x2_ASAP7_75t_L g16197 ( 
.A(n_15478),
.B(n_15239),
.Y(n_16197)
);

OR2x2_ASAP7_75t_L g16198 ( 
.A(n_15684),
.B(n_15689),
.Y(n_16198)
);

AND2x2_ASAP7_75t_L g16199 ( 
.A(n_15538),
.B(n_15243),
.Y(n_16199)
);

OR2x2_ASAP7_75t_L g16200 ( 
.A(n_15712),
.B(n_15246),
.Y(n_16200)
);

INVx1_ASAP7_75t_L g16201 ( 
.A(n_15470),
.Y(n_16201)
);

BUFx3_ASAP7_75t_L g16202 ( 
.A(n_15688),
.Y(n_16202)
);

HB1xp67_ASAP7_75t_L g16203 ( 
.A(n_16057),
.Y(n_16203)
);

INVxp67_ASAP7_75t_L g16204 ( 
.A(n_15518),
.Y(n_16204)
);

NAND2xp5_ASAP7_75t_L g16205 ( 
.A(n_15833),
.B(n_15257),
.Y(n_16205)
);

INVx2_ASAP7_75t_SL g16206 ( 
.A(n_15473),
.Y(n_16206)
);

INVx2_ASAP7_75t_L g16207 ( 
.A(n_15525),
.Y(n_16207)
);

NAND2xp5_ASAP7_75t_L g16208 ( 
.A(n_15787),
.B(n_15519),
.Y(n_16208)
);

INVx2_ASAP7_75t_L g16209 ( 
.A(n_15527),
.Y(n_16209)
);

NOR2xp67_ASAP7_75t_L g16210 ( 
.A(n_16091),
.B(n_15259),
.Y(n_16210)
);

AND2x2_ASAP7_75t_L g16211 ( 
.A(n_15517),
.B(n_15264),
.Y(n_16211)
);

AND2x2_ASAP7_75t_L g16212 ( 
.A(n_15618),
.B(n_15270),
.Y(n_16212)
);

INVx1_ASAP7_75t_L g16213 ( 
.A(n_15472),
.Y(n_16213)
);

INVx2_ASAP7_75t_L g16214 ( 
.A(n_15554),
.Y(n_16214)
);

INVx2_ASAP7_75t_L g16215 ( 
.A(n_15479),
.Y(n_16215)
);

AND2x2_ASAP7_75t_L g16216 ( 
.A(n_15628),
.B(n_15287),
.Y(n_16216)
);

AND2x2_ASAP7_75t_L g16217 ( 
.A(n_15551),
.B(n_15515),
.Y(n_16217)
);

AND2x2_ASAP7_75t_L g16218 ( 
.A(n_15516),
.B(n_15288),
.Y(n_16218)
);

OR2x2_ASAP7_75t_L g16219 ( 
.A(n_15520),
.B(n_15578),
.Y(n_16219)
);

INVx1_ASAP7_75t_L g16220 ( 
.A(n_15480),
.Y(n_16220)
);

INVx2_ASAP7_75t_SL g16221 ( 
.A(n_15482),
.Y(n_16221)
);

NAND2xp5_ASAP7_75t_L g16222 ( 
.A(n_15579),
.B(n_15290),
.Y(n_16222)
);

INVx2_ASAP7_75t_L g16223 ( 
.A(n_15486),
.Y(n_16223)
);

INVx1_ASAP7_75t_L g16224 ( 
.A(n_15562),
.Y(n_16224)
);

NAND2xp5_ASAP7_75t_L g16225 ( 
.A(n_15582),
.B(n_15293),
.Y(n_16225)
);

AOI22xp33_ASAP7_75t_L g16226 ( 
.A1(n_15506),
.A2(n_15406),
.B1(n_15400),
.B2(n_14747),
.Y(n_16226)
);

INVx1_ASAP7_75t_L g16227 ( 
.A(n_15573),
.Y(n_16227)
);

NAND2xp5_ASAP7_75t_L g16228 ( 
.A(n_15619),
.B(n_15295),
.Y(n_16228)
);

INVx1_ASAP7_75t_L g16229 ( 
.A(n_15577),
.Y(n_16229)
);

INVx1_ASAP7_75t_L g16230 ( 
.A(n_15542),
.Y(n_16230)
);

OR2x2_ASAP7_75t_L g16231 ( 
.A(n_16020),
.B(n_15296),
.Y(n_16231)
);

AND2x2_ASAP7_75t_L g16232 ( 
.A(n_15784),
.B(n_15297),
.Y(n_16232)
);

INVx1_ASAP7_75t_L g16233 ( 
.A(n_15542),
.Y(n_16233)
);

OR2x2_ASAP7_75t_L g16234 ( 
.A(n_15714),
.B(n_15299),
.Y(n_16234)
);

AND2x2_ASAP7_75t_L g16235 ( 
.A(n_15594),
.B(n_15300),
.Y(n_16235)
);

NOR2xp33_ASAP7_75t_L g16236 ( 
.A(n_15720),
.B(n_15301),
.Y(n_16236)
);

NAND2xp33_ASAP7_75t_SL g16237 ( 
.A(n_15767),
.B(n_15302),
.Y(n_16237)
);

AND2x2_ASAP7_75t_L g16238 ( 
.A(n_15463),
.B(n_15311),
.Y(n_16238)
);

INVxp67_ASAP7_75t_SL g16239 ( 
.A(n_15612),
.Y(n_16239)
);

AND2x2_ASAP7_75t_L g16240 ( 
.A(n_15634),
.B(n_15319),
.Y(n_16240)
);

INVx2_ASAP7_75t_L g16241 ( 
.A(n_15490),
.Y(n_16241)
);

AND2x4_ASAP7_75t_SL g16242 ( 
.A(n_15939),
.B(n_15332),
.Y(n_16242)
);

INVx1_ASAP7_75t_L g16243 ( 
.A(n_15493),
.Y(n_16243)
);

AND2x2_ASAP7_75t_L g16244 ( 
.A(n_15933),
.B(n_15333),
.Y(n_16244)
);

NOR2xp33_ASAP7_75t_L g16245 ( 
.A(n_15673),
.B(n_14941),
.Y(n_16245)
);

NAND2xp5_ASAP7_75t_L g16246 ( 
.A(n_15730),
.B(n_14942),
.Y(n_16246)
);

AND2x2_ASAP7_75t_L g16247 ( 
.A(n_15676),
.B(n_15365),
.Y(n_16247)
);

NAND2xp5_ASAP7_75t_L g16248 ( 
.A(n_15600),
.B(n_15408),
.Y(n_16248)
);

INVx1_ASAP7_75t_L g16249 ( 
.A(n_15494),
.Y(n_16249)
);

INVx1_ASAP7_75t_L g16250 ( 
.A(n_15496),
.Y(n_16250)
);

AND2x2_ASAP7_75t_L g16251 ( 
.A(n_15908),
.B(n_10773),
.Y(n_16251)
);

INVx2_ASAP7_75t_SL g16252 ( 
.A(n_15511),
.Y(n_16252)
);

NAND2xp5_ASAP7_75t_L g16253 ( 
.A(n_15794),
.B(n_10334),
.Y(n_16253)
);

INVx2_ASAP7_75t_L g16254 ( 
.A(n_15501),
.Y(n_16254)
);

AND2x2_ASAP7_75t_L g16255 ( 
.A(n_15559),
.B(n_10778),
.Y(n_16255)
);

HB1xp67_ASAP7_75t_L g16256 ( 
.A(n_15561),
.Y(n_16256)
);

OR2x2_ASAP7_75t_L g16257 ( 
.A(n_15580),
.B(n_10778),
.Y(n_16257)
);

NAND2xp5_ASAP7_75t_L g16258 ( 
.A(n_15798),
.B(n_10338),
.Y(n_16258)
);

AND2x2_ASAP7_75t_L g16259 ( 
.A(n_15637),
.B(n_10784),
.Y(n_16259)
);

AND2x2_ASAP7_75t_L g16260 ( 
.A(n_15931),
.B(n_10784),
.Y(n_16260)
);

NAND2xp5_ASAP7_75t_L g16261 ( 
.A(n_15581),
.B(n_10338),
.Y(n_16261)
);

AND2x2_ASAP7_75t_L g16262 ( 
.A(n_15467),
.B(n_10792),
.Y(n_16262)
);

AND2x2_ASAP7_75t_L g16263 ( 
.A(n_15604),
.B(n_10792),
.Y(n_16263)
);

INVx1_ASAP7_75t_L g16264 ( 
.A(n_15508),
.Y(n_16264)
);

AND2x4_ASAP7_75t_SL g16265 ( 
.A(n_15939),
.B(n_8752),
.Y(n_16265)
);

NAND2xp5_ASAP7_75t_L g16266 ( 
.A(n_15782),
.B(n_10339),
.Y(n_16266)
);

INVx2_ASAP7_75t_L g16267 ( 
.A(n_15680),
.Y(n_16267)
);

INVx1_ASAP7_75t_L g16268 ( 
.A(n_15528),
.Y(n_16268)
);

INVx1_ASAP7_75t_L g16269 ( 
.A(n_15535),
.Y(n_16269)
);

INVx2_ASAP7_75t_L g16270 ( 
.A(n_15680),
.Y(n_16270)
);

INVx2_ASAP7_75t_L g16271 ( 
.A(n_15521),
.Y(n_16271)
);

AND2x2_ASAP7_75t_L g16272 ( 
.A(n_15604),
.B(n_10803),
.Y(n_16272)
);

INVx1_ASAP7_75t_L g16273 ( 
.A(n_15540),
.Y(n_16273)
);

NAND2xp5_ASAP7_75t_SL g16274 ( 
.A(n_15502),
.B(n_8468),
.Y(n_16274)
);

AND2x2_ASAP7_75t_L g16275 ( 
.A(n_15465),
.B(n_10803),
.Y(n_16275)
);

AND2x2_ASAP7_75t_L g16276 ( 
.A(n_15556),
.B(n_10804),
.Y(n_16276)
);

INVxp33_ASAP7_75t_L g16277 ( 
.A(n_15938),
.Y(n_16277)
);

INVx4_ASAP7_75t_L g16278 ( 
.A(n_15816),
.Y(n_16278)
);

HB1xp67_ASAP7_75t_L g16279 ( 
.A(n_15968),
.Y(n_16279)
);

OR2x2_ASAP7_75t_L g16280 ( 
.A(n_15914),
.B(n_10804),
.Y(n_16280)
);

AND2x2_ASAP7_75t_L g16281 ( 
.A(n_15588),
.B(n_10812),
.Y(n_16281)
);

INVx2_ASAP7_75t_SL g16282 ( 
.A(n_15476),
.Y(n_16282)
);

NAND2x1_ASAP7_75t_L g16283 ( 
.A(n_15722),
.B(n_10812),
.Y(n_16283)
);

AND2x2_ASAP7_75t_L g16284 ( 
.A(n_15729),
.B(n_10814),
.Y(n_16284)
);

AND2x2_ASAP7_75t_L g16285 ( 
.A(n_15731),
.B(n_10814),
.Y(n_16285)
);

AND2x2_ASAP7_75t_L g16286 ( 
.A(n_15483),
.B(n_10819),
.Y(n_16286)
);

INVx1_ASAP7_75t_L g16287 ( 
.A(n_15552),
.Y(n_16287)
);

AND2x2_ASAP7_75t_L g16288 ( 
.A(n_15567),
.B(n_10819),
.Y(n_16288)
);

CKINVDCx14_ASAP7_75t_R g16289 ( 
.A(n_15460),
.Y(n_16289)
);

AND2x2_ASAP7_75t_L g16290 ( 
.A(n_15553),
.B(n_10825),
.Y(n_16290)
);

NAND2x1p5_ASAP7_75t_L g16291 ( 
.A(n_15471),
.B(n_8468),
.Y(n_16291)
);

AND2x2_ASAP7_75t_L g16292 ( 
.A(n_15601),
.B(n_10825),
.Y(n_16292)
);

NOR2xp33_ASAP7_75t_SL g16293 ( 
.A(n_16023),
.B(n_8468),
.Y(n_16293)
);

AND2x2_ASAP7_75t_L g16294 ( 
.A(n_15499),
.B(n_10826),
.Y(n_16294)
);

AOI21xp5_ASAP7_75t_L g16295 ( 
.A1(n_15752),
.A2(n_10834),
.B(n_10826),
.Y(n_16295)
);

INVx1_ASAP7_75t_L g16296 ( 
.A(n_15748),
.Y(n_16296)
);

AND2x2_ASAP7_75t_L g16297 ( 
.A(n_16002),
.B(n_10834),
.Y(n_16297)
);

AND2x2_ASAP7_75t_L g16298 ( 
.A(n_16040),
.B(n_10846),
.Y(n_16298)
);

INVx2_ASAP7_75t_L g16299 ( 
.A(n_15654),
.Y(n_16299)
);

AND2x2_ASAP7_75t_L g16300 ( 
.A(n_15762),
.B(n_15772),
.Y(n_16300)
);

AND2x2_ASAP7_75t_L g16301 ( 
.A(n_15776),
.B(n_10846),
.Y(n_16301)
);

AND2x2_ASAP7_75t_L g16302 ( 
.A(n_15972),
.B(n_10851),
.Y(n_16302)
);

INVx2_ASAP7_75t_L g16303 ( 
.A(n_15941),
.Y(n_16303)
);

OR2x2_ASAP7_75t_L g16304 ( 
.A(n_15635),
.B(n_10851),
.Y(n_16304)
);

INVx1_ASAP7_75t_L g16305 ( 
.A(n_15785),
.Y(n_16305)
);

AND2x2_ASAP7_75t_L g16306 ( 
.A(n_15975),
.B(n_10853),
.Y(n_16306)
);

AND2x2_ASAP7_75t_L g16307 ( 
.A(n_15892),
.B(n_10853),
.Y(n_16307)
);

AND2x2_ASAP7_75t_L g16308 ( 
.A(n_16082),
.B(n_10858),
.Y(n_16308)
);

AND2x2_ASAP7_75t_L g16309 ( 
.A(n_15647),
.B(n_10858),
.Y(n_16309)
);

AND2x2_ASAP7_75t_L g16310 ( 
.A(n_15779),
.B(n_10869),
.Y(n_16310)
);

INVx4_ASAP7_75t_L g16311 ( 
.A(n_15940),
.Y(n_16311)
);

INVx1_ASAP7_75t_L g16312 ( 
.A(n_15786),
.Y(n_16312)
);

NOR2x1_ASAP7_75t_L g16313 ( 
.A(n_15512),
.B(n_10869),
.Y(n_16313)
);

INVx1_ASAP7_75t_L g16314 ( 
.A(n_15523),
.Y(n_16314)
);

INVx2_ASAP7_75t_SL g16315 ( 
.A(n_15722),
.Y(n_16315)
);

HB1xp67_ASAP7_75t_L g16316 ( 
.A(n_16009),
.Y(n_16316)
);

INVx1_ASAP7_75t_L g16317 ( 
.A(n_15526),
.Y(n_16317)
);

INVx1_ASAP7_75t_L g16318 ( 
.A(n_15566),
.Y(n_16318)
);

NAND2xp5_ASAP7_75t_L g16319 ( 
.A(n_15742),
.B(n_10339),
.Y(n_16319)
);

HB1xp67_ASAP7_75t_L g16320 ( 
.A(n_15964),
.Y(n_16320)
);

INVx1_ASAP7_75t_L g16321 ( 
.A(n_15522),
.Y(n_16321)
);

OR2x2_ASAP7_75t_L g16322 ( 
.A(n_15745),
.B(n_10870),
.Y(n_16322)
);

AOI22xp33_ASAP7_75t_L g16323 ( 
.A1(n_15717),
.A2(n_11743),
.B1(n_8096),
.B2(n_10291),
.Y(n_16323)
);

INVx2_ASAP7_75t_L g16324 ( 
.A(n_16034),
.Y(n_16324)
);

AND2x2_ASAP7_75t_L g16325 ( 
.A(n_15944),
.B(n_10870),
.Y(n_16325)
);

INVx1_ASAP7_75t_L g16326 ( 
.A(n_15500),
.Y(n_16326)
);

AND2x2_ASAP7_75t_L g16327 ( 
.A(n_15817),
.B(n_10874),
.Y(n_16327)
);

OR2x2_ASAP7_75t_L g16328 ( 
.A(n_15750),
.B(n_10874),
.Y(n_16328)
);

AND2x2_ASAP7_75t_L g16329 ( 
.A(n_16085),
.B(n_10886),
.Y(n_16329)
);

AOI22xp33_ASAP7_75t_L g16330 ( 
.A1(n_15558),
.A2(n_8096),
.B1(n_10291),
.B2(n_9473),
.Y(n_16330)
);

AND2x2_ASAP7_75t_L g16331 ( 
.A(n_16086),
.B(n_10886),
.Y(n_16331)
);

INVx2_ASAP7_75t_L g16332 ( 
.A(n_15707),
.Y(n_16332)
);

NAND3xp33_ASAP7_75t_L g16333 ( 
.A(n_15672),
.B(n_15622),
.C(n_15583),
.Y(n_16333)
);

AND2x4_ASAP7_75t_L g16334 ( 
.A(n_15755),
.B(n_8686),
.Y(n_16334)
);

AND2x2_ASAP7_75t_L g16335 ( 
.A(n_16092),
.B(n_10889),
.Y(n_16335)
);

AND2x2_ASAP7_75t_L g16336 ( 
.A(n_15905),
.B(n_10889),
.Y(n_16336)
);

AND2x2_ASAP7_75t_L g16337 ( 
.A(n_15807),
.B(n_10891),
.Y(n_16337)
);

NAND2xp5_ASAP7_75t_L g16338 ( 
.A(n_15586),
.B(n_15595),
.Y(n_16338)
);

INVx1_ASAP7_75t_L g16339 ( 
.A(n_15607),
.Y(n_16339)
);

INVx1_ASAP7_75t_L g16340 ( 
.A(n_15610),
.Y(n_16340)
);

INVx2_ASAP7_75t_L g16341 ( 
.A(n_15652),
.Y(n_16341)
);

INVx3_ASAP7_75t_L g16342 ( 
.A(n_15477),
.Y(n_16342)
);

NAND2xp5_ASAP7_75t_L g16343 ( 
.A(n_15611),
.B(n_10340),
.Y(n_16343)
);

AND2x2_ASAP7_75t_L g16344 ( 
.A(n_15813),
.B(n_10891),
.Y(n_16344)
);

HB1xp67_ASAP7_75t_L g16345 ( 
.A(n_16065),
.Y(n_16345)
);

INVxp67_ASAP7_75t_SL g16346 ( 
.A(n_15609),
.Y(n_16346)
);

INVx1_ASAP7_75t_L g16347 ( 
.A(n_15621),
.Y(n_16347)
);

OR2x2_ASAP7_75t_L g16348 ( 
.A(n_15568),
.B(n_10893),
.Y(n_16348)
);

INVx3_ASAP7_75t_L g16349 ( 
.A(n_15655),
.Y(n_16349)
);

INVx5_ASAP7_75t_L g16350 ( 
.A(n_15936),
.Y(n_16350)
);

NOR2xp33_ASAP7_75t_L g16351 ( 
.A(n_15895),
.B(n_8468),
.Y(n_16351)
);

NOR2xp33_ASAP7_75t_L g16352 ( 
.A(n_15533),
.B(n_8468),
.Y(n_16352)
);

NAND2xp5_ASAP7_75t_L g16353 ( 
.A(n_15617),
.B(n_10340),
.Y(n_16353)
);

NAND2xp5_ASAP7_75t_L g16354 ( 
.A(n_16013),
.B(n_10341),
.Y(n_16354)
);

NAND2xp5_ASAP7_75t_L g16355 ( 
.A(n_15897),
.B(n_10341),
.Y(n_16355)
);

AND2x4_ASAP7_75t_L g16356 ( 
.A(n_15822),
.B(n_8686),
.Y(n_16356)
);

AND2x2_ASAP7_75t_L g16357 ( 
.A(n_15814),
.B(n_10893),
.Y(n_16357)
);

NOR2xp33_ASAP7_75t_L g16358 ( 
.A(n_15616),
.B(n_8468),
.Y(n_16358)
);

AND2x2_ASAP7_75t_L g16359 ( 
.A(n_15815),
.B(n_10894),
.Y(n_16359)
);

AND2x2_ASAP7_75t_L g16360 ( 
.A(n_15797),
.B(n_10894),
.Y(n_16360)
);

INVx1_ASAP7_75t_L g16361 ( 
.A(n_15534),
.Y(n_16361)
);

INVx1_ASAP7_75t_L g16362 ( 
.A(n_15536),
.Y(n_16362)
);

INVx2_ASAP7_75t_L g16363 ( 
.A(n_15630),
.Y(n_16363)
);

NOR2xp67_ASAP7_75t_L g16364 ( 
.A(n_15930),
.B(n_10895),
.Y(n_16364)
);

AND2x2_ASAP7_75t_L g16365 ( 
.A(n_15856),
.B(n_10895),
.Y(n_16365)
);

AND2x2_ASAP7_75t_L g16366 ( 
.A(n_15943),
.B(n_10900),
.Y(n_16366)
);

AND2x2_ASAP7_75t_L g16367 ( 
.A(n_15915),
.B(n_15924),
.Y(n_16367)
);

NAND2xp5_ASAP7_75t_L g16368 ( 
.A(n_15827),
.B(n_10343),
.Y(n_16368)
);

AND2x2_ASAP7_75t_L g16369 ( 
.A(n_15921),
.B(n_10900),
.Y(n_16369)
);

NAND2xp5_ASAP7_75t_SL g16370 ( 
.A(n_15591),
.B(n_8481),
.Y(n_16370)
);

INVx1_ASAP7_75t_SL g16371 ( 
.A(n_15468),
.Y(n_16371)
);

OR2x2_ASAP7_75t_L g16372 ( 
.A(n_15801),
.B(n_10902),
.Y(n_16372)
);

AND2x2_ASAP7_75t_L g16373 ( 
.A(n_15503),
.B(n_10902),
.Y(n_16373)
);

INVx2_ASAP7_75t_L g16374 ( 
.A(n_15513),
.Y(n_16374)
);

INVx1_ASAP7_75t_L g16375 ( 
.A(n_15495),
.Y(n_16375)
);

INVx1_ASAP7_75t_L g16376 ( 
.A(n_15507),
.Y(n_16376)
);

NAND2x1_ASAP7_75t_SL g16377 ( 
.A(n_16021),
.B(n_9445),
.Y(n_16377)
);

NAND2xp5_ASAP7_75t_L g16378 ( 
.A(n_15880),
.B(n_10350),
.Y(n_16378)
);

INVxp67_ASAP7_75t_L g16379 ( 
.A(n_15919),
.Y(n_16379)
);

INVx2_ASAP7_75t_L g16380 ( 
.A(n_15806),
.Y(n_16380)
);

HB1xp67_ASAP7_75t_L g16381 ( 
.A(n_15890),
.Y(n_16381)
);

INVxp67_ASAP7_75t_L g16382 ( 
.A(n_15596),
.Y(n_16382)
);

AND2x4_ASAP7_75t_L g16383 ( 
.A(n_16033),
.B(n_8686),
.Y(n_16383)
);

AND2x2_ASAP7_75t_L g16384 ( 
.A(n_16037),
.B(n_10908),
.Y(n_16384)
);

BUFx2_ASAP7_75t_L g16385 ( 
.A(n_15724),
.Y(n_16385)
);

AND2x2_ASAP7_75t_L g16386 ( 
.A(n_16078),
.B(n_15643),
.Y(n_16386)
);

INVx1_ASAP7_75t_L g16387 ( 
.A(n_15505),
.Y(n_16387)
);

OR2x2_ASAP7_75t_L g16388 ( 
.A(n_16038),
.B(n_10908),
.Y(n_16388)
);

AND2x2_ASAP7_75t_L g16389 ( 
.A(n_16074),
.B(n_10918),
.Y(n_16389)
);

INVx1_ASAP7_75t_L g16390 ( 
.A(n_15585),
.Y(n_16390)
);

INVx2_ASAP7_75t_L g16391 ( 
.A(n_15980),
.Y(n_16391)
);

INVx1_ASAP7_75t_L g16392 ( 
.A(n_15541),
.Y(n_16392)
);

NAND2xp5_ASAP7_75t_L g16393 ( 
.A(n_15898),
.B(n_10350),
.Y(n_16393)
);

INVx1_ASAP7_75t_L g16394 ( 
.A(n_15532),
.Y(n_16394)
);

INVx2_ASAP7_75t_L g16395 ( 
.A(n_15724),
.Y(n_16395)
);

INVx2_ASAP7_75t_SL g16396 ( 
.A(n_15702),
.Y(n_16396)
);

NAND2xp5_ASAP7_75t_L g16397 ( 
.A(n_15901),
.B(n_10357),
.Y(n_16397)
);

INVx2_ASAP7_75t_L g16398 ( 
.A(n_15738),
.Y(n_16398)
);

NAND2xp5_ASAP7_75t_L g16399 ( 
.A(n_15751),
.B(n_15753),
.Y(n_16399)
);

INVx1_ASAP7_75t_L g16400 ( 
.A(n_15530),
.Y(n_16400)
);

AND2x4_ASAP7_75t_L g16401 ( 
.A(n_16076),
.B(n_8686),
.Y(n_16401)
);

AND2x2_ASAP7_75t_L g16402 ( 
.A(n_15548),
.B(n_10918),
.Y(n_16402)
);

AND2x2_ASAP7_75t_L g16403 ( 
.A(n_15828),
.B(n_15877),
.Y(n_16403)
);

INVx1_ASAP7_75t_L g16404 ( 
.A(n_15539),
.Y(n_16404)
);

NAND2xp5_ASAP7_75t_L g16405 ( 
.A(n_15757),
.B(n_10357),
.Y(n_16405)
);

AND2x2_ASAP7_75t_L g16406 ( 
.A(n_15636),
.B(n_10919),
.Y(n_16406)
);

NAND2xp5_ASAP7_75t_L g16407 ( 
.A(n_15759),
.B(n_10359),
.Y(n_16407)
);

INVx1_ASAP7_75t_L g16408 ( 
.A(n_15557),
.Y(n_16408)
);

INVx1_ASAP7_75t_L g16409 ( 
.A(n_15670),
.Y(n_16409)
);

AND2x2_ASAP7_75t_L g16410 ( 
.A(n_15928),
.B(n_10919),
.Y(n_16410)
);

INVx1_ASAP7_75t_L g16411 ( 
.A(n_15692),
.Y(n_16411)
);

INVx3_ASAP7_75t_L g16412 ( 
.A(n_15846),
.Y(n_16412)
);

INVx1_ASAP7_75t_L g16413 ( 
.A(n_15703),
.Y(n_16413)
);

NOR2xp33_ASAP7_75t_L g16414 ( 
.A(n_15584),
.B(n_8481),
.Y(n_16414)
);

INVx1_ASAP7_75t_L g16415 ( 
.A(n_15974),
.Y(n_16415)
);

INVx2_ASAP7_75t_L g16416 ( 
.A(n_15738),
.Y(n_16416)
);

AND2x2_ASAP7_75t_L g16417 ( 
.A(n_15913),
.B(n_10924),
.Y(n_16417)
);

INVx2_ASAP7_75t_L g16418 ( 
.A(n_15760),
.Y(n_16418)
);

INVx1_ASAP7_75t_L g16419 ( 
.A(n_15760),
.Y(n_16419)
);

AND2x2_ASAP7_75t_SL g16420 ( 
.A(n_15572),
.B(n_7991),
.Y(n_16420)
);

NAND3xp33_ASAP7_75t_L g16421 ( 
.A(n_15906),
.B(n_9473),
.C(n_9369),
.Y(n_16421)
);

NAND2xp5_ASAP7_75t_L g16422 ( 
.A(n_15765),
.B(n_10359),
.Y(n_16422)
);

INVx1_ASAP7_75t_L g16423 ( 
.A(n_15560),
.Y(n_16423)
);

AND2x2_ASAP7_75t_L g16424 ( 
.A(n_15662),
.B(n_10924),
.Y(n_16424)
);

NAND2xp5_ASAP7_75t_SL g16425 ( 
.A(n_15629),
.B(n_8481),
.Y(n_16425)
);

HB1xp67_ASAP7_75t_L g16426 ( 
.A(n_15704),
.Y(n_16426)
);

INVx1_ASAP7_75t_L g16427 ( 
.A(n_15769),
.Y(n_16427)
);

AND2x2_ASAP7_75t_L g16428 ( 
.A(n_15570),
.B(n_15770),
.Y(n_16428)
);

AND2x2_ASAP7_75t_L g16429 ( 
.A(n_15778),
.B(n_10932),
.Y(n_16429)
);

OR2x2_ASAP7_75t_L g16430 ( 
.A(n_15589),
.B(n_15475),
.Y(n_16430)
);

HB1xp67_ASAP7_75t_L g16431 ( 
.A(n_15711),
.Y(n_16431)
);

INVx2_ASAP7_75t_L g16432 ( 
.A(n_15842),
.Y(n_16432)
);

NAND2xp5_ASAP7_75t_L g16433 ( 
.A(n_15706),
.B(n_10363),
.Y(n_16433)
);

AND2x2_ASAP7_75t_L g16434 ( 
.A(n_15773),
.B(n_10932),
.Y(n_16434)
);

HB1xp67_ASAP7_75t_L g16435 ( 
.A(n_15754),
.Y(n_16435)
);

OR2x2_ASAP7_75t_L g16436 ( 
.A(n_15747),
.B(n_10944),
.Y(n_16436)
);

NAND2xp5_ASAP7_75t_L g16437 ( 
.A(n_15888),
.B(n_10367),
.Y(n_16437)
);

OR2x2_ASAP7_75t_L g16438 ( 
.A(n_15457),
.B(n_10944),
.Y(n_16438)
);

NOR2xp33_ASAP7_75t_R g16439 ( 
.A(n_15690),
.B(n_8597),
.Y(n_16439)
);

HB1xp67_ASAP7_75t_L g16440 ( 
.A(n_15821),
.Y(n_16440)
);

NAND2xp5_ASAP7_75t_L g16441 ( 
.A(n_15631),
.B(n_10367),
.Y(n_16441)
);

NAND2xp5_ASAP7_75t_SL g16442 ( 
.A(n_15808),
.B(n_8481),
.Y(n_16442)
);

INVx2_ASAP7_75t_SL g16443 ( 
.A(n_15988),
.Y(n_16443)
);

AND2x2_ASAP7_75t_L g16444 ( 
.A(n_15633),
.B(n_10945),
.Y(n_16444)
);

INVx2_ASAP7_75t_SL g16445 ( 
.A(n_15843),
.Y(n_16445)
);

NAND2xp5_ASAP7_75t_L g16446 ( 
.A(n_15663),
.B(n_10368),
.Y(n_16446)
);

INVx1_ASAP7_75t_L g16447 ( 
.A(n_15614),
.Y(n_16447)
);

AND2x4_ASAP7_75t_SL g16448 ( 
.A(n_15946),
.B(n_8752),
.Y(n_16448)
);

OR2x2_ASAP7_75t_L g16449 ( 
.A(n_15563),
.B(n_10945),
.Y(n_16449)
);

AND2x4_ASAP7_75t_L g16450 ( 
.A(n_16087),
.B(n_8686),
.Y(n_16450)
);

INVx1_ASAP7_75t_L g16451 ( 
.A(n_15625),
.Y(n_16451)
);

INVx1_ASAP7_75t_L g16452 ( 
.A(n_15564),
.Y(n_16452)
);

AND2x2_ASAP7_75t_L g16453 ( 
.A(n_16093),
.B(n_10949),
.Y(n_16453)
);

AND2x2_ASAP7_75t_L g16454 ( 
.A(n_16094),
.B(n_10949),
.Y(n_16454)
);

INVx2_ASAP7_75t_L g16455 ( 
.A(n_15910),
.Y(n_16455)
);

INVx1_ASAP7_75t_L g16456 ( 
.A(n_15597),
.Y(n_16456)
);

AND2x2_ASAP7_75t_L g16457 ( 
.A(n_15853),
.B(n_10964),
.Y(n_16457)
);

AND2x4_ASAP7_75t_SL g16458 ( 
.A(n_15961),
.B(n_8752),
.Y(n_16458)
);

OR2x2_ASAP7_75t_L g16459 ( 
.A(n_15474),
.B(n_15603),
.Y(n_16459)
);

INVxp67_ASAP7_75t_L g16460 ( 
.A(n_15674),
.Y(n_16460)
);

INVx1_ASAP7_75t_L g16461 ( 
.A(n_15606),
.Y(n_16461)
);

INVxp67_ASAP7_75t_L g16462 ( 
.A(n_15651),
.Y(n_16462)
);

AND2x2_ASAP7_75t_L g16463 ( 
.A(n_15917),
.B(n_10964),
.Y(n_16463)
);

HB1xp67_ASAP7_75t_L g16464 ( 
.A(n_15982),
.Y(n_16464)
);

INVx1_ASAP7_75t_L g16465 ( 
.A(n_15608),
.Y(n_16465)
);

OR2x2_ASAP7_75t_L g16466 ( 
.A(n_15615),
.B(n_10971),
.Y(n_16466)
);

AND2x2_ASAP7_75t_L g16467 ( 
.A(n_15796),
.B(n_10971),
.Y(n_16467)
);

CKINVDCx20_ASAP7_75t_R g16468 ( 
.A(n_15531),
.Y(n_16468)
);

INVx2_ASAP7_75t_L g16469 ( 
.A(n_16062),
.Y(n_16469)
);

AND2x2_ASAP7_75t_L g16470 ( 
.A(n_15789),
.B(n_10977),
.Y(n_16470)
);

INVx1_ASAP7_75t_L g16471 ( 
.A(n_16055),
.Y(n_16471)
);

AND2x2_ASAP7_75t_L g16472 ( 
.A(n_15743),
.B(n_10977),
.Y(n_16472)
);

INVx1_ASAP7_75t_L g16473 ( 
.A(n_16063),
.Y(n_16473)
);

AND2x2_ASAP7_75t_L g16474 ( 
.A(n_15850),
.B(n_10995),
.Y(n_16474)
);

HB1xp67_ASAP7_75t_L g16475 ( 
.A(n_16029),
.Y(n_16475)
);

INVx1_ASAP7_75t_SL g16476 ( 
.A(n_15788),
.Y(n_16476)
);

NAND4xp25_ASAP7_75t_SL g16477 ( 
.A(n_15959),
.B(n_10998),
.C(n_10999),
.D(n_10995),
.Y(n_16477)
);

NAND2x1_ASAP7_75t_L g16478 ( 
.A(n_15824),
.B(n_10998),
.Y(n_16478)
);

INVx1_ASAP7_75t_L g16479 ( 
.A(n_15728),
.Y(n_16479)
);

INVx1_ASAP7_75t_L g16480 ( 
.A(n_15687),
.Y(n_16480)
);

INVx1_ASAP7_75t_L g16481 ( 
.A(n_15957),
.Y(n_16481)
);

NAND2xp5_ASAP7_75t_L g16482 ( 
.A(n_15696),
.B(n_10368),
.Y(n_16482)
);

INVx1_ASAP7_75t_L g16483 ( 
.A(n_15867),
.Y(n_16483)
);

AND2x2_ASAP7_75t_L g16484 ( 
.A(n_15851),
.B(n_10999),
.Y(n_16484)
);

AND2x2_ASAP7_75t_L g16485 ( 
.A(n_15852),
.B(n_11001),
.Y(n_16485)
);

AND2x2_ASAP7_75t_L g16486 ( 
.A(n_15726),
.B(n_11001),
.Y(n_16486)
);

AND2x2_ASAP7_75t_L g16487 ( 
.A(n_15764),
.B(n_15700),
.Y(n_16487)
);

OR2x2_ASAP7_75t_L g16488 ( 
.A(n_15697),
.B(n_11004),
.Y(n_16488)
);

INVxp67_ASAP7_75t_L g16489 ( 
.A(n_15732),
.Y(n_16489)
);

NAND2xp5_ASAP7_75t_L g16490 ( 
.A(n_15699),
.B(n_15705),
.Y(n_16490)
);

AOI21xp33_ASAP7_75t_L g16491 ( 
.A1(n_15590),
.A2(n_11079),
.B(n_11076),
.Y(n_16491)
);

INVx2_ASAP7_75t_L g16492 ( 
.A(n_15956),
.Y(n_16492)
);

AND2x2_ASAP7_75t_L g16493 ( 
.A(n_15965),
.B(n_11004),
.Y(n_16493)
);

BUFx12f_ASAP7_75t_L g16494 ( 
.A(n_15632),
.Y(n_16494)
);

AND2x2_ASAP7_75t_L g16495 ( 
.A(n_15990),
.B(n_11012),
.Y(n_16495)
);

INVx1_ASAP7_75t_SL g16496 ( 
.A(n_15638),
.Y(n_16496)
);

NAND2xp5_ASAP7_75t_L g16497 ( 
.A(n_15954),
.B(n_10369),
.Y(n_16497)
);

NAND2xp5_ASAP7_75t_L g16498 ( 
.A(n_15973),
.B(n_10369),
.Y(n_16498)
);

INVx2_ASAP7_75t_L g16499 ( 
.A(n_15978),
.Y(n_16499)
);

NOR2xp33_ASAP7_75t_L g16500 ( 
.A(n_15902),
.B(n_8481),
.Y(n_16500)
);

INVx1_ASAP7_75t_L g16501 ( 
.A(n_15812),
.Y(n_16501)
);

INVx1_ASAP7_75t_L g16502 ( 
.A(n_15872),
.Y(n_16502)
);

NAND2xp5_ASAP7_75t_L g16503 ( 
.A(n_16000),
.B(n_10376),
.Y(n_16503)
);

INVx1_ASAP7_75t_L g16504 ( 
.A(n_15825),
.Y(n_16504)
);

INVx1_ASAP7_75t_L g16505 ( 
.A(n_15809),
.Y(n_16505)
);

AND2x2_ASAP7_75t_L g16506 ( 
.A(n_15993),
.B(n_11012),
.Y(n_16506)
);

INVx1_ASAP7_75t_L g16507 ( 
.A(n_16001),
.Y(n_16507)
);

INVx1_ASAP7_75t_L g16508 ( 
.A(n_16007),
.Y(n_16508)
);

AND2x2_ASAP7_75t_L g16509 ( 
.A(n_16017),
.B(n_11017),
.Y(n_16509)
);

AND2x2_ASAP7_75t_L g16510 ( 
.A(n_15869),
.B(n_11017),
.Y(n_16510)
);

AND2x2_ASAP7_75t_L g16511 ( 
.A(n_15874),
.B(n_11020),
.Y(n_16511)
);

AND2x2_ASAP7_75t_L g16512 ( 
.A(n_15878),
.B(n_15879),
.Y(n_16512)
);

AND2x4_ASAP7_75t_L g16513 ( 
.A(n_16024),
.B(n_8745),
.Y(n_16513)
);

BUFx6f_ASAP7_75t_L g16514 ( 
.A(n_15719),
.Y(n_16514)
);

INVx1_ASAP7_75t_L g16515 ( 
.A(n_15802),
.Y(n_16515)
);

INVx1_ASAP7_75t_L g16516 ( 
.A(n_15803),
.Y(n_16516)
);

INVx1_ASAP7_75t_L g16517 ( 
.A(n_15804),
.Y(n_16517)
);

AOI22xp33_ASAP7_75t_L g16518 ( 
.A1(n_15945),
.A2(n_10291),
.B1(n_9473),
.B2(n_9614),
.Y(n_16518)
);

AND2x2_ASAP7_75t_L g16519 ( 
.A(n_16025),
.B(n_11020),
.Y(n_16519)
);

AND2x2_ASAP7_75t_L g16520 ( 
.A(n_15679),
.B(n_11021),
.Y(n_16520)
);

AND2x2_ASAP7_75t_L g16521 ( 
.A(n_15783),
.B(n_15805),
.Y(n_16521)
);

AND2x4_ASAP7_75t_L g16522 ( 
.A(n_16073),
.B(n_8745),
.Y(n_16522)
);

INVx1_ASAP7_75t_L g16523 ( 
.A(n_15861),
.Y(n_16523)
);

INVx2_ASAP7_75t_L g16524 ( 
.A(n_15912),
.Y(n_16524)
);

NAND2xp5_ASAP7_75t_L g16525 ( 
.A(n_15734),
.B(n_10376),
.Y(n_16525)
);

INVxp67_ASAP7_75t_SL g16526 ( 
.A(n_15775),
.Y(n_16526)
);

INVx1_ASAP7_75t_L g16527 ( 
.A(n_15863),
.Y(n_16527)
);

AND2x4_ASAP7_75t_L g16528 ( 
.A(n_16075),
.B(n_8745),
.Y(n_16528)
);

INVx1_ASAP7_75t_L g16529 ( 
.A(n_15683),
.Y(n_16529)
);

AND2x2_ASAP7_75t_L g16530 ( 
.A(n_15694),
.B(n_11021),
.Y(n_16530)
);

INVx1_ASAP7_75t_SL g16531 ( 
.A(n_15795),
.Y(n_16531)
);

INVx3_ASAP7_75t_SL g16532 ( 
.A(n_15737),
.Y(n_16532)
);

AND2x2_ASAP7_75t_L g16533 ( 
.A(n_15708),
.B(n_11022),
.Y(n_16533)
);

OR2x2_ASAP7_75t_L g16534 ( 
.A(n_15739),
.B(n_11022),
.Y(n_16534)
);

HB1xp67_ASAP7_75t_L g16535 ( 
.A(n_16039),
.Y(n_16535)
);

AND2x2_ASAP7_75t_L g16536 ( 
.A(n_15721),
.B(n_11025),
.Y(n_16536)
);

AND2x4_ASAP7_75t_L g16537 ( 
.A(n_15741),
.B(n_8745),
.Y(n_16537)
);

INVx1_ASAP7_75t_L g16538 ( 
.A(n_16011),
.Y(n_16538)
);

OR2x2_ASAP7_75t_L g16539 ( 
.A(n_15876),
.B(n_11025),
.Y(n_16539)
);

HB1xp67_ASAP7_75t_L g16540 ( 
.A(n_15763),
.Y(n_16540)
);

CKINVDCx16_ASAP7_75t_R g16541 ( 
.A(n_16067),
.Y(n_16541)
);

AND2x2_ASAP7_75t_L g16542 ( 
.A(n_15790),
.B(n_11027),
.Y(n_16542)
);

AND2x2_ASAP7_75t_L g16543 ( 
.A(n_15900),
.B(n_11027),
.Y(n_16543)
);

INVx2_ASAP7_75t_L g16544 ( 
.A(n_15777),
.Y(n_16544)
);

OR2x2_ASAP7_75t_L g16545 ( 
.A(n_15934),
.B(n_11036),
.Y(n_16545)
);

NOR4xp25_ASAP7_75t_SL g16546 ( 
.A(n_15810),
.B(n_8050),
.C(n_8092),
.D(n_7944),
.Y(n_16546)
);

AND2x2_ASAP7_75t_L g16547 ( 
.A(n_15771),
.B(n_11036),
.Y(n_16547)
);

AND2x2_ASAP7_75t_L g16548 ( 
.A(n_15819),
.B(n_11047),
.Y(n_16548)
);

AND2x2_ASAP7_75t_L g16549 ( 
.A(n_15826),
.B(n_11047),
.Y(n_16549)
);

AND2x2_ASAP7_75t_L g16550 ( 
.A(n_15834),
.B(n_11048),
.Y(n_16550)
);

NAND2xp5_ASAP7_75t_L g16551 ( 
.A(n_15849),
.B(n_10377),
.Y(n_16551)
);

INVx2_ASAP7_75t_L g16552 ( 
.A(n_15768),
.Y(n_16552)
);

OR2x2_ASAP7_75t_L g16553 ( 
.A(n_15935),
.B(n_11048),
.Y(n_16553)
);

INVx3_ASAP7_75t_L g16554 ( 
.A(n_16054),
.Y(n_16554)
);

AND2x2_ASAP7_75t_L g16555 ( 
.A(n_15835),
.B(n_8745),
.Y(n_16555)
);

INVx1_ASAP7_75t_L g16556 ( 
.A(n_15749),
.Y(n_16556)
);

INVx2_ASAP7_75t_L g16557 ( 
.A(n_15970),
.Y(n_16557)
);

AND2x2_ASAP7_75t_L g16558 ( 
.A(n_15837),
.B(n_8745),
.Y(n_16558)
);

AND2x2_ASAP7_75t_L g16559 ( 
.A(n_15845),
.B(n_15847),
.Y(n_16559)
);

AND2x2_ASAP7_75t_L g16560 ( 
.A(n_15848),
.B(n_8765),
.Y(n_16560)
);

AND2x2_ASAP7_75t_L g16561 ( 
.A(n_15854),
.B(n_8765),
.Y(n_16561)
);

NAND2xp5_ASAP7_75t_L g16562 ( 
.A(n_15627),
.B(n_10377),
.Y(n_16562)
);

INVx1_ASAP7_75t_L g16563 ( 
.A(n_15644),
.Y(n_16563)
);

HB1xp67_ASAP7_75t_L g16564 ( 
.A(n_15698),
.Y(n_16564)
);

NAND2xp5_ASAP7_75t_L g16565 ( 
.A(n_15648),
.B(n_10389),
.Y(n_16565)
);

AND2x2_ASAP7_75t_L g16566 ( 
.A(n_15858),
.B(n_8765),
.Y(n_16566)
);

INVxp67_ASAP7_75t_L g16567 ( 
.A(n_15836),
.Y(n_16567)
);

INVx1_ASAP7_75t_L g16568 ( 
.A(n_15830),
.Y(n_16568)
);

INVx1_ASAP7_75t_L g16569 ( 
.A(n_15891),
.Y(n_16569)
);

INVx3_ASAP7_75t_L g16570 ( 
.A(n_16068),
.Y(n_16570)
);

HB1xp67_ASAP7_75t_L g16571 ( 
.A(n_16010),
.Y(n_16571)
);

INVx2_ASAP7_75t_SL g16572 ( 
.A(n_16052),
.Y(n_16572)
);

INVx1_ASAP7_75t_L g16573 ( 
.A(n_15894),
.Y(n_16573)
);

INVx1_ASAP7_75t_L g16574 ( 
.A(n_15733),
.Y(n_16574)
);

INVx1_ASAP7_75t_L g16575 ( 
.A(n_15736),
.Y(n_16575)
);

NAND2xp5_ASAP7_75t_L g16576 ( 
.A(n_15950),
.B(n_15952),
.Y(n_16576)
);

INVx1_ASAP7_75t_L g16577 ( 
.A(n_15766),
.Y(n_16577)
);

AND2x2_ASAP7_75t_L g16578 ( 
.A(n_15875),
.B(n_15885),
.Y(n_16578)
);

AND2x2_ASAP7_75t_L g16579 ( 
.A(n_15984),
.B(n_15889),
.Y(n_16579)
);

AND2x2_ASAP7_75t_L g16580 ( 
.A(n_15989),
.B(n_8765),
.Y(n_16580)
);

AND2x2_ASAP7_75t_L g16581 ( 
.A(n_15992),
.B(n_8765),
.Y(n_16581)
);

AND2x2_ASAP7_75t_L g16582 ( 
.A(n_15844),
.B(n_8765),
.Y(n_16582)
);

NOR2x1_ASAP7_75t_L g16583 ( 
.A(n_15713),
.B(n_11097),
.Y(n_16583)
);

AND2x2_ASAP7_75t_L g16584 ( 
.A(n_15907),
.B(n_8767),
.Y(n_16584)
);

OR2x2_ASAP7_75t_L g16585 ( 
.A(n_15953),
.B(n_15675),
.Y(n_16585)
);

AND2x2_ASAP7_75t_L g16586 ( 
.A(n_15955),
.B(n_8767),
.Y(n_16586)
);

NAND2xp5_ASAP7_75t_L g16587 ( 
.A(n_16026),
.B(n_10389),
.Y(n_16587)
);

AND2x2_ASAP7_75t_L g16588 ( 
.A(n_15818),
.B(n_8767),
.Y(n_16588)
);

INVx1_ASAP7_75t_L g16589 ( 
.A(n_15799),
.Y(n_16589)
);

INVx1_ASAP7_75t_L g16590 ( 
.A(n_15829),
.Y(n_16590)
);

HB1xp67_ASAP7_75t_L g16591 ( 
.A(n_16012),
.Y(n_16591)
);

AND2x2_ASAP7_75t_L g16592 ( 
.A(n_15664),
.B(n_8767),
.Y(n_16592)
);

INVx1_ASAP7_75t_L g16593 ( 
.A(n_15832),
.Y(n_16593)
);

NAND2xp5_ASAP7_75t_L g16594 ( 
.A(n_16044),
.B(n_10390),
.Y(n_16594)
);

INVx2_ASAP7_75t_L g16595 ( 
.A(n_15873),
.Y(n_16595)
);

INVx1_ASAP7_75t_L g16596 ( 
.A(n_15857),
.Y(n_16596)
);

INVx1_ASAP7_75t_L g16597 ( 
.A(n_15859),
.Y(n_16597)
);

NAND2x1p5_ASAP7_75t_L g16598 ( 
.A(n_15918),
.B(n_8481),
.Y(n_16598)
);

INVx1_ASAP7_75t_L g16599 ( 
.A(n_15865),
.Y(n_16599)
);

AND2x2_ASAP7_75t_L g16600 ( 
.A(n_16014),
.B(n_8767),
.Y(n_16600)
);

NAND2xp5_ASAP7_75t_L g16601 ( 
.A(n_15838),
.B(n_10390),
.Y(n_16601)
);

AOI22xp33_ASAP7_75t_L g16602 ( 
.A1(n_15693),
.A2(n_15665),
.B1(n_15682),
.B2(n_15871),
.Y(n_16602)
);

AND2x2_ASAP7_75t_L g16603 ( 
.A(n_15916),
.B(n_8767),
.Y(n_16603)
);

INVx1_ASAP7_75t_L g16604 ( 
.A(n_15884),
.Y(n_16604)
);

INVxp67_ASAP7_75t_L g16605 ( 
.A(n_15725),
.Y(n_16605)
);

AND2x2_ASAP7_75t_L g16606 ( 
.A(n_15923),
.B(n_8804),
.Y(n_16606)
);

INVx1_ASAP7_75t_L g16607 ( 
.A(n_15718),
.Y(n_16607)
);

INVx1_ASAP7_75t_L g16608 ( 
.A(n_16015),
.Y(n_16608)
);

AND2x2_ASAP7_75t_L g16609 ( 
.A(n_15925),
.B(n_8804),
.Y(n_16609)
);

OAI211xp5_ASAP7_75t_L g16610 ( 
.A1(n_15658),
.A2(n_9473),
.B(n_9614),
.C(n_9369),
.Y(n_16610)
);

INVx1_ASAP7_75t_L g16611 ( 
.A(n_16018),
.Y(n_16611)
);

INVx1_ASAP7_75t_L g16612 ( 
.A(n_15981),
.Y(n_16612)
);

CKINVDCx14_ASAP7_75t_R g16613 ( 
.A(n_16071),
.Y(n_16613)
);

AND2x2_ASAP7_75t_L g16614 ( 
.A(n_15926),
.B(n_8804),
.Y(n_16614)
);

INVx1_ASAP7_75t_L g16615 ( 
.A(n_15881),
.Y(n_16615)
);

OR2x2_ASAP7_75t_L g16616 ( 
.A(n_16059),
.B(n_8999),
.Y(n_16616)
);

INVx2_ASAP7_75t_L g16617 ( 
.A(n_16043),
.Y(n_16617)
);

AND2x4_ASAP7_75t_L g16618 ( 
.A(n_15942),
.B(n_8804),
.Y(n_16618)
);

INVx1_ASAP7_75t_SL g16619 ( 
.A(n_15740),
.Y(n_16619)
);

NAND2x1_ASAP7_75t_SL g16620 ( 
.A(n_15996),
.B(n_9470),
.Y(n_16620)
);

AND2x4_ASAP7_75t_L g16621 ( 
.A(n_15958),
.B(n_11774),
.Y(n_16621)
);

AND2x4_ASAP7_75t_L g16622 ( 
.A(n_15977),
.B(n_11774),
.Y(n_16622)
);

INVx2_ASAP7_75t_L g16623 ( 
.A(n_16041),
.Y(n_16623)
);

AND2x2_ASAP7_75t_L g16624 ( 
.A(n_15927),
.B(n_8804),
.Y(n_16624)
);

AND2x2_ASAP7_75t_L g16625 ( 
.A(n_15932),
.B(n_8804),
.Y(n_16625)
);

OR2x2_ASAP7_75t_L g16626 ( 
.A(n_16047),
.B(n_15922),
.Y(n_16626)
);

OR2x2_ASAP7_75t_L g16627 ( 
.A(n_15709),
.B(n_8055),
.Y(n_16627)
);

INVx1_ASAP7_75t_L g16628 ( 
.A(n_15882),
.Y(n_16628)
);

AND2x2_ASAP7_75t_L g16629 ( 
.A(n_15948),
.B(n_15971),
.Y(n_16629)
);

NAND2xp5_ASAP7_75t_L g16630 ( 
.A(n_16028),
.B(n_15962),
.Y(n_16630)
);

INVx2_ASAP7_75t_L g16631 ( 
.A(n_15963),
.Y(n_16631)
);

INVx1_ASAP7_75t_L g16632 ( 
.A(n_15723),
.Y(n_16632)
);

INVx1_ASAP7_75t_L g16633 ( 
.A(n_15860),
.Y(n_16633)
);

AND2x2_ASAP7_75t_L g16634 ( 
.A(n_15976),
.B(n_8824),
.Y(n_16634)
);

AND2x2_ASAP7_75t_L g16635 ( 
.A(n_15656),
.B(n_8824),
.Y(n_16635)
);

INVx2_ASAP7_75t_L g16636 ( 
.A(n_15998),
.Y(n_16636)
);

OAI221xp5_ASAP7_75t_SL g16637 ( 
.A1(n_15761),
.A2(n_10589),
.B1(n_10598),
.B2(n_10587),
.C(n_10565),
.Y(n_16637)
);

AND2x2_ASAP7_75t_L g16638 ( 
.A(n_15979),
.B(n_8824),
.Y(n_16638)
);

AND2x4_ASAP7_75t_L g16639 ( 
.A(n_15983),
.B(n_11794),
.Y(n_16639)
);

AND2x2_ASAP7_75t_L g16640 ( 
.A(n_16077),
.B(n_15896),
.Y(n_16640)
);

AND2x2_ASAP7_75t_L g16641 ( 
.A(n_15657),
.B(n_8824),
.Y(n_16641)
);

NOR2x1_ASAP7_75t_SL g16642 ( 
.A(n_16003),
.B(n_8481),
.Y(n_16642)
);

OR2x2_ASAP7_75t_L g16643 ( 
.A(n_15758),
.B(n_8055),
.Y(n_16643)
);

INVx1_ASAP7_75t_L g16644 ( 
.A(n_15864),
.Y(n_16644)
);

NAND2xp5_ASAP7_75t_L g16645 ( 
.A(n_16006),
.B(n_10391),
.Y(n_16645)
);

NAND2xp5_ASAP7_75t_L g16646 ( 
.A(n_15855),
.B(n_10391),
.Y(n_16646)
);

NAND2xp5_ASAP7_75t_L g16647 ( 
.A(n_15862),
.B(n_10417),
.Y(n_16647)
);

INVxp67_ASAP7_75t_L g16648 ( 
.A(n_15841),
.Y(n_16648)
);

NAND2xp5_ASAP7_75t_L g16649 ( 
.A(n_15866),
.B(n_10417),
.Y(n_16649)
);

AND2x2_ASAP7_75t_L g16650 ( 
.A(n_16053),
.B(n_8824),
.Y(n_16650)
);

INVx2_ASAP7_75t_L g16651 ( 
.A(n_15756),
.Y(n_16651)
);

INVx1_ASAP7_75t_L g16652 ( 
.A(n_15947),
.Y(n_16652)
);

BUFx2_ASAP7_75t_L g16653 ( 
.A(n_15951),
.Y(n_16653)
);

HB1xp67_ASAP7_75t_L g16654 ( 
.A(n_15949),
.Y(n_16654)
);

INVx1_ASAP7_75t_SL g16655 ( 
.A(n_15909),
.Y(n_16655)
);

AND2x2_ASAP7_75t_L g16656 ( 
.A(n_16066),
.B(n_8824),
.Y(n_16656)
);

AND2x2_ASAP7_75t_L g16657 ( 
.A(n_15868),
.B(n_8844),
.Y(n_16657)
);

INVx1_ASAP7_75t_L g16658 ( 
.A(n_15839),
.Y(n_16658)
);

INVx1_ASAP7_75t_L g16659 ( 
.A(n_16385),
.Y(n_16659)
);

NAND4xp25_ASAP7_75t_L g16660 ( 
.A(n_16127),
.B(n_15904),
.C(n_15823),
.D(n_15911),
.Y(n_16660)
);

OR2x2_ASAP7_75t_L g16661 ( 
.A(n_16103),
.B(n_16072),
.Y(n_16661)
);

AND2x2_ASAP7_75t_L g16662 ( 
.A(n_16117),
.B(n_15985),
.Y(n_16662)
);

AOI21xp33_ASAP7_75t_L g16663 ( 
.A1(n_16277),
.A2(n_15701),
.B(n_16030),
.Y(n_16663)
);

INVx1_ASAP7_75t_L g16664 ( 
.A(n_16385),
.Y(n_16664)
);

INVx1_ASAP7_75t_L g16665 ( 
.A(n_16097),
.Y(n_16665)
);

NAND2xp5_ASAP7_75t_L g16666 ( 
.A(n_16252),
.B(n_15986),
.Y(n_16666)
);

INVx1_ASAP7_75t_L g16667 ( 
.A(n_16097),
.Y(n_16667)
);

NOR2xp67_ASAP7_75t_L g16668 ( 
.A(n_16350),
.B(n_16032),
.Y(n_16668)
);

INVx1_ASAP7_75t_L g16669 ( 
.A(n_16195),
.Y(n_16669)
);

AOI22xp33_ASAP7_75t_L g16670 ( 
.A1(n_16333),
.A2(n_16019),
.B1(n_16083),
.B2(n_15920),
.Y(n_16670)
);

INVx1_ASAP7_75t_L g16671 ( 
.A(n_16203),
.Y(n_16671)
);

AND2x4_ASAP7_75t_L g16672 ( 
.A(n_16346),
.B(n_16149),
.Y(n_16672)
);

INVx1_ASAP7_75t_L g16673 ( 
.A(n_16096),
.Y(n_16673)
);

NAND2xp5_ASAP7_75t_L g16674 ( 
.A(n_16126),
.B(n_15987),
.Y(n_16674)
);

HB1xp67_ASAP7_75t_L g16675 ( 
.A(n_16350),
.Y(n_16675)
);

INVx1_ASAP7_75t_SL g16676 ( 
.A(n_16112),
.Y(n_16676)
);

AND2x2_ASAP7_75t_L g16677 ( 
.A(n_16172),
.B(n_15994),
.Y(n_16677)
);

NOR2xp33_ASAP7_75t_L g16678 ( 
.A(n_16541),
.B(n_15995),
.Y(n_16678)
);

BUFx2_ASAP7_75t_L g16679 ( 
.A(n_16141),
.Y(n_16679)
);

INVx4_ASAP7_75t_L g16680 ( 
.A(n_16350),
.Y(n_16680)
);

NOR2x1_ASAP7_75t_L g16681 ( 
.A(n_16132),
.B(n_15999),
.Y(n_16681)
);

INVx1_ASAP7_75t_L g16682 ( 
.A(n_16320),
.Y(n_16682)
);

AND2x4_ASAP7_75t_L g16683 ( 
.A(n_16282),
.B(n_16031),
.Y(n_16683)
);

INVx2_ASAP7_75t_L g16684 ( 
.A(n_16130),
.Y(n_16684)
);

OR2x2_ASAP7_75t_L g16685 ( 
.A(n_16118),
.B(n_16080),
.Y(n_16685)
);

NAND2xp5_ASAP7_75t_L g16686 ( 
.A(n_16145),
.B(n_16046),
.Y(n_16686)
);

AND2x2_ASAP7_75t_L g16687 ( 
.A(n_16217),
.B(n_16049),
.Y(n_16687)
);

NAND2xp5_ASAP7_75t_L g16688 ( 
.A(n_16342),
.B(n_16060),
.Y(n_16688)
);

AND2x2_ASAP7_75t_L g16689 ( 
.A(n_16189),
.B(n_16061),
.Y(n_16689)
);

INVx1_ASAP7_75t_L g16690 ( 
.A(n_16316),
.Y(n_16690)
);

INVx1_ASAP7_75t_L g16691 ( 
.A(n_16170),
.Y(n_16691)
);

AND2x2_ASAP7_75t_L g16692 ( 
.A(n_16184),
.B(n_16386),
.Y(n_16692)
);

BUFx2_ASAP7_75t_L g16693 ( 
.A(n_16256),
.Y(n_16693)
);

INVxp67_ASAP7_75t_L g16694 ( 
.A(n_16279),
.Y(n_16694)
);

AND2x2_ASAP7_75t_L g16695 ( 
.A(n_16175),
.B(n_16098),
.Y(n_16695)
);

AND2x2_ASAP7_75t_L g16696 ( 
.A(n_16181),
.B(n_16186),
.Y(n_16696)
);

INVx1_ASAP7_75t_SL g16697 ( 
.A(n_16242),
.Y(n_16697)
);

NOR2xp67_ASAP7_75t_L g16698 ( 
.A(n_16099),
.B(n_16035),
.Y(n_16698)
);

INVx1_ASAP7_75t_L g16699 ( 
.A(n_16100),
.Y(n_16699)
);

AND2x2_ASAP7_75t_L g16700 ( 
.A(n_16162),
.B(n_16070),
.Y(n_16700)
);

NAND2xp5_ASAP7_75t_L g16701 ( 
.A(n_16315),
.B(n_16095),
.Y(n_16701)
);

AND2x2_ASAP7_75t_L g16702 ( 
.A(n_16179),
.B(n_16058),
.Y(n_16702)
);

AOI22xp33_ASAP7_75t_L g16703 ( 
.A1(n_16226),
.A2(n_16045),
.B1(n_16051),
.B2(n_16048),
.Y(n_16703)
);

NAND2xp5_ASAP7_75t_L g16704 ( 
.A(n_16247),
.B(n_16271),
.Y(n_16704)
);

NAND2x1p5_ASAP7_75t_L g16705 ( 
.A(n_16311),
.B(n_16069),
.Y(n_16705)
);

INVx1_ASAP7_75t_L g16706 ( 
.A(n_16440),
.Y(n_16706)
);

BUFx3_ASAP7_75t_L g16707 ( 
.A(n_16202),
.Y(n_16707)
);

AND2x2_ASAP7_75t_L g16708 ( 
.A(n_16160),
.B(n_16081),
.Y(n_16708)
);

NAND2xp5_ASAP7_75t_L g16709 ( 
.A(n_16114),
.B(n_15967),
.Y(n_16709)
);

AND2x2_ASAP7_75t_L g16710 ( 
.A(n_16167),
.B(n_16171),
.Y(n_16710)
);

INVx3_ASAP7_75t_L g16711 ( 
.A(n_16134),
.Y(n_16711)
);

NAND2xp5_ASAP7_75t_L g16712 ( 
.A(n_16239),
.B(n_15991),
.Y(n_16712)
);

HB1xp67_ASAP7_75t_L g16713 ( 
.A(n_16289),
.Y(n_16713)
);

AND2x2_ASAP7_75t_L g16714 ( 
.A(n_16111),
.B(n_16088),
.Y(n_16714)
);

INVx1_ASAP7_75t_L g16715 ( 
.A(n_16464),
.Y(n_16715)
);

NOR2xp33_ASAP7_75t_L g16716 ( 
.A(n_16278),
.B(n_16008),
.Y(n_16716)
);

AND2x2_ASAP7_75t_L g16717 ( 
.A(n_16123),
.B(n_16089),
.Y(n_16717)
);

AND2x2_ASAP7_75t_L g16718 ( 
.A(n_16206),
.B(n_16221),
.Y(n_16718)
);

INVx1_ASAP7_75t_L g16719 ( 
.A(n_16540),
.Y(n_16719)
);

INVx1_ASAP7_75t_L g16720 ( 
.A(n_16475),
.Y(n_16720)
);

AND2x2_ASAP7_75t_L g16721 ( 
.A(n_16168),
.B(n_15997),
.Y(n_16721)
);

AND2x4_ASAP7_75t_L g16722 ( 
.A(n_16192),
.B(n_16004),
.Y(n_16722)
);

AND2x2_ASAP7_75t_L g16723 ( 
.A(n_16177),
.B(n_16022),
.Y(n_16723)
);

CKINVDCx5p33_ASAP7_75t_R g16724 ( 
.A(n_16148),
.Y(n_16724)
);

AND2x2_ASAP7_75t_L g16725 ( 
.A(n_16131),
.B(n_16079),
.Y(n_16725)
);

AND2x2_ASAP7_75t_L g16726 ( 
.A(n_16122),
.B(n_16027),
.Y(n_16726)
);

INVx1_ASAP7_75t_SL g16727 ( 
.A(n_16532),
.Y(n_16727)
);

HB1xp67_ASAP7_75t_L g16728 ( 
.A(n_16210),
.Y(n_16728)
);

AND2x4_ASAP7_75t_L g16729 ( 
.A(n_16150),
.B(n_16016),
.Y(n_16729)
);

INVx1_ASAP7_75t_L g16730 ( 
.A(n_16535),
.Y(n_16730)
);

AND2x2_ASAP7_75t_L g16731 ( 
.A(n_16487),
.B(n_16064),
.Y(n_16731)
);

AND2x2_ASAP7_75t_L g16732 ( 
.A(n_16579),
.B(n_16084),
.Y(n_16732)
);

INVx2_ASAP7_75t_L g16733 ( 
.A(n_16377),
.Y(n_16733)
);

AOI22xp33_ASAP7_75t_L g16734 ( 
.A1(n_16494),
.A2(n_16324),
.B1(n_16154),
.B2(n_16363),
.Y(n_16734)
);

AND2x2_ASAP7_75t_L g16735 ( 
.A(n_16113),
.B(n_16084),
.Y(n_16735)
);

AND2x2_ASAP7_75t_L g16736 ( 
.A(n_16374),
.B(n_16056),
.Y(n_16736)
);

NOR2xp33_ASAP7_75t_L g16737 ( 
.A(n_16531),
.B(n_16056),
.Y(n_16737)
);

OAI21xp5_ASAP7_75t_L g16738 ( 
.A1(n_16274),
.A2(n_15660),
.B(n_10755),
.Y(n_16738)
);

INVx1_ASAP7_75t_L g16739 ( 
.A(n_16435),
.Y(n_16739)
);

AND2x2_ASAP7_75t_L g16740 ( 
.A(n_16107),
.B(n_8844),
.Y(n_16740)
);

INVxp67_ASAP7_75t_SL g16741 ( 
.A(n_16426),
.Y(n_16741)
);

INVx1_ASAP7_75t_L g16742 ( 
.A(n_16571),
.Y(n_16742)
);

INVx1_ASAP7_75t_L g16743 ( 
.A(n_16591),
.Y(n_16743)
);

OR2x2_ASAP7_75t_L g16744 ( 
.A(n_16208),
.B(n_8065),
.Y(n_16744)
);

A2O1A1Ixp33_ASAP7_75t_L g16745 ( 
.A1(n_16237),
.A2(n_11046),
.B(n_11067),
.C(n_10783),
.Y(n_16745)
);

INVx2_ASAP7_75t_SL g16746 ( 
.A(n_16178),
.Y(n_16746)
);

NAND5xp2_ASAP7_75t_L g16747 ( 
.A(n_16245),
.B(n_9209),
.C(n_7984),
.D(n_8007),
.E(n_8002),
.Y(n_16747)
);

NOR2xp33_ASAP7_75t_L g16748 ( 
.A(n_16476),
.B(n_8481),
.Y(n_16748)
);

AND2x2_ASAP7_75t_L g16749 ( 
.A(n_16559),
.B(n_8844),
.Y(n_16749)
);

OR2x2_ASAP7_75t_L g16750 ( 
.A(n_16119),
.B(n_8065),
.Y(n_16750)
);

INVx5_ASAP7_75t_L g16751 ( 
.A(n_16514),
.Y(n_16751)
);

AOI22xp5_ASAP7_75t_L g16752 ( 
.A1(n_16468),
.A2(n_8608),
.B1(n_8639),
.B2(n_8492),
.Y(n_16752)
);

INVx1_ASAP7_75t_L g16753 ( 
.A(n_16381),
.Y(n_16753)
);

AND2x2_ASAP7_75t_L g16754 ( 
.A(n_16578),
.B(n_8844),
.Y(n_16754)
);

NAND2xp5_ASAP7_75t_L g16755 ( 
.A(n_16129),
.B(n_10418),
.Y(n_16755)
);

INVx1_ASAP7_75t_L g16756 ( 
.A(n_16156),
.Y(n_16756)
);

INVx1_ASAP7_75t_L g16757 ( 
.A(n_16419),
.Y(n_16757)
);

NAND2xp5_ASAP7_75t_L g16758 ( 
.A(n_16135),
.B(n_10418),
.Y(n_16758)
);

AND2x2_ASAP7_75t_L g16759 ( 
.A(n_16104),
.B(n_8844),
.Y(n_16759)
);

INVx2_ASAP7_75t_L g16760 ( 
.A(n_16140),
.Y(n_16760)
);

AOI221xp5_ASAP7_75t_L g16761 ( 
.A1(n_16602),
.A2(n_10589),
.B1(n_10598),
.B2(n_10587),
.C(n_10565),
.Y(n_16761)
);

NAND2x1p5_ASAP7_75t_L g16762 ( 
.A(n_16619),
.B(n_8492),
.Y(n_16762)
);

INVx1_ASAP7_75t_L g16763 ( 
.A(n_16431),
.Y(n_16763)
);

AND2x2_ASAP7_75t_L g16764 ( 
.A(n_16496),
.B(n_8844),
.Y(n_16764)
);

INVx1_ASAP7_75t_SL g16765 ( 
.A(n_16430),
.Y(n_16765)
);

AND2x2_ASAP7_75t_L g16766 ( 
.A(n_16367),
.B(n_8894),
.Y(n_16766)
);

INVx1_ASAP7_75t_SL g16767 ( 
.A(n_16371),
.Y(n_16767)
);

INVx2_ASAP7_75t_L g16768 ( 
.A(n_16138),
.Y(n_16768)
);

BUFx3_ASAP7_75t_L g16769 ( 
.A(n_16305),
.Y(n_16769)
);

NAND2x1_ASAP7_75t_L g16770 ( 
.A(n_16166),
.B(n_11097),
.Y(n_16770)
);

INVx1_ASAP7_75t_L g16771 ( 
.A(n_16230),
.Y(n_16771)
);

NAND2xp5_ASAP7_75t_L g16772 ( 
.A(n_16137),
.B(n_16233),
.Y(n_16772)
);

HB1xp67_ASAP7_75t_L g16773 ( 
.A(n_16364),
.Y(n_16773)
);

AND2x2_ASAP7_75t_L g16774 ( 
.A(n_16136),
.B(n_8894),
.Y(n_16774)
);

NAND2xp5_ASAP7_75t_L g16775 ( 
.A(n_16445),
.B(n_16173),
.Y(n_16775)
);

OR2x2_ASAP7_75t_L g16776 ( 
.A(n_16125),
.B(n_9262),
.Y(n_16776)
);

AND2x2_ASAP7_75t_L g16777 ( 
.A(n_16349),
.B(n_8894),
.Y(n_16777)
);

AND2x2_ASAP7_75t_L g16778 ( 
.A(n_16183),
.B(n_8894),
.Y(n_16778)
);

NOR2xp33_ASAP7_75t_L g16779 ( 
.A(n_16204),
.B(n_8492),
.Y(n_16779)
);

OR2x2_ASAP7_75t_L g16780 ( 
.A(n_16219),
.B(n_9262),
.Y(n_16780)
);

INVx2_ASAP7_75t_L g16781 ( 
.A(n_16620),
.Y(n_16781)
);

AND2x4_ASAP7_75t_L g16782 ( 
.A(n_16182),
.B(n_8894),
.Y(n_16782)
);

OR2x2_ASAP7_75t_L g16783 ( 
.A(n_16146),
.B(n_10291),
.Y(n_16783)
);

AND2x2_ASAP7_75t_L g16784 ( 
.A(n_16428),
.B(n_8894),
.Y(n_16784)
);

INVx1_ASAP7_75t_L g16785 ( 
.A(n_16395),
.Y(n_16785)
);

OR2x2_ASAP7_75t_L g16786 ( 
.A(n_16174),
.B(n_9113),
.Y(n_16786)
);

INVx1_ASAP7_75t_L g16787 ( 
.A(n_16398),
.Y(n_16787)
);

OR2x2_ASAP7_75t_L g16788 ( 
.A(n_16142),
.B(n_9113),
.Y(n_16788)
);

BUFx3_ASAP7_75t_L g16789 ( 
.A(n_16312),
.Y(n_16789)
);

INVx1_ASAP7_75t_L g16790 ( 
.A(n_16416),
.Y(n_16790)
);

AOI22xp5_ASAP7_75t_L g16791 ( 
.A1(n_16613),
.A2(n_8608),
.B1(n_8639),
.B2(n_8492),
.Y(n_16791)
);

INVx1_ASAP7_75t_L g16792 ( 
.A(n_16418),
.Y(n_16792)
);

AND2x2_ASAP7_75t_L g16793 ( 
.A(n_16211),
.B(n_16238),
.Y(n_16793)
);

OR2x2_ASAP7_75t_L g16794 ( 
.A(n_16153),
.B(n_11101),
.Y(n_16794)
);

INVx2_ASAP7_75t_L g16795 ( 
.A(n_16642),
.Y(n_16795)
);

INVx1_ASAP7_75t_L g16796 ( 
.A(n_16564),
.Y(n_16796)
);

AND2x2_ASAP7_75t_L g16797 ( 
.A(n_16155),
.B(n_8910),
.Y(n_16797)
);

INVx2_ASAP7_75t_L g16798 ( 
.A(n_16283),
.Y(n_16798)
);

AND2x2_ASAP7_75t_L g16799 ( 
.A(n_16554),
.B(n_8910),
.Y(n_16799)
);

OR2x2_ASAP7_75t_L g16800 ( 
.A(n_16159),
.B(n_11101),
.Y(n_16800)
);

INVx2_ASAP7_75t_L g16801 ( 
.A(n_16109),
.Y(n_16801)
);

NAND3xp33_ASAP7_75t_L g16802 ( 
.A(n_16105),
.B(n_9614),
.C(n_9369),
.Y(n_16802)
);

AND2x2_ASAP7_75t_L g16803 ( 
.A(n_16570),
.B(n_8910),
.Y(n_16803)
);

AND2x2_ASAP7_75t_L g16804 ( 
.A(n_16300),
.B(n_8910),
.Y(n_16804)
);

INVx1_ASAP7_75t_L g16805 ( 
.A(n_16345),
.Y(n_16805)
);

NAND5xp2_ASAP7_75t_SL g16806 ( 
.A(n_16420),
.B(n_8564),
.C(n_8490),
.D(n_8567),
.E(n_8520),
.Y(n_16806)
);

INVx2_ASAP7_75t_SL g16807 ( 
.A(n_16265),
.Y(n_16807)
);

INVx2_ASAP7_75t_L g16808 ( 
.A(n_16412),
.Y(n_16808)
);

INVx2_ASAP7_75t_L g16809 ( 
.A(n_16267),
.Y(n_16809)
);

AND2x2_ASAP7_75t_L g16810 ( 
.A(n_16218),
.B(n_8910),
.Y(n_16810)
);

NAND4xp25_ASAP7_75t_L g16811 ( 
.A(n_16236),
.B(n_7837),
.C(n_7851),
.D(n_7806),
.Y(n_16811)
);

NAND2xp5_ASAP7_75t_L g16812 ( 
.A(n_16161),
.B(n_10419),
.Y(n_16812)
);

NAND2xp5_ASAP7_75t_L g16813 ( 
.A(n_16165),
.B(n_10419),
.Y(n_16813)
);

AND2x2_ASAP7_75t_L g16814 ( 
.A(n_16190),
.B(n_8910),
.Y(n_16814)
);

NAND2xp5_ASAP7_75t_L g16815 ( 
.A(n_16164),
.B(n_10426),
.Y(n_16815)
);

INVx2_ASAP7_75t_L g16816 ( 
.A(n_16270),
.Y(n_16816)
);

INVx1_ASAP7_75t_L g16817 ( 
.A(n_16106),
.Y(n_16817)
);

AND2x2_ASAP7_75t_L g16818 ( 
.A(n_16133),
.B(n_9026),
.Y(n_16818)
);

AOI22xp33_ASAP7_75t_L g16819 ( 
.A1(n_16383),
.A2(n_8608),
.B1(n_8639),
.B2(n_8492),
.Y(n_16819)
);

OR2x2_ASAP7_75t_L g16820 ( 
.A(n_16158),
.B(n_11108),
.Y(n_16820)
);

INVx2_ASAP7_75t_L g16821 ( 
.A(n_16164),
.Y(n_16821)
);

AOI221xp5_ASAP7_75t_L g16822 ( 
.A1(n_16102),
.A2(n_10598),
.B1(n_10599),
.B2(n_10589),
.C(n_10587),
.Y(n_16822)
);

INVx1_ASAP7_75t_L g16823 ( 
.A(n_16147),
.Y(n_16823)
);

INVx1_ASAP7_75t_L g16824 ( 
.A(n_16263),
.Y(n_16824)
);

BUFx2_ASAP7_75t_L g16825 ( 
.A(n_16654),
.Y(n_16825)
);

BUFx2_ASAP7_75t_L g16826 ( 
.A(n_16272),
.Y(n_16826)
);

NAND2xp5_ASAP7_75t_L g16827 ( 
.A(n_16296),
.B(n_10426),
.Y(n_16827)
);

NAND2xp5_ASAP7_75t_L g16828 ( 
.A(n_16396),
.B(n_10430),
.Y(n_16828)
);

HB1xp67_ASAP7_75t_L g16829 ( 
.A(n_16514),
.Y(n_16829)
);

HB1xp67_ASAP7_75t_L g16830 ( 
.A(n_16313),
.Y(n_16830)
);

AND2x2_ASAP7_75t_L g16831 ( 
.A(n_16235),
.B(n_9026),
.Y(n_16831)
);

OR2x2_ASAP7_75t_L g16832 ( 
.A(n_16157),
.B(n_11108),
.Y(n_16832)
);

NAND2x1_ASAP7_75t_L g16833 ( 
.A(n_16309),
.B(n_16259),
.Y(n_16833)
);

INVx2_ASAP7_75t_L g16834 ( 
.A(n_16207),
.Y(n_16834)
);

NAND2xp5_ASAP7_75t_L g16835 ( 
.A(n_16209),
.B(n_10430),
.Y(n_16835)
);

OR2x2_ASAP7_75t_L g16836 ( 
.A(n_16215),
.B(n_11110),
.Y(n_16836)
);

HB1xp67_ASAP7_75t_L g16837 ( 
.A(n_16232),
.Y(n_16837)
);

AND2x2_ASAP7_75t_L g16838 ( 
.A(n_16380),
.B(n_16199),
.Y(n_16838)
);

INVx1_ASAP7_75t_L g16839 ( 
.A(n_16197),
.Y(n_16839)
);

INVx1_ASAP7_75t_L g16840 ( 
.A(n_16198),
.Y(n_16840)
);

NOR2x1_ASAP7_75t_L g16841 ( 
.A(n_16231),
.B(n_11110),
.Y(n_16841)
);

INVxp67_ASAP7_75t_L g16842 ( 
.A(n_16629),
.Y(n_16842)
);

AND2x2_ASAP7_75t_L g16843 ( 
.A(n_16391),
.B(n_9026),
.Y(n_16843)
);

AND2x2_ASAP7_75t_L g16844 ( 
.A(n_16432),
.B(n_16455),
.Y(n_16844)
);

INVx1_ASAP7_75t_SL g16845 ( 
.A(n_16101),
.Y(n_16845)
);

CKINVDCx16_ASAP7_75t_R g16846 ( 
.A(n_16585),
.Y(n_16846)
);

NAND2xp5_ASAP7_75t_L g16847 ( 
.A(n_16214),
.B(n_10432),
.Y(n_16847)
);

NAND2xp5_ASAP7_75t_L g16848 ( 
.A(n_16241),
.B(n_10432),
.Y(n_16848)
);

INVxp67_ASAP7_75t_L g16849 ( 
.A(n_16653),
.Y(n_16849)
);

OR2x2_ASAP7_75t_L g16850 ( 
.A(n_16223),
.B(n_11111),
.Y(n_16850)
);

NAND2xp5_ASAP7_75t_L g16851 ( 
.A(n_16254),
.B(n_10433),
.Y(n_16851)
);

INVx1_ASAP7_75t_SL g16852 ( 
.A(n_16406),
.Y(n_16852)
);

INVx1_ASAP7_75t_L g16853 ( 
.A(n_16163),
.Y(n_16853)
);

NAND3xp33_ASAP7_75t_L g16854 ( 
.A(n_16176),
.B(n_9614),
.C(n_11111),
.Y(n_16854)
);

NAND2xp5_ASAP7_75t_L g16855 ( 
.A(n_16185),
.B(n_10433),
.Y(n_16855)
);

NOR2x1_ASAP7_75t_SL g16856 ( 
.A(n_16388),
.B(n_8492),
.Y(n_16856)
);

INVx1_ASAP7_75t_L g16857 ( 
.A(n_16120),
.Y(n_16857)
);

BUFx2_ASAP7_75t_L g16858 ( 
.A(n_16653),
.Y(n_16858)
);

INVx1_ASAP7_75t_SL g16859 ( 
.A(n_16234),
.Y(n_16859)
);

INVx1_ASAP7_75t_L g16860 ( 
.A(n_16121),
.Y(n_16860)
);

INVx3_ASAP7_75t_L g16861 ( 
.A(n_16334),
.Y(n_16861)
);

AOI22xp33_ASAP7_75t_L g16862 ( 
.A1(n_16375),
.A2(n_8608),
.B1(n_8639),
.B2(n_8492),
.Y(n_16862)
);

INVx1_ASAP7_75t_L g16863 ( 
.A(n_16110),
.Y(n_16863)
);

AND2x4_ASAP7_75t_L g16864 ( 
.A(n_16544),
.B(n_9026),
.Y(n_16864)
);

INVx1_ASAP7_75t_L g16865 ( 
.A(n_16246),
.Y(n_16865)
);

INVx2_ASAP7_75t_L g16866 ( 
.A(n_16552),
.Y(n_16866)
);

INVx2_ASAP7_75t_SL g16867 ( 
.A(n_16410),
.Y(n_16867)
);

NAND2xp5_ASAP7_75t_SL g16868 ( 
.A(n_16303),
.B(n_8492),
.Y(n_16868)
);

INVx2_ASAP7_75t_L g16869 ( 
.A(n_16557),
.Y(n_16869)
);

AND2x2_ASAP7_75t_L g16870 ( 
.A(n_16595),
.B(n_9026),
.Y(n_16870)
);

INVx1_ASAP7_75t_L g16871 ( 
.A(n_16108),
.Y(n_16871)
);

OR2x2_ASAP7_75t_L g16872 ( 
.A(n_16483),
.B(n_16451),
.Y(n_16872)
);

INVx1_ASAP7_75t_L g16873 ( 
.A(n_16116),
.Y(n_16873)
);

AND2x2_ASAP7_75t_L g16874 ( 
.A(n_16492),
.B(n_16499),
.Y(n_16874)
);

INVx1_ASAP7_75t_L g16875 ( 
.A(n_16243),
.Y(n_16875)
);

AND2x2_ASAP7_75t_L g16876 ( 
.A(n_16524),
.B(n_9026),
.Y(n_16876)
);

AND2x4_ASAP7_75t_L g16877 ( 
.A(n_16617),
.B(n_9075),
.Y(n_16877)
);

OR2x2_ASAP7_75t_L g16878 ( 
.A(n_16504),
.B(n_11121),
.Y(n_16878)
);

INVx2_ASAP7_75t_L g16879 ( 
.A(n_16291),
.Y(n_16879)
);

OR2x2_ASAP7_75t_L g16880 ( 
.A(n_16515),
.B(n_11121),
.Y(n_16880)
);

AND2x2_ASAP7_75t_L g16881 ( 
.A(n_16341),
.B(n_9075),
.Y(n_16881)
);

AND2x2_ASAP7_75t_L g16882 ( 
.A(n_16326),
.B(n_9075),
.Y(n_16882)
);

AND2x2_ASAP7_75t_L g16883 ( 
.A(n_16212),
.B(n_16216),
.Y(n_16883)
);

AND2x2_ASAP7_75t_L g16884 ( 
.A(n_16240),
.B(n_9075),
.Y(n_16884)
);

OR2x2_ASAP7_75t_L g16885 ( 
.A(n_16516),
.B(n_11139),
.Y(n_16885)
);

OR2x2_ASAP7_75t_L g16886 ( 
.A(n_16517),
.B(n_11139),
.Y(n_16886)
);

INVx5_ASAP7_75t_L g16887 ( 
.A(n_16512),
.Y(n_16887)
);

INVx1_ASAP7_75t_SL g16888 ( 
.A(n_16655),
.Y(n_16888)
);

AND2x2_ASAP7_75t_L g16889 ( 
.A(n_16260),
.B(n_9075),
.Y(n_16889)
);

INVx2_ASAP7_75t_L g16890 ( 
.A(n_16424),
.Y(n_16890)
);

OR2x2_ASAP7_75t_L g16891 ( 
.A(n_16523),
.B(n_11151),
.Y(n_16891)
);

INVx1_ASAP7_75t_L g16892 ( 
.A(n_16249),
.Y(n_16892)
);

AND2x2_ASAP7_75t_L g16893 ( 
.A(n_16318),
.B(n_16332),
.Y(n_16893)
);

OR2x6_ASAP7_75t_L g16894 ( 
.A(n_16469),
.B(n_7806),
.Y(n_16894)
);

AND2x2_ASAP7_75t_L g16895 ( 
.A(n_16361),
.B(n_9075),
.Y(n_16895)
);

INVx1_ASAP7_75t_L g16896 ( 
.A(n_16250),
.Y(n_16896)
);

AND2x4_ASAP7_75t_L g16897 ( 
.A(n_16527),
.B(n_9078),
.Y(n_16897)
);

INVx1_ASAP7_75t_L g16898 ( 
.A(n_16264),
.Y(n_16898)
);

OR2x2_ASAP7_75t_L g16899 ( 
.A(n_16529),
.B(n_11151),
.Y(n_16899)
);

NAND2x1_ASAP7_75t_L g16900 ( 
.A(n_16583),
.B(n_11160),
.Y(n_16900)
);

AOI21xp5_ASAP7_75t_L g16901 ( 
.A1(n_16338),
.A2(n_11173),
.B(n_11160),
.Y(n_16901)
);

AND2x2_ASAP7_75t_L g16902 ( 
.A(n_16362),
.B(n_9078),
.Y(n_16902)
);

OR2x2_ASAP7_75t_L g16903 ( 
.A(n_16268),
.B(n_11173),
.Y(n_16903)
);

OR2x2_ASAP7_75t_L g16904 ( 
.A(n_16269),
.B(n_11192),
.Y(n_16904)
);

OR2x2_ASAP7_75t_L g16905 ( 
.A(n_16273),
.B(n_11192),
.Y(n_16905)
);

INVx1_ASAP7_75t_L g16906 ( 
.A(n_16193),
.Y(n_16906)
);

BUFx3_ASAP7_75t_L g16907 ( 
.A(n_16409),
.Y(n_16907)
);

INVx2_ASAP7_75t_L g16908 ( 
.A(n_16308),
.Y(n_16908)
);

INVx1_ASAP7_75t_L g16909 ( 
.A(n_16201),
.Y(n_16909)
);

OR2x2_ASAP7_75t_L g16910 ( 
.A(n_16287),
.B(n_11205),
.Y(n_16910)
);

BUFx2_ASAP7_75t_L g16911 ( 
.A(n_16623),
.Y(n_16911)
);

NAND2xp5_ASAP7_75t_L g16912 ( 
.A(n_16213),
.B(n_16220),
.Y(n_16912)
);

BUFx3_ASAP7_75t_L g16913 ( 
.A(n_16411),
.Y(n_16913)
);

INVx1_ASAP7_75t_L g16914 ( 
.A(n_16224),
.Y(n_16914)
);

INVx1_ASAP7_75t_L g16915 ( 
.A(n_16227),
.Y(n_16915)
);

INVx1_ASAP7_75t_L g16916 ( 
.A(n_16229),
.Y(n_16916)
);

AND2x2_ASAP7_75t_L g16917 ( 
.A(n_16403),
.B(n_9078),
.Y(n_16917)
);

CKINVDCx5p33_ASAP7_75t_R g16918 ( 
.A(n_16382),
.Y(n_16918)
);

AND2x2_ASAP7_75t_L g16919 ( 
.A(n_16152),
.B(n_9078),
.Y(n_16919)
);

INVx6_ASAP7_75t_L g16920 ( 
.A(n_16196),
.Y(n_16920)
);

INVx1_ASAP7_75t_L g16921 ( 
.A(n_16244),
.Y(n_16921)
);

OR2x2_ASAP7_75t_L g16922 ( 
.A(n_16413),
.B(n_11205),
.Y(n_16922)
);

NAND2xp5_ASAP7_75t_L g16923 ( 
.A(n_16480),
.B(n_10440),
.Y(n_16923)
);

AOI21xp5_ASAP7_75t_L g16924 ( 
.A1(n_16477),
.A2(n_11214),
.B(n_10783),
.Y(n_16924)
);

AND2x4_ASAP7_75t_SL g16925 ( 
.A(n_16299),
.B(n_8752),
.Y(n_16925)
);

NAND4xp25_ASAP7_75t_L g16926 ( 
.A(n_16462),
.B(n_7837),
.C(n_7851),
.D(n_7806),
.Y(n_16926)
);

OR2x2_ASAP7_75t_L g16927 ( 
.A(n_16481),
.B(n_11214),
.Y(n_16927)
);

HB1xp67_ASAP7_75t_L g16928 ( 
.A(n_16608),
.Y(n_16928)
);

INVx1_ASAP7_75t_L g16929 ( 
.A(n_16115),
.Y(n_16929)
);

INVx1_ASAP7_75t_L g16930 ( 
.A(n_16124),
.Y(n_16930)
);

INVx1_ASAP7_75t_SL g16931 ( 
.A(n_16298),
.Y(n_16931)
);

INVx1_ASAP7_75t_L g16932 ( 
.A(n_16128),
.Y(n_16932)
);

INVx1_ASAP7_75t_L g16933 ( 
.A(n_16151),
.Y(n_16933)
);

AND2x2_ASAP7_75t_L g16934 ( 
.A(n_16379),
.B(n_9078),
.Y(n_16934)
);

AND2x2_ASAP7_75t_L g16935 ( 
.A(n_16572),
.B(n_9078),
.Y(n_16935)
);

AND2x2_ASAP7_75t_L g16936 ( 
.A(n_16423),
.B(n_9178),
.Y(n_16936)
);

INVx1_ASAP7_75t_L g16937 ( 
.A(n_16180),
.Y(n_16937)
);

INVx1_ASAP7_75t_L g16938 ( 
.A(n_16200),
.Y(n_16938)
);

AND2x2_ASAP7_75t_SL g16939 ( 
.A(n_16471),
.B(n_7991),
.Y(n_16939)
);

AOI221xp5_ASAP7_75t_L g16940 ( 
.A1(n_16139),
.A2(n_16491),
.B1(n_16314),
.B2(n_16340),
.C(n_16339),
.Y(n_16940)
);

AND2x2_ASAP7_75t_SL g16941 ( 
.A(n_16473),
.B(n_7991),
.Y(n_16941)
);

HB1xp67_ASAP7_75t_L g16942 ( 
.A(n_16611),
.Y(n_16942)
);

INVx1_ASAP7_75t_L g16943 ( 
.A(n_16569),
.Y(n_16943)
);

AND2x2_ASAP7_75t_L g16944 ( 
.A(n_16443),
.B(n_9178),
.Y(n_16944)
);

INVx2_ASAP7_75t_L g16945 ( 
.A(n_16650),
.Y(n_16945)
);

AND2x2_ASAP7_75t_L g16946 ( 
.A(n_16489),
.B(n_9178),
.Y(n_16946)
);

AND2x2_ASAP7_75t_L g16947 ( 
.A(n_16573),
.B(n_9178),
.Y(n_16947)
);

NAND2x1_ASAP7_75t_L g16948 ( 
.A(n_16255),
.B(n_9470),
.Y(n_16948)
);

HB1xp67_ASAP7_75t_L g16949 ( 
.A(n_16478),
.Y(n_16949)
);

NAND3xp33_ASAP7_75t_L g16950 ( 
.A(n_16293),
.B(n_8639),
.C(n_8608),
.Y(n_16950)
);

INVx1_ASAP7_75t_L g16951 ( 
.A(n_16169),
.Y(n_16951)
);

AOI21xp33_ASAP7_75t_L g16952 ( 
.A1(n_16459),
.A2(n_11367),
.B(n_11360),
.Y(n_16952)
);

INVx1_ASAP7_75t_SL g16953 ( 
.A(n_16262),
.Y(n_16953)
);

AND2x4_ASAP7_75t_L g16954 ( 
.A(n_16612),
.B(n_16415),
.Y(n_16954)
);

INVx1_ASAP7_75t_L g16955 ( 
.A(n_16304),
.Y(n_16955)
);

INVx2_ASAP7_75t_L g16956 ( 
.A(n_16656),
.Y(n_16956)
);

INVx1_ASAP7_75t_L g16957 ( 
.A(n_16143),
.Y(n_16957)
);

NAND2xp5_ASAP7_75t_L g16958 ( 
.A(n_16321),
.B(n_10440),
.Y(n_16958)
);

AND2x2_ASAP7_75t_L g16959 ( 
.A(n_16460),
.B(n_16404),
.Y(n_16959)
);

INVx1_ASAP7_75t_L g16960 ( 
.A(n_16399),
.Y(n_16960)
);

NOR2xp33_ASAP7_75t_R g16961 ( 
.A(n_16317),
.B(n_8597),
.Y(n_16961)
);

AND2x2_ASAP7_75t_L g16962 ( 
.A(n_16390),
.B(n_9178),
.Y(n_16962)
);

INVx1_ASAP7_75t_L g16963 ( 
.A(n_16310),
.Y(n_16963)
);

OR2x2_ASAP7_75t_L g16964 ( 
.A(n_16144),
.B(n_8439),
.Y(n_16964)
);

INVx2_ASAP7_75t_L g16965 ( 
.A(n_16356),
.Y(n_16965)
);

HB1xp67_ASAP7_75t_L g16966 ( 
.A(n_16286),
.Y(n_16966)
);

AND2x2_ASAP7_75t_L g16967 ( 
.A(n_16392),
.B(n_9178),
.Y(n_16967)
);

INVx1_ASAP7_75t_L g16968 ( 
.A(n_16327),
.Y(n_16968)
);

INVx1_ASAP7_75t_L g16969 ( 
.A(n_16337),
.Y(n_16969)
);

AND2x2_ASAP7_75t_L g16970 ( 
.A(n_16567),
.B(n_9180),
.Y(n_16970)
);

HB1xp67_ASAP7_75t_L g16971 ( 
.A(n_16276),
.Y(n_16971)
);

AND2x2_ASAP7_75t_L g16972 ( 
.A(n_16605),
.B(n_9180),
.Y(n_16972)
);

INVxp67_ASAP7_75t_SL g16973 ( 
.A(n_16626),
.Y(n_16973)
);

INVx2_ASAP7_75t_L g16974 ( 
.A(n_16598),
.Y(n_16974)
);

INVx1_ASAP7_75t_L g16975 ( 
.A(n_16344),
.Y(n_16975)
);

HB1xp67_ASAP7_75t_L g16976 ( 
.A(n_16281),
.Y(n_16976)
);

INVx1_ASAP7_75t_L g16977 ( 
.A(n_16357),
.Y(n_16977)
);

INVx3_ASAP7_75t_SL g16978 ( 
.A(n_16521),
.Y(n_16978)
);

AND2x2_ASAP7_75t_L g16979 ( 
.A(n_16640),
.B(n_9180),
.Y(n_16979)
);

AND2x2_ASAP7_75t_L g16980 ( 
.A(n_16376),
.B(n_9180),
.Y(n_16980)
);

NAND2xp5_ASAP7_75t_L g16981 ( 
.A(n_16359),
.B(n_10442),
.Y(n_16981)
);

INVx1_ASAP7_75t_L g16982 ( 
.A(n_16336),
.Y(n_16982)
);

INVx1_ASAP7_75t_L g16983 ( 
.A(n_16366),
.Y(n_16983)
);

INVx1_ASAP7_75t_L g16984 ( 
.A(n_16222),
.Y(n_16984)
);

AND2x2_ASAP7_75t_L g16985 ( 
.A(n_16387),
.B(n_9180),
.Y(n_16985)
);

NAND2x1p5_ASAP7_75t_L g16986 ( 
.A(n_16658),
.B(n_8608),
.Y(n_16986)
);

NAND2x1_ASAP7_75t_L g16987 ( 
.A(n_16288),
.B(n_9478),
.Y(n_16987)
);

AND2x2_ASAP7_75t_L g16988 ( 
.A(n_16408),
.B(n_9180),
.Y(n_16988)
);

INVx2_ASAP7_75t_L g16989 ( 
.A(n_16592),
.Y(n_16989)
);

NAND2xp5_ASAP7_75t_SL g16990 ( 
.A(n_16631),
.B(n_8608),
.Y(n_16990)
);

INVx2_ASAP7_75t_SL g16991 ( 
.A(n_16448),
.Y(n_16991)
);

NAND2xp5_ASAP7_75t_L g16992 ( 
.A(n_16347),
.B(n_10442),
.Y(n_16992)
);

INVx1_ASAP7_75t_L g16993 ( 
.A(n_16225),
.Y(n_16993)
);

AND2x2_ASAP7_75t_L g16994 ( 
.A(n_16400),
.B(n_9210),
.Y(n_16994)
);

OR2x2_ASAP7_75t_L g16995 ( 
.A(n_16228),
.B(n_8439),
.Y(n_16995)
);

INVx1_ASAP7_75t_L g16996 ( 
.A(n_16369),
.Y(n_16996)
);

INVx1_ASAP7_75t_L g16997 ( 
.A(n_16187),
.Y(n_16997)
);

NAND2xp5_ASAP7_75t_L g16998 ( 
.A(n_16652),
.B(n_10449),
.Y(n_16998)
);

AND2x4_ASAP7_75t_SL g16999 ( 
.A(n_16651),
.B(n_8752),
.Y(n_16999)
);

AND2x2_ASAP7_75t_L g17000 ( 
.A(n_16447),
.B(n_9210),
.Y(n_17000)
);

AND2x2_ASAP7_75t_L g17001 ( 
.A(n_16461),
.B(n_9210),
.Y(n_17001)
);

INVx6_ASAP7_75t_L g17002 ( 
.A(n_16284),
.Y(n_17002)
);

OAI33xp33_ASAP7_75t_L g17003 ( 
.A1(n_16248),
.A2(n_10638),
.A3(n_10619),
.B1(n_10642),
.B2(n_10635),
.B3(n_10599),
.Y(n_17003)
);

BUFx2_ASAP7_75t_L g17004 ( 
.A(n_16294),
.Y(n_17004)
);

OR2x2_ASAP7_75t_L g17005 ( 
.A(n_16636),
.B(n_8439),
.Y(n_17005)
);

OR2x2_ASAP7_75t_L g17006 ( 
.A(n_16188),
.B(n_8456),
.Y(n_17006)
);

NAND2xp5_ASAP7_75t_L g17007 ( 
.A(n_16427),
.B(n_10449),
.Y(n_17007)
);

OR2x2_ASAP7_75t_L g17008 ( 
.A(n_16191),
.B(n_8456),
.Y(n_17008)
);

AOI22xp33_ASAP7_75t_L g17009 ( 
.A1(n_16522),
.A2(n_8639),
.B1(n_8838),
.B2(n_8608),
.Y(n_17009)
);

OR2x2_ASAP7_75t_L g17010 ( 
.A(n_16194),
.B(n_8456),
.Y(n_17010)
);

INVx1_ASAP7_75t_L g17011 ( 
.A(n_16205),
.Y(n_17011)
);

AND2x2_ASAP7_75t_L g17012 ( 
.A(n_16465),
.B(n_9210),
.Y(n_17012)
);

AND2x2_ASAP7_75t_L g17013 ( 
.A(n_16394),
.B(n_9210),
.Y(n_17013)
);

NOR2xp33_ASAP7_75t_R g17014 ( 
.A(n_16574),
.B(n_8597),
.Y(n_17014)
);

INVx3_ASAP7_75t_L g17015 ( 
.A(n_16528),
.Y(n_17015)
);

OR2x2_ASAP7_75t_L g17016 ( 
.A(n_16490),
.B(n_8575),
.Y(n_17016)
);

INVx1_ASAP7_75t_L g17017 ( 
.A(n_16576),
.Y(n_17017)
);

AND2x4_ASAP7_75t_L g17018 ( 
.A(n_16526),
.B(n_9210),
.Y(n_17018)
);

NAND2xp5_ASAP7_75t_L g17019 ( 
.A(n_16575),
.B(n_16577),
.Y(n_17019)
);

NAND2xp5_ASAP7_75t_L g17020 ( 
.A(n_16589),
.B(n_10454),
.Y(n_17020)
);

INVxp67_ASAP7_75t_L g17021 ( 
.A(n_16373),
.Y(n_17021)
);

AND4x1_ASAP7_75t_L g17022 ( 
.A(n_16452),
.B(n_7741),
.C(n_8691),
.D(n_8689),
.Y(n_17022)
);

AND2x2_ASAP7_75t_L g17023 ( 
.A(n_16641),
.B(n_9215),
.Y(n_17023)
);

NAND4xp25_ASAP7_75t_L g17024 ( 
.A(n_16630),
.B(n_7837),
.C(n_7851),
.D(n_7806),
.Y(n_17024)
);

NAND2xp5_ASAP7_75t_L g17025 ( 
.A(n_16590),
.B(n_10454),
.Y(n_17025)
);

NOR3xp33_ASAP7_75t_SL g17026 ( 
.A(n_16456),
.B(n_8691),
.C(n_8689),
.Y(n_17026)
);

NAND2xp5_ASAP7_75t_L g17027 ( 
.A(n_16593),
.B(n_10455),
.Y(n_17027)
);

AOI31xp33_ASAP7_75t_SL g17028 ( 
.A1(n_16648),
.A2(n_16351),
.A3(n_16414),
.B(n_16358),
.Y(n_17028)
);

OR2x2_ASAP7_75t_L g17029 ( 
.A(n_16438),
.B(n_8575),
.Y(n_17029)
);

INVx2_ASAP7_75t_L g17030 ( 
.A(n_16290),
.Y(n_17030)
);

INVx1_ASAP7_75t_L g17031 ( 
.A(n_16436),
.Y(n_17031)
);

OR2x2_ASAP7_75t_L g17032 ( 
.A(n_16257),
.B(n_16596),
.Y(n_17032)
);

NAND2xp5_ASAP7_75t_L g17033 ( 
.A(n_16597),
.B(n_10455),
.Y(n_17033)
);

AND2x4_ASAP7_75t_L g17034 ( 
.A(n_16599),
.B(n_9215),
.Y(n_17034)
);

AND2x2_ASAP7_75t_L g17035 ( 
.A(n_16275),
.B(n_9215),
.Y(n_17035)
);

AOI221xp5_ASAP7_75t_L g17036 ( 
.A1(n_16563),
.A2(n_10635),
.B1(n_10638),
.B2(n_10619),
.C(n_10599),
.Y(n_17036)
);

NAND2xp5_ASAP7_75t_L g17037 ( 
.A(n_16604),
.B(n_10456),
.Y(n_17037)
);

AND2x2_ASAP7_75t_L g17038 ( 
.A(n_16384),
.B(n_9215),
.Y(n_17038)
);

AND2x2_ASAP7_75t_L g17039 ( 
.A(n_16479),
.B(n_9215),
.Y(n_17039)
);

OR2x2_ASAP7_75t_L g17040 ( 
.A(n_16348),
.B(n_8682),
.Y(n_17040)
);

INVxp67_ASAP7_75t_L g17041 ( 
.A(n_16297),
.Y(n_17041)
);

INVx1_ASAP7_75t_L g17042 ( 
.A(n_16285),
.Y(n_17042)
);

INVx2_ASAP7_75t_L g17043 ( 
.A(n_16580),
.Y(n_17043)
);

INVx1_ASAP7_75t_L g17044 ( 
.A(n_16307),
.Y(n_17044)
);

AND2x2_ASAP7_75t_L g17045 ( 
.A(n_16444),
.B(n_9215),
.Y(n_17045)
);

AND2x2_ASAP7_75t_L g17046 ( 
.A(n_16502),
.B(n_9225),
.Y(n_17046)
);

NAND3xp33_ASAP7_75t_SL g17047 ( 
.A(n_16546),
.B(n_8613),
.C(n_8483),
.Y(n_17047)
);

OR2x2_ASAP7_75t_L g17048 ( 
.A(n_16643),
.B(n_16446),
.Y(n_17048)
);

AND2x4_ASAP7_75t_L g17049 ( 
.A(n_16505),
.B(n_9225),
.Y(n_17049)
);

NAND2xp5_ASAP7_75t_L g17050 ( 
.A(n_16507),
.B(n_10456),
.Y(n_17050)
);

AOI221xp5_ASAP7_75t_L g17051 ( 
.A1(n_16568),
.A2(n_10638),
.B1(n_10642),
.B2(n_10635),
.C(n_10619),
.Y(n_17051)
);

INVx1_ASAP7_75t_L g17052 ( 
.A(n_16325),
.Y(n_17052)
);

NOR3xp33_ASAP7_75t_L g17053 ( 
.A(n_16501),
.B(n_8269),
.C(n_8219),
.Y(n_17053)
);

AOI221xp5_ASAP7_75t_L g17054 ( 
.A1(n_16607),
.A2(n_10654),
.B1(n_10683),
.B2(n_10650),
.C(n_10642),
.Y(n_17054)
);

AND2x2_ASAP7_75t_SL g17055 ( 
.A(n_16508),
.B(n_8183),
.Y(n_17055)
);

BUFx3_ASAP7_75t_L g17056 ( 
.A(n_16615),
.Y(n_17056)
);

OAI211xp5_ASAP7_75t_SL g17057 ( 
.A1(n_16556),
.A2(n_10654),
.B(n_10683),
.C(n_10650),
.Y(n_17057)
);

INVx2_ASAP7_75t_L g17058 ( 
.A(n_16581),
.Y(n_17058)
);

AND2x2_ASAP7_75t_L g17059 ( 
.A(n_16638),
.B(n_9225),
.Y(n_17059)
);

NAND2xp5_ASAP7_75t_L g17060 ( 
.A(n_16402),
.B(n_10458),
.Y(n_17060)
);

NAND2xp5_ASAP7_75t_L g17061 ( 
.A(n_16457),
.B(n_16467),
.Y(n_17061)
);

INVxp67_ASAP7_75t_SL g17062 ( 
.A(n_16466),
.Y(n_17062)
);

CKINVDCx16_ASAP7_75t_R g17063 ( 
.A(n_16632),
.Y(n_17063)
);

INVx1_ASAP7_75t_L g17064 ( 
.A(n_16280),
.Y(n_17064)
);

AND2x2_ASAP7_75t_L g17065 ( 
.A(n_16657),
.B(n_9225),
.Y(n_17065)
);

INVx2_ASAP7_75t_L g17066 ( 
.A(n_16582),
.Y(n_17066)
);

INVx1_ASAP7_75t_L g17067 ( 
.A(n_16488),
.Y(n_17067)
);

NAND2x1_ASAP7_75t_L g17068 ( 
.A(n_16434),
.B(n_9478),
.Y(n_17068)
);

AND2x4_ASAP7_75t_L g17069 ( 
.A(n_16538),
.B(n_16633),
.Y(n_17069)
);

AND2x2_ASAP7_75t_L g17070 ( 
.A(n_16513),
.B(n_9225),
.Y(n_17070)
);

AND2x2_ASAP7_75t_L g17071 ( 
.A(n_16292),
.B(n_9225),
.Y(n_17071)
);

OAI21xp5_ASAP7_75t_SL g17072 ( 
.A1(n_16635),
.A2(n_9209),
.B(n_8862),
.Y(n_17072)
);

OR2x2_ASAP7_75t_L g17073 ( 
.A(n_16627),
.B(n_8682),
.Y(n_17073)
);

CKINVDCx20_ASAP7_75t_R g17074 ( 
.A(n_16644),
.Y(n_17074)
);

BUFx3_ASAP7_75t_L g17075 ( 
.A(n_16628),
.Y(n_17075)
);

INVx1_ASAP7_75t_L g17076 ( 
.A(n_16534),
.Y(n_17076)
);

INVx2_ASAP7_75t_L g17077 ( 
.A(n_16584),
.Y(n_17077)
);

NAND2xp5_ASAP7_75t_L g17078 ( 
.A(n_16474),
.B(n_10458),
.Y(n_17078)
);

NAND2x1p5_ASAP7_75t_L g17079 ( 
.A(n_16370),
.B(n_16322),
.Y(n_17079)
);

NAND2xp33_ASAP7_75t_SL g17080 ( 
.A(n_16519),
.B(n_8639),
.Y(n_17080)
);

OAI21xp5_ASAP7_75t_SL g17081 ( 
.A1(n_16458),
.A2(n_8862),
.B(n_8183),
.Y(n_17081)
);

NAND2xp5_ASAP7_75t_L g17082 ( 
.A(n_16484),
.B(n_10466),
.Y(n_17082)
);

NAND2xp5_ASAP7_75t_L g17083 ( 
.A(n_16485),
.B(n_10466),
.Y(n_17083)
);

INVx1_ASAP7_75t_L g17084 ( 
.A(n_16429),
.Y(n_17084)
);

OR2x2_ASAP7_75t_L g17085 ( 
.A(n_16328),
.B(n_8238),
.Y(n_17085)
);

INVx2_ASAP7_75t_L g17086 ( 
.A(n_16586),
.Y(n_17086)
);

AND2x2_ASAP7_75t_L g17087 ( 
.A(n_16537),
.B(n_9276),
.Y(n_17087)
);

INVx2_ASAP7_75t_L g17088 ( 
.A(n_16588),
.Y(n_17088)
);

AND2x2_ASAP7_75t_L g17089 ( 
.A(n_16251),
.B(n_9276),
.Y(n_17089)
);

AND2x2_ASAP7_75t_L g17090 ( 
.A(n_16450),
.B(n_9276),
.Y(n_17090)
);

AND2x2_ASAP7_75t_L g17091 ( 
.A(n_16463),
.B(n_9276),
.Y(n_17091)
);

INVx1_ASAP7_75t_L g17092 ( 
.A(n_16453),
.Y(n_17092)
);

AOI22xp33_ASAP7_75t_L g17093 ( 
.A1(n_16401),
.A2(n_8838),
.B1(n_8883),
.B2(n_8639),
.Y(n_17093)
);

INVx1_ASAP7_75t_L g17094 ( 
.A(n_16454),
.Y(n_17094)
);

NAND2xp5_ASAP7_75t_L g17095 ( 
.A(n_16472),
.B(n_10468),
.Y(n_17095)
);

INVx1_ASAP7_75t_L g17096 ( 
.A(n_16449),
.Y(n_17096)
);

INVx1_ASAP7_75t_L g17097 ( 
.A(n_16301),
.Y(n_17097)
);

INVx1_ASAP7_75t_L g17098 ( 
.A(n_16302),
.Y(n_17098)
);

INVxp67_ASAP7_75t_L g17099 ( 
.A(n_16306),
.Y(n_17099)
);

OR2x2_ASAP7_75t_L g17100 ( 
.A(n_16372),
.B(n_9482),
.Y(n_17100)
);

OR2x2_ASAP7_75t_L g17101 ( 
.A(n_16539),
.B(n_9482),
.Y(n_17101)
);

INVx1_ASAP7_75t_L g17102 ( 
.A(n_16360),
.Y(n_17102)
);

INVx2_ASAP7_75t_L g17103 ( 
.A(n_16555),
.Y(n_17103)
);

AND2x2_ASAP7_75t_L g17104 ( 
.A(n_16618),
.B(n_9276),
.Y(n_17104)
);

OR2x2_ASAP7_75t_L g17105 ( 
.A(n_16616),
.B(n_9482),
.Y(n_17105)
);

INVx2_ASAP7_75t_L g17106 ( 
.A(n_16558),
.Y(n_17106)
);

NAND2xp5_ASAP7_75t_L g17107 ( 
.A(n_16365),
.B(n_16510),
.Y(n_17107)
);

INVx2_ASAP7_75t_L g17108 ( 
.A(n_16560),
.Y(n_17108)
);

OR2x2_ASAP7_75t_L g17109 ( 
.A(n_16545),
.B(n_9485),
.Y(n_17109)
);

OR2x2_ASAP7_75t_L g17110 ( 
.A(n_16553),
.B(n_9485),
.Y(n_17110)
);

INVx1_ASAP7_75t_L g17111 ( 
.A(n_16253),
.Y(n_17111)
);

NAND2xp5_ASAP7_75t_L g17112 ( 
.A(n_16511),
.B(n_16329),
.Y(n_17112)
);

INVx2_ASAP7_75t_L g17113 ( 
.A(n_16561),
.Y(n_17113)
);

NAND2xp5_ASAP7_75t_L g17114 ( 
.A(n_16331),
.B(n_10468),
.Y(n_17114)
);

INVx1_ASAP7_75t_L g17115 ( 
.A(n_16258),
.Y(n_17115)
);

INVx2_ASAP7_75t_L g17116 ( 
.A(n_16566),
.Y(n_17116)
);

AND2x2_ASAP7_75t_L g17117 ( 
.A(n_16417),
.B(n_9276),
.Y(n_17117)
);

NOR2xp33_ASAP7_75t_L g17118 ( 
.A(n_16355),
.B(n_8838),
.Y(n_17118)
);

INVx1_ASAP7_75t_L g17119 ( 
.A(n_16437),
.Y(n_17119)
);

CKINVDCx5p33_ASAP7_75t_R g17120 ( 
.A(n_16500),
.Y(n_17120)
);

NAND2xp5_ASAP7_75t_L g17121 ( 
.A(n_16335),
.B(n_10469),
.Y(n_17121)
);

INVx1_ASAP7_75t_L g17122 ( 
.A(n_16261),
.Y(n_17122)
);

NAND2x1p5_ASAP7_75t_L g17123 ( 
.A(n_16425),
.B(n_8838),
.Y(n_17123)
);

INVx2_ASAP7_75t_L g17124 ( 
.A(n_16600),
.Y(n_17124)
);

INVx1_ASAP7_75t_L g17125 ( 
.A(n_16493),
.Y(n_17125)
);

OR2x2_ASAP7_75t_L g17126 ( 
.A(n_16441),
.B(n_9485),
.Y(n_17126)
);

OR2x2_ASAP7_75t_L g17127 ( 
.A(n_16354),
.B(n_9488),
.Y(n_17127)
);

AND2x2_ASAP7_75t_L g17128 ( 
.A(n_16389),
.B(n_16603),
.Y(n_17128)
);

INVx2_ASAP7_75t_L g17129 ( 
.A(n_16606),
.Y(n_17129)
);

INVx1_ASAP7_75t_L g17130 ( 
.A(n_16495),
.Y(n_17130)
);

INVx1_ASAP7_75t_L g17131 ( 
.A(n_16506),
.Y(n_17131)
);

INVx2_ASAP7_75t_L g17132 ( 
.A(n_16609),
.Y(n_17132)
);

INVx2_ASAP7_75t_L g17133 ( 
.A(n_16614),
.Y(n_17133)
);

OAI221xp5_ASAP7_75t_L g17134 ( 
.A1(n_16352),
.A2(n_8410),
.B1(n_8499),
.B2(n_8269),
.C(n_8219),
.Y(n_17134)
);

INVx1_ASAP7_75t_L g17135 ( 
.A(n_16509),
.Y(n_17135)
);

AND2x2_ASAP7_75t_L g17136 ( 
.A(n_16624),
.B(n_9290),
.Y(n_17136)
);

NOR2x1_ASAP7_75t_L g17137 ( 
.A(n_16645),
.B(n_10469),
.Y(n_17137)
);

INVx2_ASAP7_75t_L g17138 ( 
.A(n_16625),
.Y(n_17138)
);

AND2x2_ASAP7_75t_L g17139 ( 
.A(n_16634),
.B(n_9290),
.Y(n_17139)
);

INVx2_ASAP7_75t_L g17140 ( 
.A(n_16520),
.Y(n_17140)
);

AND2x2_ASAP7_75t_L g17141 ( 
.A(n_16470),
.B(n_9290),
.Y(n_17141)
);

NAND2xp5_ASAP7_75t_L g17142 ( 
.A(n_16547),
.B(n_10470),
.Y(n_17142)
);

AOI31xp33_ASAP7_75t_L g17143 ( 
.A1(n_16343),
.A2(n_7984),
.A3(n_8002),
.B(n_7942),
.Y(n_17143)
);

AND2x2_ASAP7_75t_L g17144 ( 
.A(n_16543),
.B(n_9290),
.Y(n_17144)
);

NAND2x1p5_ASAP7_75t_L g17145 ( 
.A(n_16486),
.B(n_8838),
.Y(n_17145)
);

AND2x2_ASAP7_75t_L g17146 ( 
.A(n_16530),
.B(n_9290),
.Y(n_17146)
);

INVx1_ASAP7_75t_L g17147 ( 
.A(n_16319),
.Y(n_17147)
);

INVxp67_ASAP7_75t_L g17148 ( 
.A(n_16368),
.Y(n_17148)
);

INVx1_ASAP7_75t_L g17149 ( 
.A(n_16433),
.Y(n_17149)
);

AND2x2_ASAP7_75t_L g17150 ( 
.A(n_16533),
.B(n_16536),
.Y(n_17150)
);

NAND2xp5_ASAP7_75t_L g17151 ( 
.A(n_16601),
.B(n_10470),
.Y(n_17151)
);

INVx1_ASAP7_75t_L g17152 ( 
.A(n_16405),
.Y(n_17152)
);

INVx2_ASAP7_75t_L g17153 ( 
.A(n_16542),
.Y(n_17153)
);

INVx2_ASAP7_75t_L g17154 ( 
.A(n_16548),
.Y(n_17154)
);

OR2x2_ASAP7_75t_L g17155 ( 
.A(n_16378),
.B(n_9488),
.Y(n_17155)
);

AND2x2_ASAP7_75t_L g17156 ( 
.A(n_16549),
.B(n_9290),
.Y(n_17156)
);

NOR3xp33_ASAP7_75t_L g17157 ( 
.A(n_16353),
.B(n_8269),
.C(n_8219),
.Y(n_17157)
);

INVx1_ASAP7_75t_L g17158 ( 
.A(n_16407),
.Y(n_17158)
);

AOI211x1_ASAP7_75t_SL g17159 ( 
.A1(n_16393),
.A2(n_10654),
.B(n_10683),
.C(n_10650),
.Y(n_17159)
);

INVx1_ASAP7_75t_L g17160 ( 
.A(n_16422),
.Y(n_17160)
);

INVx1_ASAP7_75t_L g17161 ( 
.A(n_16397),
.Y(n_17161)
);

AND2x2_ASAP7_75t_L g17162 ( 
.A(n_16550),
.B(n_9292),
.Y(n_17162)
);

AOI22xp33_ASAP7_75t_L g17163 ( 
.A1(n_16421),
.A2(n_8883),
.B1(n_8934),
.B2(n_8838),
.Y(n_17163)
);

INVx1_ASAP7_75t_SL g17164 ( 
.A(n_16266),
.Y(n_17164)
);

INVx1_ASAP7_75t_L g17165 ( 
.A(n_16482),
.Y(n_17165)
);

INVx1_ASAP7_75t_SL g17166 ( 
.A(n_16497),
.Y(n_17166)
);

AND2x4_ASAP7_75t_L g17167 ( 
.A(n_16498),
.B(n_9292),
.Y(n_17167)
);

INVx1_ASAP7_75t_L g17168 ( 
.A(n_16525),
.Y(n_17168)
);

AOI221xp5_ASAP7_75t_L g17169 ( 
.A1(n_16637),
.A2(n_10698),
.B1(n_10701),
.B2(n_10694),
.C(n_10685),
.Y(n_17169)
);

AND2x2_ASAP7_75t_L g17170 ( 
.A(n_16503),
.B(n_9292),
.Y(n_17170)
);

INVx1_ASAP7_75t_SL g17171 ( 
.A(n_16551),
.Y(n_17171)
);

AND2x2_ASAP7_75t_L g17172 ( 
.A(n_16562),
.B(n_9292),
.Y(n_17172)
);

INVx1_ASAP7_75t_L g17173 ( 
.A(n_16565),
.Y(n_17173)
);

AND2x2_ASAP7_75t_L g17174 ( 
.A(n_16646),
.B(n_9292),
.Y(n_17174)
);

CKINVDCx5p33_ASAP7_75t_R g17175 ( 
.A(n_16647),
.Y(n_17175)
);

NAND3xp33_ASAP7_75t_L g17176 ( 
.A(n_16649),
.B(n_8883),
.C(n_8838),
.Y(n_17176)
);

INVx2_ASAP7_75t_SL g17177 ( 
.A(n_16587),
.Y(n_17177)
);

AND2x2_ASAP7_75t_L g17178 ( 
.A(n_16594),
.B(n_16439),
.Y(n_17178)
);

NAND2xp5_ASAP7_75t_L g17179 ( 
.A(n_16295),
.B(n_16442),
.Y(n_17179)
);

AND2x2_ASAP7_75t_L g17180 ( 
.A(n_16621),
.B(n_9292),
.Y(n_17180)
);

AND2x2_ASAP7_75t_L g17181 ( 
.A(n_16621),
.B(n_8219),
.Y(n_17181)
);

NAND3xp33_ASAP7_75t_L g17182 ( 
.A(n_16330),
.B(n_8883),
.C(n_8838),
.Y(n_17182)
);

NAND2xp5_ASAP7_75t_L g17183 ( 
.A(n_16622),
.B(n_10471),
.Y(n_17183)
);

OR2x2_ASAP7_75t_L g17184 ( 
.A(n_16610),
.B(n_9488),
.Y(n_17184)
);

INVx1_ASAP7_75t_SL g17185 ( 
.A(n_16622),
.Y(n_17185)
);

INVx2_ASAP7_75t_L g17186 ( 
.A(n_16639),
.Y(n_17186)
);

AND2x4_ASAP7_75t_L g17187 ( 
.A(n_16751),
.B(n_16639),
.Y(n_17187)
);

INVx2_ASAP7_75t_L g17188 ( 
.A(n_16680),
.Y(n_17188)
);

NAND2x1_ASAP7_75t_L g17189 ( 
.A(n_16920),
.B(n_16323),
.Y(n_17189)
);

INVx2_ASAP7_75t_SL g17190 ( 
.A(n_16751),
.Y(n_17190)
);

NAND2xp5_ASAP7_75t_L g17191 ( 
.A(n_16713),
.B(n_16518),
.Y(n_17191)
);

INVx1_ASAP7_75t_L g17192 ( 
.A(n_16675),
.Y(n_17192)
);

INVx1_ASAP7_75t_L g17193 ( 
.A(n_16728),
.Y(n_17193)
);

INVx1_ASAP7_75t_L g17194 ( 
.A(n_16858),
.Y(n_17194)
);

INVx6_ASAP7_75t_L g17195 ( 
.A(n_16751),
.Y(n_17195)
);

INVx2_ASAP7_75t_L g17196 ( 
.A(n_16679),
.Y(n_17196)
);

AND2x4_ASAP7_75t_L g17197 ( 
.A(n_16887),
.B(n_11794),
.Y(n_17197)
);

AOI32xp33_ASAP7_75t_L g17198 ( 
.A1(n_16676),
.A2(n_11099),
.A3(n_11134),
.B1(n_11096),
.B2(n_11071),
.Y(n_17198)
);

AND2x2_ASAP7_75t_L g17199 ( 
.A(n_16692),
.B(n_10484),
.Y(n_17199)
);

OR2x6_ASAP7_75t_L g17200 ( 
.A(n_16672),
.B(n_7837),
.Y(n_17200)
);

OAI211xp5_ASAP7_75t_L g17201 ( 
.A1(n_16738),
.A2(n_10694),
.B(n_10698),
.C(n_10685),
.Y(n_17201)
);

INVx1_ASAP7_75t_L g17202 ( 
.A(n_16830),
.Y(n_17202)
);

INVx1_ASAP7_75t_L g17203 ( 
.A(n_16825),
.Y(n_17203)
);

NOR2x1_ASAP7_75t_L g17204 ( 
.A(n_16665),
.B(n_10471),
.Y(n_17204)
);

NOR2xp33_ASAP7_75t_L g17205 ( 
.A(n_16846),
.B(n_8883),
.Y(n_17205)
);

NOR2x1p5_ASAP7_75t_L g17206 ( 
.A(n_16741),
.B(n_8269),
.Y(n_17206)
);

INVx1_ASAP7_75t_L g17207 ( 
.A(n_16773),
.Y(n_17207)
);

OR2x2_ASAP7_75t_L g17208 ( 
.A(n_16821),
.B(n_9492),
.Y(n_17208)
);

AND2x2_ASAP7_75t_L g17209 ( 
.A(n_16695),
.B(n_10484),
.Y(n_17209)
);

INVx1_ASAP7_75t_L g17210 ( 
.A(n_16667),
.Y(n_17210)
);

OAI33xp33_ASAP7_75t_L g17211 ( 
.A1(n_16659),
.A2(n_10701),
.A3(n_10694),
.B1(n_10704),
.B2(n_10698),
.B3(n_10685),
.Y(n_17211)
);

O2A1O1Ixp5_ASAP7_75t_R g17212 ( 
.A1(n_16704),
.A2(n_7320),
.B(n_7332),
.C(n_7319),
.Y(n_17212)
);

OR2x2_ASAP7_75t_L g17213 ( 
.A(n_16765),
.B(n_16978),
.Y(n_17213)
);

OAI33xp33_ASAP7_75t_L g17214 ( 
.A1(n_16664),
.A2(n_10714),
.A3(n_10704),
.B1(n_10705),
.B2(n_10701),
.B3(n_9507),
.Y(n_17214)
);

INVx1_ASAP7_75t_L g17215 ( 
.A(n_16887),
.Y(n_17215)
);

INVx2_ASAP7_75t_L g17216 ( 
.A(n_16887),
.Y(n_17216)
);

INVx2_ASAP7_75t_L g17217 ( 
.A(n_16920),
.Y(n_17217)
);

AOI32xp33_ASAP7_75t_L g17218 ( 
.A1(n_16697),
.A2(n_11099),
.A3(n_11134),
.B1(n_11096),
.B2(n_11071),
.Y(n_17218)
);

INVx1_ASAP7_75t_L g17219 ( 
.A(n_16693),
.Y(n_17219)
);

INVx2_ASAP7_75t_L g17220 ( 
.A(n_16718),
.Y(n_17220)
);

OA222x2_ASAP7_75t_L g17221 ( 
.A1(n_16849),
.A2(n_16682),
.B1(n_16690),
.B2(n_16753),
.C1(n_16684),
.C2(n_16673),
.Y(n_17221)
);

INVx1_ASAP7_75t_L g17222 ( 
.A(n_16837),
.Y(n_17222)
);

INVx2_ASAP7_75t_L g17223 ( 
.A(n_17002),
.Y(n_17223)
);

INVx1_ASAP7_75t_SL g17224 ( 
.A(n_16661),
.Y(n_17224)
);

NAND2xp5_ASAP7_75t_L g17225 ( 
.A(n_16793),
.B(n_10481),
.Y(n_17225)
);

INVx1_ASAP7_75t_SL g17226 ( 
.A(n_17004),
.Y(n_17226)
);

AOI211xp5_ASAP7_75t_L g17227 ( 
.A1(n_16663),
.A2(n_11872),
.B(n_11877),
.C(n_11797),
.Y(n_17227)
);

OAI22xp5_ASAP7_75t_L g17228 ( 
.A1(n_16734),
.A2(n_8934),
.B1(n_8939),
.B2(n_8883),
.Y(n_17228)
);

INVx1_ASAP7_75t_L g17229 ( 
.A(n_16826),
.Y(n_17229)
);

INVx1_ASAP7_75t_L g17230 ( 
.A(n_16966),
.Y(n_17230)
);

NAND2x1p5_ASAP7_75t_L g17231 ( 
.A(n_16727),
.B(n_16711),
.Y(n_17231)
);

AND2x2_ASAP7_75t_SL g17232 ( 
.A(n_16911),
.B(n_8883),
.Y(n_17232)
);

OA222x2_ASAP7_75t_L g17233 ( 
.A1(n_16733),
.A2(n_9507),
.B1(n_9493),
.B2(n_9511),
.C1(n_9504),
.C2(n_9492),
.Y(n_17233)
);

AOI22xp5_ASAP7_75t_L g17234 ( 
.A1(n_16767),
.A2(n_8934),
.B1(n_8939),
.B2(n_8883),
.Y(n_17234)
);

AND2x2_ASAP7_75t_L g17235 ( 
.A(n_16696),
.B(n_10486),
.Y(n_17235)
);

INVx1_ASAP7_75t_L g17236 ( 
.A(n_16971),
.Y(n_17236)
);

AOI21xp33_ASAP7_75t_SL g17237 ( 
.A1(n_17063),
.A2(n_11872),
.B(n_11797),
.Y(n_17237)
);

INVxp67_ASAP7_75t_SL g17238 ( 
.A(n_16668),
.Y(n_17238)
);

INVxp67_ASAP7_75t_L g17239 ( 
.A(n_16928),
.Y(n_17239)
);

NAND2xp5_ASAP7_75t_L g17240 ( 
.A(n_16710),
.B(n_10481),
.Y(n_17240)
);

OAI32xp33_ASAP7_75t_L g17241 ( 
.A1(n_16829),
.A2(n_9504),
.A3(n_9507),
.B1(n_9493),
.B2(n_9492),
.Y(n_17241)
);

NAND2xp5_ASAP7_75t_L g17242 ( 
.A(n_16838),
.B(n_10492),
.Y(n_17242)
);

NAND2x1_ASAP7_75t_L g17243 ( 
.A(n_17002),
.B(n_9493),
.Y(n_17243)
);

INVx1_ASAP7_75t_L g17244 ( 
.A(n_16976),
.Y(n_17244)
);

OAI221xp5_ASAP7_75t_SL g17245 ( 
.A1(n_16670),
.A2(n_10714),
.B1(n_10705),
.B2(n_10704),
.C(n_9516),
.Y(n_17245)
);

INVx3_ASAP7_75t_L g17246 ( 
.A(n_16833),
.Y(n_17246)
);

INVxp67_ASAP7_75t_L g17247 ( 
.A(n_16942),
.Y(n_17247)
);

AND2x2_ASAP7_75t_L g17248 ( 
.A(n_16714),
.B(n_10486),
.Y(n_17248)
);

INVx1_ASAP7_75t_L g17249 ( 
.A(n_16949),
.Y(n_17249)
);

INVx2_ASAP7_75t_SL g17250 ( 
.A(n_16883),
.Y(n_17250)
);

INVx2_ASAP7_75t_L g17251 ( 
.A(n_16707),
.Y(n_17251)
);

INVx1_ASAP7_75t_L g17252 ( 
.A(n_16662),
.Y(n_17252)
);

INVx1_ASAP7_75t_L g17253 ( 
.A(n_16677),
.Y(n_17253)
);

OAI22xp5_ASAP7_75t_L g17254 ( 
.A1(n_16703),
.A2(n_8939),
.B1(n_9081),
.B2(n_8934),
.Y(n_17254)
);

INVx1_ASAP7_75t_L g17255 ( 
.A(n_16687),
.Y(n_17255)
);

OR2x2_ASAP7_75t_L g17256 ( 
.A(n_16852),
.B(n_9504),
.Y(n_17256)
);

NAND2xp5_ASAP7_75t_L g17257 ( 
.A(n_16746),
.B(n_10492),
.Y(n_17257)
);

INVx1_ASAP7_75t_L g17258 ( 
.A(n_16708),
.Y(n_17258)
);

INVx1_ASAP7_75t_L g17259 ( 
.A(n_16874),
.Y(n_17259)
);

OAI22xp33_ASAP7_75t_SL g17260 ( 
.A1(n_16762),
.A2(n_9516),
.B1(n_9520),
.B2(n_9511),
.Y(n_17260)
);

INVx1_ASAP7_75t_L g17261 ( 
.A(n_16689),
.Y(n_17261)
);

OAI32xp33_ASAP7_75t_L g17262 ( 
.A1(n_16772),
.A2(n_9520),
.A3(n_9523),
.B1(n_9516),
.B2(n_9511),
.Y(n_17262)
);

NOR2x1_ASAP7_75t_L g17263 ( 
.A(n_16681),
.B(n_10494),
.Y(n_17263)
);

INVx1_ASAP7_75t_L g17264 ( 
.A(n_16973),
.Y(n_17264)
);

NAND2xp5_ASAP7_75t_L g17265 ( 
.A(n_16867),
.B(n_10494),
.Y(n_17265)
);

AND2x4_ASAP7_75t_L g17266 ( 
.A(n_16698),
.B(n_11877),
.Y(n_17266)
);

INVx1_ASAP7_75t_SL g17267 ( 
.A(n_16845),
.Y(n_17267)
);

INVx1_ASAP7_75t_SL g17268 ( 
.A(n_16888),
.Y(n_17268)
);

AOI211xp5_ASAP7_75t_L g17269 ( 
.A1(n_17028),
.A2(n_11878),
.B(n_11407),
.C(n_11411),
.Y(n_17269)
);

INVxp67_ASAP7_75t_L g17270 ( 
.A(n_16678),
.Y(n_17270)
);

AND2x4_ASAP7_75t_SL g17271 ( 
.A(n_16722),
.B(n_8752),
.Y(n_17271)
);

INVxp67_ASAP7_75t_L g17272 ( 
.A(n_16737),
.Y(n_17272)
);

OR2x2_ASAP7_75t_L g17273 ( 
.A(n_16953),
.B(n_9520),
.Y(n_17273)
);

OAI22xp5_ASAP7_75t_L g17274 ( 
.A1(n_16724),
.A2(n_8939),
.B1(n_9081),
.B2(n_8934),
.Y(n_17274)
);

NOR2xp33_ASAP7_75t_L g17275 ( 
.A(n_16694),
.B(n_8934),
.Y(n_17275)
);

AOI32xp33_ASAP7_75t_L g17276 ( 
.A1(n_16716),
.A2(n_11143),
.A3(n_11197),
.B1(n_11169),
.B2(n_10714),
.Y(n_17276)
);

NOR3xp33_ASAP7_75t_L g17277 ( 
.A(n_16660),
.B(n_8410),
.C(n_8269),
.Y(n_17277)
);

AO22x1_ASAP7_75t_L g17278 ( 
.A1(n_17062),
.A2(n_16796),
.B1(n_16683),
.B2(n_16763),
.Y(n_17278)
);

INVx1_ASAP7_75t_L g17279 ( 
.A(n_16691),
.Y(n_17279)
);

NAND2xp5_ASAP7_75t_L g17280 ( 
.A(n_16706),
.B(n_10501),
.Y(n_17280)
);

OAI21xp33_ASAP7_75t_L g17281 ( 
.A1(n_16811),
.A2(n_10705),
.B(n_8499),
.Y(n_17281)
);

AND2x2_ASAP7_75t_L g17282 ( 
.A(n_16844),
.B(n_10506),
.Y(n_17282)
);

OAI33xp33_ASAP7_75t_L g17283 ( 
.A1(n_16805),
.A2(n_9545),
.A3(n_9528),
.B1(n_9553),
.B2(n_9531),
.B3(n_9523),
.Y(n_17283)
);

OR2x2_ASAP7_75t_L g17284 ( 
.A(n_16931),
.B(n_16872),
.Y(n_17284)
);

NAND2xp5_ASAP7_75t_L g17285 ( 
.A(n_16715),
.B(n_10501),
.Y(n_17285)
);

INVxp67_ASAP7_75t_L g17286 ( 
.A(n_16732),
.Y(n_17286)
);

INVx2_ASAP7_75t_L g17287 ( 
.A(n_16856),
.Y(n_17287)
);

AND2x2_ASAP7_75t_L g17288 ( 
.A(n_16808),
.B(n_10506),
.Y(n_17288)
);

INVx1_ASAP7_75t_L g17289 ( 
.A(n_17186),
.Y(n_17289)
);

AND2x2_ASAP7_75t_L g17290 ( 
.A(n_16717),
.B(n_10511),
.Y(n_17290)
);

INVx2_ASAP7_75t_L g17291 ( 
.A(n_16907),
.Y(n_17291)
);

NAND2xp5_ASAP7_75t_L g17292 ( 
.A(n_16719),
.B(n_16739),
.Y(n_17292)
);

AOI322xp5_ASAP7_75t_L g17293 ( 
.A1(n_16940),
.A2(n_9545),
.A3(n_9528),
.B1(n_9553),
.B2(n_9566),
.C1(n_9531),
.C2(n_9523),
.Y(n_17293)
);

INVx1_ASAP7_75t_L g17294 ( 
.A(n_16742),
.Y(n_17294)
);

INVx1_ASAP7_75t_L g17295 ( 
.A(n_16743),
.Y(n_17295)
);

AND2x2_ASAP7_75t_L g17296 ( 
.A(n_16700),
.B(n_10511),
.Y(n_17296)
);

AOI22xp5_ASAP7_75t_L g17297 ( 
.A1(n_17074),
.A2(n_16842),
.B1(n_16918),
.B2(n_16764),
.Y(n_17297)
);

INVxp67_ASAP7_75t_L g17298 ( 
.A(n_16735),
.Y(n_17298)
);

OR2x2_ASAP7_75t_L g17299 ( 
.A(n_16768),
.B(n_16890),
.Y(n_17299)
);

INVx2_ASAP7_75t_SL g17300 ( 
.A(n_17055),
.Y(n_17300)
);

INVx1_ASAP7_75t_L g17301 ( 
.A(n_17150),
.Y(n_17301)
);

AOI22xp33_ASAP7_75t_L g17302 ( 
.A1(n_16806),
.A2(n_8934),
.B1(n_9081),
.B2(n_8939),
.Y(n_17302)
);

AND2x2_ASAP7_75t_L g17303 ( 
.A(n_16893),
.B(n_8410),
.Y(n_17303)
);

INVx1_ASAP7_75t_L g17304 ( 
.A(n_16669),
.Y(n_17304)
);

INVx2_ASAP7_75t_L g17305 ( 
.A(n_16913),
.Y(n_17305)
);

AOI22xp5_ASAP7_75t_L g17306 ( 
.A1(n_16777),
.A2(n_8939),
.B1(n_9081),
.B2(n_8934),
.Y(n_17306)
);

OAI32xp33_ASAP7_75t_L g17307 ( 
.A1(n_16671),
.A2(n_9545),
.A3(n_9553),
.B1(n_9531),
.B2(n_9528),
.Y(n_17307)
);

INVx1_ASAP7_75t_L g17308 ( 
.A(n_16666),
.Y(n_17308)
);

NOR2xp67_ASAP7_75t_L g17309 ( 
.A(n_17047),
.B(n_8410),
.Y(n_17309)
);

AND2x2_ASAP7_75t_L g17310 ( 
.A(n_16726),
.B(n_8410),
.Y(n_17310)
);

INVxp67_ASAP7_75t_L g17311 ( 
.A(n_16736),
.Y(n_17311)
);

AOI21x1_ASAP7_75t_L g17312 ( 
.A1(n_16720),
.A2(n_10093),
.B(n_10064),
.Y(n_17312)
);

INVx1_ASAP7_75t_L g17313 ( 
.A(n_16674),
.Y(n_17313)
);

OR2x2_ASAP7_75t_L g17314 ( 
.A(n_16730),
.B(n_16859),
.Y(n_17314)
);

INVx1_ASAP7_75t_L g17315 ( 
.A(n_16775),
.Y(n_17315)
);

INVx1_ASAP7_75t_L g17316 ( 
.A(n_16686),
.Y(n_17316)
);

NAND2xp5_ASAP7_75t_L g17317 ( 
.A(n_16839),
.B(n_10504),
.Y(n_17317)
);

OAI22xp33_ASAP7_75t_L g17318 ( 
.A1(n_16791),
.A2(n_9568),
.B1(n_9569),
.B2(n_9566),
.Y(n_17318)
);

NAND2xp5_ASAP7_75t_L g17319 ( 
.A(n_16824),
.B(n_10504),
.Y(n_17319)
);

INVx1_ASAP7_75t_L g17320 ( 
.A(n_16769),
.Y(n_17320)
);

INVx1_ASAP7_75t_L g17321 ( 
.A(n_16789),
.Y(n_17321)
);

OR2x2_ASAP7_75t_L g17322 ( 
.A(n_16685),
.B(n_9566),
.Y(n_17322)
);

AOI21xp5_ASAP7_75t_L g17323 ( 
.A1(n_17019),
.A2(n_11169),
.B(n_11143),
.Y(n_17323)
);

INVx2_ASAP7_75t_SL g17324 ( 
.A(n_16894),
.Y(n_17324)
);

INVx1_ASAP7_75t_L g17325 ( 
.A(n_16688),
.Y(n_17325)
);

OR2x2_ASAP7_75t_L g17326 ( 
.A(n_16809),
.B(n_9568),
.Y(n_17326)
);

NAND4xp75_ASAP7_75t_L g17327 ( 
.A(n_16840),
.B(n_8386),
.C(n_7921),
.D(n_8035),
.Y(n_17327)
);

INVx1_ASAP7_75t_L g17328 ( 
.A(n_16760),
.Y(n_17328)
);

NAND4xp75_ASAP7_75t_L g17329 ( 
.A(n_16699),
.B(n_8386),
.C(n_7921),
.D(n_8035),
.Y(n_17329)
);

INVx1_ASAP7_75t_L g17330 ( 
.A(n_17061),
.Y(n_17330)
);

OR2x2_ASAP7_75t_L g17331 ( 
.A(n_16816),
.B(n_9568),
.Y(n_17331)
);

INVx1_ASAP7_75t_L g17332 ( 
.A(n_16701),
.Y(n_17332)
);

INVx1_ASAP7_75t_L g17333 ( 
.A(n_17112),
.Y(n_17333)
);

OAI22xp33_ASAP7_75t_L g17334 ( 
.A1(n_16752),
.A2(n_16894),
.B1(n_16834),
.B2(n_16801),
.Y(n_17334)
);

NAND2xp5_ASAP7_75t_L g17335 ( 
.A(n_17015),
.B(n_10507),
.Y(n_17335)
);

NOR3xp33_ASAP7_75t_L g17336 ( 
.A(n_16756),
.B(n_16933),
.C(n_16951),
.Y(n_17336)
);

INVx1_ASAP7_75t_L g17337 ( 
.A(n_16785),
.Y(n_17337)
);

INVx1_ASAP7_75t_L g17338 ( 
.A(n_16787),
.Y(n_17338)
);

INVx1_ASAP7_75t_L g17339 ( 
.A(n_16790),
.Y(n_17339)
);

OAI22xp5_ASAP7_75t_L g17340 ( 
.A1(n_17021),
.A2(n_9081),
.B1(n_9226),
.B2(n_8939),
.Y(n_17340)
);

AOI22xp5_ASAP7_75t_L g17341 ( 
.A1(n_16799),
.A2(n_9081),
.B1(n_9226),
.B2(n_8939),
.Y(n_17341)
);

AND2x4_ASAP7_75t_L g17342 ( 
.A(n_16861),
.B(n_16937),
.Y(n_17342)
);

INVx1_ASAP7_75t_L g17343 ( 
.A(n_16792),
.Y(n_17343)
);

INVxp33_ASAP7_75t_L g17344 ( 
.A(n_16705),
.Y(n_17344)
);

INVx1_ASAP7_75t_L g17345 ( 
.A(n_16757),
.Y(n_17345)
);

OAI32xp33_ASAP7_75t_L g17346 ( 
.A1(n_16912),
.A2(n_9585),
.A3(n_9569),
.B1(n_10211),
.B2(n_10200),
.Y(n_17346)
);

INVx2_ASAP7_75t_L g17347 ( 
.A(n_16798),
.Y(n_17347)
);

INVxp67_ASAP7_75t_L g17348 ( 
.A(n_16702),
.Y(n_17348)
);

NOR2xp33_ASAP7_75t_L g17349 ( 
.A(n_17041),
.B(n_9081),
.Y(n_17349)
);

NAND2xp5_ASAP7_75t_L g17350 ( 
.A(n_16908),
.B(n_10507),
.Y(n_17350)
);

INVx1_ASAP7_75t_L g17351 ( 
.A(n_17107),
.Y(n_17351)
);

OAI33xp33_ASAP7_75t_L g17352 ( 
.A1(n_16771),
.A2(n_16817),
.A3(n_16892),
.B1(n_16898),
.B2(n_16896),
.B3(n_16875),
.Y(n_17352)
);

AOI22xp5_ASAP7_75t_L g17353 ( 
.A1(n_16803),
.A2(n_9226),
.B1(n_9245),
.B2(n_9081),
.Y(n_17353)
);

AOI33xp33_ASAP7_75t_L g17354 ( 
.A1(n_16921),
.A2(n_9585),
.A3(n_9569),
.B1(n_10211),
.B2(n_10214),
.B3(n_10200),
.Y(n_17354)
);

HB1xp67_ASAP7_75t_L g17355 ( 
.A(n_16795),
.Y(n_17355)
);

INVx1_ASAP7_75t_L g17356 ( 
.A(n_16721),
.Y(n_17356)
);

OAI33xp33_ASAP7_75t_L g17357 ( 
.A1(n_16853),
.A2(n_9585),
.A3(n_10214),
.B1(n_10216),
.B2(n_10211),
.B3(n_10200),
.Y(n_17357)
);

BUFx2_ASAP7_75t_L g17358 ( 
.A(n_17079),
.Y(n_17358)
);

NAND2xp5_ASAP7_75t_L g17359 ( 
.A(n_17030),
.B(n_10510),
.Y(n_17359)
);

NAND2xp5_ASAP7_75t_SL g17360 ( 
.A(n_16729),
.B(n_9226),
.Y(n_17360)
);

INVx1_ASAP7_75t_L g17361 ( 
.A(n_16723),
.Y(n_17361)
);

O2A1O1Ixp5_ASAP7_75t_L g17362 ( 
.A1(n_16900),
.A2(n_10216),
.B(n_10220),
.C(n_10214),
.Y(n_17362)
);

AND2x2_ASAP7_75t_L g17363 ( 
.A(n_17128),
.B(n_8499),
.Y(n_17363)
);

INVx1_ASAP7_75t_L g17364 ( 
.A(n_16725),
.Y(n_17364)
);

INVx1_ASAP7_75t_L g17365 ( 
.A(n_16963),
.Y(n_17365)
);

INVx1_ASAP7_75t_L g17366 ( 
.A(n_16968),
.Y(n_17366)
);

INVx1_ASAP7_75t_L g17367 ( 
.A(n_16969),
.Y(n_17367)
);

NAND5xp2_ASAP7_75t_L g17368 ( 
.A(n_16959),
.B(n_7942),
.C(n_8007),
.D(n_8002),
.E(n_7984),
.Y(n_17368)
);

INVx1_ASAP7_75t_L g17369 ( 
.A(n_16975),
.Y(n_17369)
);

INVx2_ASAP7_75t_L g17370 ( 
.A(n_16781),
.Y(n_17370)
);

INVx3_ASAP7_75t_L g17371 ( 
.A(n_17018),
.Y(n_17371)
);

INVx1_ASAP7_75t_L g17372 ( 
.A(n_16977),
.Y(n_17372)
);

NAND2xp5_ASAP7_75t_L g17373 ( 
.A(n_17140),
.B(n_10510),
.Y(n_17373)
);

NAND2xp5_ASAP7_75t_L g17374 ( 
.A(n_17153),
.B(n_10524),
.Y(n_17374)
);

INVx1_ASAP7_75t_SL g17375 ( 
.A(n_17032),
.Y(n_17375)
);

INVx2_ASAP7_75t_L g17376 ( 
.A(n_16986),
.Y(n_17376)
);

INVx1_ASAP7_75t_L g17377 ( 
.A(n_16982),
.Y(n_17377)
);

NOR2x1p5_ASAP7_75t_SL g17378 ( 
.A(n_16878),
.B(n_10216),
.Y(n_17378)
);

AND2x2_ASAP7_75t_L g17379 ( 
.A(n_16989),
.B(n_8499),
.Y(n_17379)
);

OAI32xp33_ASAP7_75t_L g17380 ( 
.A1(n_17185),
.A2(n_16995),
.A3(n_16964),
.B1(n_16712),
.B2(n_17006),
.Y(n_17380)
);

INVx2_ASAP7_75t_L g17381 ( 
.A(n_17154),
.Y(n_17381)
);

INVx1_ASAP7_75t_L g17382 ( 
.A(n_16983),
.Y(n_17382)
);

INVx3_ASAP7_75t_L g17383 ( 
.A(n_16954),
.Y(n_17383)
);

OR2x2_ASAP7_75t_L g17384 ( 
.A(n_16866),
.B(n_9845),
.Y(n_17384)
);

AOI22xp33_ASAP7_75t_L g17385 ( 
.A1(n_16945),
.A2(n_9226),
.B1(n_9261),
.B2(n_9245),
.Y(n_17385)
);

AOI22xp5_ASAP7_75t_L g17386 ( 
.A1(n_16935),
.A2(n_9245),
.B1(n_9261),
.B2(n_9226),
.Y(n_17386)
);

NOR2x1p5_ASAP7_75t_SL g17387 ( 
.A(n_16880),
.B(n_10220),
.Y(n_17387)
);

OR2x2_ASAP7_75t_L g17388 ( 
.A(n_16869),
.B(n_9845),
.Y(n_17388)
);

INVx2_ASAP7_75t_SL g17389 ( 
.A(n_16939),
.Y(n_17389)
);

INVx1_ASAP7_75t_L g17390 ( 
.A(n_16996),
.Y(n_17390)
);

INVx2_ASAP7_75t_L g17391 ( 
.A(n_17180),
.Y(n_17391)
);

AND2x2_ASAP7_75t_L g17392 ( 
.A(n_16956),
.B(n_8499),
.Y(n_17392)
);

NOR3xp33_ASAP7_75t_L g17393 ( 
.A(n_16857),
.B(n_8563),
.C(n_8551),
.Y(n_17393)
);

NOR2xp33_ASAP7_75t_L g17394 ( 
.A(n_17052),
.B(n_17092),
.Y(n_17394)
);

NAND2xp5_ASAP7_75t_L g17395 ( 
.A(n_17094),
.B(n_10524),
.Y(n_17395)
);

NAND2xp5_ASAP7_75t_L g17396 ( 
.A(n_16938),
.B(n_10535),
.Y(n_17396)
);

BUFx2_ASAP7_75t_L g17397 ( 
.A(n_16841),
.Y(n_17397)
);

NAND2xp5_ASAP7_75t_SL g17398 ( 
.A(n_16941),
.B(n_9226),
.Y(n_17398)
);

NOR2x1_ASAP7_75t_R g17399 ( 
.A(n_17056),
.B(n_5627),
.Y(n_17399)
);

O2A1O1Ixp33_ASAP7_75t_SL g17400 ( 
.A1(n_17179),
.A2(n_7921),
.B(n_8035),
.C(n_7916),
.Y(n_17400)
);

INVx1_ASAP7_75t_L g17401 ( 
.A(n_17042),
.Y(n_17401)
);

O2A1O1Ixp5_ASAP7_75t_R g17402 ( 
.A1(n_16709),
.A2(n_16755),
.B(n_16758),
.C(n_16827),
.Y(n_17402)
);

INVx1_ASAP7_75t_L g17403 ( 
.A(n_17044),
.Y(n_17403)
);

AND2x2_ASAP7_75t_L g17404 ( 
.A(n_17043),
.B(n_17058),
.Y(n_17404)
);

INVx1_ASAP7_75t_L g17405 ( 
.A(n_17084),
.Y(n_17405)
);

OAI33xp33_ASAP7_75t_L g17406 ( 
.A1(n_16906),
.A2(n_10220),
.A3(n_10229),
.B1(n_10251),
.B2(n_10241),
.B3(n_10228),
.Y(n_17406)
);

A2O1A1Ixp33_ASAP7_75t_R g17407 ( 
.A1(n_16944),
.A2(n_8520),
.B(n_8567),
.C(n_8490),
.Y(n_17407)
);

OAI22xp33_ASAP7_75t_L g17408 ( 
.A1(n_16926),
.A2(n_9245),
.B1(n_9261),
.B2(n_9226),
.Y(n_17408)
);

OR2x2_ASAP7_75t_L g17409 ( 
.A(n_17005),
.B(n_9845),
.Y(n_17409)
);

INVx1_ASAP7_75t_L g17410 ( 
.A(n_16965),
.Y(n_17410)
);

INVx1_ASAP7_75t_L g17411 ( 
.A(n_17064),
.Y(n_17411)
);

INVxp33_ASAP7_75t_L g17412 ( 
.A(n_16748),
.Y(n_17412)
);

AOI22xp5_ASAP7_75t_L g17413 ( 
.A1(n_16759),
.A2(n_9261),
.B1(n_9245),
.B2(n_8563),
.Y(n_17413)
);

INVx1_ASAP7_75t_L g17414 ( 
.A(n_17097),
.Y(n_17414)
);

OAI32xp33_ASAP7_75t_L g17415 ( 
.A1(n_17008),
.A2(n_10228),
.A3(n_10251),
.B1(n_10241),
.B2(n_10229),
.Y(n_17415)
);

OR2x2_ASAP7_75t_L g17416 ( 
.A(n_16750),
.B(n_9865),
.Y(n_17416)
);

OR2x2_ASAP7_75t_L g17417 ( 
.A(n_17098),
.B(n_9865),
.Y(n_17417)
);

INVx1_ASAP7_75t_L g17418 ( 
.A(n_17102),
.Y(n_17418)
);

OAI33xp33_ASAP7_75t_L g17419 ( 
.A1(n_16909),
.A2(n_10229),
.A3(n_10241),
.B1(n_10254),
.B2(n_10251),
.B3(n_10228),
.Y(n_17419)
);

INVx1_ASAP7_75t_SL g17420 ( 
.A(n_16999),
.Y(n_17420)
);

XOR2x2_ASAP7_75t_L g17421 ( 
.A(n_16991),
.B(n_7851),
.Y(n_17421)
);

INVx1_ASAP7_75t_L g17422 ( 
.A(n_17125),
.Y(n_17422)
);

INVx1_ASAP7_75t_L g17423 ( 
.A(n_17130),
.Y(n_17423)
);

OAI33xp33_ASAP7_75t_L g17424 ( 
.A1(n_16914),
.A2(n_10258),
.A3(n_10259),
.B1(n_10292),
.B2(n_10269),
.B3(n_10254),
.Y(n_17424)
);

AOI22xp5_ASAP7_75t_L g17425 ( 
.A1(n_16778),
.A2(n_16917),
.B1(n_16864),
.B2(n_16877),
.Y(n_17425)
);

AND2x2_ASAP7_75t_L g17426 ( 
.A(n_17066),
.B(n_8551),
.Y(n_17426)
);

INVx2_ASAP7_75t_L g17427 ( 
.A(n_16774),
.Y(n_17427)
);

INVx1_ASAP7_75t_L g17428 ( 
.A(n_17131),
.Y(n_17428)
);

INVx1_ASAP7_75t_L g17429 ( 
.A(n_17135),
.Y(n_17429)
);

INVx1_ASAP7_75t_L g17430 ( 
.A(n_17031),
.Y(n_17430)
);

NOR2xp33_ASAP7_75t_SL g17431 ( 
.A(n_16807),
.B(n_9245),
.Y(n_17431)
);

INVx1_ASAP7_75t_L g17432 ( 
.A(n_16943),
.Y(n_17432)
);

INVx1_ASAP7_75t_L g17433 ( 
.A(n_17067),
.Y(n_17433)
);

INVx1_ASAP7_75t_L g17434 ( 
.A(n_17076),
.Y(n_17434)
);

OAI221xp5_ASAP7_75t_SL g17435 ( 
.A1(n_17081),
.A2(n_10259),
.B1(n_10269),
.B2(n_10258),
.C(n_10254),
.Y(n_17435)
);

INVxp67_ASAP7_75t_L g17436 ( 
.A(n_16731),
.Y(n_17436)
);

AOI21xp5_ASAP7_75t_L g17437 ( 
.A1(n_16990),
.A2(n_11197),
.B(n_11069),
.Y(n_17437)
);

INVx1_ASAP7_75t_L g17438 ( 
.A(n_16794),
.Y(n_17438)
);

AOI22xp33_ASAP7_75t_L g17439 ( 
.A1(n_17077),
.A2(n_9261),
.B1(n_9245),
.B2(n_9234),
.Y(n_17439)
);

AND2x2_ASAP7_75t_L g17440 ( 
.A(n_17086),
.B(n_8551),
.Y(n_17440)
);

INVx1_ASAP7_75t_L g17441 ( 
.A(n_16800),
.Y(n_17441)
);

AND2x2_ASAP7_75t_L g17442 ( 
.A(n_17088),
.B(n_8551),
.Y(n_17442)
);

INVx1_ASAP7_75t_L g17443 ( 
.A(n_16832),
.Y(n_17443)
);

NAND2xp5_ASAP7_75t_L g17444 ( 
.A(n_17103),
.B(n_10535),
.Y(n_17444)
);

A2O1A1Ixp33_ASAP7_75t_L g17445 ( 
.A1(n_16779),
.A2(n_11293),
.B(n_11284),
.C(n_11323),
.Y(n_17445)
);

AOI32xp33_ASAP7_75t_L g17446 ( 
.A1(n_16934),
.A2(n_10954),
.A3(n_10970),
.B1(n_10953),
.B2(n_10920),
.Y(n_17446)
);

BUFx3_ASAP7_75t_L g17447 ( 
.A(n_17075),
.Y(n_17447)
);

OAI33xp33_ASAP7_75t_L g17448 ( 
.A1(n_16915),
.A2(n_10259),
.A3(n_10269),
.B1(n_10293),
.B2(n_10292),
.B3(n_10258),
.Y(n_17448)
);

INVx1_ASAP7_75t_L g17449 ( 
.A(n_16780),
.Y(n_17449)
);

INVx1_ASAP7_75t_L g17450 ( 
.A(n_16916),
.Y(n_17450)
);

INVx1_ASAP7_75t_L g17451 ( 
.A(n_16744),
.Y(n_17451)
);

INVxp67_ASAP7_75t_L g17452 ( 
.A(n_17106),
.Y(n_17452)
);

AOI22xp5_ASAP7_75t_L g17453 ( 
.A1(n_16881),
.A2(n_9261),
.B1(n_9245),
.B2(n_8563),
.Y(n_17453)
);

INVx1_ASAP7_75t_L g17454 ( 
.A(n_16836),
.Y(n_17454)
);

INVx1_ASAP7_75t_L g17455 ( 
.A(n_16850),
.Y(n_17455)
);

INVx1_ASAP7_75t_L g17456 ( 
.A(n_16903),
.Y(n_17456)
);

OR2x2_ASAP7_75t_L g17457 ( 
.A(n_17129),
.B(n_9865),
.Y(n_17457)
);

INVx2_ASAP7_75t_L g17458 ( 
.A(n_16740),
.Y(n_17458)
);

OR2x2_ASAP7_75t_L g17459 ( 
.A(n_17132),
.B(n_9875),
.Y(n_17459)
);

OAI33xp33_ASAP7_75t_L g17460 ( 
.A1(n_16929),
.A2(n_10301),
.A3(n_10292),
.B1(n_10309),
.B2(n_10304),
.B3(n_10293),
.Y(n_17460)
);

INVx2_ASAP7_75t_L g17461 ( 
.A(n_16749),
.Y(n_17461)
);

OR2x2_ASAP7_75t_L g17462 ( 
.A(n_17133),
.B(n_9875),
.Y(n_17462)
);

AOI21xp33_ASAP7_75t_L g17463 ( 
.A1(n_16860),
.A2(n_11367),
.B(n_11360),
.Y(n_17463)
);

OR2x2_ASAP7_75t_L g17464 ( 
.A(n_17138),
.B(n_16788),
.Y(n_17464)
);

XOR2x2_ASAP7_75t_L g17465 ( 
.A(n_16863),
.B(n_7855),
.Y(n_17465)
);

AOI322xp5_ASAP7_75t_L g17466 ( 
.A1(n_16871),
.A2(n_10304),
.A3(n_10293),
.B1(n_10309),
.B2(n_10314),
.C1(n_10313),
.C2(n_10301),
.Y(n_17466)
);

NAND2xp5_ASAP7_75t_L g17467 ( 
.A(n_17108),
.B(n_10536),
.Y(n_17467)
);

INVx1_ASAP7_75t_SL g17468 ( 
.A(n_16925),
.Y(n_17468)
);

OR2x2_ASAP7_75t_L g17469 ( 
.A(n_17113),
.B(n_17116),
.Y(n_17469)
);

INVx2_ASAP7_75t_SL g17470 ( 
.A(n_16782),
.Y(n_17470)
);

XNOR2xp5_ASAP7_75t_L g17471 ( 
.A(n_17024),
.B(n_8183),
.Y(n_17471)
);

OR2x6_ASAP7_75t_L g17472 ( 
.A(n_16865),
.B(n_7855),
.Y(n_17472)
);

OAI222xp33_ASAP7_75t_L g17473 ( 
.A1(n_17184),
.A2(n_10313),
.B1(n_10304),
.B2(n_10314),
.C1(n_10309),
.C2(n_10301),
.Y(n_17473)
);

INVx1_ASAP7_75t_L g17474 ( 
.A(n_16904),
.Y(n_17474)
);

INVx2_ASAP7_75t_L g17475 ( 
.A(n_16754),
.Y(n_17475)
);

INVx1_ASAP7_75t_L g17476 ( 
.A(n_16905),
.Y(n_17476)
);

INVx1_ASAP7_75t_L g17477 ( 
.A(n_16910),
.Y(n_17477)
);

NAND4xp25_ASAP7_75t_L g17478 ( 
.A(n_17124),
.B(n_7894),
.C(n_7905),
.D(n_7855),
.Y(n_17478)
);

BUFx2_ASAP7_75t_L g17479 ( 
.A(n_17099),
.Y(n_17479)
);

OAI22xp33_ASAP7_75t_L g17480 ( 
.A1(n_17143),
.A2(n_16823),
.B1(n_17010),
.B2(n_16776),
.Y(n_17480)
);

OR2x2_ASAP7_75t_L g17481 ( 
.A(n_16955),
.B(n_9875),
.Y(n_17481)
);

NAND2xp5_ASAP7_75t_L g17482 ( 
.A(n_17096),
.B(n_10536),
.Y(n_17482)
);

OR2x2_ASAP7_75t_L g17483 ( 
.A(n_17048),
.B(n_8715),
.Y(n_17483)
);

OAI322xp33_ASAP7_75t_L g17484 ( 
.A1(n_16984),
.A2(n_10328),
.A3(n_10314),
.B1(n_10332),
.B2(n_10345),
.C1(n_10326),
.C2(n_10313),
.Y(n_17484)
);

INVx1_ASAP7_75t_L g17485 ( 
.A(n_17178),
.Y(n_17485)
);

HB1xp67_ASAP7_75t_L g17486 ( 
.A(n_16770),
.Y(n_17486)
);

INVx1_ASAP7_75t_L g17487 ( 
.A(n_16820),
.Y(n_17487)
);

NAND4xp75_ASAP7_75t_L g17488 ( 
.A(n_16873),
.B(n_8386),
.C(n_8053),
.D(n_8138),
.Y(n_17488)
);

OAI22xp5_ASAP7_75t_L g17489 ( 
.A1(n_16862),
.A2(n_9261),
.B1(n_8563),
.B2(n_8668),
.Y(n_17489)
);

INVx1_ASAP7_75t_L g17490 ( 
.A(n_16815),
.Y(n_17490)
);

BUFx12f_ASAP7_75t_L g17491 ( 
.A(n_17069),
.Y(n_17491)
);

NAND2xp5_ASAP7_75t_L g17492 ( 
.A(n_16882),
.B(n_17177),
.Y(n_17492)
);

NAND2xp5_ASAP7_75t_L g17493 ( 
.A(n_16895),
.B(n_10537),
.Y(n_17493)
);

INVx1_ASAP7_75t_L g17494 ( 
.A(n_16885),
.Y(n_17494)
);

OR2x2_ASAP7_75t_L g17495 ( 
.A(n_17029),
.B(n_8715),
.Y(n_17495)
);

AND2x2_ASAP7_75t_L g17496 ( 
.A(n_16902),
.B(n_8551),
.Y(n_17496)
);

INVx1_ASAP7_75t_L g17497 ( 
.A(n_16886),
.Y(n_17497)
);

INVx1_ASAP7_75t_SL g17498 ( 
.A(n_17164),
.Y(n_17498)
);

INVx1_ASAP7_75t_L g17499 ( 
.A(n_16891),
.Y(n_17499)
);

NAND2xp5_ASAP7_75t_L g17500 ( 
.A(n_17166),
.B(n_10537),
.Y(n_17500)
);

INVxp67_ASAP7_75t_SL g17501 ( 
.A(n_16879),
.Y(n_17501)
);

INVx2_ASAP7_75t_L g17502 ( 
.A(n_16818),
.Y(n_17502)
);

NAND4xp75_ASAP7_75t_L g17503 ( 
.A(n_16993),
.B(n_8386),
.C(n_8053),
.D(n_8138),
.Y(n_17503)
);

OAI33xp33_ASAP7_75t_L g17504 ( 
.A1(n_16930),
.A2(n_10345),
.A3(n_10328),
.B1(n_10351),
.B2(n_10332),
.B3(n_10326),
.Y(n_17504)
);

INVx1_ASAP7_75t_L g17505 ( 
.A(n_16899),
.Y(n_17505)
);

NAND2xp5_ASAP7_75t_L g17506 ( 
.A(n_17171),
.B(n_16936),
.Y(n_17506)
);

OAI33xp33_ASAP7_75t_L g17507 ( 
.A1(n_16932),
.A2(n_10345),
.A3(n_10328),
.B1(n_10351),
.B2(n_10332),
.B3(n_10326),
.Y(n_17507)
);

AOI322xp5_ASAP7_75t_L g17508 ( 
.A1(n_16957),
.A2(n_10360),
.A3(n_10354),
.B1(n_10373),
.B2(n_10374),
.C1(n_10355),
.C2(n_10351),
.Y(n_17508)
);

HB1xp67_ASAP7_75t_L g17509 ( 
.A(n_16974),
.Y(n_17509)
);

NAND2x1p5_ASAP7_75t_L g17510 ( 
.A(n_16960),
.B(n_9261),
.Y(n_17510)
);

O2A1O1Ixp5_ASAP7_75t_R g17511 ( 
.A1(n_16828),
.A2(n_16813),
.B(n_16835),
.C(n_16812),
.Y(n_17511)
);

NOR2x1_ASAP7_75t_L g17512 ( 
.A(n_16997),
.B(n_10542),
.Y(n_17512)
);

NOR2x1p5_ASAP7_75t_L g17513 ( 
.A(n_17120),
.B(n_8563),
.Y(n_17513)
);

INVx1_ASAP7_75t_SL g17514 ( 
.A(n_16922),
.Y(n_17514)
);

AOI22xp5_ASAP7_75t_L g17515 ( 
.A1(n_16797),
.A2(n_8672),
.B1(n_8683),
.B2(n_8668),
.Y(n_17515)
);

INVx1_ASAP7_75t_L g17516 ( 
.A(n_16927),
.Y(n_17516)
);

INVx2_ASAP7_75t_L g17517 ( 
.A(n_16810),
.Y(n_17517)
);

OAI22xp5_ASAP7_75t_L g17518 ( 
.A1(n_16786),
.A2(n_8672),
.B1(n_8683),
.B2(n_8668),
.Y(n_17518)
);

AND2x4_ASAP7_75t_L g17519 ( 
.A(n_17111),
.B(n_11878),
.Y(n_17519)
);

INVx2_ASAP7_75t_L g17520 ( 
.A(n_16814),
.Y(n_17520)
);

NOR2xp67_ASAP7_75t_L g17521 ( 
.A(n_17148),
.B(n_8668),
.Y(n_17521)
);

OAI22xp33_ASAP7_75t_L g17522 ( 
.A1(n_16783),
.A2(n_8672),
.B1(n_8683),
.B2(n_8668),
.Y(n_17522)
);

OAI33xp33_ASAP7_75t_L g17523 ( 
.A1(n_17011),
.A2(n_10373),
.A3(n_10355),
.B1(n_10374),
.B2(n_10360),
.B3(n_10354),
.Y(n_17523)
);

OR2x2_ASAP7_75t_L g17524 ( 
.A(n_17040),
.B(n_8715),
.Y(n_17524)
);

NOR2xp33_ASAP7_75t_L g17525 ( 
.A(n_17017),
.B(n_17175),
.Y(n_17525)
);

BUFx2_ASAP7_75t_L g17526 ( 
.A(n_16843),
.Y(n_17526)
);

OR2x2_ASAP7_75t_L g17527 ( 
.A(n_17073),
.B(n_8806),
.Y(n_17527)
);

INVx1_ASAP7_75t_L g17528 ( 
.A(n_16847),
.Y(n_17528)
);

XNOR2x2_ASAP7_75t_L g17529 ( 
.A(n_17115),
.B(n_17152),
.Y(n_17529)
);

INVx3_ASAP7_75t_L g17530 ( 
.A(n_17034),
.Y(n_17530)
);

INVx2_ASAP7_75t_L g17531 ( 
.A(n_16831),
.Y(n_17531)
);

AOI22xp5_ASAP7_75t_L g17532 ( 
.A1(n_16897),
.A2(n_8683),
.B1(n_8688),
.B2(n_8672),
.Y(n_17532)
);

OR2x2_ASAP7_75t_L g17533 ( 
.A(n_17016),
.B(n_8806),
.Y(n_17533)
);

AND2x4_ASAP7_75t_L g17534 ( 
.A(n_17122),
.B(n_11401),
.Y(n_17534)
);

INVx2_ASAP7_75t_L g17535 ( 
.A(n_16884),
.Y(n_17535)
);

OAI22xp5_ASAP7_75t_L g17536 ( 
.A1(n_17026),
.A2(n_8683),
.B1(n_8688),
.B2(n_8672),
.Y(n_17536)
);

INVx2_ASAP7_75t_SL g17537 ( 
.A(n_16784),
.Y(n_17537)
);

INVx1_ASAP7_75t_L g17538 ( 
.A(n_16848),
.Y(n_17538)
);

INVx1_ASAP7_75t_L g17539 ( 
.A(n_16851),
.Y(n_17539)
);

NAND2xp5_ASAP7_75t_L g17540 ( 
.A(n_16970),
.B(n_10542),
.Y(n_17540)
);

INVx1_ASAP7_75t_L g17541 ( 
.A(n_16923),
.Y(n_17541)
);

AND2x2_ASAP7_75t_L g17542 ( 
.A(n_16972),
.B(n_8688),
.Y(n_17542)
);

INVx1_ASAP7_75t_L g17543 ( 
.A(n_16998),
.Y(n_17543)
);

INVx1_ASAP7_75t_L g17544 ( 
.A(n_17020),
.Y(n_17544)
);

INVx1_ASAP7_75t_L g17545 ( 
.A(n_17025),
.Y(n_17545)
);

NAND2x2_ASAP7_75t_L g17546 ( 
.A(n_17027),
.B(n_7855),
.Y(n_17546)
);

AOI22xp33_ASAP7_75t_L g17547 ( 
.A1(n_17049),
.A2(n_8048),
.B1(n_10355),
.B2(n_10354),
.Y(n_17547)
);

NAND2xp5_ASAP7_75t_L g17548 ( 
.A(n_16985),
.B(n_10543),
.Y(n_17548)
);

INVxp67_ASAP7_75t_L g17549 ( 
.A(n_17161),
.Y(n_17549)
);

INVx2_ASAP7_75t_L g17550 ( 
.A(n_17145),
.Y(n_17550)
);

NOR2x1_ASAP7_75t_L g17551 ( 
.A(n_17158),
.B(n_10543),
.Y(n_17551)
);

INVx1_ASAP7_75t_L g17552 ( 
.A(n_17033),
.Y(n_17552)
);

NAND2xp5_ASAP7_75t_SL g17553 ( 
.A(n_17022),
.B(n_17014),
.Y(n_17553)
);

INVx2_ASAP7_75t_L g17554 ( 
.A(n_17045),
.Y(n_17554)
);

OAI22xp5_ASAP7_75t_L g17555 ( 
.A1(n_17072),
.A2(n_8754),
.B1(n_8774),
.B2(n_8688),
.Y(n_17555)
);

INVx2_ASAP7_75t_L g17556 ( 
.A(n_16889),
.Y(n_17556)
);

INVx2_ASAP7_75t_SL g17557 ( 
.A(n_16946),
.Y(n_17557)
);

INVx1_ASAP7_75t_L g17558 ( 
.A(n_17037),
.Y(n_17558)
);

INVx2_ASAP7_75t_L g17559 ( 
.A(n_16766),
.Y(n_17559)
);

AOI22xp5_ASAP7_75t_L g17560 ( 
.A1(n_16870),
.A2(n_8754),
.B1(n_8774),
.B2(n_8688),
.Y(n_17560)
);

INVx2_ASAP7_75t_SL g17561 ( 
.A(n_16804),
.Y(n_17561)
);

OR2x2_ASAP7_75t_L g17562 ( 
.A(n_17119),
.B(n_8806),
.Y(n_17562)
);

O2A1O1Ixp33_ASAP7_75t_L g17563 ( 
.A1(n_17149),
.A2(n_10373),
.B(n_10374),
.C(n_10360),
.Y(n_17563)
);

INVx1_ASAP7_75t_L g17564 ( 
.A(n_16855),
.Y(n_17564)
);

INVx1_ASAP7_75t_L g17565 ( 
.A(n_16958),
.Y(n_17565)
);

AND2x4_ASAP7_75t_L g17566 ( 
.A(n_17147),
.B(n_11401),
.Y(n_17566)
);

NAND2xp5_ASAP7_75t_L g17567 ( 
.A(n_16988),
.B(n_16962),
.Y(n_17567)
);

OR3x2_ASAP7_75t_L g17568 ( 
.A(n_17160),
.B(n_8359),
.C(n_8952),
.Y(n_17568)
);

NOR2xp33_ASAP7_75t_L g17569 ( 
.A(n_17165),
.B(n_8754),
.Y(n_17569)
);

OR2x2_ASAP7_75t_L g17570 ( 
.A(n_17060),
.B(n_10547),
.Y(n_17570)
);

OR2x6_ASAP7_75t_L g17571 ( 
.A(n_17168),
.B(n_7894),
.Y(n_17571)
);

HB1xp67_ASAP7_75t_L g17572 ( 
.A(n_17137),
.Y(n_17572)
);

INVxp67_ASAP7_75t_SL g17573 ( 
.A(n_16868),
.Y(n_17573)
);

INVx1_ASAP7_75t_L g17574 ( 
.A(n_16992),
.Y(n_17574)
);

AND2x2_ASAP7_75t_L g17575 ( 
.A(n_16967),
.B(n_8754),
.Y(n_17575)
);

NAND2xp5_ASAP7_75t_L g17576 ( 
.A(n_16994),
.B(n_10547),
.Y(n_17576)
);

OAI22xp33_ASAP7_75t_L g17577 ( 
.A1(n_17182),
.A2(n_8774),
.B1(n_8829),
.B2(n_8754),
.Y(n_17577)
);

AND2x2_ASAP7_75t_L g17578 ( 
.A(n_17013),
.B(n_8774),
.Y(n_17578)
);

OR2x2_ASAP7_75t_L g17579 ( 
.A(n_16981),
.B(n_10550),
.Y(n_17579)
);

INVx1_ASAP7_75t_L g17580 ( 
.A(n_17007),
.Y(n_17580)
);

HB1xp67_ASAP7_75t_L g17581 ( 
.A(n_16980),
.Y(n_17581)
);

HB1xp67_ASAP7_75t_L g17582 ( 
.A(n_17000),
.Y(n_17582)
);

INVx1_ASAP7_75t_L g17583 ( 
.A(n_17050),
.Y(n_17583)
);

INVx1_ASAP7_75t_L g17584 ( 
.A(n_17173),
.Y(n_17584)
);

INVx1_ASAP7_75t_L g17585 ( 
.A(n_17078),
.Y(n_17585)
);

AND2x2_ASAP7_75t_L g17586 ( 
.A(n_16979),
.B(n_8774),
.Y(n_17586)
);

OAI31xp67_ASAP7_75t_L g17587 ( 
.A1(n_16747),
.A2(n_10392),
.A3(n_10399),
.B(n_10381),
.Y(n_17587)
);

INVx1_ASAP7_75t_L g17588 ( 
.A(n_17082),
.Y(n_17588)
);

AND2x4_ASAP7_75t_L g17589 ( 
.A(n_16947),
.B(n_11407),
.Y(n_17589)
);

INVx1_ASAP7_75t_L g17590 ( 
.A(n_17083),
.Y(n_17590)
);

OAI31xp33_ASAP7_75t_L g17591 ( 
.A1(n_16745),
.A2(n_10392),
.A3(n_10399),
.B(n_10381),
.Y(n_17591)
);

NAND2xp5_ASAP7_75t_L g17592 ( 
.A(n_17001),
.B(n_10550),
.Y(n_17592)
);

INVx2_ASAP7_75t_L g17593 ( 
.A(n_16919),
.Y(n_17593)
);

OR2x2_ASAP7_75t_L g17594 ( 
.A(n_17142),
.B(n_10556),
.Y(n_17594)
);

INVx2_ASAP7_75t_L g17595 ( 
.A(n_17123),
.Y(n_17595)
);

INVx2_ASAP7_75t_L g17596 ( 
.A(n_17035),
.Y(n_17596)
);

INVx1_ASAP7_75t_L g17597 ( 
.A(n_17095),
.Y(n_17597)
);

INVx2_ASAP7_75t_L g17598 ( 
.A(n_17071),
.Y(n_17598)
);

INVx1_ASAP7_75t_L g17599 ( 
.A(n_17114),
.Y(n_17599)
);

INVx1_ASAP7_75t_L g17600 ( 
.A(n_17121),
.Y(n_17600)
);

OA222x2_ASAP7_75t_L g17601 ( 
.A1(n_17085),
.A2(n_10438),
.B1(n_10392),
.B2(n_10445),
.C1(n_10399),
.C2(n_10381),
.Y(n_17601)
);

OAI322xp33_ASAP7_75t_L g17602 ( 
.A1(n_17118),
.A2(n_10445),
.A3(n_10447),
.B1(n_10438),
.B2(n_8708),
.C1(n_8483),
.C2(n_8613),
.Y(n_17602)
);

INVx1_ASAP7_75t_L g17603 ( 
.A(n_17151),
.Y(n_17603)
);

AND2x4_ASAP7_75t_L g17604 ( 
.A(n_17012),
.B(n_11411),
.Y(n_17604)
);

INVx1_ASAP7_75t_L g17605 ( 
.A(n_17183),
.Y(n_17605)
);

INVx1_ASAP7_75t_L g17606 ( 
.A(n_17039),
.Y(n_17606)
);

NAND2xp5_ASAP7_75t_L g17607 ( 
.A(n_17046),
.B(n_10556),
.Y(n_17607)
);

INVx1_ASAP7_75t_L g17608 ( 
.A(n_16876),
.Y(n_17608)
);

INVx1_ASAP7_75t_L g17609 ( 
.A(n_17170),
.Y(n_17609)
);

AND2x4_ASAP7_75t_L g17610 ( 
.A(n_17070),
.B(n_11440),
.Y(n_17610)
);

NAND2xp5_ASAP7_75t_L g17611 ( 
.A(n_17172),
.B(n_10558),
.Y(n_17611)
);

NAND2xp5_ASAP7_75t_L g17612 ( 
.A(n_17174),
.B(n_10558),
.Y(n_17612)
);

AND2x2_ASAP7_75t_L g17613 ( 
.A(n_17144),
.B(n_8829),
.Y(n_17613)
);

NAND2xp5_ASAP7_75t_L g17614 ( 
.A(n_17167),
.B(n_10560),
.Y(n_17614)
);

AOI322xp5_ASAP7_75t_L g17615 ( 
.A1(n_17163),
.A2(n_10445),
.A3(n_10447),
.B1(n_10438),
.B2(n_8978),
.C1(n_8708),
.C2(n_8725),
.Y(n_17615)
);

AND2x2_ASAP7_75t_L g17616 ( 
.A(n_17038),
.B(n_8829),
.Y(n_17616)
);

OAI22xp33_ASAP7_75t_L g17617 ( 
.A1(n_16854),
.A2(n_8980),
.B1(n_9022),
.B2(n_8829),
.Y(n_17617)
);

INVxp67_ASAP7_75t_SL g17618 ( 
.A(n_16901),
.Y(n_17618)
);

OR2x2_ASAP7_75t_L g17619 ( 
.A(n_17155),
.B(n_10560),
.Y(n_17619)
);

NAND2xp5_ASAP7_75t_L g17620 ( 
.A(n_17091),
.B(n_10562),
.Y(n_17620)
);

NAND2xp5_ASAP7_75t_L g17621 ( 
.A(n_17246),
.B(n_17089),
.Y(n_17621)
);

INVx2_ASAP7_75t_L g17622 ( 
.A(n_17195),
.Y(n_17622)
);

INVx1_ASAP7_75t_L g17623 ( 
.A(n_17486),
.Y(n_17623)
);

NAND2xp5_ASAP7_75t_L g17624 ( 
.A(n_17250),
.B(n_17117),
.Y(n_17624)
);

NAND4xp25_ASAP7_75t_L g17625 ( 
.A(n_17297),
.B(n_17053),
.C(n_17023),
.D(n_16924),
.Y(n_17625)
);

NAND2x1p5_ASAP7_75t_L g17626 ( 
.A(n_17268),
.B(n_17181),
.Y(n_17626)
);

NAND2xp5_ASAP7_75t_L g17627 ( 
.A(n_17383),
.B(n_17146),
.Y(n_17627)
);

NAND3xp33_ASAP7_75t_L g17628 ( 
.A(n_17194),
.B(n_17080),
.C(n_17176),
.Y(n_17628)
);

INVx1_ASAP7_75t_L g17629 ( 
.A(n_17397),
.Y(n_17629)
);

AND2x2_ASAP7_75t_L g17630 ( 
.A(n_17220),
.B(n_17087),
.Y(n_17630)
);

NAND2xp5_ASAP7_75t_L g17631 ( 
.A(n_17238),
.B(n_17156),
.Y(n_17631)
);

OAI21xp33_ASAP7_75t_SL g17632 ( 
.A1(n_17263),
.A2(n_17104),
.B(n_17090),
.Y(n_17632)
);

AND2x2_ASAP7_75t_L g17633 ( 
.A(n_17231),
.B(n_17059),
.Y(n_17633)
);

AND2x2_ASAP7_75t_L g17634 ( 
.A(n_17226),
.B(n_17065),
.Y(n_17634)
);

NAND2xp5_ASAP7_75t_L g17635 ( 
.A(n_17278),
.B(n_17162),
.Y(n_17635)
);

OR2x2_ASAP7_75t_L g17636 ( 
.A(n_17224),
.B(n_17126),
.Y(n_17636)
);

INVx1_ASAP7_75t_L g17637 ( 
.A(n_17215),
.Y(n_17637)
);

NAND2xp5_ASAP7_75t_L g17638 ( 
.A(n_17342),
.B(n_17141),
.Y(n_17638)
);

NOR3xp33_ASAP7_75t_L g17639 ( 
.A(n_17358),
.B(n_16952),
.C(n_17157),
.Y(n_17639)
);

AOI211xp5_ASAP7_75t_SL g17640 ( 
.A1(n_17334),
.A2(n_17100),
.B(n_17101),
.C(n_17109),
.Y(n_17640)
);

INVx1_ASAP7_75t_L g17641 ( 
.A(n_17195),
.Y(n_17641)
);

HB1xp67_ASAP7_75t_L g17642 ( 
.A(n_17216),
.Y(n_17642)
);

AOI22xp33_ASAP7_75t_L g17643 ( 
.A1(n_17491),
.A2(n_16802),
.B1(n_17139),
.B2(n_17136),
.Y(n_17643)
);

NOR2x1_ASAP7_75t_L g17644 ( 
.A(n_17187),
.B(n_16948),
.Y(n_17644)
);

NAND2xp5_ASAP7_75t_L g17645 ( 
.A(n_17342),
.B(n_16961),
.Y(n_17645)
);

INVx1_ASAP7_75t_L g17646 ( 
.A(n_17572),
.Y(n_17646)
);

INVx1_ASAP7_75t_SL g17647 ( 
.A(n_17213),
.Y(n_17647)
);

INVx1_ASAP7_75t_L g17648 ( 
.A(n_17355),
.Y(n_17648)
);

INVx1_ASAP7_75t_L g17649 ( 
.A(n_17190),
.Y(n_17649)
);

OR2x2_ASAP7_75t_L g17650 ( 
.A(n_17284),
.B(n_17110),
.Y(n_17650)
);

AOI322xp5_ASAP7_75t_L g17651 ( 
.A1(n_17267),
.A2(n_16761),
.A3(n_16819),
.B1(n_17093),
.B2(n_17009),
.C1(n_16987),
.C2(n_17068),
.Y(n_17651)
);

INVx2_ASAP7_75t_L g17652 ( 
.A(n_17187),
.Y(n_17652)
);

INVx1_ASAP7_75t_SL g17653 ( 
.A(n_17375),
.Y(n_17653)
);

NAND2xp5_ASAP7_75t_L g17654 ( 
.A(n_17258),
.B(n_17127),
.Y(n_17654)
);

INVx1_ASAP7_75t_L g17655 ( 
.A(n_17192),
.Y(n_17655)
);

OR2x2_ASAP7_75t_L g17656 ( 
.A(n_17299),
.B(n_17469),
.Y(n_17656)
);

AND2x2_ASAP7_75t_L g17657 ( 
.A(n_17404),
.B(n_17105),
.Y(n_17657)
);

INVx1_ASAP7_75t_L g17658 ( 
.A(n_17219),
.Y(n_17658)
);

NAND2xp5_ASAP7_75t_L g17659 ( 
.A(n_17301),
.B(n_17159),
.Y(n_17659)
);

INVx2_ASAP7_75t_SL g17660 ( 
.A(n_17206),
.Y(n_17660)
);

NAND2xp5_ASAP7_75t_L g17661 ( 
.A(n_17196),
.B(n_16950),
.Y(n_17661)
);

AOI33xp33_ASAP7_75t_L g17662 ( 
.A1(n_17203),
.A2(n_16822),
.A3(n_17036),
.B1(n_17054),
.B2(n_17051),
.B3(n_17169),
.Y(n_17662)
);

INVx1_ASAP7_75t_SL g17663 ( 
.A(n_17314),
.Y(n_17663)
);

OR2x2_ASAP7_75t_L g17664 ( 
.A(n_17217),
.B(n_17134),
.Y(n_17664)
);

OR2x2_ASAP7_75t_L g17665 ( 
.A(n_17259),
.B(n_9586),
.Y(n_17665)
);

INVxp67_ASAP7_75t_L g17666 ( 
.A(n_17581),
.Y(n_17666)
);

AND2x2_ASAP7_75t_L g17667 ( 
.A(n_17221),
.B(n_17251),
.Y(n_17667)
);

INVx1_ASAP7_75t_SL g17668 ( 
.A(n_17526),
.Y(n_17668)
);

NOR2xp33_ASAP7_75t_L g17669 ( 
.A(n_17344),
.B(n_17003),
.Y(n_17669)
);

INVxp67_ASAP7_75t_L g17670 ( 
.A(n_17582),
.Y(n_17670)
);

OR2x2_ASAP7_75t_L g17671 ( 
.A(n_17230),
.B(n_9586),
.Y(n_17671)
);

INVx1_ASAP7_75t_L g17672 ( 
.A(n_17249),
.Y(n_17672)
);

INVx5_ASAP7_75t_L g17673 ( 
.A(n_17188),
.Y(n_17673)
);

NOR2x1_ASAP7_75t_L g17674 ( 
.A(n_17447),
.B(n_17264),
.Y(n_17674)
);

INVxp67_ASAP7_75t_SL g17675 ( 
.A(n_17239),
.Y(n_17675)
);

BUFx2_ASAP7_75t_L g17676 ( 
.A(n_17200),
.Y(n_17676)
);

INVx1_ASAP7_75t_L g17677 ( 
.A(n_17236),
.Y(n_17677)
);

NAND2xp5_ASAP7_75t_L g17678 ( 
.A(n_17286),
.B(n_10562),
.Y(n_17678)
);

NAND2xp5_ASAP7_75t_L g17679 ( 
.A(n_17348),
.B(n_10564),
.Y(n_17679)
);

NAND2x1p5_ASAP7_75t_L g17680 ( 
.A(n_17498),
.B(n_7894),
.Y(n_17680)
);

OR3x1_ASAP7_75t_L g17681 ( 
.A(n_17380),
.B(n_17057),
.C(n_10575),
.Y(n_17681)
);

AOI31xp33_ASAP7_75t_L g17682 ( 
.A1(n_17247),
.A2(n_7984),
.A3(n_8002),
.B(n_7942),
.Y(n_17682)
);

INVx2_ASAP7_75t_SL g17683 ( 
.A(n_17200),
.Y(n_17683)
);

NAND2xp5_ASAP7_75t_L g17684 ( 
.A(n_17244),
.B(n_17252),
.Y(n_17684)
);

OR2x2_ASAP7_75t_L g17685 ( 
.A(n_17223),
.B(n_9586),
.Y(n_17685)
);

INVx1_ASAP7_75t_L g17686 ( 
.A(n_17229),
.Y(n_17686)
);

INVx1_ASAP7_75t_SL g17687 ( 
.A(n_17464),
.Y(n_17687)
);

AOI22xp33_ASAP7_75t_L g17688 ( 
.A1(n_17291),
.A2(n_17305),
.B1(n_17321),
.B2(n_17320),
.Y(n_17688)
);

AND2x2_ASAP7_75t_L g17689 ( 
.A(n_17253),
.B(n_11376),
.Y(n_17689)
);

AND2x2_ASAP7_75t_L g17690 ( 
.A(n_17255),
.B(n_11376),
.Y(n_17690)
);

INVxp67_ASAP7_75t_L g17691 ( 
.A(n_17509),
.Y(n_17691)
);

NOR2xp33_ASAP7_75t_L g17692 ( 
.A(n_17298),
.B(n_8829),
.Y(n_17692)
);

NAND2xp5_ASAP7_75t_L g17693 ( 
.A(n_17210),
.B(n_10564),
.Y(n_17693)
);

OR2x2_ASAP7_75t_L g17694 ( 
.A(n_17193),
.B(n_9588),
.Y(n_17694)
);

NAND2xp33_ASAP7_75t_SL g17695 ( 
.A(n_17300),
.B(n_8980),
.Y(n_17695)
);

INVx2_ASAP7_75t_L g17696 ( 
.A(n_17421),
.Y(n_17696)
);

INVx1_ASAP7_75t_L g17697 ( 
.A(n_17222),
.Y(n_17697)
);

INVx1_ASAP7_75t_L g17698 ( 
.A(n_17261),
.Y(n_17698)
);

AND2x2_ASAP7_75t_L g17699 ( 
.A(n_17371),
.B(n_11440),
.Y(n_17699)
);

INVx1_ASAP7_75t_L g17700 ( 
.A(n_17289),
.Y(n_17700)
);

NAND5xp2_ASAP7_75t_SL g17701 ( 
.A(n_17336),
.B(n_8564),
.C(n_8567),
.D(n_8520),
.E(n_8490),
.Y(n_17701)
);

NAND2xp33_ASAP7_75t_SL g17702 ( 
.A(n_17389),
.B(n_8980),
.Y(n_17702)
);

NOR2xp33_ASAP7_75t_R g17703 ( 
.A(n_17364),
.B(n_7894),
.Y(n_17703)
);

AND2x2_ASAP7_75t_L g17704 ( 
.A(n_17530),
.B(n_11465),
.Y(n_17704)
);

INVx2_ASAP7_75t_SL g17705 ( 
.A(n_17271),
.Y(n_17705)
);

NAND2xp5_ASAP7_75t_L g17706 ( 
.A(n_17501),
.B(n_10575),
.Y(n_17706)
);

INVx1_ASAP7_75t_SL g17707 ( 
.A(n_17514),
.Y(n_17707)
);

AOI22xp5_ASAP7_75t_L g17708 ( 
.A1(n_17436),
.A2(n_9022),
.B1(n_9065),
.B2(n_8980),
.Y(n_17708)
);

INVxp67_ASAP7_75t_L g17709 ( 
.A(n_17394),
.Y(n_17709)
);

INVx1_ASAP7_75t_L g17710 ( 
.A(n_17479),
.Y(n_17710)
);

AND2x2_ASAP7_75t_L g17711 ( 
.A(n_17381),
.B(n_17311),
.Y(n_17711)
);

NOR2xp33_ASAP7_75t_L g17712 ( 
.A(n_17352),
.B(n_8980),
.Y(n_17712)
);

AND2x2_ASAP7_75t_L g17713 ( 
.A(n_17410),
.B(n_11465),
.Y(n_17713)
);

INVx2_ASAP7_75t_L g17714 ( 
.A(n_17287),
.Y(n_17714)
);

NAND2xp5_ASAP7_75t_L g17715 ( 
.A(n_17537),
.B(n_10578),
.Y(n_17715)
);

AND2x4_ASAP7_75t_L g17716 ( 
.A(n_17561),
.B(n_9022),
.Y(n_17716)
);

INVx1_ASAP7_75t_L g17717 ( 
.A(n_17292),
.Y(n_17717)
);

INVx2_ASAP7_75t_L g17718 ( 
.A(n_17243),
.Y(n_17718)
);

AND2x2_ASAP7_75t_L g17719 ( 
.A(n_17461),
.B(n_11520),
.Y(n_17719)
);

INVx1_ASAP7_75t_L g17720 ( 
.A(n_17207),
.Y(n_17720)
);

AND2x2_ASAP7_75t_L g17721 ( 
.A(n_17475),
.B(n_11520),
.Y(n_17721)
);

NAND2xp5_ASAP7_75t_L g17722 ( 
.A(n_17324),
.B(n_10578),
.Y(n_17722)
);

NAND2xp5_ASAP7_75t_L g17723 ( 
.A(n_17347),
.B(n_10581),
.Y(n_17723)
);

AND2x2_ASAP7_75t_SL g17724 ( 
.A(n_17449),
.B(n_17506),
.Y(n_17724)
);

INVx1_ASAP7_75t_L g17725 ( 
.A(n_17204),
.Y(n_17725)
);

AND2x2_ASAP7_75t_L g17726 ( 
.A(n_17502),
.B(n_17559),
.Y(n_17726)
);

INVx2_ASAP7_75t_L g17727 ( 
.A(n_17232),
.Y(n_17727)
);

NAND2xp5_ASAP7_75t_L g17728 ( 
.A(n_17470),
.B(n_10581),
.Y(n_17728)
);

NAND2xp5_ASAP7_75t_L g17729 ( 
.A(n_17452),
.B(n_10584),
.Y(n_17729)
);

INVx2_ASAP7_75t_SL g17730 ( 
.A(n_17513),
.Y(n_17730)
);

NAND2xp5_ASAP7_75t_L g17731 ( 
.A(n_17557),
.B(n_10584),
.Y(n_17731)
);

OR2x2_ASAP7_75t_L g17732 ( 
.A(n_17328),
.B(n_9588),
.Y(n_17732)
);

INVx1_ASAP7_75t_L g17733 ( 
.A(n_17202),
.Y(n_17733)
);

AND2x2_ASAP7_75t_L g17734 ( 
.A(n_17427),
.B(n_11542),
.Y(n_17734)
);

INVx2_ASAP7_75t_L g17735 ( 
.A(n_17458),
.Y(n_17735)
);

HB1xp67_ASAP7_75t_L g17736 ( 
.A(n_17521),
.Y(n_17736)
);

NAND2xp5_ASAP7_75t_L g17737 ( 
.A(n_17205),
.B(n_17356),
.Y(n_17737)
);

INVx1_ASAP7_75t_L g17738 ( 
.A(n_17279),
.Y(n_17738)
);

INVx1_ASAP7_75t_L g17739 ( 
.A(n_17304),
.Y(n_17739)
);

INVx1_ASAP7_75t_L g17740 ( 
.A(n_17430),
.Y(n_17740)
);

NAND2xp5_ASAP7_75t_L g17741 ( 
.A(n_17361),
.B(n_10586),
.Y(n_17741)
);

OR2x2_ASAP7_75t_L g17742 ( 
.A(n_17517),
.B(n_9588),
.Y(n_17742)
);

OAI211xp5_ASAP7_75t_SL g17743 ( 
.A1(n_17270),
.A2(n_9065),
.B(n_9205),
.C(n_9022),
.Y(n_17743)
);

HB1xp67_ASAP7_75t_L g17744 ( 
.A(n_17472),
.Y(n_17744)
);

OR2x2_ASAP7_75t_L g17745 ( 
.A(n_17520),
.B(n_9589),
.Y(n_17745)
);

NAND2xp5_ASAP7_75t_L g17746 ( 
.A(n_17531),
.B(n_10586),
.Y(n_17746)
);

NOR2xp67_ASAP7_75t_SL g17747 ( 
.A(n_17411),
.B(n_7582),
.Y(n_17747)
);

NOR3xp33_ASAP7_75t_L g17748 ( 
.A(n_17191),
.B(n_9065),
.C(n_9022),
.Y(n_17748)
);

INVx1_ASAP7_75t_L g17749 ( 
.A(n_17294),
.Y(n_17749)
);

BUFx3_ASAP7_75t_L g17750 ( 
.A(n_17391),
.Y(n_17750)
);

NAND2xp5_ASAP7_75t_L g17751 ( 
.A(n_17535),
.B(n_10596),
.Y(n_17751)
);

AND2x4_ASAP7_75t_L g17752 ( 
.A(n_17554),
.B(n_9065),
.Y(n_17752)
);

NOR2x1_ASAP7_75t_L g17753 ( 
.A(n_17438),
.B(n_10596),
.Y(n_17753)
);

OR2x2_ASAP7_75t_L g17754 ( 
.A(n_17593),
.B(n_9589),
.Y(n_17754)
);

HB1xp67_ASAP7_75t_L g17755 ( 
.A(n_17472),
.Y(n_17755)
);

INVx1_ASAP7_75t_L g17756 ( 
.A(n_17295),
.Y(n_17756)
);

NAND3xp33_ASAP7_75t_L g17757 ( 
.A(n_17272),
.B(n_10447),
.C(n_9205),
.Y(n_17757)
);

OR2x2_ASAP7_75t_L g17758 ( 
.A(n_17596),
.B(n_9589),
.Y(n_17758)
);

INVx1_ASAP7_75t_L g17759 ( 
.A(n_17492),
.Y(n_17759)
);

AND2x2_ASAP7_75t_L g17760 ( 
.A(n_17598),
.B(n_11542),
.Y(n_17760)
);

AO21x2_ASAP7_75t_L g17761 ( 
.A1(n_17345),
.A2(n_11293),
.B(n_11284),
.Y(n_17761)
);

INVx1_ASAP7_75t_L g17762 ( 
.A(n_17529),
.Y(n_17762)
);

AND2x2_ASAP7_75t_L g17763 ( 
.A(n_17556),
.B(n_11561),
.Y(n_17763)
);

AND3x1_ASAP7_75t_L g17764 ( 
.A(n_17370),
.B(n_9205),
.C(n_9065),
.Y(n_17764)
);

NOR2xp33_ASAP7_75t_L g17765 ( 
.A(n_17478),
.B(n_9205),
.Y(n_17765)
);

OR2x2_ASAP7_75t_L g17766 ( 
.A(n_17483),
.B(n_9594),
.Y(n_17766)
);

AND2x2_ASAP7_75t_L g17767 ( 
.A(n_17606),
.B(n_11561),
.Y(n_17767)
);

OR2x2_ASAP7_75t_L g17768 ( 
.A(n_17433),
.B(n_9594),
.Y(n_17768)
);

NAND2xp5_ASAP7_75t_L g17769 ( 
.A(n_17441),
.B(n_10597),
.Y(n_17769)
);

NAND4xp25_ASAP7_75t_L g17770 ( 
.A(n_17525),
.B(n_7905),
.C(n_9172),
.D(n_9014),
.Y(n_17770)
);

OR2x6_ASAP7_75t_L g17771 ( 
.A(n_17434),
.B(n_7905),
.Y(n_17771)
);

AND2x4_ASAP7_75t_L g17772 ( 
.A(n_17608),
.B(n_9205),
.Y(n_17772)
);

INVx1_ASAP7_75t_L g17773 ( 
.A(n_17337),
.Y(n_17773)
);

OR2x2_ASAP7_75t_L g17774 ( 
.A(n_17338),
.B(n_9594),
.Y(n_17774)
);

NOR2xp33_ASAP7_75t_R g17775 ( 
.A(n_17339),
.B(n_7905),
.Y(n_17775)
);

AND2x2_ASAP7_75t_SL g17776 ( 
.A(n_17451),
.B(n_9014),
.Y(n_17776)
);

AND2x2_ASAP7_75t_L g17777 ( 
.A(n_17485),
.B(n_11579),
.Y(n_17777)
);

AND2x2_ASAP7_75t_L g17778 ( 
.A(n_17468),
.B(n_11579),
.Y(n_17778)
);

NOR2x1_ASAP7_75t_L g17779 ( 
.A(n_17494),
.B(n_10597),
.Y(n_17779)
);

OR2x2_ASAP7_75t_L g17780 ( 
.A(n_17343),
.B(n_9603),
.Y(n_17780)
);

INVx1_ASAP7_75t_L g17781 ( 
.A(n_17618),
.Y(n_17781)
);

NAND2xp33_ASAP7_75t_R g17782 ( 
.A(n_17402),
.B(n_8386),
.Y(n_17782)
);

AND2x2_ASAP7_75t_L g17783 ( 
.A(n_17420),
.B(n_11588),
.Y(n_17783)
);

AND2x2_ASAP7_75t_L g17784 ( 
.A(n_17609),
.B(n_11588),
.Y(n_17784)
);

NAND3xp33_ASAP7_75t_L g17785 ( 
.A(n_17189),
.B(n_9611),
.C(n_9603),
.Y(n_17785)
);

AND3x1_ASAP7_75t_L g17786 ( 
.A(n_17275),
.B(n_8053),
.C(n_7916),
.Y(n_17786)
);

NAND3xp33_ASAP7_75t_L g17787 ( 
.A(n_17431),
.B(n_9611),
.C(n_9603),
.Y(n_17787)
);

NAND2xp33_ASAP7_75t_SL g17788 ( 
.A(n_17412),
.B(n_9035),
.Y(n_17788)
);

INVx1_ASAP7_75t_L g17789 ( 
.A(n_17497),
.Y(n_17789)
);

OR2x2_ASAP7_75t_L g17790 ( 
.A(n_17365),
.B(n_9611),
.Y(n_17790)
);

OR2x2_ASAP7_75t_L g17791 ( 
.A(n_17366),
.B(n_9622),
.Y(n_17791)
);

NAND2xp5_ASAP7_75t_L g17792 ( 
.A(n_17499),
.B(n_10600),
.Y(n_17792)
);

INVx2_ASAP7_75t_L g17793 ( 
.A(n_17465),
.Y(n_17793)
);

INVx1_ASAP7_75t_L g17794 ( 
.A(n_17505),
.Y(n_17794)
);

OR2x2_ASAP7_75t_L g17795 ( 
.A(n_17367),
.B(n_9622),
.Y(n_17795)
);

NAND2xp5_ASAP7_75t_L g17796 ( 
.A(n_17516),
.B(n_10600),
.Y(n_17796)
);

INVx1_ASAP7_75t_L g17797 ( 
.A(n_17443),
.Y(n_17797)
);

CKINVDCx20_ASAP7_75t_R g17798 ( 
.A(n_17330),
.Y(n_17798)
);

INVx1_ASAP7_75t_L g17799 ( 
.A(n_17369),
.Y(n_17799)
);

OR2x4_ASAP7_75t_L g17800 ( 
.A(n_17315),
.B(n_8903),
.Y(n_17800)
);

AND2x2_ASAP7_75t_L g17801 ( 
.A(n_17425),
.B(n_11637),
.Y(n_17801)
);

AND2x2_ASAP7_75t_L g17802 ( 
.A(n_17313),
.B(n_11637),
.Y(n_17802)
);

AND2x2_ASAP7_75t_L g17803 ( 
.A(n_17333),
.B(n_11696),
.Y(n_17803)
);

NOR2xp33_ASAP7_75t_L g17804 ( 
.A(n_17372),
.B(n_10603),
.Y(n_17804)
);

AND2x2_ASAP7_75t_L g17805 ( 
.A(n_17351),
.B(n_11696),
.Y(n_17805)
);

AND2x2_ASAP7_75t_SL g17806 ( 
.A(n_17487),
.B(n_9014),
.Y(n_17806)
);

OAI21xp5_ASAP7_75t_L g17807 ( 
.A1(n_17309),
.A2(n_11713),
.B(n_10871),
.Y(n_17807)
);

OR2x2_ASAP7_75t_L g17808 ( 
.A(n_17377),
.B(n_17382),
.Y(n_17808)
);

AND2x2_ASAP7_75t_L g17809 ( 
.A(n_17332),
.B(n_11713),
.Y(n_17809)
);

INVx1_ASAP7_75t_L g17810 ( 
.A(n_17390),
.Y(n_17810)
);

NAND2xp5_ASAP7_75t_L g17811 ( 
.A(n_17405),
.B(n_10603),
.Y(n_17811)
);

OR2x2_ASAP7_75t_L g17812 ( 
.A(n_17401),
.B(n_9622),
.Y(n_17812)
);

AOI31xp33_ASAP7_75t_L g17813 ( 
.A1(n_17403),
.A2(n_7942),
.A3(n_8007),
.B(n_8002),
.Y(n_17813)
);

NAND2xp5_ASAP7_75t_L g17814 ( 
.A(n_17414),
.B(n_10606),
.Y(n_17814)
);

AND2x2_ASAP7_75t_L g17815 ( 
.A(n_17308),
.B(n_17571),
.Y(n_17815)
);

AND2x2_ASAP7_75t_L g17816 ( 
.A(n_17571),
.B(n_11323),
.Y(n_17816)
);

INVx2_ASAP7_75t_SL g17817 ( 
.A(n_17546),
.Y(n_17817)
);

INVxp67_ASAP7_75t_L g17818 ( 
.A(n_17399),
.Y(n_17818)
);

AND2x2_ASAP7_75t_L g17819 ( 
.A(n_17316),
.B(n_11343),
.Y(n_17819)
);

NOR2xp33_ASAP7_75t_L g17820 ( 
.A(n_17418),
.B(n_17422),
.Y(n_17820)
);

AND2x4_ASAP7_75t_L g17821 ( 
.A(n_17423),
.B(n_17428),
.Y(n_17821)
);

INVx2_ASAP7_75t_L g17822 ( 
.A(n_17266),
.Y(n_17822)
);

OR2x2_ASAP7_75t_L g17823 ( 
.A(n_17429),
.B(n_9625),
.Y(n_17823)
);

INVx3_ASAP7_75t_SL g17824 ( 
.A(n_17325),
.Y(n_17824)
);

NAND2xp5_ASAP7_75t_L g17825 ( 
.A(n_17456),
.B(n_10606),
.Y(n_17825)
);

NAND2xp5_ASAP7_75t_L g17826 ( 
.A(n_17474),
.B(n_10607),
.Y(n_17826)
);

NAND3xp33_ASAP7_75t_L g17827 ( 
.A(n_17432),
.B(n_9638),
.C(n_9625),
.Y(n_17827)
);

INVx1_ASAP7_75t_L g17828 ( 
.A(n_17573),
.Y(n_17828)
);

OR2x2_ASAP7_75t_L g17829 ( 
.A(n_17562),
.B(n_9625),
.Y(n_17829)
);

INVx2_ASAP7_75t_SL g17830 ( 
.A(n_17303),
.Y(n_17830)
);

AND2x2_ASAP7_75t_L g17831 ( 
.A(n_17476),
.B(n_11343),
.Y(n_17831)
);

AND2x2_ASAP7_75t_L g17832 ( 
.A(n_17477),
.B(n_11348),
.Y(n_17832)
);

NAND2xp5_ASAP7_75t_L g17833 ( 
.A(n_17454),
.B(n_10607),
.Y(n_17833)
);

INVx1_ASAP7_75t_L g17834 ( 
.A(n_17455),
.Y(n_17834)
);

OR2x2_ASAP7_75t_L g17835 ( 
.A(n_17567),
.B(n_9638),
.Y(n_17835)
);

INVx2_ASAP7_75t_L g17836 ( 
.A(n_17266),
.Y(n_17836)
);

AND2x2_ASAP7_75t_L g17837 ( 
.A(n_17310),
.B(n_11348),
.Y(n_17837)
);

AND2x2_ASAP7_75t_L g17838 ( 
.A(n_17549),
.B(n_10852),
.Y(n_17838)
);

INVx1_ASAP7_75t_L g17839 ( 
.A(n_17335),
.Y(n_17839)
);

NOR3xp33_ASAP7_75t_L g17840 ( 
.A(n_17480),
.B(n_9939),
.C(n_9906),
.Y(n_17840)
);

NAND2xp5_ASAP7_75t_SL g17841 ( 
.A(n_17234),
.B(n_10852),
.Y(n_17841)
);

OAI211xp5_ASAP7_75t_L g17842 ( 
.A1(n_17553),
.A2(n_7582),
.B(n_7809),
.C(n_10871),
.Y(n_17842)
);

NAND2xp5_ASAP7_75t_L g17843 ( 
.A(n_17450),
.B(n_10614),
.Y(n_17843)
);

NAND2xp5_ASAP7_75t_L g17844 ( 
.A(n_17595),
.B(n_10614),
.Y(n_17844)
);

AND2x2_ASAP7_75t_L g17845 ( 
.A(n_17379),
.B(n_10877),
.Y(n_17845)
);

AND2x2_ASAP7_75t_L g17846 ( 
.A(n_17392),
.B(n_10877),
.Y(n_17846)
);

NAND3xp33_ASAP7_75t_SL g17847 ( 
.A(n_17376),
.B(n_8725),
.C(n_8667),
.Y(n_17847)
);

NAND2xp5_ASAP7_75t_L g17848 ( 
.A(n_17349),
.B(n_10615),
.Y(n_17848)
);

INVxp67_ASAP7_75t_L g17849 ( 
.A(n_17257),
.Y(n_17849)
);

INVx1_ASAP7_75t_L g17850 ( 
.A(n_17240),
.Y(n_17850)
);

HB1xp67_ASAP7_75t_L g17851 ( 
.A(n_17510),
.Y(n_17851)
);

NAND2xp5_ASAP7_75t_L g17852 ( 
.A(n_17490),
.B(n_10615),
.Y(n_17852)
);

NAND2xp5_ASAP7_75t_L g17853 ( 
.A(n_17528),
.B(n_10616),
.Y(n_17853)
);

NOR2xp33_ASAP7_75t_L g17854 ( 
.A(n_17584),
.B(n_10616),
.Y(n_17854)
);

INVx1_ASAP7_75t_L g17855 ( 
.A(n_17225),
.Y(n_17855)
);

AOI21xp33_ASAP7_75t_L g17856 ( 
.A1(n_17599),
.A2(n_10105),
.B(n_10015),
.Y(n_17856)
);

NAND3xp33_ASAP7_75t_L g17857 ( 
.A(n_17245),
.B(n_9647),
.C(n_9638),
.Y(n_17857)
);

NAND2xp5_ASAP7_75t_L g17858 ( 
.A(n_17538),
.B(n_10617),
.Y(n_17858)
);

NAND2xp5_ASAP7_75t_L g17859 ( 
.A(n_17539),
.B(n_10617),
.Y(n_17859)
);

INVxp67_ASAP7_75t_L g17860 ( 
.A(n_17280),
.Y(n_17860)
);

NAND2xp5_ASAP7_75t_L g17861 ( 
.A(n_17585),
.B(n_10620),
.Y(n_17861)
);

NAND2xp5_ASAP7_75t_L g17862 ( 
.A(n_17588),
.B(n_10620),
.Y(n_17862)
);

NAND2xp5_ASAP7_75t_L g17863 ( 
.A(n_17590),
.B(n_17597),
.Y(n_17863)
);

OR2x2_ASAP7_75t_L g17864 ( 
.A(n_17533),
.B(n_9647),
.Y(n_17864)
);

OAI211xp5_ASAP7_75t_SL g17865 ( 
.A1(n_17511),
.A2(n_7809),
.B(n_9653),
.C(n_9647),
.Y(n_17865)
);

AND2x2_ASAP7_75t_L g17866 ( 
.A(n_17426),
.B(n_10884),
.Y(n_17866)
);

NOR2xp33_ASAP7_75t_L g17867 ( 
.A(n_17600),
.B(n_10621),
.Y(n_17867)
);

INVx1_ASAP7_75t_SL g17868 ( 
.A(n_17360),
.Y(n_17868)
);

NAND2xp5_ASAP7_75t_L g17869 ( 
.A(n_17543),
.B(n_10621),
.Y(n_17869)
);

OR2x2_ASAP7_75t_L g17870 ( 
.A(n_17527),
.B(n_9653),
.Y(n_17870)
);

AOI22xp33_ASAP7_75t_L g17871 ( 
.A1(n_17277),
.A2(n_8386),
.B1(n_8762),
.B2(n_8760),
.Y(n_17871)
);

NAND2xp5_ASAP7_75t_L g17872 ( 
.A(n_17544),
.B(n_10623),
.Y(n_17872)
);

AND2x2_ASAP7_75t_L g17873 ( 
.A(n_17440),
.B(n_10884),
.Y(n_17873)
);

OR2x2_ASAP7_75t_L g17874 ( 
.A(n_17524),
.B(n_9653),
.Y(n_17874)
);

AND2x2_ASAP7_75t_L g17875 ( 
.A(n_17442),
.B(n_10015),
.Y(n_17875)
);

AOI321xp33_ASAP7_75t_L g17876 ( 
.A1(n_17398),
.A2(n_9172),
.A3(n_9014),
.B1(n_8092),
.B2(n_8050),
.C(n_8749),
.Y(n_17876)
);

INVxp67_ASAP7_75t_L g17877 ( 
.A(n_17285),
.Y(n_17877)
);

INVx1_ASAP7_75t_L g17878 ( 
.A(n_17242),
.Y(n_17878)
);

NAND4xp25_ASAP7_75t_L g17879 ( 
.A(n_17569),
.B(n_9172),
.C(n_9014),
.D(n_7153),
.Y(n_17879)
);

AND2x4_ASAP7_75t_L g17880 ( 
.A(n_17603),
.B(n_8138),
.Y(n_17880)
);

OR2x2_ASAP7_75t_L g17881 ( 
.A(n_17495),
.B(n_9673),
.Y(n_17881)
);

OR2x2_ASAP7_75t_L g17882 ( 
.A(n_17208),
.B(n_17256),
.Y(n_17882)
);

OR2x6_ASAP7_75t_L g17883 ( 
.A(n_17545),
.B(n_8477),
.Y(n_17883)
);

AND2x2_ASAP7_75t_L g17884 ( 
.A(n_17363),
.B(n_10105),
.Y(n_17884)
);

AND2x2_ASAP7_75t_SL g17885 ( 
.A(n_17550),
.B(n_9014),
.Y(n_17885)
);

NOR2xp33_ASAP7_75t_L g17886 ( 
.A(n_17552),
.B(n_10623),
.Y(n_17886)
);

AND2x2_ASAP7_75t_L g17887 ( 
.A(n_17471),
.B(n_10920),
.Y(n_17887)
);

NOR2x1_ASAP7_75t_L g17888 ( 
.A(n_17558),
.B(n_10627),
.Y(n_17888)
);

NAND2xp33_ASAP7_75t_R g17889 ( 
.A(n_17541),
.B(n_8572),
.Y(n_17889)
);

NOR2xp33_ASAP7_75t_R g17890 ( 
.A(n_17564),
.B(n_9048),
.Y(n_17890)
);

OR2x2_ASAP7_75t_L g17891 ( 
.A(n_17273),
.B(n_9673),
.Y(n_17891)
);

OR2x2_ASAP7_75t_L g17892 ( 
.A(n_17322),
.B(n_9673),
.Y(n_17892)
);

INVx1_ASAP7_75t_L g17893 ( 
.A(n_17265),
.Y(n_17893)
);

INVx2_ASAP7_75t_L g17894 ( 
.A(n_17568),
.Y(n_17894)
);

INVx1_ASAP7_75t_L g17895 ( 
.A(n_17444),
.Y(n_17895)
);

OAI211xp5_ASAP7_75t_SL g17896 ( 
.A1(n_17565),
.A2(n_7809),
.B(n_9685),
.C(n_9682),
.Y(n_17896)
);

NOR2x1_ASAP7_75t_L g17897 ( 
.A(n_17574),
.B(n_17580),
.Y(n_17897)
);

NAND2xp5_ASAP7_75t_L g17898 ( 
.A(n_17583),
.B(n_17605),
.Y(n_17898)
);

AND2x2_ASAP7_75t_L g17899 ( 
.A(n_17542),
.B(n_10953),
.Y(n_17899)
);

HB1xp67_ASAP7_75t_L g17900 ( 
.A(n_17512),
.Y(n_17900)
);

OR2x2_ASAP7_75t_L g17901 ( 
.A(n_17467),
.B(n_9682),
.Y(n_17901)
);

INVx1_ASAP7_75t_L g17902 ( 
.A(n_17359),
.Y(n_17902)
);

INVx1_ASAP7_75t_L g17903 ( 
.A(n_17373),
.Y(n_17903)
);

AND2x2_ASAP7_75t_L g17904 ( 
.A(n_17496),
.B(n_10954),
.Y(n_17904)
);

INVx2_ASAP7_75t_L g17905 ( 
.A(n_17326),
.Y(n_17905)
);

AND2x4_ASAP7_75t_L g17906 ( 
.A(n_17551),
.B(n_8164),
.Y(n_17906)
);

INVx2_ASAP7_75t_L g17907 ( 
.A(n_17331),
.Y(n_17907)
);

INVx2_ASAP7_75t_L g17908 ( 
.A(n_17586),
.Y(n_17908)
);

INVx4_ASAP7_75t_L g17909 ( 
.A(n_17384),
.Y(n_17909)
);

INVx1_ASAP7_75t_L g17910 ( 
.A(n_17374),
.Y(n_17910)
);

INVxp67_ASAP7_75t_L g17911 ( 
.A(n_17500),
.Y(n_17911)
);

AND2x2_ASAP7_75t_L g17912 ( 
.A(n_17575),
.B(n_17578),
.Y(n_17912)
);

OR2x2_ASAP7_75t_L g17913 ( 
.A(n_17457),
.B(n_9682),
.Y(n_17913)
);

INVx1_ASAP7_75t_L g17914 ( 
.A(n_17350),
.Y(n_17914)
);

OR2x2_ASAP7_75t_L g17915 ( 
.A(n_17459),
.B(n_9685),
.Y(n_17915)
);

OR2x2_ASAP7_75t_L g17916 ( 
.A(n_17462),
.B(n_9685),
.Y(n_17916)
);

INVx1_ASAP7_75t_L g17917 ( 
.A(n_17396),
.Y(n_17917)
);

INVx2_ASAP7_75t_L g17918 ( 
.A(n_17613),
.Y(n_17918)
);

INVx1_ASAP7_75t_L g17919 ( 
.A(n_17319),
.Y(n_17919)
);

INVx1_ASAP7_75t_SL g17920 ( 
.A(n_17388),
.Y(n_17920)
);

HB1xp67_ASAP7_75t_L g17921 ( 
.A(n_17481),
.Y(n_17921)
);

AND2x4_ASAP7_75t_SL g17922 ( 
.A(n_17296),
.B(n_9048),
.Y(n_17922)
);

AND2x2_ASAP7_75t_L g17923 ( 
.A(n_17616),
.B(n_10970),
.Y(n_17923)
);

INVx1_ASAP7_75t_L g17924 ( 
.A(n_17317),
.Y(n_17924)
);

NAND2xp5_ASAP7_75t_L g17925 ( 
.A(n_17395),
.B(n_10627),
.Y(n_17925)
);

NAND2x1p5_ASAP7_75t_L g17926 ( 
.A(n_17288),
.B(n_8667),
.Y(n_17926)
);

INVx1_ASAP7_75t_SL g17927 ( 
.A(n_17482),
.Y(n_17927)
);

NAND2xp5_ASAP7_75t_L g17928 ( 
.A(n_17540),
.B(n_10630),
.Y(n_17928)
);

NAND2xp5_ASAP7_75t_L g17929 ( 
.A(n_17548),
.B(n_10630),
.Y(n_17929)
);

AND2x4_ASAP7_75t_L g17930 ( 
.A(n_17378),
.B(n_8164),
.Y(n_17930)
);

NAND2xp33_ASAP7_75t_SL g17931 ( 
.A(n_17417),
.B(n_9035),
.Y(n_17931)
);

NAND2xp5_ASAP7_75t_L g17932 ( 
.A(n_17576),
.B(n_10639),
.Y(n_17932)
);

INVx1_ASAP7_75t_L g17933 ( 
.A(n_17387),
.Y(n_17933)
);

AND2x2_ASAP7_75t_L g17934 ( 
.A(n_17439),
.B(n_7114),
.Y(n_17934)
);

AND2x4_ASAP7_75t_L g17935 ( 
.A(n_17199),
.B(n_8164),
.Y(n_17935)
);

INVx1_ASAP7_75t_L g17936 ( 
.A(n_17579),
.Y(n_17936)
);

INVx1_ASAP7_75t_L g17937 ( 
.A(n_17570),
.Y(n_17937)
);

NAND2xp5_ASAP7_75t_L g17938 ( 
.A(n_17592),
.B(n_10639),
.Y(n_17938)
);

NAND2xp5_ASAP7_75t_L g17939 ( 
.A(n_17607),
.B(n_10643),
.Y(n_17939)
);

AND2x4_ASAP7_75t_L g17940 ( 
.A(n_17235),
.B(n_8172),
.Y(n_17940)
);

NAND2xp33_ASAP7_75t_L g17941 ( 
.A(n_17393),
.B(n_9054),
.Y(n_17941)
);

INVxp67_ASAP7_75t_SL g17942 ( 
.A(n_17619),
.Y(n_17942)
);

AND2x4_ASAP7_75t_L g17943 ( 
.A(n_17209),
.B(n_17282),
.Y(n_17943)
);

INVx3_ASAP7_75t_L g17944 ( 
.A(n_17610),
.Y(n_17944)
);

OAI211xp5_ASAP7_75t_SL g17945 ( 
.A1(n_17281),
.A2(n_7809),
.B(n_9689),
.C(n_9687),
.Y(n_17945)
);

INVx1_ASAP7_75t_L g17946 ( 
.A(n_17594),
.Y(n_17946)
);

NAND2xp5_ASAP7_75t_SL g17947 ( 
.A(n_17254),
.B(n_8172),
.Y(n_17947)
);

NAND2xp5_ASAP7_75t_L g17948 ( 
.A(n_17611),
.B(n_10643),
.Y(n_17948)
);

NAND2xp5_ASAP7_75t_L g17949 ( 
.A(n_17612),
.B(n_10649),
.Y(n_17949)
);

AND2x2_ASAP7_75t_L g17950 ( 
.A(n_17290),
.B(n_7114),
.Y(n_17950)
);

OR2x4_ASAP7_75t_L g17951 ( 
.A(n_17212),
.B(n_8903),
.Y(n_17951)
);

BUFx2_ASAP7_75t_L g17952 ( 
.A(n_17493),
.Y(n_17952)
);

AND2x2_ASAP7_75t_L g17953 ( 
.A(n_17248),
.B(n_7132),
.Y(n_17953)
);

INVx1_ASAP7_75t_L g17954 ( 
.A(n_17614),
.Y(n_17954)
);

AND2x2_ASAP7_75t_L g17955 ( 
.A(n_17620),
.B(n_7132),
.Y(n_17955)
);

INVx1_ASAP7_75t_L g17956 ( 
.A(n_17409),
.Y(n_17956)
);

AOI22xp5_ASAP7_75t_L g17957 ( 
.A1(n_17228),
.A2(n_8172),
.B1(n_8304),
.B2(n_8255),
.Y(n_17957)
);

NOR2x1_ASAP7_75t_R g17958 ( 
.A(n_17407),
.B(n_5627),
.Y(n_17958)
);

INVx2_ASAP7_75t_SL g17959 ( 
.A(n_17416),
.Y(n_17959)
);

NAND2xp5_ASAP7_75t_L g17960 ( 
.A(n_17408),
.B(n_17269),
.Y(n_17960)
);

HB1xp67_ASAP7_75t_L g17961 ( 
.A(n_17274),
.Y(n_17961)
);

NAND4xp25_ASAP7_75t_SL g17962 ( 
.A(n_17276),
.B(n_17218),
.C(n_17302),
.D(n_17227),
.Y(n_17962)
);

INVx1_ASAP7_75t_L g17963 ( 
.A(n_17602),
.Y(n_17963)
);

AND2x2_ASAP7_75t_L g17964 ( 
.A(n_17385),
.B(n_7132),
.Y(n_17964)
);

INVx2_ASAP7_75t_SL g17965 ( 
.A(n_17197),
.Y(n_17965)
);

NAND2xp5_ASAP7_75t_L g17966 ( 
.A(n_17323),
.B(n_10649),
.Y(n_17966)
);

INVx1_ASAP7_75t_L g17967 ( 
.A(n_17312),
.Y(n_17967)
);

INVx1_ASAP7_75t_L g17968 ( 
.A(n_17362),
.Y(n_17968)
);

BUFx2_ASAP7_75t_SL g17969 ( 
.A(n_17197),
.Y(n_17969)
);

INVx2_ASAP7_75t_SL g17970 ( 
.A(n_17604),
.Y(n_17970)
);

INVx1_ASAP7_75t_L g17971 ( 
.A(n_17260),
.Y(n_17971)
);

NOR2xp33_ASAP7_75t_L g17972 ( 
.A(n_17435),
.B(n_10652),
.Y(n_17972)
);

INVx2_ASAP7_75t_L g17973 ( 
.A(n_17329),
.Y(n_17973)
);

OR2x2_ASAP7_75t_L g17974 ( 
.A(n_17340),
.B(n_9687),
.Y(n_17974)
);

AND2x2_ASAP7_75t_L g17975 ( 
.A(n_17386),
.B(n_7132),
.Y(n_17975)
);

BUFx3_ASAP7_75t_L g17976 ( 
.A(n_17604),
.Y(n_17976)
);

OR2x2_ASAP7_75t_L g17977 ( 
.A(n_17368),
.B(n_9687),
.Y(n_17977)
);

NOR2xp33_ASAP7_75t_R g17978 ( 
.A(n_17587),
.B(n_9048),
.Y(n_17978)
);

NAND2xp5_ASAP7_75t_L g17979 ( 
.A(n_17237),
.B(n_10652),
.Y(n_17979)
);

NAND2xp5_ASAP7_75t_L g17980 ( 
.A(n_17198),
.B(n_10653),
.Y(n_17980)
);

NAND3xp33_ASAP7_75t_SL g17981 ( 
.A(n_17591),
.B(n_17446),
.C(n_17615),
.Y(n_17981)
);

NAND2xp5_ASAP7_75t_L g17982 ( 
.A(n_17617),
.B(n_17577),
.Y(n_17982)
);

INVx1_ASAP7_75t_L g17983 ( 
.A(n_17307),
.Y(n_17983)
);

INVx2_ASAP7_75t_L g17984 ( 
.A(n_17327),
.Y(n_17984)
);

AND2x2_ASAP7_75t_L g17985 ( 
.A(n_17610),
.B(n_7167),
.Y(n_17985)
);

NAND2xp5_ASAP7_75t_L g17986 ( 
.A(n_17488),
.B(n_10653),
.Y(n_17986)
);

NAND2xp5_ASAP7_75t_SL g17987 ( 
.A(n_17522),
.B(n_8255),
.Y(n_17987)
);

AND2x2_ASAP7_75t_L g17988 ( 
.A(n_17306),
.B(n_7167),
.Y(n_17988)
);

OR2x2_ASAP7_75t_L g17989 ( 
.A(n_17536),
.B(n_9689),
.Y(n_17989)
);

AND2x2_ASAP7_75t_L g17990 ( 
.A(n_17341),
.B(n_7167),
.Y(n_17990)
);

AOI211xp5_ASAP7_75t_L g17991 ( 
.A1(n_17463),
.A2(n_9906),
.B(n_9956),
.C(n_9939),
.Y(n_17991)
);

AND2x2_ASAP7_75t_L g17992 ( 
.A(n_17353),
.B(n_7167),
.Y(n_17992)
);

NOR4xp25_ASAP7_75t_SL g17993 ( 
.A(n_17400),
.B(n_10658),
.C(n_10662),
.D(n_10657),
.Y(n_17993)
);

BUFx3_ASAP7_75t_L g17994 ( 
.A(n_17589),
.Y(n_17994)
);

O2A1O1Ixp33_ASAP7_75t_L g17995 ( 
.A1(n_17445),
.A2(n_9689),
.B(n_9715),
.C(n_9705),
.Y(n_17995)
);

INVx1_ASAP7_75t_L g17996 ( 
.A(n_17503),
.Y(n_17996)
);

AOI31xp33_ASAP7_75t_SL g17997 ( 
.A1(n_17437),
.A2(n_9705),
.A3(n_9716),
.B(n_9715),
.Y(n_17997)
);

AOI32xp33_ASAP7_75t_L g17998 ( 
.A1(n_17519),
.A2(n_11069),
.A3(n_8776),
.B1(n_9099),
.B2(n_9071),
.Y(n_17998)
);

OAI33xp33_ASAP7_75t_L g17999 ( 
.A1(n_17318),
.A2(n_10674),
.A3(n_10658),
.B1(n_10675),
.B2(n_10662),
.B3(n_10657),
.Y(n_17999)
);

NAND2xp5_ASAP7_75t_L g18000 ( 
.A(n_17589),
.B(n_10674),
.Y(n_18000)
);

NOR3xp33_ASAP7_75t_L g18001 ( 
.A(n_17201),
.B(n_9956),
.C(n_10193),
.Y(n_18001)
);

NAND2xp33_ASAP7_75t_R g18002 ( 
.A(n_17519),
.B(n_8572),
.Y(n_18002)
);

INVx2_ASAP7_75t_L g18003 ( 
.A(n_17566),
.Y(n_18003)
);

NOR2xp33_ASAP7_75t_R g18004 ( 
.A(n_17566),
.B(n_9048),
.Y(n_18004)
);

NAND5xp2_ASAP7_75t_L g18005 ( 
.A(n_17563),
.B(n_7942),
.C(n_8208),
.D(n_8114),
.E(n_8007),
.Y(n_18005)
);

INVx1_ASAP7_75t_L g18006 ( 
.A(n_17241),
.Y(n_18006)
);

NOR2xp33_ASAP7_75t_L g18007 ( 
.A(n_17453),
.B(n_10675),
.Y(n_18007)
);

INVx1_ASAP7_75t_SL g18008 ( 
.A(n_17534),
.Y(n_18008)
);

AND2x2_ASAP7_75t_L g18009 ( 
.A(n_17413),
.B(n_7170),
.Y(n_18009)
);

AND2x2_ASAP7_75t_L g18010 ( 
.A(n_17601),
.B(n_7170),
.Y(n_18010)
);

INVx1_ASAP7_75t_L g18011 ( 
.A(n_17262),
.Y(n_18011)
);

AND2x2_ASAP7_75t_L g18012 ( 
.A(n_17560),
.B(n_7170),
.Y(n_18012)
);

AOI21xp33_ASAP7_75t_SL g18013 ( 
.A1(n_17518),
.A2(n_8304),
.B(n_8255),
.Y(n_18013)
);

OR2x2_ASAP7_75t_L g18014 ( 
.A(n_17555),
.B(n_9705),
.Y(n_18014)
);

NOR4xp25_ASAP7_75t_SL g18015 ( 
.A(n_17233),
.B(n_10678),
.C(n_10679),
.D(n_10676),
.Y(n_18015)
);

INVx1_ASAP7_75t_L g18016 ( 
.A(n_17346),
.Y(n_18016)
);

NAND2x1p5_ASAP7_75t_L g18017 ( 
.A(n_17534),
.B(n_8776),
.Y(n_18017)
);

NOR2xp33_ASAP7_75t_L g18018 ( 
.A(n_17283),
.B(n_10676),
.Y(n_18018)
);

AND2x2_ASAP7_75t_L g18019 ( 
.A(n_17515),
.B(n_7170),
.Y(n_18019)
);

INVx2_ASAP7_75t_L g18020 ( 
.A(n_17532),
.Y(n_18020)
);

NOR2xp33_ASAP7_75t_R g18021 ( 
.A(n_17547),
.B(n_9048),
.Y(n_18021)
);

INVx1_ASAP7_75t_L g18022 ( 
.A(n_17354),
.Y(n_18022)
);

INVx2_ASAP7_75t_L g18023 ( 
.A(n_17489),
.Y(n_18023)
);

NAND2xp33_ASAP7_75t_R g18024 ( 
.A(n_17473),
.B(n_8572),
.Y(n_18024)
);

NAND2xp5_ASAP7_75t_L g18025 ( 
.A(n_17293),
.B(n_17415),
.Y(n_18025)
);

AND2x6_ASAP7_75t_L g18026 ( 
.A(n_17357),
.B(n_9172),
.Y(n_18026)
);

NOR2xp33_ASAP7_75t_L g18027 ( 
.A(n_17523),
.B(n_10678),
.Y(n_18027)
);

OR2x2_ASAP7_75t_L g18028 ( 
.A(n_17406),
.B(n_9715),
.Y(n_18028)
);

AND2x2_ASAP7_75t_L g18029 ( 
.A(n_17466),
.B(n_17508),
.Y(n_18029)
);

INVx1_ASAP7_75t_L g18030 ( 
.A(n_17969),
.Y(n_18030)
);

AND2x2_ASAP7_75t_L g18031 ( 
.A(n_17633),
.B(n_7179),
.Y(n_18031)
);

INVx1_ASAP7_75t_L g18032 ( 
.A(n_17644),
.Y(n_18032)
);

OR2x2_ASAP7_75t_L g18033 ( 
.A(n_17762),
.B(n_9994),
.Y(n_18033)
);

NOR2xp33_ASAP7_75t_L g18034 ( 
.A(n_17652),
.B(n_17214),
.Y(n_18034)
);

AOI22xp33_ASAP7_75t_L g18035 ( 
.A1(n_17750),
.A2(n_17419),
.B1(n_17448),
.B2(n_17424),
.Y(n_18035)
);

INVx1_ASAP7_75t_L g18036 ( 
.A(n_17900),
.Y(n_18036)
);

OR2x2_ASAP7_75t_L g18037 ( 
.A(n_17668),
.B(n_9994),
.Y(n_18037)
);

NAND2xp5_ASAP7_75t_L g18038 ( 
.A(n_17673),
.B(n_10679),
.Y(n_18038)
);

AND2x2_ASAP7_75t_L g18039 ( 
.A(n_17667),
.B(n_7179),
.Y(n_18039)
);

INVx4_ASAP7_75t_L g18040 ( 
.A(n_17673),
.Y(n_18040)
);

INVx1_ASAP7_75t_L g18041 ( 
.A(n_17642),
.Y(n_18041)
);

AND2x2_ASAP7_75t_L g18042 ( 
.A(n_17726),
.B(n_7179),
.Y(n_18042)
);

INVx2_ASAP7_75t_L g18043 ( 
.A(n_18010),
.Y(n_18043)
);

NOR2xp33_ASAP7_75t_L g18044 ( 
.A(n_17691),
.B(n_17460),
.Y(n_18044)
);

NAND2xp5_ASAP7_75t_L g18045 ( 
.A(n_17673),
.B(n_17724),
.Y(n_18045)
);

INVx1_ASAP7_75t_L g18046 ( 
.A(n_17933),
.Y(n_18046)
);

OR2x2_ASAP7_75t_L g18047 ( 
.A(n_17656),
.B(n_9994),
.Y(n_18047)
);

INVxp67_ASAP7_75t_L g18048 ( 
.A(n_17638),
.Y(n_18048)
);

INVx1_ASAP7_75t_SL g18049 ( 
.A(n_17687),
.Y(n_18049)
);

AOI22xp33_ASAP7_75t_L g18050 ( 
.A1(n_17701),
.A2(n_17504),
.B1(n_17507),
.B2(n_17211),
.Y(n_18050)
);

OA21x2_ASAP7_75t_L g18051 ( 
.A1(n_17725),
.A2(n_9860),
.B(n_9847),
.Y(n_18051)
);

INVx1_ASAP7_75t_SL g18052 ( 
.A(n_17653),
.Y(n_18052)
);

AND2x2_ASAP7_75t_L g18053 ( 
.A(n_17634),
.B(n_7179),
.Y(n_18053)
);

OR2x6_ASAP7_75t_L g18054 ( 
.A(n_17666),
.B(n_5627),
.Y(n_18054)
);

HB1xp67_ASAP7_75t_L g18055 ( 
.A(n_17680),
.Y(n_18055)
);

INVx1_ASAP7_75t_L g18056 ( 
.A(n_17641),
.Y(n_18056)
);

NAND2xp5_ASAP7_75t_L g18057 ( 
.A(n_17622),
.B(n_10680),
.Y(n_18057)
);

NAND2xp5_ASAP7_75t_L g18058 ( 
.A(n_17649),
.B(n_17663),
.Y(n_18058)
);

INVx1_ASAP7_75t_SL g18059 ( 
.A(n_17707),
.Y(n_18059)
);

AND2x2_ASAP7_75t_L g18060 ( 
.A(n_17630),
.B(n_7183),
.Y(n_18060)
);

HB1xp67_ASAP7_75t_L g18061 ( 
.A(n_17965),
.Y(n_18061)
);

INVx1_ASAP7_75t_L g18062 ( 
.A(n_17626),
.Y(n_18062)
);

AOI22xp33_ASAP7_75t_L g18063 ( 
.A1(n_17710),
.A2(n_17484),
.B1(n_8353),
.B2(n_8426),
.Y(n_18063)
);

NOR2xp33_ASAP7_75t_L g18064 ( 
.A(n_17632),
.B(n_17670),
.Y(n_18064)
);

INVx1_ASAP7_75t_SL g18065 ( 
.A(n_17650),
.Y(n_18065)
);

OR2x2_ASAP7_75t_L g18066 ( 
.A(n_17635),
.B(n_10003),
.Y(n_18066)
);

INVx1_ASAP7_75t_L g18067 ( 
.A(n_17657),
.Y(n_18067)
);

BUFx2_ASAP7_75t_R g18068 ( 
.A(n_17824),
.Y(n_18068)
);

AND2x2_ASAP7_75t_L g18069 ( 
.A(n_17735),
.B(n_7183),
.Y(n_18069)
);

AND2x2_ASAP7_75t_L g18070 ( 
.A(n_17711),
.B(n_7183),
.Y(n_18070)
);

HB1xp67_ASAP7_75t_L g18071 ( 
.A(n_17681),
.Y(n_18071)
);

INVx2_ASAP7_75t_L g18072 ( 
.A(n_17930),
.Y(n_18072)
);

HB1xp67_ASAP7_75t_L g18073 ( 
.A(n_18017),
.Y(n_18073)
);

AND2x2_ASAP7_75t_L g18074 ( 
.A(n_17647),
.B(n_17674),
.Y(n_18074)
);

NAND2xp5_ASAP7_75t_L g18075 ( 
.A(n_17623),
.B(n_10680),
.Y(n_18075)
);

INVx1_ASAP7_75t_L g18076 ( 
.A(n_17631),
.Y(n_18076)
);

AND2x2_ASAP7_75t_L g18077 ( 
.A(n_17675),
.B(n_7183),
.Y(n_18077)
);

INVx1_ASAP7_75t_L g18078 ( 
.A(n_17944),
.Y(n_18078)
);

INVx3_ASAP7_75t_L g18079 ( 
.A(n_17976),
.Y(n_18079)
);

INVx1_ASAP7_75t_L g18080 ( 
.A(n_17627),
.Y(n_18080)
);

AND2x2_ASAP7_75t_L g18081 ( 
.A(n_17828),
.B(n_8581),
.Y(n_18081)
);

AND2x2_ASAP7_75t_L g18082 ( 
.A(n_17648),
.B(n_8581),
.Y(n_18082)
);

AND2x2_ASAP7_75t_L g18083 ( 
.A(n_17658),
.B(n_8581),
.Y(n_18083)
);

AND2x4_ASAP7_75t_L g18084 ( 
.A(n_17686),
.B(n_8304),
.Y(n_18084)
);

AND2x4_ASAP7_75t_L g18085 ( 
.A(n_17683),
.B(n_8353),
.Y(n_18085)
);

INVx4_ASAP7_75t_L g18086 ( 
.A(n_17821),
.Y(n_18086)
);

INVx2_ASAP7_75t_L g18087 ( 
.A(n_17994),
.Y(n_18087)
);

INVx1_ASAP7_75t_L g18088 ( 
.A(n_17744),
.Y(n_18088)
);

INVx1_ASAP7_75t_L g18089 ( 
.A(n_17755),
.Y(n_18089)
);

INVx1_ASAP7_75t_L g18090 ( 
.A(n_17736),
.Y(n_18090)
);

AND2x2_ASAP7_75t_L g18091 ( 
.A(n_17643),
.B(n_9172),
.Y(n_18091)
);

INVx1_ASAP7_75t_L g18092 ( 
.A(n_17624),
.Y(n_18092)
);

OAI22xp5_ASAP7_75t_L g18093 ( 
.A1(n_17688),
.A2(n_10687),
.B1(n_10688),
.B2(n_10684),
.Y(n_18093)
);

NAND2xp5_ASAP7_75t_L g18094 ( 
.A(n_17714),
.B(n_10684),
.Y(n_18094)
);

INVx2_ASAP7_75t_L g18095 ( 
.A(n_17906),
.Y(n_18095)
);

OAI21xp5_ASAP7_75t_L g18096 ( 
.A1(n_17709),
.A2(n_10429),
.B(n_10346),
.Y(n_18096)
);

INVx1_ASAP7_75t_L g18097 ( 
.A(n_17676),
.Y(n_18097)
);

AND2x2_ASAP7_75t_L g18098 ( 
.A(n_17815),
.B(n_9172),
.Y(n_18098)
);

BUFx3_ASAP7_75t_L g18099 ( 
.A(n_17655),
.Y(n_18099)
);

INVx1_ASAP7_75t_L g18100 ( 
.A(n_17921),
.Y(n_18100)
);

OR2x2_ASAP7_75t_L g18101 ( 
.A(n_17621),
.B(n_17636),
.Y(n_18101)
);

NAND2xp5_ASAP7_75t_L g18102 ( 
.A(n_17637),
.B(n_10687),
.Y(n_18102)
);

AND2x2_ASAP7_75t_L g18103 ( 
.A(n_17912),
.B(n_17698),
.Y(n_18103)
);

INVx1_ASAP7_75t_L g18104 ( 
.A(n_17822),
.Y(n_18104)
);

AOI222xp33_ASAP7_75t_L g18105 ( 
.A1(n_17981),
.A2(n_9729),
.B1(n_9716),
.B2(n_9748),
.C1(n_9743),
.C2(n_9725),
.Y(n_18105)
);

AND2x2_ASAP7_75t_L g18106 ( 
.A(n_17720),
.B(n_17771),
.Y(n_18106)
);

INVx1_ASAP7_75t_L g18107 ( 
.A(n_17836),
.Y(n_18107)
);

AND2x2_ASAP7_75t_L g18108 ( 
.A(n_17771),
.B(n_8909),
.Y(n_18108)
);

HB1xp67_ASAP7_75t_L g18109 ( 
.A(n_17718),
.Y(n_18109)
);

INVx2_ASAP7_75t_L g18110 ( 
.A(n_17970),
.Y(n_18110)
);

INVx2_ASAP7_75t_L g18111 ( 
.A(n_17882),
.Y(n_18111)
);

AOI22xp33_ASAP7_75t_L g18112 ( 
.A1(n_17963),
.A2(n_8426),
.B1(n_8465),
.B2(n_8353),
.Y(n_18112)
);

AND2x2_ASAP7_75t_L g18113 ( 
.A(n_17908),
.B(n_17918),
.Y(n_18113)
);

INVx3_ASAP7_75t_SL g18114 ( 
.A(n_17808),
.Y(n_18114)
);

OR2x2_ASAP7_75t_L g18115 ( 
.A(n_17645),
.B(n_10003),
.Y(n_18115)
);

NAND2xp5_ASAP7_75t_L g18116 ( 
.A(n_17640),
.B(n_10688),
.Y(n_18116)
);

INVx1_ASAP7_75t_L g18117 ( 
.A(n_17967),
.Y(n_18117)
);

AND2x2_ASAP7_75t_L g18118 ( 
.A(n_17672),
.B(n_8909),
.Y(n_18118)
);

HB1xp67_ASAP7_75t_L g18119 ( 
.A(n_17800),
.Y(n_18119)
);

AND2x2_ASAP7_75t_L g18120 ( 
.A(n_17677),
.B(n_8909),
.Y(n_18120)
);

INVx1_ASAP7_75t_L g18121 ( 
.A(n_17684),
.Y(n_18121)
);

OAI21xp33_ASAP7_75t_SL g18122 ( 
.A1(n_17651),
.A2(n_10429),
.B(n_10346),
.Y(n_18122)
);

AOI21xp5_ASAP7_75t_L g18123 ( 
.A1(n_17788),
.A2(n_9725),
.B(n_9716),
.Y(n_18123)
);

AND2x2_ASAP7_75t_L g18124 ( 
.A(n_17697),
.B(n_8909),
.Y(n_18124)
);

NAND2xp5_ASAP7_75t_L g18125 ( 
.A(n_18008),
.B(n_10689),
.Y(n_18125)
);

AND2x4_ASAP7_75t_L g18126 ( 
.A(n_17830),
.B(n_8426),
.Y(n_18126)
);

INVx1_ASAP7_75t_L g18127 ( 
.A(n_18003),
.Y(n_18127)
);

AND2x2_ASAP7_75t_L g18128 ( 
.A(n_17759),
.B(n_8909),
.Y(n_18128)
);

INVx1_ASAP7_75t_L g18129 ( 
.A(n_17629),
.Y(n_18129)
);

OAI22xp5_ASAP7_75t_L g18130 ( 
.A1(n_17798),
.A2(n_10693),
.B1(n_10708),
.B2(n_10689),
.Y(n_18130)
);

INVx1_ASAP7_75t_SL g18131 ( 
.A(n_17703),
.Y(n_18131)
);

INVx2_ASAP7_75t_L g18132 ( 
.A(n_17926),
.Y(n_18132)
);

NAND2xp5_ASAP7_75t_L g18133 ( 
.A(n_17943),
.B(n_10693),
.Y(n_18133)
);

NOR2xp33_ASAP7_75t_L g18134 ( 
.A(n_17797),
.B(n_8978),
.Y(n_18134)
);

INVx1_ASAP7_75t_SL g18135 ( 
.A(n_17775),
.Y(n_18135)
);

NOR2x1_ASAP7_75t_L g18136 ( 
.A(n_17909),
.B(n_10708),
.Y(n_18136)
);

AND2x2_ASAP7_75t_L g18137 ( 
.A(n_17705),
.B(n_8909),
.Y(n_18137)
);

INVx1_ASAP7_75t_L g18138 ( 
.A(n_17654),
.Y(n_18138)
);

INVx2_ASAP7_75t_L g18139 ( 
.A(n_17885),
.Y(n_18139)
);

INVx2_ASAP7_75t_L g18140 ( 
.A(n_17806),
.Y(n_18140)
);

AND2x2_ASAP7_75t_L g18141 ( 
.A(n_17733),
.B(n_8909),
.Y(n_18141)
);

NAND2xp5_ASAP7_75t_L g18142 ( 
.A(n_17646),
.B(n_10710),
.Y(n_18142)
);

AND2x2_ASAP7_75t_L g18143 ( 
.A(n_17700),
.B(n_8909),
.Y(n_18143)
);

AND2x2_ASAP7_75t_L g18144 ( 
.A(n_17696),
.B(n_8909),
.Y(n_18144)
);

INVx2_ASAP7_75t_L g18145 ( 
.A(n_17776),
.Y(n_18145)
);

INVx1_ASAP7_75t_L g18146 ( 
.A(n_17789),
.Y(n_18146)
);

AND2x4_ASAP7_75t_L g18147 ( 
.A(n_17834),
.B(n_17794),
.Y(n_18147)
);

INVx1_ASAP7_75t_SL g18148 ( 
.A(n_17695),
.Y(n_18148)
);

HB1xp67_ASAP7_75t_L g18149 ( 
.A(n_17851),
.Y(n_18149)
);

INVx1_ASAP7_75t_SL g18150 ( 
.A(n_17702),
.Y(n_18150)
);

AND2x2_ASAP7_75t_L g18151 ( 
.A(n_17817),
.B(n_8957),
.Y(n_18151)
);

AND2x2_ASAP7_75t_L g18152 ( 
.A(n_18029),
.B(n_8957),
.Y(n_18152)
);

NAND3xp33_ASAP7_75t_L g18153 ( 
.A(n_17669),
.B(n_9729),
.C(n_9725),
.Y(n_18153)
);

AND2x2_ASAP7_75t_L g18154 ( 
.A(n_17793),
.B(n_8957),
.Y(n_18154)
);

AND2x2_ASAP7_75t_L g18155 ( 
.A(n_17717),
.B(n_8957),
.Y(n_18155)
);

INVx1_ASAP7_75t_L g18156 ( 
.A(n_17968),
.Y(n_18156)
);

NAND2xp5_ASAP7_75t_L g18157 ( 
.A(n_17983),
.B(n_10710),
.Y(n_18157)
);

INVx1_ASAP7_75t_SL g18158 ( 
.A(n_17920),
.Y(n_18158)
);

INVx1_ASAP7_75t_L g18159 ( 
.A(n_17781),
.Y(n_18159)
);

NAND2xp5_ASAP7_75t_L g18160 ( 
.A(n_18006),
.B(n_10711),
.Y(n_18160)
);

INVx1_ASAP7_75t_L g18161 ( 
.A(n_17971),
.Y(n_18161)
);

OR2x2_ASAP7_75t_L g18162 ( 
.A(n_17847),
.B(n_10003),
.Y(n_18162)
);

INVx2_ASAP7_75t_L g18163 ( 
.A(n_17716),
.Y(n_18163)
);

CKINVDCx16_ASAP7_75t_R g18164 ( 
.A(n_17897),
.Y(n_18164)
);

INVx1_ASAP7_75t_L g18165 ( 
.A(n_17942),
.Y(n_18165)
);

INVx1_ASAP7_75t_L g18166 ( 
.A(n_17712),
.Y(n_18166)
);

AND2x2_ASAP7_75t_L g18167 ( 
.A(n_17894),
.B(n_8957),
.Y(n_18167)
);

INVx1_ASAP7_75t_L g18168 ( 
.A(n_17740),
.Y(n_18168)
);

INVx1_ASAP7_75t_L g18169 ( 
.A(n_17738),
.Y(n_18169)
);

INVx1_ASAP7_75t_SL g18170 ( 
.A(n_17868),
.Y(n_18170)
);

AO21x2_ASAP7_75t_L g18171 ( 
.A1(n_17799),
.A2(n_10711),
.B(n_10213),
.Y(n_18171)
);

INVx2_ASAP7_75t_L g18172 ( 
.A(n_17752),
.Y(n_18172)
);

AOI22xp33_ASAP7_75t_L g18173 ( 
.A1(n_17639),
.A2(n_8509),
.B1(n_8512),
.B2(n_8465),
.Y(n_18173)
);

AND2x2_ASAP7_75t_L g18174 ( 
.A(n_17820),
.B(n_8957),
.Y(n_18174)
);

NAND2xp5_ASAP7_75t_L g18175 ( 
.A(n_18011),
.B(n_7995),
.Y(n_18175)
);

NAND2xp5_ASAP7_75t_L g18176 ( 
.A(n_18016),
.B(n_7995),
.Y(n_18176)
);

AND2x2_ASAP7_75t_L g18177 ( 
.A(n_17739),
.B(n_8957),
.Y(n_18177)
);

AND2x2_ASAP7_75t_L g18178 ( 
.A(n_17749),
.B(n_17756),
.Y(n_18178)
);

INVx1_ASAP7_75t_L g18179 ( 
.A(n_17810),
.Y(n_18179)
);

AOI22xp5_ASAP7_75t_L g18180 ( 
.A1(n_17747),
.A2(n_10010),
.B1(n_10017),
.B2(n_10007),
.Y(n_18180)
);

INVx2_ASAP7_75t_L g18181 ( 
.A(n_17935),
.Y(n_18181)
);

OR2x2_ASAP7_75t_L g18182 ( 
.A(n_18025),
.B(n_10007),
.Y(n_18182)
);

INVx1_ASAP7_75t_L g18183 ( 
.A(n_17661),
.Y(n_18183)
);

INVx1_ASAP7_75t_L g18184 ( 
.A(n_17905),
.Y(n_18184)
);

INVx1_ASAP7_75t_L g18185 ( 
.A(n_17907),
.Y(n_18185)
);

INVx2_ASAP7_75t_L g18186 ( 
.A(n_17940),
.Y(n_18186)
);

INVx1_ASAP7_75t_SL g18187 ( 
.A(n_17890),
.Y(n_18187)
);

INVx2_ASAP7_75t_SL g18188 ( 
.A(n_17922),
.Y(n_18188)
);

INVx1_ASAP7_75t_SL g18189 ( 
.A(n_17931),
.Y(n_18189)
);

OR2x2_ASAP7_75t_L g18190 ( 
.A(n_17625),
.B(n_10007),
.Y(n_18190)
);

INVx1_ASAP7_75t_L g18191 ( 
.A(n_17961),
.Y(n_18191)
);

OR2x2_ASAP7_75t_L g18192 ( 
.A(n_17737),
.B(n_10010),
.Y(n_18192)
);

AND2x4_ASAP7_75t_L g18193 ( 
.A(n_17818),
.B(n_8465),
.Y(n_18193)
);

INVx1_ASAP7_75t_SL g18194 ( 
.A(n_17927),
.Y(n_18194)
);

INVx1_ASAP7_75t_L g18195 ( 
.A(n_17753),
.Y(n_18195)
);

AND2x2_ASAP7_75t_L g18196 ( 
.A(n_18022),
.B(n_8957),
.Y(n_18196)
);

AOI22xp33_ASAP7_75t_L g18197 ( 
.A1(n_18026),
.A2(n_17962),
.B1(n_17840),
.B2(n_17770),
.Y(n_18197)
);

AOI22x1_ASAP7_75t_L g18198 ( 
.A1(n_17973),
.A2(n_17984),
.B1(n_17996),
.B2(n_17660),
.Y(n_18198)
);

AO21x2_ASAP7_75t_L g18199 ( 
.A1(n_17773),
.A2(n_10213),
.B(n_10193),
.Y(n_18199)
);

INVx2_ASAP7_75t_L g18200 ( 
.A(n_17950),
.Y(n_18200)
);

INVx1_ASAP7_75t_SL g18201 ( 
.A(n_17664),
.Y(n_18201)
);

NAND2xp5_ASAP7_75t_L g18202 ( 
.A(n_17959),
.B(n_17956),
.Y(n_18202)
);

BUFx3_ASAP7_75t_L g18203 ( 
.A(n_17952),
.Y(n_18203)
);

AND2x4_ASAP7_75t_SL g18204 ( 
.A(n_17727),
.B(n_9048),
.Y(n_18204)
);

OR2x2_ASAP7_75t_L g18205 ( 
.A(n_17728),
.B(n_10010),
.Y(n_18205)
);

NAND2xp5_ASAP7_75t_L g18206 ( 
.A(n_17730),
.B(n_7995),
.Y(n_18206)
);

BUFx2_ASAP7_75t_L g18207 ( 
.A(n_18004),
.Y(n_18207)
);

NOR2xp33_ASAP7_75t_L g18208 ( 
.A(n_17865),
.B(n_9071),
.Y(n_18208)
);

NOR2x1_ASAP7_75t_L g18209 ( 
.A(n_17628),
.B(n_8847),
.Y(n_18209)
);

BUFx2_ASAP7_75t_L g18210 ( 
.A(n_17779),
.Y(n_18210)
);

BUFx3_ASAP7_75t_L g18211 ( 
.A(n_18020),
.Y(n_18211)
);

NAND2x1p5_ASAP7_75t_L g18212 ( 
.A(n_17936),
.B(n_9099),
.Y(n_18212)
);

AOI22xp33_ASAP7_75t_L g18213 ( 
.A1(n_18026),
.A2(n_8512),
.B1(n_8643),
.B2(n_8509),
.Y(n_18213)
);

NOR2xp33_ASAP7_75t_L g18214 ( 
.A(n_17911),
.B(n_9247),
.Y(n_18214)
);

NOR2xp33_ASAP7_75t_L g18215 ( 
.A(n_17958),
.B(n_9247),
.Y(n_18215)
);

OR2x2_ASAP7_75t_L g18216 ( 
.A(n_17659),
.B(n_10017),
.Y(n_18216)
);

INVx1_ASAP7_75t_L g18217 ( 
.A(n_17706),
.Y(n_18217)
);

NAND3xp33_ASAP7_75t_SL g18218 ( 
.A(n_17863),
.B(n_9289),
.C(n_9288),
.Y(n_18218)
);

INVx1_ASAP7_75t_L g18219 ( 
.A(n_17715),
.Y(n_18219)
);

INVx1_ASAP7_75t_L g18220 ( 
.A(n_17731),
.Y(n_18220)
);

NOR2xp33_ASAP7_75t_L g18221 ( 
.A(n_17849),
.B(n_17860),
.Y(n_18221)
);

NOR2xp33_ASAP7_75t_L g18222 ( 
.A(n_17877),
.B(n_9288),
.Y(n_18222)
);

AND2x2_ASAP7_75t_L g18223 ( 
.A(n_17778),
.B(n_8957),
.Y(n_18223)
);

AND2x4_ASAP7_75t_L g18224 ( 
.A(n_18023),
.B(n_8509),
.Y(n_18224)
);

BUFx3_ASAP7_75t_L g18225 ( 
.A(n_17937),
.Y(n_18225)
);

INVx1_ASAP7_75t_L g18226 ( 
.A(n_17746),
.Y(n_18226)
);

INVx1_ASAP7_75t_L g18227 ( 
.A(n_17751),
.Y(n_18227)
);

AOI22xp33_ASAP7_75t_L g18228 ( 
.A1(n_18026),
.A2(n_8643),
.B1(n_8671),
.B2(n_8512),
.Y(n_18228)
);

INVxp67_ASAP7_75t_SL g18229 ( 
.A(n_17888),
.Y(n_18229)
);

AND2x2_ASAP7_75t_L g18230 ( 
.A(n_17783),
.B(n_8564),
.Y(n_18230)
);

AO21x2_ASAP7_75t_L g18231 ( 
.A1(n_17898),
.A2(n_8705),
.B(n_8600),
.Y(n_18231)
);

INVx2_ASAP7_75t_SL g18232 ( 
.A(n_17772),
.Y(n_18232)
);

INVx4_ASAP7_75t_L g18233 ( 
.A(n_17946),
.Y(n_18233)
);

INVx1_ASAP7_75t_SL g18234 ( 
.A(n_17960),
.Y(n_18234)
);

OR2x2_ASAP7_75t_L g18235 ( 
.A(n_17835),
.B(n_10017),
.Y(n_18235)
);

INVx2_ASAP7_75t_L g18236 ( 
.A(n_17953),
.Y(n_18236)
);

AND2x2_ASAP7_75t_L g18237 ( 
.A(n_17692),
.B(n_7606),
.Y(n_18237)
);

AOI22xp5_ASAP7_75t_L g18238 ( 
.A1(n_17765),
.A2(n_10021),
.B1(n_10024),
.B2(n_10020),
.Y(n_18238)
);

NOR2x1_ASAP7_75t_L g18239 ( 
.A(n_17917),
.B(n_8847),
.Y(n_18239)
);

BUFx3_ASAP7_75t_L g18240 ( 
.A(n_17839),
.Y(n_18240)
);

OR2x2_ASAP7_75t_L g18241 ( 
.A(n_17742),
.B(n_10020),
.Y(n_18241)
);

INVx1_ASAP7_75t_L g18242 ( 
.A(n_17722),
.Y(n_18242)
);

AND2x2_ASAP7_75t_L g18243 ( 
.A(n_17801),
.B(n_7606),
.Y(n_18243)
);

NOR2xp33_ASAP7_75t_L g18244 ( 
.A(n_17850),
.B(n_9289),
.Y(n_18244)
);

HB1xp67_ASAP7_75t_L g18245 ( 
.A(n_17889),
.Y(n_18245)
);

NOR2x1_ASAP7_75t_L g18246 ( 
.A(n_17919),
.B(n_8847),
.Y(n_18246)
);

AND2x2_ASAP7_75t_L g18247 ( 
.A(n_17855),
.B(n_9847),
.Y(n_18247)
);

BUFx3_ASAP7_75t_L g18248 ( 
.A(n_17878),
.Y(n_18248)
);

AOI22xp33_ASAP7_75t_L g18249 ( 
.A1(n_17748),
.A2(n_8671),
.B1(n_8714),
.B2(n_8643),
.Y(n_18249)
);

OR2x2_ASAP7_75t_L g18250 ( 
.A(n_17745),
.B(n_10020),
.Y(n_18250)
);

INVx4_ASAP7_75t_L g18251 ( 
.A(n_17924),
.Y(n_18251)
);

INVx2_ASAP7_75t_L g18252 ( 
.A(n_17985),
.Y(n_18252)
);

INVx2_ASAP7_75t_L g18253 ( 
.A(n_17704),
.Y(n_18253)
);

INVx1_ASAP7_75t_L g18254 ( 
.A(n_17723),
.Y(n_18254)
);

BUFx3_ASAP7_75t_L g18255 ( 
.A(n_17893),
.Y(n_18255)
);

NOR2x1_ASAP7_75t_L g18256 ( 
.A(n_17895),
.B(n_8847),
.Y(n_18256)
);

INVx1_ASAP7_75t_L g18257 ( 
.A(n_17678),
.Y(n_18257)
);

INVx1_ASAP7_75t_L g18258 ( 
.A(n_17693),
.Y(n_18258)
);

OR2x6_ASAP7_75t_L g18259 ( 
.A(n_17902),
.B(n_5627),
.Y(n_18259)
);

OR2x2_ASAP7_75t_L g18260 ( 
.A(n_17754),
.B(n_10021),
.Y(n_18260)
);

INVx1_ASAP7_75t_SL g18261 ( 
.A(n_17685),
.Y(n_18261)
);

INVx1_ASAP7_75t_L g18262 ( 
.A(n_17729),
.Y(n_18262)
);

NOR2xp33_ASAP7_75t_L g18263 ( 
.A(n_17954),
.B(n_9054),
.Y(n_18263)
);

OAI22xp5_ASAP7_75t_L g18264 ( 
.A1(n_17951),
.A2(n_8714),
.B1(n_8796),
.B2(n_8671),
.Y(n_18264)
);

INVx1_ASAP7_75t_SL g18265 ( 
.A(n_17713),
.Y(n_18265)
);

AOI22xp33_ASAP7_75t_L g18266 ( 
.A1(n_17978),
.A2(n_8714),
.B1(n_8833),
.B2(n_8796),
.Y(n_18266)
);

INVx1_ASAP7_75t_L g18267 ( 
.A(n_17833),
.Y(n_18267)
);

OR2x2_ASAP7_75t_L g18268 ( 
.A(n_17758),
.B(n_10021),
.Y(n_18268)
);

AND2x2_ASAP7_75t_L g18269 ( 
.A(n_17777),
.B(n_9860),
.Y(n_18269)
);

INVx1_ASAP7_75t_L g18270 ( 
.A(n_17769),
.Y(n_18270)
);

INVxp67_ASAP7_75t_SL g18271 ( 
.A(n_17679),
.Y(n_18271)
);

INVx1_ASAP7_75t_L g18272 ( 
.A(n_17792),
.Y(n_18272)
);

INVx1_ASAP7_75t_L g18273 ( 
.A(n_17796),
.Y(n_18273)
);

INVx1_ASAP7_75t_L g18274 ( 
.A(n_17825),
.Y(n_18274)
);

OR2x2_ASAP7_75t_L g18275 ( 
.A(n_17977),
.B(n_10024),
.Y(n_18275)
);

HB1xp67_ASAP7_75t_L g18276 ( 
.A(n_17782),
.Y(n_18276)
);

INVx2_ASAP7_75t_L g18277 ( 
.A(n_17699),
.Y(n_18277)
);

INVxp67_ASAP7_75t_SL g18278 ( 
.A(n_17811),
.Y(n_18278)
);

CKINVDCx16_ASAP7_75t_R g18279 ( 
.A(n_17903),
.Y(n_18279)
);

AND2x2_ASAP7_75t_L g18280 ( 
.A(n_17955),
.B(n_9874),
.Y(n_18280)
);

INVx1_ASAP7_75t_L g18281 ( 
.A(n_17826),
.Y(n_18281)
);

AOI22xp5_ASAP7_75t_L g18282 ( 
.A1(n_17842),
.A2(n_10058),
.B1(n_10072),
.B2(n_10024),
.Y(n_18282)
);

INVx2_ASAP7_75t_L g18283 ( 
.A(n_17891),
.Y(n_18283)
);

NAND2xp5_ASAP7_75t_L g18284 ( 
.A(n_17662),
.B(n_7995),
.Y(n_18284)
);

INVx2_ASAP7_75t_L g18285 ( 
.A(n_17892),
.Y(n_18285)
);

AND2x2_ASAP7_75t_L g18286 ( 
.A(n_17880),
.B(n_9874),
.Y(n_18286)
);

INVx1_ASAP7_75t_L g18287 ( 
.A(n_17814),
.Y(n_18287)
);

INVx4_ASAP7_75t_L g18288 ( 
.A(n_17910),
.Y(n_18288)
);

OR2x2_ASAP7_75t_L g18289 ( 
.A(n_17980),
.B(n_10058),
.Y(n_18289)
);

INVx2_ASAP7_75t_L g18290 ( 
.A(n_17719),
.Y(n_18290)
);

INVx2_ASAP7_75t_L g18291 ( 
.A(n_17721),
.Y(n_18291)
);

NAND2xp5_ASAP7_75t_L g18292 ( 
.A(n_18018),
.B(n_7995),
.Y(n_18292)
);

CKINVDCx16_ASAP7_75t_R g18293 ( 
.A(n_17914),
.Y(n_18293)
);

AND2x2_ASAP7_75t_L g18294 ( 
.A(n_17784),
.B(n_7028),
.Y(n_18294)
);

AND3x1_ASAP7_75t_L g18295 ( 
.A(n_17982),
.B(n_9743),
.C(n_9729),
.Y(n_18295)
);

INVx1_ASAP7_75t_SL g18296 ( 
.A(n_17694),
.Y(n_18296)
);

OAI22xp5_ASAP7_75t_L g18297 ( 
.A1(n_17708),
.A2(n_8833),
.B1(n_8892),
.B2(n_8796),
.Y(n_18297)
);

AND2x2_ASAP7_75t_L g18298 ( 
.A(n_17689),
.B(n_7028),
.Y(n_18298)
);

INVx2_ASAP7_75t_L g18299 ( 
.A(n_17734),
.Y(n_18299)
);

OR2x2_ASAP7_75t_L g18300 ( 
.A(n_17844),
.B(n_10058),
.Y(n_18300)
);

INVx1_ASAP7_75t_SL g18301 ( 
.A(n_17671),
.Y(n_18301)
);

NAND2xp5_ASAP7_75t_L g18302 ( 
.A(n_18027),
.B(n_8014),
.Y(n_18302)
);

AND2x2_ASAP7_75t_L g18303 ( 
.A(n_17690),
.B(n_7028),
.Y(n_18303)
);

AOI22xp33_ASAP7_75t_L g18304 ( 
.A1(n_17896),
.A2(n_8892),
.B1(n_8904),
.B2(n_8833),
.Y(n_18304)
);

AND2x2_ASAP7_75t_L g18305 ( 
.A(n_17767),
.B(n_7028),
.Y(n_18305)
);

OA21x2_ASAP7_75t_L g18306 ( 
.A1(n_17843),
.A2(n_10460),
.B(n_10443),
.Y(n_18306)
);

OR2x2_ASAP7_75t_L g18307 ( 
.A(n_17665),
.B(n_10072),
.Y(n_18307)
);

AND2x2_ASAP7_75t_L g18308 ( 
.A(n_17803),
.B(n_7028),
.Y(n_18308)
);

INVxp67_ASAP7_75t_L g18309 ( 
.A(n_17854),
.Y(n_18309)
);

AND2x4_ASAP7_75t_L g18310 ( 
.A(n_17741),
.B(n_8892),
.Y(n_18310)
);

INVx1_ASAP7_75t_SL g18311 ( 
.A(n_17838),
.Y(n_18311)
);

OR2x2_ASAP7_75t_L g18312 ( 
.A(n_18028),
.B(n_10072),
.Y(n_18312)
);

OAI22xp5_ASAP7_75t_L g18313 ( 
.A1(n_17757),
.A2(n_8913),
.B1(n_8932),
.B2(n_8904),
.Y(n_18313)
);

INVx1_ASAP7_75t_L g18314 ( 
.A(n_17804),
.Y(n_18314)
);

INVx1_ASAP7_75t_L g18315 ( 
.A(n_17861),
.Y(n_18315)
);

INVx2_ASAP7_75t_L g18316 ( 
.A(n_17760),
.Y(n_18316)
);

AND2x2_ASAP7_75t_L g18317 ( 
.A(n_17805),
.B(n_17887),
.Y(n_18317)
);

OR2x2_ASAP7_75t_L g18318 ( 
.A(n_17732),
.B(n_10077),
.Y(n_18318)
);

INVx1_ASAP7_75t_SL g18319 ( 
.A(n_17809),
.Y(n_18319)
);

AND2x4_ASAP7_75t_L g18320 ( 
.A(n_17763),
.B(n_17802),
.Y(n_18320)
);

OAI22xp5_ASAP7_75t_L g18321 ( 
.A1(n_17786),
.A2(n_8913),
.B1(n_8932),
.B2(n_8904),
.Y(n_18321)
);

INVxp67_ASAP7_75t_L g18322 ( 
.A(n_17867),
.Y(n_18322)
);

NAND2xp5_ASAP7_75t_L g18323 ( 
.A(n_17886),
.B(n_17819),
.Y(n_18323)
);

AND2x2_ASAP7_75t_L g18324 ( 
.A(n_17831),
.B(n_17832),
.Y(n_18324)
);

INVx1_ASAP7_75t_SL g18325 ( 
.A(n_18021),
.Y(n_18325)
);

INVx1_ASAP7_75t_L g18326 ( 
.A(n_17862),
.Y(n_18326)
);

NAND2xp5_ASAP7_75t_L g18327 ( 
.A(n_17948),
.B(n_8014),
.Y(n_18327)
);

INVx1_ASAP7_75t_L g18328 ( 
.A(n_17852),
.Y(n_18328)
);

INVx1_ASAP7_75t_SL g18329 ( 
.A(n_17768),
.Y(n_18329)
);

INVx1_ASAP7_75t_SL g18330 ( 
.A(n_17790),
.Y(n_18330)
);

AOI22xp33_ASAP7_75t_L g18331 ( 
.A1(n_17934),
.A2(n_8932),
.B1(n_8951),
.B2(n_8913),
.Y(n_18331)
);

NOR2xp67_ASAP7_75t_SL g18332 ( 
.A(n_17774),
.B(n_5751),
.Y(n_18332)
);

AOI222xp33_ASAP7_75t_L g18333 ( 
.A1(n_17941),
.A2(n_9750),
.B1(n_9748),
.B2(n_9763),
.C1(n_9759),
.C2(n_9743),
.Y(n_18333)
);

INVx2_ASAP7_75t_L g18334 ( 
.A(n_17913),
.Y(n_18334)
);

AND2x2_ASAP7_75t_L g18335 ( 
.A(n_17993),
.B(n_18012),
.Y(n_18335)
);

NAND2xp5_ASAP7_75t_L g18336 ( 
.A(n_17949),
.B(n_8014),
.Y(n_18336)
);

OR2x2_ASAP7_75t_L g18337 ( 
.A(n_17791),
.B(n_10077),
.Y(n_18337)
);

INVx2_ASAP7_75t_L g18338 ( 
.A(n_17915),
.Y(n_18338)
);

INVx1_ASAP7_75t_SL g18339 ( 
.A(n_17795),
.Y(n_18339)
);

INVx1_ASAP7_75t_SL g18340 ( 
.A(n_17812),
.Y(n_18340)
);

AND2x2_ASAP7_75t_L g18341 ( 
.A(n_18019),
.B(n_7028),
.Y(n_18341)
);

AND2x2_ASAP7_75t_L g18342 ( 
.A(n_17964),
.B(n_7029),
.Y(n_18342)
);

NAND2xp5_ASAP7_75t_L g18343 ( 
.A(n_17928),
.B(n_8014),
.Y(n_18343)
);

INVx1_ASAP7_75t_SL g18344 ( 
.A(n_17823),
.Y(n_18344)
);

NOR2xp33_ASAP7_75t_L g18345 ( 
.A(n_17853),
.B(n_9109),
.Y(n_18345)
);

INVx1_ASAP7_75t_L g18346 ( 
.A(n_17858),
.Y(n_18346)
);

INVx2_ASAP7_75t_L g18347 ( 
.A(n_17916),
.Y(n_18347)
);

AND2x4_ASAP7_75t_L g18348 ( 
.A(n_17859),
.B(n_8951),
.Y(n_18348)
);

NOR2xp33_ASAP7_75t_L g18349 ( 
.A(n_17869),
.B(n_9109),
.Y(n_18349)
);

INVx1_ASAP7_75t_SL g18350 ( 
.A(n_17780),
.Y(n_18350)
);

BUFx3_ASAP7_75t_L g18351 ( 
.A(n_17872),
.Y(n_18351)
);

OAI21xp33_ASAP7_75t_L g18352 ( 
.A1(n_17879),
.A2(n_9750),
.B(n_9748),
.Y(n_18352)
);

INVx1_ASAP7_75t_L g18353 ( 
.A(n_17925),
.Y(n_18353)
);

HB1xp67_ASAP7_75t_L g18354 ( 
.A(n_18002),
.Y(n_18354)
);

INVx1_ASAP7_75t_L g18355 ( 
.A(n_17929),
.Y(n_18355)
);

INVx1_ASAP7_75t_SL g18356 ( 
.A(n_17816),
.Y(n_18356)
);

INVx1_ASAP7_75t_SL g18357 ( 
.A(n_17966),
.Y(n_18357)
);

INVx1_ASAP7_75t_SL g18358 ( 
.A(n_17986),
.Y(n_18358)
);

INVx4_ASAP7_75t_L g18359 ( 
.A(n_17988),
.Y(n_18359)
);

NAND2xp5_ASAP7_75t_L g18360 ( 
.A(n_17932),
.B(n_8014),
.Y(n_18360)
);

NAND2xp5_ASAP7_75t_L g18361 ( 
.A(n_17938),
.B(n_8251),
.Y(n_18361)
);

AND2x4_ASAP7_75t_L g18362 ( 
.A(n_17990),
.B(n_8951),
.Y(n_18362)
);

INVx2_ASAP7_75t_L g18363 ( 
.A(n_17829),
.Y(n_18363)
);

INVx1_ASAP7_75t_L g18364 ( 
.A(n_17939),
.Y(n_18364)
);

INVx2_ASAP7_75t_L g18365 ( 
.A(n_17766),
.Y(n_18365)
);

INVx1_ASAP7_75t_SL g18366 ( 
.A(n_17979),
.Y(n_18366)
);

AND2x2_ASAP7_75t_L g18367 ( 
.A(n_17992),
.B(n_7029),
.Y(n_18367)
);

AOI21xp5_ASAP7_75t_L g18368 ( 
.A1(n_18045),
.A2(n_17841),
.B(n_18015),
.Y(n_18368)
);

AOI22xp5_ASAP7_75t_L g18369 ( 
.A1(n_18062),
.A2(n_18065),
.B1(n_18059),
.B2(n_18052),
.Y(n_18369)
);

AND2x2_ASAP7_75t_L g18370 ( 
.A(n_18039),
.B(n_17975),
.Y(n_18370)
);

INVx1_ASAP7_75t_L g18371 ( 
.A(n_18068),
.Y(n_18371)
);

OR2x2_ASAP7_75t_L g18372 ( 
.A(n_18164),
.B(n_18086),
.Y(n_18372)
);

INVx1_ASAP7_75t_SL g18373 ( 
.A(n_18114),
.Y(n_18373)
);

INVx1_ASAP7_75t_L g18374 ( 
.A(n_18040),
.Y(n_18374)
);

NAND3xp33_ASAP7_75t_L g18375 ( 
.A(n_18064),
.B(n_17998),
.C(n_17972),
.Y(n_18375)
);

O2A1O1Ixp33_ASAP7_75t_L g18376 ( 
.A1(n_18276),
.A2(n_17997),
.B(n_17945),
.C(n_17848),
.Y(n_18376)
);

INVx1_ASAP7_75t_L g18377 ( 
.A(n_18061),
.Y(n_18377)
);

AOI21xp5_ASAP7_75t_L g18378 ( 
.A1(n_18202),
.A2(n_17987),
.B(n_17947),
.Y(n_18378)
);

AND2x2_ASAP7_75t_SL g18379 ( 
.A(n_18074),
.B(n_17764),
.Y(n_18379)
);

INVxp67_ASAP7_75t_SL g18380 ( 
.A(n_18055),
.Y(n_18380)
);

AOI32xp33_ASAP7_75t_L g18381 ( 
.A1(n_18049),
.A2(n_18007),
.A3(n_18009),
.B1(n_17743),
.B2(n_18001),
.Y(n_18381)
);

OAI22xp33_ASAP7_75t_L g18382 ( 
.A1(n_18189),
.A2(n_17957),
.B1(n_17785),
.B2(n_17989),
.Y(n_18382)
);

INVx2_ASAP7_75t_L g18383 ( 
.A(n_18043),
.Y(n_18383)
);

AOI22xp5_ASAP7_75t_L g18384 ( 
.A1(n_18097),
.A2(n_17999),
.B1(n_17827),
.B2(n_18024),
.Y(n_18384)
);

INVx1_ASAP7_75t_L g18385 ( 
.A(n_18210),
.Y(n_18385)
);

INVx1_ASAP7_75t_L g18386 ( 
.A(n_18149),
.Y(n_18386)
);

NAND2xp5_ASAP7_75t_L g18387 ( 
.A(n_18067),
.B(n_18013),
.Y(n_18387)
);

AND2x2_ASAP7_75t_L g18388 ( 
.A(n_18103),
.B(n_17845),
.Y(n_18388)
);

INVx1_ASAP7_75t_L g18389 ( 
.A(n_18109),
.Y(n_18389)
);

INVx1_ASAP7_75t_L g18390 ( 
.A(n_18058),
.Y(n_18390)
);

OAI22xp5_ASAP7_75t_L g18391 ( 
.A1(n_18197),
.A2(n_17991),
.B1(n_17871),
.B2(n_17864),
.Y(n_18391)
);

INVx1_ASAP7_75t_L g18392 ( 
.A(n_18119),
.Y(n_18392)
);

INVx1_ASAP7_75t_L g18393 ( 
.A(n_18071),
.Y(n_18393)
);

AOI21xp33_ASAP7_75t_SL g18394 ( 
.A1(n_18279),
.A2(n_17901),
.B(n_18000),
.Y(n_18394)
);

NAND2xp5_ASAP7_75t_L g18395 ( 
.A(n_18030),
.B(n_17807),
.Y(n_18395)
);

AOI22xp5_ASAP7_75t_L g18396 ( 
.A1(n_18170),
.A2(n_17846),
.B1(n_17873),
.B2(n_17866),
.Y(n_18396)
);

AOI22xp5_ASAP7_75t_L g18397 ( 
.A1(n_18088),
.A2(n_17837),
.B1(n_17899),
.B2(n_17904),
.Y(n_18397)
);

INVxp67_ASAP7_75t_L g18398 ( 
.A(n_18073),
.Y(n_18398)
);

NAND2x1_ASAP7_75t_L g18399 ( 
.A(n_18195),
.B(n_17923),
.Y(n_18399)
);

INVx2_ASAP7_75t_SL g18400 ( 
.A(n_18212),
.Y(n_18400)
);

AND2x2_ASAP7_75t_L g18401 ( 
.A(n_18113),
.B(n_17875),
.Y(n_18401)
);

OR2x2_ASAP7_75t_L g18402 ( 
.A(n_18191),
.B(n_18005),
.Y(n_18402)
);

OAI221xp5_ASAP7_75t_L g18403 ( 
.A1(n_18122),
.A2(n_17876),
.B1(n_17881),
.B2(n_17874),
.C(n_17870),
.Y(n_18403)
);

OAI21xp33_ASAP7_75t_L g18404 ( 
.A1(n_18091),
.A2(n_18014),
.B(n_17682),
.Y(n_18404)
);

HB1xp67_ASAP7_75t_L g18405 ( 
.A(n_18032),
.Y(n_18405)
);

OA22x2_ASAP7_75t_L g18406 ( 
.A1(n_18072),
.A2(n_17884),
.B1(n_17883),
.B2(n_17761),
.Y(n_18406)
);

AOI21xp33_ASAP7_75t_SL g18407 ( 
.A1(n_18293),
.A2(n_18041),
.B(n_18100),
.Y(n_18407)
);

INVx1_ASAP7_75t_L g18408 ( 
.A(n_18101),
.Y(n_18408)
);

INVx1_ASAP7_75t_L g18409 ( 
.A(n_18245),
.Y(n_18409)
);

HB1xp67_ASAP7_75t_L g18410 ( 
.A(n_18354),
.Y(n_18410)
);

AOI21xp33_ASAP7_75t_L g18411 ( 
.A1(n_18089),
.A2(n_17974),
.B(n_17813),
.Y(n_18411)
);

NAND2xp5_ASAP7_75t_L g18412 ( 
.A(n_18079),
.B(n_17856),
.Y(n_18412)
);

INVx1_ASAP7_75t_L g18413 ( 
.A(n_18229),
.Y(n_18413)
);

NAND2xp5_ASAP7_75t_L g18414 ( 
.A(n_18078),
.B(n_17857),
.Y(n_18414)
);

OAI211xp5_ASAP7_75t_L g18415 ( 
.A1(n_18198),
.A2(n_17995),
.B(n_17787),
.C(n_17883),
.Y(n_18415)
);

NAND2xp5_ASAP7_75t_L g18416 ( 
.A(n_18110),
.B(n_8230),
.Y(n_18416)
);

NOR2xp33_ASAP7_75t_L g18417 ( 
.A(n_18233),
.B(n_9115),
.Y(n_18417)
);

NAND2x1p5_ASAP7_75t_L g18418 ( 
.A(n_18158),
.B(n_18203),
.Y(n_18418)
);

NAND2x1_ASAP7_75t_L g18419 ( 
.A(n_18136),
.B(n_8600),
.Y(n_18419)
);

AND2x4_ASAP7_75t_L g18420 ( 
.A(n_18111),
.B(n_10443),
.Y(n_18420)
);

OR2x2_ASAP7_75t_L g18421 ( 
.A(n_18087),
.B(n_9750),
.Y(n_18421)
);

INVx1_ASAP7_75t_L g18422 ( 
.A(n_18082),
.Y(n_18422)
);

INVx1_ASAP7_75t_L g18423 ( 
.A(n_18083),
.Y(n_18423)
);

NAND2xp5_ASAP7_75t_L g18424 ( 
.A(n_18127),
.B(n_8230),
.Y(n_18424)
);

AOI21xp5_ASAP7_75t_L g18425 ( 
.A1(n_18165),
.A2(n_9763),
.B(n_9759),
.Y(n_18425)
);

OAI222xp33_ASAP7_75t_L g18426 ( 
.A1(n_18234),
.A2(n_9199),
.B1(n_9084),
.B2(n_9216),
.C1(n_9131),
.C2(n_9047),
.Y(n_18426)
);

AOI322xp5_ASAP7_75t_L g18427 ( 
.A1(n_18152),
.A2(n_9774),
.A3(n_9763),
.B1(n_9782),
.B2(n_9795),
.C1(n_9770),
.C2(n_9759),
.Y(n_18427)
);

OAI221xp5_ASAP7_75t_L g18428 ( 
.A1(n_18112),
.A2(n_9131),
.B1(n_9199),
.B2(n_9084),
.C(n_9047),
.Y(n_18428)
);

BUFx2_ASAP7_75t_L g18429 ( 
.A(n_18295),
.Y(n_18429)
);

NAND2xp5_ASAP7_75t_L g18430 ( 
.A(n_18081),
.B(n_8230),
.Y(n_18430)
);

INVx1_ASAP7_75t_L g18431 ( 
.A(n_18056),
.Y(n_18431)
);

OAI22xp5_ASAP7_75t_L g18432 ( 
.A1(n_18266),
.A2(n_10081),
.B1(n_10083),
.B2(n_10077),
.Y(n_18432)
);

INVx2_ASAP7_75t_L g18433 ( 
.A(n_18099),
.Y(n_18433)
);

OAI21xp5_ASAP7_75t_SL g18434 ( 
.A1(n_18201),
.A2(n_8114),
.B(n_8007),
.Y(n_18434)
);

INVx1_ASAP7_75t_L g18435 ( 
.A(n_18116),
.Y(n_18435)
);

AOI21xp33_ASAP7_75t_L g18436 ( 
.A1(n_18090),
.A2(n_18161),
.B(n_18048),
.Y(n_18436)
);

NAND2xp5_ASAP7_75t_L g18437 ( 
.A(n_18104),
.B(n_8233),
.Y(n_18437)
);

CKINVDCx5p33_ASAP7_75t_R g18438 ( 
.A(n_18211),
.Y(n_18438)
);

INVx1_ASAP7_75t_L g18439 ( 
.A(n_18335),
.Y(n_18439)
);

INVx1_ASAP7_75t_L g18440 ( 
.A(n_18324),
.Y(n_18440)
);

OR2x2_ASAP7_75t_L g18441 ( 
.A(n_18107),
.B(n_9770),
.Y(n_18441)
);

INVx1_ASAP7_75t_L g18442 ( 
.A(n_18106),
.Y(n_18442)
);

INVx1_ASAP7_75t_L g18443 ( 
.A(n_18077),
.Y(n_18443)
);

INVx1_ASAP7_75t_L g18444 ( 
.A(n_18033),
.Y(n_18444)
);

AOI21xp33_ASAP7_75t_SL g18445 ( 
.A1(n_18036),
.A2(n_10467),
.B(n_10460),
.Y(n_18445)
);

AOI22xp5_ASAP7_75t_L g18446 ( 
.A1(n_18208),
.A2(n_9774),
.B1(n_9782),
.B2(n_9770),
.Y(n_18446)
);

O2A1O1Ixp33_ASAP7_75t_L g18447 ( 
.A1(n_18156),
.A2(n_8705),
.B(n_8739),
.C(n_8600),
.Y(n_18447)
);

INVx2_ASAP7_75t_L g18448 ( 
.A(n_18031),
.Y(n_18448)
);

INVx1_ASAP7_75t_L g18449 ( 
.A(n_18038),
.Y(n_18449)
);

INVx1_ASAP7_75t_L g18450 ( 
.A(n_18129),
.Y(n_18450)
);

AND2x2_ASAP7_75t_L g18451 ( 
.A(n_18098),
.B(n_10467),
.Y(n_18451)
);

INVx1_ASAP7_75t_L g18452 ( 
.A(n_18046),
.Y(n_18452)
);

AOI21xp5_ASAP7_75t_R g18453 ( 
.A1(n_18147),
.A2(n_7701),
.B(n_7706),
.Y(n_18453)
);

AOI22xp5_ASAP7_75t_L g18454 ( 
.A1(n_18215),
.A2(n_9782),
.B1(n_9795),
.B2(n_9774),
.Y(n_18454)
);

OAI22xp5_ASAP7_75t_L g18455 ( 
.A1(n_18050),
.A2(n_10083),
.B1(n_10084),
.B2(n_10081),
.Y(n_18455)
);

AOI21xp33_ASAP7_75t_L g18456 ( 
.A1(n_18034),
.A2(n_9800),
.B(n_9795),
.Y(n_18456)
);

NAND2xp5_ASAP7_75t_L g18457 ( 
.A(n_18296),
.B(n_8233),
.Y(n_18457)
);

NAND2xp5_ASAP7_75t_L g18458 ( 
.A(n_18301),
.B(n_8233),
.Y(n_18458)
);

AOI22xp5_ASAP7_75t_L g18459 ( 
.A1(n_18194),
.A2(n_9809),
.B1(n_9814),
.B2(n_9800),
.Y(n_18459)
);

INVx1_ASAP7_75t_L g18460 ( 
.A(n_18140),
.Y(n_18460)
);

INVx1_ASAP7_75t_L g18461 ( 
.A(n_18145),
.Y(n_18461)
);

INVx2_ASAP7_75t_L g18462 ( 
.A(n_18225),
.Y(n_18462)
);

NOR2xp33_ASAP7_75t_SL g18463 ( 
.A(n_18288),
.B(n_8705),
.Y(n_18463)
);

AOI211xp5_ASAP7_75t_L g18464 ( 
.A1(n_18044),
.A2(n_10479),
.B(n_9084),
.C(n_9131),
.Y(n_18464)
);

OR2x2_ASAP7_75t_L g18465 ( 
.A(n_18184),
.B(n_9800),
.Y(n_18465)
);

NAND2xp5_ASAP7_75t_L g18466 ( 
.A(n_18185),
.B(n_10081),
.Y(n_18466)
);

NOR2x1_ASAP7_75t_L g18467 ( 
.A(n_18251),
.B(n_8847),
.Y(n_18467)
);

INVx1_ASAP7_75t_L g18468 ( 
.A(n_18178),
.Y(n_18468)
);

OAI22xp33_ASAP7_75t_SL g18469 ( 
.A1(n_18312),
.A2(n_9814),
.B1(n_9823),
.B2(n_9809),
.Y(n_18469)
);

NAND4xp25_ASAP7_75t_L g18470 ( 
.A(n_18035),
.B(n_18134),
.C(n_18080),
.D(n_18221),
.Y(n_18470)
);

INVx1_ASAP7_75t_L g18471 ( 
.A(n_18139),
.Y(n_18471)
);

OAI22xp5_ASAP7_75t_L g18472 ( 
.A1(n_18213),
.A2(n_10084),
.B1(n_10088),
.B2(n_10083),
.Y(n_18472)
);

NAND2xp5_ASAP7_75t_L g18473 ( 
.A(n_18329),
.B(n_10084),
.Y(n_18473)
);

AOI22xp5_ASAP7_75t_L g18474 ( 
.A1(n_18076),
.A2(n_9814),
.B1(n_9823),
.B2(n_9809),
.Y(n_18474)
);

INVx1_ASAP7_75t_L g18475 ( 
.A(n_18317),
.Y(n_18475)
);

INVx1_ASAP7_75t_L g18476 ( 
.A(n_18146),
.Y(n_18476)
);

AOI22xp5_ASAP7_75t_L g18477 ( 
.A1(n_18092),
.A2(n_18053),
.B1(n_18183),
.B2(n_18196),
.Y(n_18477)
);

INVxp67_ASAP7_75t_L g18478 ( 
.A(n_18200),
.Y(n_18478)
);

A2O1A1Ixp33_ASAP7_75t_L g18479 ( 
.A1(n_18263),
.A2(n_10479),
.B(n_10096),
.C(n_10127),
.Y(n_18479)
);

INVx1_ASAP7_75t_L g18480 ( 
.A(n_18236),
.Y(n_18480)
);

NOR4xp25_ASAP7_75t_L g18481 ( 
.A(n_18358),
.B(n_9837),
.C(n_9841),
.D(n_9823),
.Y(n_18481)
);

AND2x2_ASAP7_75t_L g18482 ( 
.A(n_18252),
.B(n_7029),
.Y(n_18482)
);

OR2x2_ASAP7_75t_L g18483 ( 
.A(n_18265),
.B(n_9837),
.Y(n_18483)
);

NAND2x1p5_ASAP7_75t_L g18484 ( 
.A(n_18135),
.B(n_8656),
.Y(n_18484)
);

HB1xp67_ASAP7_75t_L g18485 ( 
.A(n_18132),
.Y(n_18485)
);

AOI322xp5_ASAP7_75t_L g18486 ( 
.A1(n_18284),
.A2(n_9841),
.A3(n_9837),
.B1(n_10096),
.B2(n_10127),
.C1(n_10128),
.C2(n_10088),
.Y(n_18486)
);

AND2x2_ASAP7_75t_L g18487 ( 
.A(n_18070),
.B(n_7029),
.Y(n_18487)
);

INVxp67_ASAP7_75t_L g18488 ( 
.A(n_18095),
.Y(n_18488)
);

BUFx3_ASAP7_75t_L g18489 ( 
.A(n_18248),
.Y(n_18489)
);

NAND2xp5_ASAP7_75t_L g18490 ( 
.A(n_18330),
.B(n_10088),
.Y(n_18490)
);

INVx1_ASAP7_75t_L g18491 ( 
.A(n_18159),
.Y(n_18491)
);

INVx1_ASAP7_75t_L g18492 ( 
.A(n_18125),
.Y(n_18492)
);

NAND2xp5_ASAP7_75t_L g18493 ( 
.A(n_18339),
.B(n_10096),
.Y(n_18493)
);

AOI211x1_ASAP7_75t_L g18494 ( 
.A1(n_18332),
.A2(n_8852),
.B(n_8782),
.C(n_8359),
.Y(n_18494)
);

AOI22xp33_ASAP7_75t_L g18495 ( 
.A1(n_18193),
.A2(n_9047),
.B1(n_9216),
.B2(n_9199),
.Y(n_18495)
);

OAI22xp5_ASAP7_75t_L g18496 ( 
.A1(n_18228),
.A2(n_10127),
.B1(n_10128),
.B2(n_9841),
.Y(n_18496)
);

AOI221xp5_ASAP7_75t_L g18497 ( 
.A1(n_18218),
.A2(n_10128),
.B1(n_8739),
.B2(n_9064),
.C(n_8728),
.Y(n_18497)
);

NAND2xp5_ASAP7_75t_L g18498 ( 
.A(n_18340),
.B(n_8251),
.Y(n_18498)
);

OAI32xp33_ASAP7_75t_L g18499 ( 
.A1(n_18182),
.A2(n_8329),
.A3(n_8381),
.B1(n_8208),
.B2(n_8114),
.Y(n_18499)
);

AOI21xp33_ASAP7_75t_L g18500 ( 
.A1(n_18166),
.A2(n_8739),
.B(n_8760),
.Y(n_18500)
);

INVx2_ASAP7_75t_L g18501 ( 
.A(n_18126),
.Y(n_18501)
);

INVx1_ASAP7_75t_L g18502 ( 
.A(n_18320),
.Y(n_18502)
);

INVx1_ASAP7_75t_L g18503 ( 
.A(n_18363),
.Y(n_18503)
);

INVx1_ASAP7_75t_L g18504 ( 
.A(n_18365),
.Y(n_18504)
);

INVx2_ASAP7_75t_L g18505 ( 
.A(n_18230),
.Y(n_18505)
);

INVx3_ASAP7_75t_L g18506 ( 
.A(n_18084),
.Y(n_18506)
);

AOI22xp5_ASAP7_75t_L g18507 ( 
.A1(n_18060),
.A2(n_9304),
.B1(n_9216),
.B2(n_8728),
.Y(n_18507)
);

INVx1_ASAP7_75t_L g18508 ( 
.A(n_18323),
.Y(n_18508)
);

NAND2xp5_ASAP7_75t_L g18509 ( 
.A(n_18344),
.B(n_8251),
.Y(n_18509)
);

OR2x2_ASAP7_75t_L g18510 ( 
.A(n_18319),
.B(n_9115),
.Y(n_18510)
);

OAI21xp33_ASAP7_75t_L g18511 ( 
.A1(n_18214),
.A2(n_18222),
.B(n_18131),
.Y(n_18511)
);

INVx1_ASAP7_75t_L g18512 ( 
.A(n_18117),
.Y(n_18512)
);

INVx1_ASAP7_75t_L g18513 ( 
.A(n_18168),
.Y(n_18513)
);

INVx2_ASAP7_75t_SL g18514 ( 
.A(n_18204),
.Y(n_18514)
);

OAI22xp5_ASAP7_75t_L g18515 ( 
.A1(n_18173),
.A2(n_9304),
.B1(n_8749),
.B2(n_8841),
.Y(n_18515)
);

AOI21xp33_ASAP7_75t_SL g18516 ( 
.A1(n_18232),
.A2(n_10141),
.B(n_10136),
.Y(n_18516)
);

NAND2xp5_ASAP7_75t_SL g18517 ( 
.A(n_18085),
.B(n_9304),
.Y(n_18517)
);

OAI22xp33_ASAP7_75t_L g18518 ( 
.A1(n_18292),
.A2(n_9177),
.B1(n_9222),
.B2(n_9132),
.Y(n_18518)
);

AOI211xp5_ASAP7_75t_L g18519 ( 
.A1(n_18311),
.A2(n_8723),
.B(n_8656),
.C(n_10136),
.Y(n_18519)
);

AND2x2_ASAP7_75t_L g18520 ( 
.A(n_18069),
.B(n_7029),
.Y(n_18520)
);

INVx1_ASAP7_75t_L g18521 ( 
.A(n_18169),
.Y(n_18521)
);

INVx1_ASAP7_75t_L g18522 ( 
.A(n_18179),
.Y(n_18522)
);

O2A1O1Ixp33_ASAP7_75t_SL g18523 ( 
.A1(n_18148),
.A2(n_9177),
.B(n_9222),
.C(n_9132),
.Y(n_18523)
);

INVx1_ASAP7_75t_L g18524 ( 
.A(n_18160),
.Y(n_18524)
);

AND2x2_ASAP7_75t_L g18525 ( 
.A(n_18042),
.B(n_7029),
.Y(n_18525)
);

OAI221xp5_ASAP7_75t_L g18526 ( 
.A1(n_18063),
.A2(n_8114),
.B1(n_8381),
.B2(n_8329),
.C(n_8208),
.Y(n_18526)
);

INVx1_ASAP7_75t_L g18527 ( 
.A(n_18157),
.Y(n_18527)
);

NOR2x1_ASAP7_75t_L g18528 ( 
.A(n_18255),
.B(n_8893),
.Y(n_18528)
);

AOI21xp33_ASAP7_75t_L g18529 ( 
.A1(n_18325),
.A2(n_8762),
.B(n_8760),
.Y(n_18529)
);

INVxp67_ASAP7_75t_L g18530 ( 
.A(n_18207),
.Y(n_18530)
);

OAI32xp33_ASAP7_75t_L g18531 ( 
.A1(n_18175),
.A2(n_8329),
.A3(n_8381),
.B1(n_8208),
.B2(n_8114),
.Y(n_18531)
);

INVx1_ASAP7_75t_L g18532 ( 
.A(n_18283),
.Y(n_18532)
);

INVx1_ASAP7_75t_L g18533 ( 
.A(n_18334),
.Y(n_18533)
);

AOI21xp5_ASAP7_75t_L g18534 ( 
.A1(n_18278),
.A2(n_8068),
.B(n_8252),
.Y(n_18534)
);

NAND3xp33_ASAP7_75t_L g18535 ( 
.A(n_18121),
.B(n_9249),
.C(n_9232),
.Y(n_18535)
);

NAND2xp5_ASAP7_75t_L g18536 ( 
.A(n_18350),
.B(n_8252),
.Y(n_18536)
);

INVxp67_ASAP7_75t_L g18537 ( 
.A(n_18181),
.Y(n_18537)
);

AOI21xp33_ASAP7_75t_SL g18538 ( 
.A1(n_18188),
.A2(n_10163),
.B(n_10141),
.Y(n_18538)
);

AND2x2_ASAP7_75t_SL g18539 ( 
.A(n_18359),
.B(n_7633),
.Y(n_18539)
);

NAND2xp5_ASAP7_75t_L g18540 ( 
.A(n_18261),
.B(n_18224),
.Y(n_18540)
);

INVx1_ASAP7_75t_L g18541 ( 
.A(n_18338),
.Y(n_18541)
);

INVx1_ASAP7_75t_L g18542 ( 
.A(n_18347),
.Y(n_18542)
);

OAI21xp33_ASAP7_75t_SL g18543 ( 
.A1(n_18209),
.A2(n_10163),
.B(n_8723),
.Y(n_18543)
);

OAI22xp33_ASAP7_75t_L g18544 ( 
.A1(n_18302),
.A2(n_9249),
.B1(n_9268),
.B2(n_9232),
.Y(n_18544)
);

AOI21xp5_ASAP7_75t_R g18545 ( 
.A1(n_18130),
.A2(n_7701),
.B(n_7706),
.Y(n_18545)
);

AOI21xp5_ASAP7_75t_L g18546 ( 
.A1(n_18271),
.A2(n_8068),
.B(n_8252),
.Y(n_18546)
);

INVx2_ASAP7_75t_L g18547 ( 
.A(n_18171),
.Y(n_18547)
);

OR2x2_ASAP7_75t_L g18548 ( 
.A(n_18356),
.B(n_9268),
.Y(n_18548)
);

OR2x2_ASAP7_75t_L g18549 ( 
.A(n_18150),
.B(n_8893),
.Y(n_18549)
);

NOR3xp33_ASAP7_75t_L g18550 ( 
.A(n_18138),
.B(n_8723),
.C(n_8656),
.Y(n_18550)
);

OAI21xp5_ASAP7_75t_L g18551 ( 
.A1(n_18244),
.A2(n_8821),
.B(n_8477),
.Y(n_18551)
);

INVx1_ASAP7_75t_L g18552 ( 
.A(n_18186),
.Y(n_18552)
);

NOR4xp25_ASAP7_75t_SL g18553 ( 
.A(n_18314),
.B(n_8841),
.C(n_8916),
.D(n_7944),
.Y(n_18553)
);

OAI22xp5_ASAP7_75t_L g18554 ( 
.A1(n_18331),
.A2(n_18304),
.B1(n_18190),
.B2(n_18187),
.Y(n_18554)
);

OAI21xp5_ASAP7_75t_L g18555 ( 
.A1(n_18176),
.A2(n_8821),
.B(n_8477),
.Y(n_18555)
);

NOR2xp33_ASAP7_75t_L g18556 ( 
.A(n_18163),
.B(n_9053),
.Y(n_18556)
);

OR2x2_ASAP7_75t_L g18557 ( 
.A(n_18290),
.B(n_8893),
.Y(n_18557)
);

NOR2xp33_ASAP7_75t_L g18558 ( 
.A(n_18357),
.B(n_9053),
.Y(n_18558)
);

INVx1_ASAP7_75t_L g18559 ( 
.A(n_18285),
.Y(n_18559)
);

INVx1_ASAP7_75t_L g18560 ( 
.A(n_18253),
.Y(n_18560)
);

AOI31xp33_ASAP7_75t_L g18561 ( 
.A1(n_18322),
.A2(n_8329),
.A3(n_8381),
.B(n_8208),
.Y(n_18561)
);

INVx2_ASAP7_75t_L g18562 ( 
.A(n_18308),
.Y(n_18562)
);

BUFx2_ASAP7_75t_L g18563 ( 
.A(n_18054),
.Y(n_18563)
);

AOI22xp5_ASAP7_75t_L g18564 ( 
.A1(n_18144),
.A2(n_8916),
.B1(n_8893),
.B2(n_8895),
.Y(n_18564)
);

OAI22xp5_ASAP7_75t_SL g18565 ( 
.A1(n_18366),
.A2(n_8329),
.B1(n_8427),
.B2(n_8381),
.Y(n_18565)
);

AOI22xp5_ASAP7_75t_L g18566 ( 
.A1(n_18154),
.A2(n_8893),
.B1(n_8895),
.B2(n_8790),
.Y(n_18566)
);

INVxp67_ASAP7_75t_SL g18567 ( 
.A(n_18142),
.Y(n_18567)
);

AOI21xp33_ASAP7_75t_L g18568 ( 
.A1(n_18216),
.A2(n_8762),
.B(n_8760),
.Y(n_18568)
);

INVx1_ASAP7_75t_L g18569 ( 
.A(n_18277),
.Y(n_18569)
);

OAI21xp5_ASAP7_75t_SL g18570 ( 
.A1(n_18137),
.A2(n_8435),
.B(n_8427),
.Y(n_18570)
);

AND2x2_ASAP7_75t_L g18571 ( 
.A(n_18240),
.B(n_9057),
.Y(n_18571)
);

AOI21xp5_ASAP7_75t_L g18572 ( 
.A1(n_18206),
.A2(n_8068),
.B(n_8790),
.Y(n_18572)
);

INVx1_ASAP7_75t_L g18573 ( 
.A(n_18291),
.Y(n_18573)
);

OAI22xp5_ASAP7_75t_L g18574 ( 
.A1(n_18153),
.A2(n_8435),
.B1(n_8525),
.B2(n_8427),
.Y(n_18574)
);

OAI22xp33_ASAP7_75t_L g18575 ( 
.A1(n_18066),
.A2(n_8435),
.B1(n_8525),
.B2(n_8427),
.Y(n_18575)
);

OAI21xp33_ASAP7_75t_L g18576 ( 
.A1(n_18151),
.A2(n_18167),
.B(n_18174),
.Y(n_18576)
);

INVx1_ASAP7_75t_L g18577 ( 
.A(n_18299),
.Y(n_18577)
);

OAI22xp5_ASAP7_75t_L g18578 ( 
.A1(n_18249),
.A2(n_8435),
.B1(n_8525),
.B2(n_8427),
.Y(n_18578)
);

O2A1O1Ixp33_ASAP7_75t_SL g18579 ( 
.A1(n_18075),
.A2(n_7482),
.B(n_7497),
.C(n_7491),
.Y(n_18579)
);

INVxp67_ASAP7_75t_L g18580 ( 
.A(n_18316),
.Y(n_18580)
);

INVx1_ASAP7_75t_L g18581 ( 
.A(n_18094),
.Y(n_18581)
);

INVx2_ASAP7_75t_L g18582 ( 
.A(n_18231),
.Y(n_18582)
);

AOI21xp5_ASAP7_75t_L g18583 ( 
.A1(n_18309),
.A2(n_8794),
.B(n_8790),
.Y(n_18583)
);

NAND2xp5_ASAP7_75t_L g18584 ( 
.A(n_18172),
.B(n_8760),
.Y(n_18584)
);

INVx1_ASAP7_75t_SL g18585 ( 
.A(n_18037),
.Y(n_18585)
);

OAI211xp5_ASAP7_75t_L g18586 ( 
.A1(n_18242),
.A2(n_8359),
.B(n_8852),
.C(n_8782),
.Y(n_18586)
);

OAI21xp33_ASAP7_75t_SL g18587 ( 
.A1(n_18256),
.A2(n_7962),
.B(n_7959),
.Y(n_18587)
);

AOI22xp33_ASAP7_75t_SL g18588 ( 
.A1(n_18243),
.A2(n_9064),
.B1(n_7101),
.B2(n_7210),
.Y(n_18588)
);

AOI22xp33_ASAP7_75t_L g18589 ( 
.A1(n_18362),
.A2(n_8657),
.B1(n_8895),
.B2(n_8785),
.Y(n_18589)
);

AND2x2_ASAP7_75t_L g18590 ( 
.A(n_18054),
.B(n_9057),
.Y(n_18590)
);

OAI22xp5_ASAP7_75t_L g18591 ( 
.A1(n_18162),
.A2(n_8525),
.B1(n_8609),
.B2(n_8435),
.Y(n_18591)
);

AND2x2_ASAP7_75t_L g18592 ( 
.A(n_18118),
.B(n_9057),
.Y(n_18592)
);

AND2x4_ASAP7_75t_L g18593 ( 
.A(n_18351),
.B(n_8036),
.Y(n_18593)
);

NOR2x1_ASAP7_75t_L g18594 ( 
.A(n_18217),
.B(n_8790),
.Y(n_18594)
);

HB1xp67_ASAP7_75t_L g18595 ( 
.A(n_18259),
.Y(n_18595)
);

AOI22xp5_ASAP7_75t_L g18596 ( 
.A1(n_18128),
.A2(n_8895),
.B1(n_8794),
.B2(n_8790),
.Y(n_18596)
);

INVx1_ASAP7_75t_L g18597 ( 
.A(n_18102),
.Y(n_18597)
);

NAND2xp5_ASAP7_75t_L g18598 ( 
.A(n_18345),
.B(n_8762),
.Y(n_18598)
);

INVx1_ASAP7_75t_L g18599 ( 
.A(n_18057),
.Y(n_18599)
);

NAND2xp5_ASAP7_75t_L g18600 ( 
.A(n_18349),
.B(n_8762),
.Y(n_18600)
);

OAI22xp5_ASAP7_75t_SL g18601 ( 
.A1(n_18219),
.A2(n_8525),
.B1(n_8747),
.B2(n_8609),
.Y(n_18601)
);

OAI21xp5_ASAP7_75t_L g18602 ( 
.A1(n_18155),
.A2(n_8821),
.B(n_8549),
.Y(n_18602)
);

NAND2xp5_ASAP7_75t_L g18603 ( 
.A(n_18120),
.B(n_8785),
.Y(n_18603)
);

INVx1_ASAP7_75t_L g18604 ( 
.A(n_18133),
.Y(n_18604)
);

A2O1A1Ixp33_ASAP7_75t_L g18605 ( 
.A1(n_18124),
.A2(n_8067),
.B(n_8052),
.C(n_8324),
.Y(n_18605)
);

NAND2xp5_ASAP7_75t_L g18606 ( 
.A(n_18141),
.B(n_8785),
.Y(n_18606)
);

NOR3xp33_ASAP7_75t_L g18607 ( 
.A(n_18355),
.B(n_8462),
.C(n_8215),
.Y(n_18607)
);

OAI22xp5_ASAP7_75t_L g18608 ( 
.A1(n_18275),
.A2(n_8609),
.B1(n_8768),
.B2(n_8747),
.Y(n_18608)
);

AOI21xp5_ASAP7_75t_L g18609 ( 
.A1(n_18259),
.A2(n_8794),
.B(n_8785),
.Y(n_18609)
);

INVx1_ASAP7_75t_L g18610 ( 
.A(n_18220),
.Y(n_18610)
);

AOI22xp5_ASAP7_75t_L g18611 ( 
.A1(n_18143),
.A2(n_8895),
.B1(n_8794),
.B2(n_7535),
.Y(n_18611)
);

INVx1_ASAP7_75t_L g18612 ( 
.A(n_18267),
.Y(n_18612)
);

NOR3xp33_ASAP7_75t_L g18613 ( 
.A(n_18364),
.B(n_8462),
.C(n_8215),
.Y(n_18613)
);

NAND2xp5_ASAP7_75t_L g18614 ( 
.A(n_18254),
.B(n_18226),
.Y(n_18614)
);

OAI32xp33_ASAP7_75t_L g18615 ( 
.A1(n_18115),
.A2(n_8747),
.A3(n_8781),
.B1(n_8768),
.B2(n_8609),
.Y(n_18615)
);

INVx1_ASAP7_75t_SL g18616 ( 
.A(n_18047),
.Y(n_18616)
);

NAND2xp5_ASAP7_75t_L g18617 ( 
.A(n_18227),
.B(n_8785),
.Y(n_18617)
);

NAND3xp33_ASAP7_75t_L g18618 ( 
.A(n_18270),
.B(n_7053),
.C(n_7020),
.Y(n_18618)
);

INVx1_ASAP7_75t_L g18619 ( 
.A(n_18272),
.Y(n_18619)
);

INVxp67_ASAP7_75t_SL g18620 ( 
.A(n_18273),
.Y(n_18620)
);

NOR2xp67_ASAP7_75t_SL g18621 ( 
.A(n_18262),
.B(n_5751),
.Y(n_18621)
);

NAND2xp5_ASAP7_75t_L g18622 ( 
.A(n_18274),
.B(n_8794),
.Y(n_18622)
);

INVx2_ASAP7_75t_L g18623 ( 
.A(n_18294),
.Y(n_18623)
);

OAI22xp5_ASAP7_75t_L g18624 ( 
.A1(n_18264),
.A2(n_8609),
.B1(n_8768),
.B2(n_8747),
.Y(n_18624)
);

NAND2xp5_ASAP7_75t_L g18625 ( 
.A(n_18281),
.B(n_8285),
.Y(n_18625)
);

INVx1_ASAP7_75t_L g18626 ( 
.A(n_18258),
.Y(n_18626)
);

NAND2xp5_ASAP7_75t_L g18627 ( 
.A(n_18287),
.B(n_8285),
.Y(n_18627)
);

AND2x2_ASAP7_75t_L g18628 ( 
.A(n_18177),
.B(n_8299),
.Y(n_18628)
);

INVx1_ASAP7_75t_L g18629 ( 
.A(n_18257),
.Y(n_18629)
);

OR2x2_ASAP7_75t_L g18630 ( 
.A(n_18192),
.B(n_8903),
.Y(n_18630)
);

INVx1_ASAP7_75t_L g18631 ( 
.A(n_18315),
.Y(n_18631)
);

INVx1_ASAP7_75t_L g18632 ( 
.A(n_18326),
.Y(n_18632)
);

NAND2xp5_ASAP7_75t_L g18633 ( 
.A(n_18328),
.B(n_8285),
.Y(n_18633)
);

NAND2xp5_ASAP7_75t_L g18634 ( 
.A(n_18346),
.B(n_8285),
.Y(n_18634)
);

INVx2_ASAP7_75t_L g18635 ( 
.A(n_18298),
.Y(n_18635)
);

OAI22xp33_ASAP7_75t_SL g18636 ( 
.A1(n_18289),
.A2(n_8747),
.B1(n_8781),
.B2(n_8768),
.Y(n_18636)
);

OAI332xp33_ASAP7_75t_L g18637 ( 
.A1(n_18353),
.A2(n_8737),
.A3(n_8694),
.B1(n_8718),
.B2(n_8493),
.B3(n_7254),
.C1(n_7307),
.C2(n_7234),
.Y(n_18637)
);

INVx1_ASAP7_75t_L g18638 ( 
.A(n_18108),
.Y(n_18638)
);

INVx2_ASAP7_75t_L g18639 ( 
.A(n_18303),
.Y(n_18639)
);

INVx1_ASAP7_75t_L g18640 ( 
.A(n_18348),
.Y(n_18640)
);

OAI22xp5_ASAP7_75t_L g18641 ( 
.A1(n_18305),
.A2(n_18223),
.B1(n_18342),
.B2(n_18336),
.Y(n_18641)
);

AND2x2_ASAP7_75t_L g18642 ( 
.A(n_18341),
.B(n_8299),
.Y(n_18642)
);

NAND2xp5_ASAP7_75t_L g18643 ( 
.A(n_18310),
.B(n_8315),
.Y(n_18643)
);

INVx1_ASAP7_75t_L g18644 ( 
.A(n_18093),
.Y(n_18644)
);

OAI21xp5_ASAP7_75t_L g18645 ( 
.A1(n_18247),
.A2(n_8549),
.B(n_8462),
.Y(n_18645)
);

NOR2x1_ASAP7_75t_L g18646 ( 
.A(n_18239),
.B(n_8546),
.Y(n_18646)
);

INVx1_ASAP7_75t_SL g18647 ( 
.A(n_18300),
.Y(n_18647)
);

OAI221xp5_ASAP7_75t_L g18648 ( 
.A1(n_18327),
.A2(n_8781),
.B1(n_8834),
.B2(n_8800),
.C(n_8768),
.Y(n_18648)
);

AND2x4_ASAP7_75t_L g18649 ( 
.A(n_18367),
.B(n_8036),
.Y(n_18649)
);

INVx1_ASAP7_75t_L g18650 ( 
.A(n_18205),
.Y(n_18650)
);

INVx2_ASAP7_75t_L g18651 ( 
.A(n_18318),
.Y(n_18651)
);

AOI33xp33_ASAP7_75t_L g18652 ( 
.A1(n_18237),
.A2(n_7497),
.A3(n_7491),
.B1(n_7482),
.B2(n_7036),
.B3(n_7633),
.Y(n_18652)
);

NAND2xp5_ASAP7_75t_L g18653 ( 
.A(n_18269),
.B(n_8315),
.Y(n_18653)
);

NAND2xp5_ASAP7_75t_L g18654 ( 
.A(n_18371),
.B(n_18286),
.Y(n_18654)
);

INVx1_ASAP7_75t_SL g18655 ( 
.A(n_18372),
.Y(n_18655)
);

AOI21xp5_ASAP7_75t_L g18656 ( 
.A1(n_18380),
.A2(n_18361),
.B(n_18360),
.Y(n_18656)
);

AND2x2_ASAP7_75t_L g18657 ( 
.A(n_18439),
.B(n_18280),
.Y(n_18657)
);

NAND2xp5_ASAP7_75t_L g18658 ( 
.A(n_18386),
.B(n_18373),
.Y(n_18658)
);

NAND2xp5_ASAP7_75t_L g18659 ( 
.A(n_18377),
.B(n_18321),
.Y(n_18659)
);

OAI22xp33_ASAP7_75t_L g18660 ( 
.A1(n_18369),
.A2(n_18343),
.B1(n_18235),
.B2(n_18307),
.Y(n_18660)
);

OAI32xp33_ASAP7_75t_L g18661 ( 
.A1(n_18418),
.A2(n_18250),
.A3(n_18268),
.B1(n_18260),
.B2(n_18241),
.Y(n_18661)
);

NAND2xp5_ASAP7_75t_L g18662 ( 
.A(n_18389),
.B(n_18400),
.Y(n_18662)
);

AOI22xp33_ASAP7_75t_L g18663 ( 
.A1(n_18392),
.A2(n_18352),
.B1(n_18297),
.B2(n_18199),
.Y(n_18663)
);

HB1xp67_ASAP7_75t_L g18664 ( 
.A(n_18406),
.Y(n_18664)
);

INVxp67_ASAP7_75t_L g18665 ( 
.A(n_18405),
.Y(n_18665)
);

OAI22xp5_ASAP7_75t_L g18666 ( 
.A1(n_18398),
.A2(n_18337),
.B1(n_18282),
.B2(n_18238),
.Y(n_18666)
);

INVx1_ASAP7_75t_L g18667 ( 
.A(n_18485),
.Y(n_18667)
);

INVxp67_ASAP7_75t_L g18668 ( 
.A(n_18388),
.Y(n_18668)
);

AOI21xp5_ASAP7_75t_L g18669 ( 
.A1(n_18368),
.A2(n_18246),
.B(n_18123),
.Y(n_18669)
);

NAND2xp5_ASAP7_75t_L g18670 ( 
.A(n_18374),
.B(n_18313),
.Y(n_18670)
);

AOI22x1_ASAP7_75t_L g18671 ( 
.A1(n_18429),
.A2(n_18105),
.B1(n_18096),
.B2(n_18333),
.Y(n_18671)
);

NOR3xp33_ASAP7_75t_SL g18672 ( 
.A(n_18438),
.B(n_18180),
.C(n_18306),
.Y(n_18672)
);

NOR2xp33_ASAP7_75t_L g18673 ( 
.A(n_18537),
.B(n_18051),
.Y(n_18673)
);

AOI332xp33_ASAP7_75t_L g18674 ( 
.A1(n_18393),
.A2(n_8795),
.A3(n_8779),
.B1(n_8803),
.B2(n_8798),
.B3(n_8820),
.C1(n_8786),
.C2(n_8777),
.Y(n_18674)
);

INVx2_ASAP7_75t_SL g18675 ( 
.A(n_18379),
.Y(n_18675)
);

NAND2xp5_ASAP7_75t_L g18676 ( 
.A(n_18442),
.B(n_18401),
.Y(n_18676)
);

OAI321xp33_ASAP7_75t_L g18677 ( 
.A1(n_18381),
.A2(n_8781),
.A3(n_8800),
.B1(n_8944),
.B2(n_8868),
.C(n_8834),
.Y(n_18677)
);

AOI22xp5_ASAP7_75t_L g18678 ( 
.A1(n_18408),
.A2(n_7535),
.B1(n_7408),
.B2(n_8546),
.Y(n_18678)
);

NAND2xp5_ASAP7_75t_SL g18679 ( 
.A(n_18407),
.B(n_7020),
.Y(n_18679)
);

NOR2xp33_ASAP7_75t_L g18680 ( 
.A(n_18478),
.B(n_9053),
.Y(n_18680)
);

AOI22xp33_ASAP7_75t_SL g18681 ( 
.A1(n_18489),
.A2(n_9064),
.B1(n_7101),
.B2(n_7210),
.Y(n_18681)
);

NAND2xp5_ASAP7_75t_SL g18682 ( 
.A(n_18539),
.B(n_7020),
.Y(n_18682)
);

NAND2xp5_ASAP7_75t_SL g18683 ( 
.A(n_18463),
.B(n_7020),
.Y(n_18683)
);

NAND2xp5_ASAP7_75t_L g18684 ( 
.A(n_18383),
.B(n_8315),
.Y(n_18684)
);

O2A1O1Ixp33_ASAP7_75t_SL g18685 ( 
.A1(n_18399),
.A2(n_7482),
.B(n_7497),
.C(n_7491),
.Y(n_18685)
);

OAI31xp33_ASAP7_75t_L g18686 ( 
.A1(n_18415),
.A2(n_8800),
.A3(n_8834),
.B(n_8781),
.Y(n_18686)
);

NOR2xp33_ASAP7_75t_L g18687 ( 
.A(n_18440),
.B(n_9053),
.Y(n_18687)
);

A2O1A1Ixp33_ASAP7_75t_L g18688 ( 
.A1(n_18376),
.A2(n_8067),
.B(n_8052),
.C(n_8215),
.Y(n_18688)
);

NAND3xp33_ASAP7_75t_L g18689 ( 
.A(n_18375),
.B(n_7053),
.C(n_7020),
.Y(n_18689)
);

INVxp33_ASAP7_75t_L g18690 ( 
.A(n_18370),
.Y(n_18690)
);

OAI22xp5_ASAP7_75t_L g18691 ( 
.A1(n_18545),
.A2(n_8800),
.B1(n_8868),
.B2(n_8834),
.Y(n_18691)
);

INVx1_ASAP7_75t_L g18692 ( 
.A(n_18410),
.Y(n_18692)
);

OAI21xp5_ASAP7_75t_L g18693 ( 
.A1(n_18378),
.A2(n_18530),
.B(n_18488),
.Y(n_18693)
);

INVx3_ASAP7_75t_L g18694 ( 
.A(n_18506),
.Y(n_18694)
);

INVxp67_ASAP7_75t_L g18695 ( 
.A(n_18552),
.Y(n_18695)
);

INVx2_ASAP7_75t_L g18696 ( 
.A(n_18462),
.Y(n_18696)
);

INVx1_ASAP7_75t_L g18697 ( 
.A(n_18548),
.Y(n_18697)
);

INVx1_ASAP7_75t_L g18698 ( 
.A(n_18468),
.Y(n_18698)
);

OAI21xp33_ASAP7_75t_L g18699 ( 
.A1(n_18470),
.A2(n_18511),
.B(n_18390),
.Y(n_18699)
);

INVx2_ASAP7_75t_L g18700 ( 
.A(n_18510),
.Y(n_18700)
);

NAND2xp5_ASAP7_75t_L g18701 ( 
.A(n_18444),
.B(n_8315),
.Y(n_18701)
);

AND2x2_ASAP7_75t_L g18702 ( 
.A(n_18505),
.B(n_8299),
.Y(n_18702)
);

INVx1_ASAP7_75t_L g18703 ( 
.A(n_18475),
.Y(n_18703)
);

AOI21xp33_ASAP7_75t_SL g18704 ( 
.A1(n_18382),
.A2(n_8834),
.B(n_8800),
.Y(n_18704)
);

INVx1_ASAP7_75t_L g18705 ( 
.A(n_18503),
.Y(n_18705)
);

AOI32xp33_ASAP7_75t_L g18706 ( 
.A1(n_18460),
.A2(n_8476),
.A3(n_8549),
.B1(n_8283),
.B2(n_8638),
.Y(n_18706)
);

INVx1_ASAP7_75t_L g18707 ( 
.A(n_18504),
.Y(n_18707)
);

OAI21xp33_ASAP7_75t_L g18708 ( 
.A1(n_18471),
.A2(n_8493),
.B(n_8694),
.Y(n_18708)
);

INVxp67_ASAP7_75t_L g18709 ( 
.A(n_18540),
.Y(n_18709)
);

INVx1_ASAP7_75t_L g18710 ( 
.A(n_18532),
.Y(n_18710)
);

INVx2_ASAP7_75t_L g18711 ( 
.A(n_18419),
.Y(n_18711)
);

NAND2xp5_ASAP7_75t_SL g18712 ( 
.A(n_18385),
.B(n_7020),
.Y(n_18712)
);

INVx1_ASAP7_75t_SL g18713 ( 
.A(n_18585),
.Y(n_18713)
);

OAI221xp5_ASAP7_75t_L g18714 ( 
.A1(n_18384),
.A2(n_18404),
.B1(n_18397),
.B2(n_18396),
.C(n_18403),
.Y(n_18714)
);

OAI322xp33_ASAP7_75t_L g18715 ( 
.A1(n_18580),
.A2(n_8493),
.A3(n_8694),
.B1(n_8718),
.B2(n_8737),
.C1(n_8944),
.C2(n_8868),
.Y(n_18715)
);

INVx2_ASAP7_75t_L g18716 ( 
.A(n_18433),
.Y(n_18716)
);

INVx1_ASAP7_75t_L g18717 ( 
.A(n_18533),
.Y(n_18717)
);

NAND2xp5_ASAP7_75t_L g18718 ( 
.A(n_18422),
.B(n_8322),
.Y(n_18718)
);

INVx1_ASAP7_75t_L g18719 ( 
.A(n_18541),
.Y(n_18719)
);

AOI22xp5_ASAP7_75t_L g18720 ( 
.A1(n_18480),
.A2(n_7535),
.B1(n_8546),
.B2(n_7101),
.Y(n_18720)
);

AOI21xp5_ASAP7_75t_L g18721 ( 
.A1(n_18395),
.A2(n_8245),
.B(n_8235),
.Y(n_18721)
);

OAI322xp33_ASAP7_75t_L g18722 ( 
.A1(n_18402),
.A2(n_8737),
.A3(n_8718),
.B1(n_8868),
.B2(n_9072),
.C1(n_9024),
.C2(n_8944),
.Y(n_18722)
);

AND2x2_ASAP7_75t_L g18723 ( 
.A(n_18502),
.B(n_8299),
.Y(n_18723)
);

AND2x2_ASAP7_75t_L g18724 ( 
.A(n_18448),
.B(n_8299),
.Y(n_18724)
);

AND2x2_ASAP7_75t_L g18725 ( 
.A(n_18562),
.B(n_8299),
.Y(n_18725)
);

AOI22xp33_ASAP7_75t_L g18726 ( 
.A1(n_18461),
.A2(n_18559),
.B1(n_18542),
.B2(n_18560),
.Y(n_18726)
);

NOR3xp33_ASAP7_75t_SL g18727 ( 
.A(n_18436),
.B(n_18414),
.C(n_18412),
.Y(n_18727)
);

NAND2xp5_ASAP7_75t_L g18728 ( 
.A(n_18506),
.B(n_8322),
.Y(n_18728)
);

INVx1_ASAP7_75t_L g18729 ( 
.A(n_18431),
.Y(n_18729)
);

INVx1_ASAP7_75t_L g18730 ( 
.A(n_18443),
.Y(n_18730)
);

NOR3xp33_ASAP7_75t_L g18731 ( 
.A(n_18394),
.B(n_5120),
.C(n_5066),
.Y(n_18731)
);

NAND2xp33_ASAP7_75t_SL g18732 ( 
.A(n_18621),
.B(n_7535),
.Y(n_18732)
);

AOI22xp33_ASAP7_75t_SL g18733 ( 
.A1(n_18409),
.A2(n_7101),
.B1(n_7210),
.B2(n_7020),
.Y(n_18733)
);

OR2x2_ASAP7_75t_L g18734 ( 
.A(n_18423),
.B(n_8299),
.Y(n_18734)
);

INVxp67_ASAP7_75t_L g18735 ( 
.A(n_18417),
.Y(n_18735)
);

AOI221xp5_ASAP7_75t_L g18736 ( 
.A1(n_18411),
.A2(n_8440),
.B1(n_8431),
.B2(n_8048),
.C(n_7497),
.Y(n_18736)
);

NAND2xp5_ASAP7_75t_L g18737 ( 
.A(n_18616),
.B(n_8322),
.Y(n_18737)
);

OAI32xp33_ASAP7_75t_L g18738 ( 
.A1(n_18413),
.A2(n_9024),
.A3(n_9072),
.B1(n_8944),
.B2(n_8868),
.Y(n_18738)
);

OAI22xp5_ASAP7_75t_L g18739 ( 
.A1(n_18453),
.A2(n_8944),
.B1(n_9072),
.B2(n_9024),
.Y(n_18739)
);

INVx2_ASAP7_75t_L g18740 ( 
.A(n_18630),
.Y(n_18740)
);

OAI22xp33_ASAP7_75t_L g18741 ( 
.A1(n_18477),
.A2(n_9072),
.B1(n_9134),
.B2(n_9024),
.Y(n_18741)
);

O2A1O1Ixp5_ASAP7_75t_L g18742 ( 
.A1(n_18547),
.A2(n_8852),
.B(n_8332),
.C(n_8952),
.Y(n_18742)
);

AND2x2_ASAP7_75t_L g18743 ( 
.A(n_18623),
.B(n_8299),
.Y(n_18743)
);

NAND2x1p5_ASAP7_75t_L g18744 ( 
.A(n_18450),
.B(n_5382),
.Y(n_18744)
);

XNOR2x2_ASAP7_75t_L g18745 ( 
.A(n_18647),
.B(n_8513),
.Y(n_18745)
);

AND2x2_ASAP7_75t_L g18746 ( 
.A(n_18635),
.B(n_8299),
.Y(n_18746)
);

OAI22xp5_ASAP7_75t_L g18747 ( 
.A1(n_18569),
.A2(n_9024),
.B1(n_9134),
.B2(n_9072),
.Y(n_18747)
);

INVx1_ASAP7_75t_L g18748 ( 
.A(n_18639),
.Y(n_18748)
);

INVx2_ASAP7_75t_L g18749 ( 
.A(n_18482),
.Y(n_18749)
);

NAND2xp5_ASAP7_75t_L g18750 ( 
.A(n_18573),
.B(n_8322),
.Y(n_18750)
);

NAND2xp5_ASAP7_75t_L g18751 ( 
.A(n_18577),
.B(n_8048),
.Y(n_18751)
);

INVx1_ASAP7_75t_L g18752 ( 
.A(n_18387),
.Y(n_18752)
);

AOI22xp5_ASAP7_75t_L g18753 ( 
.A1(n_18556),
.A2(n_18558),
.B1(n_18508),
.B2(n_18514),
.Y(n_18753)
);

AND2x2_ASAP7_75t_L g18754 ( 
.A(n_18501),
.B(n_8533),
.Y(n_18754)
);

INVx1_ASAP7_75t_L g18755 ( 
.A(n_18491),
.Y(n_18755)
);

INVx1_ASAP7_75t_L g18756 ( 
.A(n_18452),
.Y(n_18756)
);

INVx1_ASAP7_75t_L g18757 ( 
.A(n_18476),
.Y(n_18757)
);

NAND2x1p5_ASAP7_75t_L g18758 ( 
.A(n_18563),
.B(n_5382),
.Y(n_18758)
);

INVx1_ASAP7_75t_L g18759 ( 
.A(n_18513),
.Y(n_18759)
);

OAI21xp5_ASAP7_75t_L g18760 ( 
.A1(n_18391),
.A2(n_8549),
.B(n_8283),
.Y(n_18760)
);

NOR4xp25_ASAP7_75t_SL g18761 ( 
.A(n_18435),
.B(n_8777),
.C(n_8786),
.D(n_8779),
.Y(n_18761)
);

INVx1_ASAP7_75t_L g18762 ( 
.A(n_18521),
.Y(n_18762)
);

NOR2xp33_ASAP7_75t_SL g18763 ( 
.A(n_18620),
.B(n_18576),
.Y(n_18763)
);

NAND2xp5_ASAP7_75t_L g18764 ( 
.A(n_18522),
.B(n_8048),
.Y(n_18764)
);

OR2x2_ASAP7_75t_L g18765 ( 
.A(n_18535),
.B(n_18512),
.Y(n_18765)
);

AOI22xp5_ASAP7_75t_L g18766 ( 
.A1(n_18554),
.A2(n_7535),
.B1(n_8546),
.B2(n_7101),
.Y(n_18766)
);

NAND2xp5_ASAP7_75t_L g18767 ( 
.A(n_18651),
.B(n_8048),
.Y(n_18767)
);

AOI22xp33_ASAP7_75t_SL g18768 ( 
.A1(n_18571),
.A2(n_7101),
.B1(n_7210),
.B2(n_7020),
.Y(n_18768)
);

INVx1_ASAP7_75t_L g18769 ( 
.A(n_18595),
.Y(n_18769)
);

OR2x2_ASAP7_75t_L g18770 ( 
.A(n_18640),
.B(n_8533),
.Y(n_18770)
);

AOI211xp5_ASAP7_75t_SL g18771 ( 
.A1(n_18638),
.A2(n_7087),
.B(n_7104),
.C(n_7067),
.Y(n_18771)
);

AOI222xp33_ASAP7_75t_L g18772 ( 
.A1(n_18644),
.A2(n_8067),
.B1(n_8052),
.B2(n_8516),
.C1(n_8513),
.C2(n_8301),
.Y(n_18772)
);

OA22x2_ASAP7_75t_L g18773 ( 
.A1(n_18610),
.A2(n_7491),
.B1(n_8433),
.B2(n_8476),
.Y(n_18773)
);

NAND2xp33_ASAP7_75t_SL g18774 ( 
.A(n_18553),
.B(n_7535),
.Y(n_18774)
);

A2O1A1Ixp33_ASAP7_75t_L g18775 ( 
.A1(n_18464),
.A2(n_8324),
.B(n_8433),
.C(n_8476),
.Y(n_18775)
);

NAND2xp5_ASAP7_75t_L g18776 ( 
.A(n_18650),
.B(n_8709),
.Y(n_18776)
);

INVxp33_ASAP7_75t_L g18777 ( 
.A(n_18614),
.Y(n_18777)
);

INVx2_ASAP7_75t_L g18778 ( 
.A(n_18441),
.Y(n_18778)
);

OAI32xp33_ASAP7_75t_L g18779 ( 
.A1(n_18483),
.A2(n_9282),
.A3(n_9287),
.B1(n_9212),
.B2(n_9134),
.Y(n_18779)
);

INVx1_ASAP7_75t_L g18780 ( 
.A(n_18449),
.Y(n_18780)
);

INVx2_ASAP7_75t_L g18781 ( 
.A(n_18465),
.Y(n_18781)
);

NAND3xp33_ASAP7_75t_L g18782 ( 
.A(n_18629),
.B(n_7101),
.C(n_7020),
.Y(n_18782)
);

INVx1_ASAP7_75t_L g18783 ( 
.A(n_18582),
.Y(n_18783)
);

NAND2xp5_ASAP7_75t_L g18784 ( 
.A(n_18492),
.B(n_8709),
.Y(n_18784)
);

INVx1_ASAP7_75t_L g18785 ( 
.A(n_18523),
.Y(n_18785)
);

AND2x4_ASAP7_75t_L g18786 ( 
.A(n_18524),
.B(n_8036),
.Y(n_18786)
);

INVx1_ASAP7_75t_L g18787 ( 
.A(n_18567),
.Y(n_18787)
);

INVx2_ASAP7_75t_SL g18788 ( 
.A(n_18421),
.Y(n_18788)
);

INVx1_ASAP7_75t_L g18789 ( 
.A(n_18612),
.Y(n_18789)
);

AND2x2_ASAP7_75t_L g18790 ( 
.A(n_18619),
.B(n_8533),
.Y(n_18790)
);

AOI221x1_ASAP7_75t_L g18791 ( 
.A1(n_18626),
.A2(n_18632),
.B1(n_18631),
.B2(n_18527),
.C(n_18604),
.Y(n_18791)
);

INVx1_ASAP7_75t_L g18792 ( 
.A(n_18641),
.Y(n_18792)
);

OAI22xp5_ASAP7_75t_L g18793 ( 
.A1(n_18526),
.A2(n_9134),
.B1(n_9282),
.B2(n_9212),
.Y(n_18793)
);

NAND3xp33_ASAP7_75t_L g18794 ( 
.A(n_18599),
.B(n_18581),
.C(n_18597),
.Y(n_18794)
);

INVx1_ASAP7_75t_L g18795 ( 
.A(n_18466),
.Y(n_18795)
);

NAND2xp5_ASAP7_75t_L g18796 ( 
.A(n_18518),
.B(n_18544),
.Y(n_18796)
);

NOR3xp33_ASAP7_75t_L g18797 ( 
.A(n_18416),
.B(n_5120),
.C(n_5066),
.Y(n_18797)
);

AOI22xp5_ASAP7_75t_L g18798 ( 
.A1(n_18455),
.A2(n_8546),
.B1(n_7101),
.B2(n_7210),
.Y(n_18798)
);

INVx2_ASAP7_75t_L g18799 ( 
.A(n_18484),
.Y(n_18799)
);

INVx2_ASAP7_75t_L g18800 ( 
.A(n_18549),
.Y(n_18800)
);

INVx1_ASAP7_75t_L g18801 ( 
.A(n_18473),
.Y(n_18801)
);

NAND2xp5_ASAP7_75t_SL g18802 ( 
.A(n_18456),
.B(n_18543),
.Y(n_18802)
);

INVx2_ASAP7_75t_L g18803 ( 
.A(n_18557),
.Y(n_18803)
);

INVx1_ASAP7_75t_L g18804 ( 
.A(n_18490),
.Y(n_18804)
);

INVxp67_ASAP7_75t_L g18805 ( 
.A(n_18424),
.Y(n_18805)
);

NOR2x1_ASAP7_75t_SL g18806 ( 
.A(n_18437),
.B(n_5751),
.Y(n_18806)
);

INVx2_ASAP7_75t_L g18807 ( 
.A(n_18628),
.Y(n_18807)
);

HB1xp67_ASAP7_75t_L g18808 ( 
.A(n_18457),
.Y(n_18808)
);

AND2x2_ASAP7_75t_L g18809 ( 
.A(n_18520),
.B(n_8533),
.Y(n_18809)
);

NAND2xp5_ASAP7_75t_L g18810 ( 
.A(n_18487),
.B(n_18525),
.Y(n_18810)
);

OAI21xp5_ASAP7_75t_SL g18811 ( 
.A1(n_18493),
.A2(n_9212),
.B(n_9134),
.Y(n_18811)
);

AOI22xp5_ASAP7_75t_L g18812 ( 
.A1(n_18517),
.A2(n_7101),
.B1(n_7210),
.B2(n_7020),
.Y(n_18812)
);

INVx1_ASAP7_75t_L g18813 ( 
.A(n_18498),
.Y(n_18813)
);

AND2x2_ASAP7_75t_L g18814 ( 
.A(n_18642),
.B(n_8533),
.Y(n_18814)
);

NAND2xp5_ASAP7_75t_SL g18815 ( 
.A(n_18618),
.B(n_7101),
.Y(n_18815)
);

NAND2xp5_ASAP7_75t_SL g18816 ( 
.A(n_18636),
.B(n_7210),
.Y(n_18816)
);

AOI21xp5_ASAP7_75t_L g18817 ( 
.A1(n_18458),
.A2(n_8245),
.B(n_8235),
.Y(n_18817)
);

AOI22xp33_ASAP7_75t_SL g18818 ( 
.A1(n_18592),
.A2(n_7218),
.B1(n_7345),
.B2(n_7210),
.Y(n_18818)
);

INVx2_ASAP7_75t_L g18819 ( 
.A(n_18590),
.Y(n_18819)
);

OAI22xp33_ASAP7_75t_L g18820 ( 
.A1(n_18446),
.A2(n_9282),
.B1(n_9287),
.B2(n_9212),
.Y(n_18820)
);

INVx1_ASAP7_75t_L g18821 ( 
.A(n_18509),
.Y(n_18821)
);

AOI21xp5_ASAP7_75t_L g18822 ( 
.A1(n_18536),
.A2(n_8245),
.B(n_8235),
.Y(n_18822)
);

AOI22xp5_ASAP7_75t_L g18823 ( 
.A1(n_18434),
.A2(n_18570),
.B1(n_18430),
.B2(n_18584),
.Y(n_18823)
);

OR2x2_ASAP7_75t_L g18824 ( 
.A(n_18625),
.B(n_8533),
.Y(n_18824)
);

AOI21xp5_ASAP7_75t_L g18825 ( 
.A1(n_18622),
.A2(n_8732),
.B(n_8709),
.Y(n_18825)
);

OAI32xp33_ASAP7_75t_L g18826 ( 
.A1(n_18627),
.A2(n_18634),
.A3(n_18633),
.B1(n_18617),
.B2(n_18600),
.Y(n_18826)
);

OAI21xp5_ASAP7_75t_L g18827 ( 
.A1(n_18598),
.A2(n_18425),
.B(n_18603),
.Y(n_18827)
);

INVx2_ASAP7_75t_L g18828 ( 
.A(n_18451),
.Y(n_18828)
);

AOI22xp5_ASAP7_75t_L g18829 ( 
.A1(n_18591),
.A2(n_7218),
.B1(n_7345),
.B2(n_7210),
.Y(n_18829)
);

INVx2_ASAP7_75t_L g18830 ( 
.A(n_18643),
.Y(n_18830)
);

INVx2_ASAP7_75t_SL g18831 ( 
.A(n_18606),
.Y(n_18831)
);

INVx1_ASAP7_75t_L g18832 ( 
.A(n_18653),
.Y(n_18832)
);

AOI21xp33_ASAP7_75t_SL g18833 ( 
.A1(n_18481),
.A2(n_18500),
.B(n_18428),
.Y(n_18833)
);

INVxp67_ASAP7_75t_L g18834 ( 
.A(n_18594),
.Y(n_18834)
);

INVx1_ASAP7_75t_L g18835 ( 
.A(n_18579),
.Y(n_18835)
);

AOI21xp5_ASAP7_75t_L g18836 ( 
.A1(n_18572),
.A2(n_18467),
.B(n_18528),
.Y(n_18836)
);

INVx1_ASAP7_75t_L g18837 ( 
.A(n_18646),
.Y(n_18837)
);

INVx1_ASAP7_75t_L g18838 ( 
.A(n_18469),
.Y(n_18838)
);

OR2x2_ASAP7_75t_L g18839 ( 
.A(n_18515),
.B(n_8533),
.Y(n_18839)
);

AND2x2_ASAP7_75t_L g18840 ( 
.A(n_18652),
.B(n_8533),
.Y(n_18840)
);

NAND2xp5_ASAP7_75t_L g18841 ( 
.A(n_18637),
.B(n_8709),
.Y(n_18841)
);

INVx1_ASAP7_75t_SL g18842 ( 
.A(n_18565),
.Y(n_18842)
);

INVx1_ASAP7_75t_L g18843 ( 
.A(n_18459),
.Y(n_18843)
);

NOR2xp33_ASAP7_75t_L g18844 ( 
.A(n_18531),
.B(n_9053),
.Y(n_18844)
);

OAI22xp33_ASAP7_75t_SL g18845 ( 
.A1(n_18648),
.A2(n_9282),
.B1(n_9287),
.B2(n_9212),
.Y(n_18845)
);

OAI21xp5_ASAP7_75t_L g18846 ( 
.A1(n_18507),
.A2(n_8283),
.B(n_8303),
.Y(n_18846)
);

AND2x2_ASAP7_75t_L g18847 ( 
.A(n_18495),
.B(n_8533),
.Y(n_18847)
);

OAI21x1_ASAP7_75t_L g18848 ( 
.A1(n_18583),
.A2(n_8332),
.B(n_8952),
.Y(n_18848)
);

NAND2xp5_ASAP7_75t_L g18849 ( 
.A(n_18497),
.B(n_8709),
.Y(n_18849)
);

INVxp67_ASAP7_75t_L g18850 ( 
.A(n_18624),
.Y(n_18850)
);

INVx1_ASAP7_75t_L g18851 ( 
.A(n_18474),
.Y(n_18851)
);

AND2x2_ASAP7_75t_L g18852 ( 
.A(n_18588),
.B(n_18649),
.Y(n_18852)
);

OAI22xp5_ASAP7_75t_L g18853 ( 
.A1(n_18454),
.A2(n_9282),
.B1(n_9287),
.B2(n_9130),
.Y(n_18853)
);

INVx1_ASAP7_75t_L g18854 ( 
.A(n_18564),
.Y(n_18854)
);

AOI221xp5_ASAP7_75t_L g18855 ( 
.A1(n_18499),
.A2(n_8440),
.B1(n_8431),
.B2(n_7104),
.C(n_7144),
.Y(n_18855)
);

OAI32xp33_ASAP7_75t_L g18856 ( 
.A1(n_18587),
.A2(n_9287),
.A3(n_7494),
.B1(n_7528),
.B2(n_7440),
.Y(n_18856)
);

NOR3xp33_ASAP7_75t_L g18857 ( 
.A(n_18529),
.B(n_5120),
.C(n_5066),
.Y(n_18857)
);

NAND2xp5_ASAP7_75t_L g18858 ( 
.A(n_18494),
.B(n_8732),
.Y(n_18858)
);

XNOR2xp5_ASAP7_75t_L g18859 ( 
.A(n_18601),
.B(n_8283),
.Y(n_18859)
);

OR2x2_ASAP7_75t_L g18860 ( 
.A(n_18649),
.B(n_8545),
.Y(n_18860)
);

OAI22xp5_ASAP7_75t_L g18861 ( 
.A1(n_18611),
.A2(n_9296),
.B1(n_9130),
.B2(n_7857),
.Y(n_18861)
);

AND2x2_ASAP7_75t_L g18862 ( 
.A(n_18555),
.B(n_8545),
.Y(n_18862)
);

AOI322xp5_ASAP7_75t_L g18863 ( 
.A1(n_18575),
.A2(n_7254),
.A3(n_7234),
.B1(n_7307),
.B2(n_7356),
.C1(n_7339),
.C2(n_7220),
.Y(n_18863)
);

AOI21xp33_ASAP7_75t_SL g18864 ( 
.A1(n_18561),
.A2(n_5499),
.B(n_5426),
.Y(n_18864)
);

INVx1_ASAP7_75t_L g18865 ( 
.A(n_18479),
.Y(n_18865)
);

HB1xp67_ASAP7_75t_L g18866 ( 
.A(n_18426),
.Y(n_18866)
);

NAND2xp5_ASAP7_75t_L g18867 ( 
.A(n_18550),
.B(n_8732),
.Y(n_18867)
);

NAND3xp33_ASAP7_75t_L g18868 ( 
.A(n_18519),
.B(n_7218),
.C(n_7210),
.Y(n_18868)
);

NAND2xp5_ASAP7_75t_L g18869 ( 
.A(n_18607),
.B(n_8732),
.Y(n_18869)
);

AOI222xp33_ASAP7_75t_L g18870 ( 
.A1(n_18602),
.A2(n_8513),
.B1(n_8516),
.B2(n_8301),
.C1(n_8403),
.C2(n_8399),
.Y(n_18870)
);

OAI21xp33_ASAP7_75t_L g18871 ( 
.A1(n_18586),
.A2(n_9296),
.B(n_9130),
.Y(n_18871)
);

NAND2xp5_ASAP7_75t_L g18872 ( 
.A(n_18613),
.B(n_8732),
.Y(n_18872)
);

NAND2xp5_ASAP7_75t_L g18873 ( 
.A(n_18538),
.B(n_8748),
.Y(n_18873)
);

INVx1_ASAP7_75t_L g18874 ( 
.A(n_18546),
.Y(n_18874)
);

INVx3_ASAP7_75t_L g18875 ( 
.A(n_18420),
.Y(n_18875)
);

AND2x4_ASAP7_75t_L g18876 ( 
.A(n_18645),
.B(n_8036),
.Y(n_18876)
);

NAND2xp5_ASAP7_75t_L g18877 ( 
.A(n_18447),
.B(n_8748),
.Y(n_18877)
);

NAND2xp5_ASAP7_75t_L g18878 ( 
.A(n_18516),
.B(n_8748),
.Y(n_18878)
);

INVx1_ASAP7_75t_L g18879 ( 
.A(n_18534),
.Y(n_18879)
);

OAI22xp5_ASAP7_75t_L g18880 ( 
.A1(n_18566),
.A2(n_9296),
.B1(n_7857),
.B2(n_7867),
.Y(n_18880)
);

INVx1_ASAP7_75t_L g18881 ( 
.A(n_18432),
.Y(n_18881)
);

INVx1_ASAP7_75t_L g18882 ( 
.A(n_18596),
.Y(n_18882)
);

NAND2xp5_ASAP7_75t_L g18883 ( 
.A(n_18608),
.B(n_8748),
.Y(n_18883)
);

NAND2xp5_ASAP7_75t_L g18884 ( 
.A(n_18445),
.B(n_8748),
.Y(n_18884)
);

NAND2xp5_ASAP7_75t_L g18885 ( 
.A(n_18574),
.B(n_8431),
.Y(n_18885)
);

INVx1_ASAP7_75t_L g18886 ( 
.A(n_18472),
.Y(n_18886)
);

HB1xp67_ASAP7_75t_L g18887 ( 
.A(n_18420),
.Y(n_18887)
);

NAND2xp5_ASAP7_75t_L g18888 ( 
.A(n_18496),
.B(n_8431),
.Y(n_18888)
);

NAND2x1p5_ASAP7_75t_L g18889 ( 
.A(n_18593),
.B(n_5382),
.Y(n_18889)
);

NAND2xp5_ASAP7_75t_SL g18890 ( 
.A(n_18568),
.B(n_7218),
.Y(n_18890)
);

NAND2xp5_ASAP7_75t_L g18891 ( 
.A(n_18578),
.B(n_8431),
.Y(n_18891)
);

INVx1_ASAP7_75t_L g18892 ( 
.A(n_18609),
.Y(n_18892)
);

OAI21xp33_ASAP7_75t_L g18893 ( 
.A1(n_18615),
.A2(n_18551),
.B(n_18486),
.Y(n_18893)
);

INVx1_ASAP7_75t_L g18894 ( 
.A(n_18605),
.Y(n_18894)
);

INVx1_ASAP7_75t_L g18895 ( 
.A(n_18593),
.Y(n_18895)
);

AOI21xp33_ASAP7_75t_L g18896 ( 
.A1(n_18589),
.A2(n_8036),
.B(n_8440),
.Y(n_18896)
);

OAI221xp5_ASAP7_75t_L g18897 ( 
.A1(n_18427),
.A2(n_8379),
.B1(n_8253),
.B2(n_7494),
.C(n_7528),
.Y(n_18897)
);

AOI221xp5_ASAP7_75t_L g18898 ( 
.A1(n_18407),
.A2(n_8440),
.B1(n_7144),
.B2(n_7149),
.C(n_7087),
.Y(n_18898)
);

NAND2xp5_ASAP7_75t_L g18899 ( 
.A(n_18371),
.B(n_8440),
.Y(n_18899)
);

NOR2xp33_ASAP7_75t_L g18900 ( 
.A(n_18371),
.B(n_9053),
.Y(n_18900)
);

NAND2xp5_ASAP7_75t_SL g18901 ( 
.A(n_18372),
.B(n_7218),
.Y(n_18901)
);

OAI21xp33_ASAP7_75t_L g18902 ( 
.A1(n_18371),
.A2(n_6838),
.B(n_7436),
.Y(n_18902)
);

OAI322xp33_ASAP7_75t_L g18903 ( 
.A1(n_18439),
.A2(n_7967),
.A3(n_7930),
.B1(n_7978),
.B2(n_8010),
.C1(n_7953),
.C2(n_7917),
.Y(n_18903)
);

INVx1_ASAP7_75t_L g18904 ( 
.A(n_18372),
.Y(n_18904)
);

INVx1_ASAP7_75t_SL g18905 ( 
.A(n_18372),
.Y(n_18905)
);

AOI21xp5_ASAP7_75t_L g18906 ( 
.A1(n_18380),
.A2(n_8516),
.B(n_8513),
.Y(n_18906)
);

OAI22xp5_ASAP7_75t_L g18907 ( 
.A1(n_18369),
.A2(n_7857),
.B1(n_7867),
.B2(n_7795),
.Y(n_18907)
);

OAI22xp5_ASAP7_75t_L g18908 ( 
.A1(n_18369),
.A2(n_7857),
.B1(n_7867),
.B2(n_7795),
.Y(n_18908)
);

INVx1_ASAP7_75t_L g18909 ( 
.A(n_18372),
.Y(n_18909)
);

NOR2xp33_ASAP7_75t_L g18910 ( 
.A(n_18371),
.B(n_7720),
.Y(n_18910)
);

INVx1_ASAP7_75t_L g18911 ( 
.A(n_18694),
.Y(n_18911)
);

NAND2xp5_ASAP7_75t_L g18912 ( 
.A(n_18694),
.B(n_8383),
.Y(n_18912)
);

INVx1_ASAP7_75t_L g18913 ( 
.A(n_18676),
.Y(n_18913)
);

AOI22xp33_ASAP7_75t_L g18914 ( 
.A1(n_18675),
.A2(n_18667),
.B1(n_18769),
.B2(n_18692),
.Y(n_18914)
);

NAND2xp5_ASAP7_75t_L g18915 ( 
.A(n_18655),
.B(n_8383),
.Y(n_18915)
);

AOI22xp33_ASAP7_75t_L g18916 ( 
.A1(n_18904),
.A2(n_7345),
.B1(n_7353),
.B2(n_7218),
.Y(n_18916)
);

AND3x1_ASAP7_75t_L g18917 ( 
.A(n_18763),
.B(n_7831),
.C(n_7812),
.Y(n_18917)
);

INVx1_ASAP7_75t_L g18918 ( 
.A(n_18887),
.Y(n_18918)
);

NAND2xp5_ASAP7_75t_L g18919 ( 
.A(n_18905),
.B(n_18668),
.Y(n_18919)
);

OAI21xp33_ASAP7_75t_L g18920 ( 
.A1(n_18690),
.A2(n_6838),
.B(n_7436),
.Y(n_18920)
);

NAND2xp5_ASAP7_75t_L g18921 ( 
.A(n_18664),
.B(n_8383),
.Y(n_18921)
);

AND2x2_ASAP7_75t_L g18922 ( 
.A(n_18909),
.B(n_8545),
.Y(n_18922)
);

NAND2xp5_ASAP7_75t_L g18923 ( 
.A(n_18748),
.B(n_8399),
.Y(n_18923)
);

INVx1_ASAP7_75t_L g18924 ( 
.A(n_18662),
.Y(n_18924)
);

INVxp67_ASAP7_75t_L g18925 ( 
.A(n_18900),
.Y(n_18925)
);

OR2x2_ASAP7_75t_L g18926 ( 
.A(n_18658),
.B(n_8545),
.Y(n_18926)
);

AND2x2_ASAP7_75t_L g18927 ( 
.A(n_18657),
.B(n_8545),
.Y(n_18927)
);

INVx1_ASAP7_75t_L g18928 ( 
.A(n_18875),
.Y(n_18928)
);

INVx2_ASAP7_75t_L g18929 ( 
.A(n_18875),
.Y(n_18929)
);

NOR2xp33_ASAP7_75t_L g18930 ( 
.A(n_18665),
.B(n_7720),
.Y(n_18930)
);

NAND2xp5_ASAP7_75t_L g18931 ( 
.A(n_18713),
.B(n_8399),
.Y(n_18931)
);

INVx1_ASAP7_75t_SL g18932 ( 
.A(n_18765),
.Y(n_18932)
);

NOR2xp33_ASAP7_75t_L g18933 ( 
.A(n_18695),
.B(n_7720),
.Y(n_18933)
);

INVx1_ASAP7_75t_L g18934 ( 
.A(n_18703),
.Y(n_18934)
);

HB1xp67_ASAP7_75t_L g18935 ( 
.A(n_18785),
.Y(n_18935)
);

INVx1_ASAP7_75t_L g18936 ( 
.A(n_18654),
.Y(n_18936)
);

AND2x2_ASAP7_75t_L g18937 ( 
.A(n_18698),
.B(n_8545),
.Y(n_18937)
);

INVx1_ASAP7_75t_L g18938 ( 
.A(n_18705),
.Y(n_18938)
);

NAND2xp5_ASAP7_75t_L g18939 ( 
.A(n_18726),
.B(n_8403),
.Y(n_18939)
);

INVx1_ASAP7_75t_L g18940 ( 
.A(n_18707),
.Y(n_18940)
);

INVx1_ASAP7_75t_L g18941 ( 
.A(n_18710),
.Y(n_18941)
);

INVx1_ASAP7_75t_L g18942 ( 
.A(n_18717),
.Y(n_18942)
);

INVx1_ASAP7_75t_L g18943 ( 
.A(n_18719),
.Y(n_18943)
);

NAND2xp5_ASAP7_75t_L g18944 ( 
.A(n_18910),
.B(n_8403),
.Y(n_18944)
);

INVx1_ASAP7_75t_L g18945 ( 
.A(n_18810),
.Y(n_18945)
);

NAND2xp5_ASAP7_75t_L g18946 ( 
.A(n_18730),
.B(n_8084),
.Y(n_18946)
);

NAND2xp5_ASAP7_75t_L g18947 ( 
.A(n_18740),
.B(n_8084),
.Y(n_18947)
);

NAND2xp5_ASAP7_75t_L g18948 ( 
.A(n_18788),
.B(n_8084),
.Y(n_18948)
);

INVx2_ASAP7_75t_L g18949 ( 
.A(n_18696),
.Y(n_18949)
);

AND2x2_ASAP7_75t_L g18950 ( 
.A(n_18716),
.B(n_8545),
.Y(n_18950)
);

NAND2xp5_ASAP7_75t_L g18951 ( 
.A(n_18792),
.B(n_18687),
.Y(n_18951)
);

AND2x2_ASAP7_75t_L g18952 ( 
.A(n_18693),
.B(n_8545),
.Y(n_18952)
);

OR2x2_ASAP7_75t_L g18953 ( 
.A(n_18700),
.B(n_8545),
.Y(n_18953)
);

NAND2xp5_ASAP7_75t_L g18954 ( 
.A(n_18709),
.B(n_8084),
.Y(n_18954)
);

INVx1_ASAP7_75t_L g18955 ( 
.A(n_18866),
.Y(n_18955)
);

NOR2xp33_ASAP7_75t_L g18956 ( 
.A(n_18777),
.B(n_7720),
.Y(n_18956)
);

INVx1_ASAP7_75t_L g18957 ( 
.A(n_18659),
.Y(n_18957)
);

NAND2xp5_ASAP7_75t_L g18958 ( 
.A(n_18673),
.B(n_8084),
.Y(n_18958)
);

NAND2xp5_ASAP7_75t_L g18959 ( 
.A(n_18729),
.B(n_7917),
.Y(n_18959)
);

INVx1_ASAP7_75t_L g18960 ( 
.A(n_18697),
.Y(n_18960)
);

AOI22xp33_ASAP7_75t_L g18961 ( 
.A1(n_18708),
.A2(n_7345),
.B1(n_7353),
.B2(n_7218),
.Y(n_18961)
);

INVx1_ASAP7_75t_SL g18962 ( 
.A(n_18774),
.Y(n_18962)
);

NAND2xp5_ASAP7_75t_L g18963 ( 
.A(n_18755),
.B(n_7917),
.Y(n_18963)
);

NOR2xp33_ASAP7_75t_L g18964 ( 
.A(n_18714),
.B(n_7720),
.Y(n_18964)
);

INVx1_ASAP7_75t_L g18965 ( 
.A(n_18756),
.Y(n_18965)
);

INVx1_ASAP7_75t_SL g18966 ( 
.A(n_18757),
.Y(n_18966)
);

INVx1_ASAP7_75t_L g18967 ( 
.A(n_18759),
.Y(n_18967)
);

INVx2_ASAP7_75t_L g18968 ( 
.A(n_18758),
.Y(n_18968)
);

AND2x2_ASAP7_75t_L g18969 ( 
.A(n_18749),
.B(n_8629),
.Y(n_18969)
);

AND2x2_ASAP7_75t_L g18970 ( 
.A(n_18680),
.B(n_8629),
.Y(n_18970)
);

NAND2xp5_ASAP7_75t_L g18971 ( 
.A(n_18762),
.B(n_7917),
.Y(n_18971)
);

INVx1_ASAP7_75t_L g18972 ( 
.A(n_18789),
.Y(n_18972)
);

HB1xp67_ASAP7_75t_L g18973 ( 
.A(n_18744),
.Y(n_18973)
);

NAND2xp5_ASAP7_75t_L g18974 ( 
.A(n_18778),
.B(n_7930),
.Y(n_18974)
);

INVx1_ASAP7_75t_L g18975 ( 
.A(n_18781),
.Y(n_18975)
);

NOR2xp33_ASAP7_75t_L g18976 ( 
.A(n_18699),
.B(n_7720),
.Y(n_18976)
);

INVx1_ASAP7_75t_L g18977 ( 
.A(n_18828),
.Y(n_18977)
);

HB1xp67_ASAP7_75t_L g18978 ( 
.A(n_18835),
.Y(n_18978)
);

INVx2_ASAP7_75t_L g18979 ( 
.A(n_18889),
.Y(n_18979)
);

AND2x2_ASAP7_75t_L g18980 ( 
.A(n_18727),
.B(n_8629),
.Y(n_18980)
);

NAND2xp5_ASAP7_75t_L g18981 ( 
.A(n_18669),
.B(n_7930),
.Y(n_18981)
);

INVx1_ASAP7_75t_L g18982 ( 
.A(n_18852),
.Y(n_18982)
);

NAND2xp5_ASAP7_75t_SL g18983 ( 
.A(n_18660),
.B(n_18704),
.Y(n_18983)
);

NAND2xp5_ASAP7_75t_L g18984 ( 
.A(n_18663),
.B(n_18838),
.Y(n_18984)
);

OR2x2_ASAP7_75t_L g18985 ( 
.A(n_18807),
.B(n_8629),
.Y(n_18985)
);

INVxp67_ASAP7_75t_L g18986 ( 
.A(n_18808),
.Y(n_18986)
);

INVx1_ASAP7_75t_L g18987 ( 
.A(n_18711),
.Y(n_18987)
);

NOR2xp33_ASAP7_75t_L g18988 ( 
.A(n_18661),
.B(n_7747),
.Y(n_18988)
);

NAND2xp5_ASAP7_75t_L g18989 ( 
.A(n_18819),
.B(n_7953),
.Y(n_18989)
);

NAND2xp5_ASAP7_75t_L g18990 ( 
.A(n_18801),
.B(n_7953),
.Y(n_18990)
);

INVx1_ASAP7_75t_L g18991 ( 
.A(n_18671),
.Y(n_18991)
);

CKINVDCx16_ASAP7_75t_R g18992 ( 
.A(n_18753),
.Y(n_18992)
);

NOR2xp33_ASAP7_75t_L g18993 ( 
.A(n_18689),
.B(n_7747),
.Y(n_18993)
);

NAND2xp5_ASAP7_75t_L g18994 ( 
.A(n_18804),
.B(n_7967),
.Y(n_18994)
);

INVx2_ASAP7_75t_L g18995 ( 
.A(n_18770),
.Y(n_18995)
);

NAND2x1_ASAP7_75t_L g18996 ( 
.A(n_18799),
.B(n_8572),
.Y(n_18996)
);

INVx1_ASAP7_75t_L g18997 ( 
.A(n_18666),
.Y(n_18997)
);

AND2x2_ASAP7_75t_L g18998 ( 
.A(n_18787),
.B(n_8629),
.Y(n_18998)
);

NOR2x1_ASAP7_75t_L g18999 ( 
.A(n_18794),
.B(n_8320),
.Y(n_18999)
);

NAND2xp5_ASAP7_75t_L g19000 ( 
.A(n_18842),
.B(n_7967),
.Y(n_19000)
);

AND2x2_ASAP7_75t_L g19001 ( 
.A(n_18752),
.B(n_8629),
.Y(n_19001)
);

HB1xp67_ASAP7_75t_L g19002 ( 
.A(n_18712),
.Y(n_19002)
);

AND2x2_ASAP7_75t_L g19003 ( 
.A(n_18723),
.B(n_8629),
.Y(n_19003)
);

NAND2xp5_ASAP7_75t_L g19004 ( 
.A(n_18790),
.B(n_18881),
.Y(n_19004)
);

NAND2xp5_ASAP7_75t_SL g19005 ( 
.A(n_18686),
.B(n_18733),
.Y(n_19005)
);

AOI22xp33_ASAP7_75t_L g19006 ( 
.A1(n_18844),
.A2(n_7345),
.B1(n_7353),
.B2(n_7218),
.Y(n_19006)
);

INVxp67_ASAP7_75t_SL g19007 ( 
.A(n_18679),
.Y(n_19007)
);

OAI21xp5_ASAP7_75t_SL g19008 ( 
.A1(n_18850),
.A2(n_18735),
.B(n_18791),
.Y(n_19008)
);

BUFx2_ASAP7_75t_L g19009 ( 
.A(n_18732),
.Y(n_19009)
);

AND2x2_ASAP7_75t_L g19010 ( 
.A(n_18754),
.B(n_8629),
.Y(n_19010)
);

INVx1_ASAP7_75t_L g19011 ( 
.A(n_18895),
.Y(n_19011)
);

NAND2xp5_ASAP7_75t_L g19012 ( 
.A(n_18886),
.B(n_18672),
.Y(n_19012)
);

NAND2xp5_ASAP7_75t_L g19013 ( 
.A(n_18780),
.B(n_7967),
.Y(n_19013)
);

NAND2xp5_ASAP7_75t_L g19014 ( 
.A(n_18783),
.B(n_7978),
.Y(n_19014)
);

AND2x2_ASAP7_75t_L g19015 ( 
.A(n_18725),
.B(n_8629),
.Y(n_19015)
);

AOI22xp33_ASAP7_75t_L g19016 ( 
.A1(n_18840),
.A2(n_7345),
.B1(n_7353),
.B2(n_7218),
.Y(n_19016)
);

AOI222xp33_ASAP7_75t_L g19017 ( 
.A1(n_18802),
.A2(n_8516),
.B1(n_8324),
.B2(n_8301),
.C1(n_8205),
.C2(n_8209),
.Y(n_19017)
);

OR2x2_ASAP7_75t_L g19018 ( 
.A(n_18901),
.B(n_8751),
.Y(n_19018)
);

AND2x2_ASAP7_75t_L g19019 ( 
.A(n_18743),
.B(n_8751),
.Y(n_19019)
);

OR2x2_ASAP7_75t_L g19020 ( 
.A(n_18670),
.B(n_8751),
.Y(n_19020)
);

NAND2xp5_ASAP7_75t_L g19021 ( 
.A(n_18843),
.B(n_7978),
.Y(n_19021)
);

AND2x2_ASAP7_75t_L g19022 ( 
.A(n_18746),
.B(n_8751),
.Y(n_19022)
);

NOR2x1p5_ASAP7_75t_L g19023 ( 
.A(n_18796),
.B(n_5751),
.Y(n_19023)
);

AOI22xp33_ASAP7_75t_L g19024 ( 
.A1(n_18731),
.A2(n_7345),
.B1(n_7353),
.B2(n_7218),
.Y(n_19024)
);

AND2x2_ASAP7_75t_L g19025 ( 
.A(n_18702),
.B(n_8751),
.Y(n_19025)
);

INVx1_ASAP7_75t_L g19026 ( 
.A(n_18865),
.Y(n_19026)
);

AND2x2_ASAP7_75t_L g19027 ( 
.A(n_18724),
.B(n_8751),
.Y(n_19027)
);

AOI22xp5_ASAP7_75t_L g19028 ( 
.A1(n_18907),
.A2(n_18908),
.B1(n_18902),
.B2(n_18893),
.Y(n_19028)
);

OAI22xp5_ASAP7_75t_L g19029 ( 
.A1(n_18818),
.A2(n_7149),
.B1(n_7067),
.B2(n_7795),
.Y(n_19029)
);

OAI222xp33_ASAP7_75t_L g19030 ( 
.A1(n_18823),
.A2(n_8253),
.B1(n_8379),
.B2(n_9025),
.C1(n_9087),
.C2(n_9069),
.Y(n_19030)
);

OR2x2_ASAP7_75t_L g19031 ( 
.A(n_18734),
.B(n_8751),
.Y(n_19031)
);

INVx1_ASAP7_75t_L g19032 ( 
.A(n_18795),
.Y(n_19032)
);

NAND2x1p5_ASAP7_75t_L g19033 ( 
.A(n_18851),
.B(n_5382),
.Y(n_19033)
);

INVx1_ASAP7_75t_L g19034 ( 
.A(n_18874),
.Y(n_19034)
);

INVxp67_ASAP7_75t_L g19035 ( 
.A(n_18899),
.Y(n_19035)
);

INVx1_ASAP7_75t_SL g19036 ( 
.A(n_18813),
.Y(n_19036)
);

NAND2x1_ASAP7_75t_L g19037 ( 
.A(n_18837),
.B(n_8572),
.Y(n_19037)
);

INVx2_ASAP7_75t_L g19038 ( 
.A(n_18860),
.Y(n_19038)
);

INVx1_ASAP7_75t_SL g19039 ( 
.A(n_18821),
.Y(n_19039)
);

NOR2xp33_ASAP7_75t_L g19040 ( 
.A(n_18833),
.B(n_7747),
.Y(n_19040)
);

INVx1_ASAP7_75t_L g19041 ( 
.A(n_18879),
.Y(n_19041)
);

NAND2xp5_ASAP7_75t_L g19042 ( 
.A(n_18656),
.B(n_7978),
.Y(n_19042)
);

HB1xp67_ASAP7_75t_L g19043 ( 
.A(n_18834),
.Y(n_19043)
);

INVx2_ASAP7_75t_L g19044 ( 
.A(n_18814),
.Y(n_19044)
);

INVx1_ASAP7_75t_L g19045 ( 
.A(n_18800),
.Y(n_19045)
);

INVx1_ASAP7_75t_L g19046 ( 
.A(n_18830),
.Y(n_19046)
);

INVx1_ASAP7_75t_SL g19047 ( 
.A(n_18832),
.Y(n_19047)
);

NAND2xp5_ASAP7_75t_L g19048 ( 
.A(n_18806),
.B(n_8010),
.Y(n_19048)
);

INVx1_ASAP7_75t_L g19049 ( 
.A(n_18894),
.Y(n_19049)
);

NOR2x1_ASAP7_75t_L g19050 ( 
.A(n_18892),
.B(n_8320),
.Y(n_19050)
);

INVx1_ASAP7_75t_L g19051 ( 
.A(n_18803),
.Y(n_19051)
);

INVx1_ASAP7_75t_L g19052 ( 
.A(n_18854),
.Y(n_19052)
);

INVx1_ASAP7_75t_L g19053 ( 
.A(n_18882),
.Y(n_19053)
);

OR2x2_ASAP7_75t_L g19054 ( 
.A(n_18839),
.B(n_18682),
.Y(n_19054)
);

AOI22xp33_ASAP7_75t_L g19055 ( 
.A1(n_18871),
.A2(n_7353),
.B1(n_7355),
.B2(n_7345),
.Y(n_19055)
);

INVx1_ASAP7_75t_L g19056 ( 
.A(n_18805),
.Y(n_19056)
);

AND2x2_ASAP7_75t_L g19057 ( 
.A(n_18809),
.B(n_8751),
.Y(n_19057)
);

INVx2_ASAP7_75t_L g19058 ( 
.A(n_18824),
.Y(n_19058)
);

OR2x2_ASAP7_75t_L g19059 ( 
.A(n_18841),
.B(n_8751),
.Y(n_19059)
);

INVx2_ASAP7_75t_L g19060 ( 
.A(n_18862),
.Y(n_19060)
);

NAND2xp5_ASAP7_75t_SL g19061 ( 
.A(n_18768),
.B(n_18864),
.Y(n_19061)
);

INVx1_ASAP7_75t_L g19062 ( 
.A(n_18831),
.Y(n_19062)
);

AND2x2_ASAP7_75t_L g19063 ( 
.A(n_18771),
.B(n_8805),
.Y(n_19063)
);

NAND2xp5_ASAP7_75t_L g19064 ( 
.A(n_18816),
.B(n_8010),
.Y(n_19064)
);

AOI22xp5_ASAP7_75t_L g19065 ( 
.A1(n_18782),
.A2(n_7353),
.B1(n_7355),
.B2(n_7345),
.Y(n_19065)
);

NAND2xp5_ASAP7_75t_L g19066 ( 
.A(n_18683),
.B(n_8010),
.Y(n_19066)
);

NOR2xp67_ASAP7_75t_L g19067 ( 
.A(n_18836),
.B(n_9025),
.Y(n_19067)
);

INVx1_ASAP7_75t_SL g19068 ( 
.A(n_18751),
.Y(n_19068)
);

INVx1_ASAP7_75t_L g19069 ( 
.A(n_18827),
.Y(n_19069)
);

INVx1_ASAP7_75t_L g19070 ( 
.A(n_18826),
.Y(n_19070)
);

INVx1_ASAP7_75t_L g19071 ( 
.A(n_18685),
.Y(n_19071)
);

HB1xp67_ASAP7_75t_L g19072 ( 
.A(n_18764),
.Y(n_19072)
);

INVx1_ASAP7_75t_SL g19073 ( 
.A(n_18784),
.Y(n_19073)
);

INVx1_ASAP7_75t_L g19074 ( 
.A(n_18815),
.Y(n_19074)
);

NAND2xp5_ASAP7_75t_L g19075 ( 
.A(n_18797),
.B(n_8023),
.Y(n_19075)
);

AND2x2_ASAP7_75t_L g19076 ( 
.A(n_18847),
.B(n_8805),
.Y(n_19076)
);

NOR2xp33_ASAP7_75t_L g19077 ( 
.A(n_18890),
.B(n_7747),
.Y(n_19077)
);

NOR2xp33_ASAP7_75t_L g19078 ( 
.A(n_18856),
.B(n_18750),
.Y(n_19078)
);

NAND2xp5_ASAP7_75t_L g19079 ( 
.A(n_18857),
.B(n_8023),
.Y(n_19079)
);

OAI22xp33_ASAP7_75t_L g19080 ( 
.A1(n_18766),
.A2(n_7353),
.B1(n_7355),
.B2(n_7345),
.Y(n_19080)
);

NAND2xp5_ASAP7_75t_L g19081 ( 
.A(n_18684),
.B(n_8023),
.Y(n_19081)
);

INVx2_ASAP7_75t_L g19082 ( 
.A(n_18859),
.Y(n_19082)
);

NAND2xp5_ASAP7_75t_L g19083 ( 
.A(n_18718),
.B(n_8023),
.Y(n_19083)
);

AND2x2_ASAP7_75t_L g19084 ( 
.A(n_18760),
.B(n_8805),
.Y(n_19084)
);

INVx1_ASAP7_75t_L g19085 ( 
.A(n_18776),
.Y(n_19085)
);

NOR2xp33_ASAP7_75t_L g19086 ( 
.A(n_18737),
.B(n_7747),
.Y(n_19086)
);

NAND2xp5_ASAP7_75t_L g19087 ( 
.A(n_18701),
.B(n_8032),
.Y(n_19087)
);

INVxp67_ASAP7_75t_L g19088 ( 
.A(n_18728),
.Y(n_19088)
);

INVx1_ASAP7_75t_L g19089 ( 
.A(n_18877),
.Y(n_19089)
);

NAND2xp5_ASAP7_75t_L g19090 ( 
.A(n_18767),
.B(n_8032),
.Y(n_19090)
);

NOR2xp33_ASAP7_75t_L g19091 ( 
.A(n_18849),
.B(n_7747),
.Y(n_19091)
);

INVx1_ASAP7_75t_L g19092 ( 
.A(n_18858),
.Y(n_19092)
);

INVx1_ASAP7_75t_L g19093 ( 
.A(n_18868),
.Y(n_19093)
);

NAND2xp5_ASAP7_75t_L g19094 ( 
.A(n_18898),
.B(n_8032),
.Y(n_19094)
);

AND2x4_ASAP7_75t_L g19095 ( 
.A(n_18829),
.B(n_8969),
.Y(n_19095)
);

NAND2xp5_ASAP7_75t_L g19096 ( 
.A(n_18811),
.B(n_8032),
.Y(n_19096)
);

INVx2_ASAP7_75t_L g19097 ( 
.A(n_18884),
.Y(n_19097)
);

AOI22xp33_ASAP7_75t_L g19098 ( 
.A1(n_18897),
.A2(n_7355),
.B1(n_7366),
.B2(n_7353),
.Y(n_19098)
);

NAND2xp5_ASAP7_75t_L g19099 ( 
.A(n_18845),
.B(n_8033),
.Y(n_19099)
);

INVx1_ASAP7_75t_SL g19100 ( 
.A(n_18873),
.Y(n_19100)
);

AOI22xp33_ASAP7_75t_SL g19101 ( 
.A1(n_18861),
.A2(n_7355),
.B1(n_7366),
.B2(n_7353),
.Y(n_19101)
);

AND2x2_ASAP7_75t_L g19102 ( 
.A(n_18761),
.B(n_8805),
.Y(n_19102)
);

INVx1_ASAP7_75t_L g19103 ( 
.A(n_18878),
.Y(n_19103)
);

NOR2xp33_ASAP7_75t_L g19104 ( 
.A(n_18880),
.B(n_5499),
.Y(n_19104)
);

AOI22xp33_ASAP7_75t_L g19105 ( 
.A1(n_18876),
.A2(n_7366),
.B1(n_7367),
.B2(n_7355),
.Y(n_19105)
);

INVx1_ASAP7_75t_L g19106 ( 
.A(n_18869),
.Y(n_19106)
);

INVx2_ASAP7_75t_L g19107 ( 
.A(n_18876),
.Y(n_19107)
);

NAND2xp5_ASAP7_75t_L g19108 ( 
.A(n_18863),
.B(n_8033),
.Y(n_19108)
);

INVx1_ASAP7_75t_L g19109 ( 
.A(n_18872),
.Y(n_19109)
);

NAND2xp5_ASAP7_75t_SL g19110 ( 
.A(n_18677),
.B(n_7355),
.Y(n_19110)
);

NAND2xp5_ASAP7_75t_L g19111 ( 
.A(n_18906),
.B(n_8033),
.Y(n_19111)
);

INVx1_ASAP7_75t_L g19112 ( 
.A(n_18867),
.Y(n_19112)
);

OR2x2_ASAP7_75t_L g19113 ( 
.A(n_18885),
.B(n_8805),
.Y(n_19113)
);

NOR2xp33_ASAP7_75t_L g19114 ( 
.A(n_18883),
.B(n_5699),
.Y(n_19114)
);

INVx1_ASAP7_75t_L g19115 ( 
.A(n_18888),
.Y(n_19115)
);

INVx1_ASAP7_75t_SL g19116 ( 
.A(n_18891),
.Y(n_19116)
);

OR2x2_ASAP7_75t_L g19117 ( 
.A(n_18853),
.B(n_8805),
.Y(n_19117)
);

INVx1_ASAP7_75t_L g19118 ( 
.A(n_18745),
.Y(n_19118)
);

INVx2_ASAP7_75t_L g19119 ( 
.A(n_18848),
.Y(n_19119)
);

CKINVDCx16_ASAP7_75t_R g19120 ( 
.A(n_18747),
.Y(n_19120)
);

AND2x4_ASAP7_75t_L g19121 ( 
.A(n_18846),
.B(n_8969),
.Y(n_19121)
);

NAND2xp5_ASAP7_75t_L g19122 ( 
.A(n_18855),
.B(n_8033),
.Y(n_19122)
);

INVx1_ASAP7_75t_L g19123 ( 
.A(n_18721),
.Y(n_19123)
);

NAND2xp33_ASAP7_75t_L g19124 ( 
.A(n_18688),
.B(n_18775),
.Y(n_19124)
);

AOI22xp33_ASAP7_75t_L g19125 ( 
.A1(n_18741),
.A2(n_7366),
.B1(n_7367),
.B2(n_7355),
.Y(n_19125)
);

NAND2xp5_ASAP7_75t_L g19126 ( 
.A(n_18820),
.B(n_8062),
.Y(n_19126)
);

AND2x2_ASAP7_75t_L g19127 ( 
.A(n_18812),
.B(n_8805),
.Y(n_19127)
);

OAI22xp33_ASAP7_75t_L g19128 ( 
.A1(n_18798),
.A2(n_7366),
.B1(n_7367),
.B2(n_7355),
.Y(n_19128)
);

NAND2xp5_ASAP7_75t_L g19129 ( 
.A(n_18817),
.B(n_8062),
.Y(n_19129)
);

NOR2xp67_ASAP7_75t_L g19130 ( 
.A(n_18822),
.B(n_9025),
.Y(n_19130)
);

INVx1_ASAP7_75t_L g19131 ( 
.A(n_18903),
.Y(n_19131)
);

OR2x2_ASAP7_75t_L g19132 ( 
.A(n_18793),
.B(n_8805),
.Y(n_19132)
);

AOI22xp33_ASAP7_75t_L g19133 ( 
.A1(n_18722),
.A2(n_7366),
.B1(n_7367),
.B2(n_7355),
.Y(n_19133)
);

OR2x2_ASAP7_75t_L g19134 ( 
.A(n_18691),
.B(n_8805),
.Y(n_19134)
);

NAND2xp5_ASAP7_75t_L g19135 ( 
.A(n_18736),
.B(n_8062),
.Y(n_19135)
);

AOI22xp33_ASAP7_75t_L g19136 ( 
.A1(n_18773),
.A2(n_7367),
.B1(n_7375),
.B2(n_7366),
.Y(n_19136)
);

NOR2xp33_ASAP7_75t_L g19137 ( 
.A(n_18896),
.B(n_5699),
.Y(n_19137)
);

NAND3xp33_ASAP7_75t_SL g19138 ( 
.A(n_18674),
.B(n_7178),
.C(n_7115),
.Y(n_19138)
);

AND2x2_ASAP7_75t_L g19139 ( 
.A(n_18681),
.B(n_8873),
.Y(n_19139)
);

AND2x2_ASAP7_75t_L g19140 ( 
.A(n_18739),
.B(n_18779),
.Y(n_19140)
);

AOI22xp33_ASAP7_75t_L g19141 ( 
.A1(n_18715),
.A2(n_7367),
.B1(n_7375),
.B2(n_7366),
.Y(n_19141)
);

INVx1_ASAP7_75t_L g19142 ( 
.A(n_18825),
.Y(n_19142)
);

INVx2_ASAP7_75t_L g19143 ( 
.A(n_18742),
.Y(n_19143)
);

NOR2xp33_ASAP7_75t_L g19144 ( 
.A(n_18738),
.B(n_9069),
.Y(n_19144)
);

NOR2xp33_ASAP7_75t_L g19145 ( 
.A(n_18678),
.B(n_9069),
.Y(n_19145)
);

INVx1_ASAP7_75t_L g19146 ( 
.A(n_18720),
.Y(n_19146)
);

AND2x2_ASAP7_75t_L g19147 ( 
.A(n_18786),
.B(n_8873),
.Y(n_19147)
);

NAND2x1_ASAP7_75t_SL g19148 ( 
.A(n_18786),
.B(n_8777),
.Y(n_19148)
);

INVx1_ASAP7_75t_L g19149 ( 
.A(n_18772),
.Y(n_19149)
);

INVx1_ASAP7_75t_L g19150 ( 
.A(n_18870),
.Y(n_19150)
);

AND2x2_ASAP7_75t_L g19151 ( 
.A(n_18706),
.B(n_8873),
.Y(n_19151)
);

NAND2xp5_ASAP7_75t_L g19152 ( 
.A(n_18694),
.B(n_8062),
.Y(n_19152)
);

AOI22xp33_ASAP7_75t_SL g19153 ( 
.A1(n_18694),
.A2(n_7367),
.B1(n_7375),
.B2(n_7366),
.Y(n_19153)
);

NAND2xp5_ASAP7_75t_L g19154 ( 
.A(n_18694),
.B(n_8069),
.Y(n_19154)
);

AOI22xp33_ASAP7_75t_L g19155 ( 
.A1(n_18675),
.A2(n_7367),
.B1(n_7375),
.B2(n_7366),
.Y(n_19155)
);

AND2x2_ASAP7_75t_L g19156 ( 
.A(n_18667),
.B(n_8873),
.Y(n_19156)
);

NAND2xp5_ASAP7_75t_L g19157 ( 
.A(n_18694),
.B(n_8069),
.Y(n_19157)
);

AOI21xp5_ASAP7_75t_L g19158 ( 
.A1(n_18676),
.A2(n_8320),
.B(n_8301),
.Y(n_19158)
);

NAND2xp5_ASAP7_75t_L g19159 ( 
.A(n_18694),
.B(n_8069),
.Y(n_19159)
);

INVx1_ASAP7_75t_L g19160 ( 
.A(n_18694),
.Y(n_19160)
);

INVx2_ASAP7_75t_L g19161 ( 
.A(n_18694),
.Y(n_19161)
);

AND2x2_ASAP7_75t_L g19162 ( 
.A(n_18667),
.B(n_8873),
.Y(n_19162)
);

NOR2xp33_ASAP7_75t_L g19163 ( 
.A(n_18694),
.B(n_9087),
.Y(n_19163)
);

NAND2xp5_ASAP7_75t_L g19164 ( 
.A(n_18694),
.B(n_8069),
.Y(n_19164)
);

AND2x2_ASAP7_75t_L g19165 ( 
.A(n_18667),
.B(n_8873),
.Y(n_19165)
);

INVx1_ASAP7_75t_L g19166 ( 
.A(n_18694),
.Y(n_19166)
);

INVx1_ASAP7_75t_L g19167 ( 
.A(n_18694),
.Y(n_19167)
);

INVx1_ASAP7_75t_L g19168 ( 
.A(n_18911),
.Y(n_19168)
);

OAI221xp5_ASAP7_75t_L g19169 ( 
.A1(n_19008),
.A2(n_8379),
.B1(n_8253),
.B2(n_7494),
.C(n_7528),
.Y(n_19169)
);

NAND2xp5_ASAP7_75t_L g19170 ( 
.A(n_18955),
.B(n_8078),
.Y(n_19170)
);

AND2x2_ASAP7_75t_L g19171 ( 
.A(n_19161),
.B(n_7120),
.Y(n_19171)
);

INVx1_ASAP7_75t_L g19172 ( 
.A(n_19160),
.Y(n_19172)
);

NOR3xp33_ASAP7_75t_L g19173 ( 
.A(n_18992),
.B(n_5120),
.C(n_5066),
.Y(n_19173)
);

NOR4xp25_ASAP7_75t_SL g19174 ( 
.A(n_18983),
.B(n_8786),
.C(n_8795),
.D(n_8779),
.Y(n_19174)
);

NOR2xp33_ASAP7_75t_SL g19175 ( 
.A(n_18935),
.B(n_5066),
.Y(n_19175)
);

NOR3xp33_ASAP7_75t_SL g19176 ( 
.A(n_18919),
.B(n_7126),
.C(n_7111),
.Y(n_19176)
);

NAND2xp33_ASAP7_75t_R g19177 ( 
.A(n_19166),
.B(n_8832),
.Y(n_19177)
);

NAND2xp5_ASAP7_75t_L g19178 ( 
.A(n_19167),
.B(n_8078),
.Y(n_19178)
);

HB1xp67_ASAP7_75t_L g19179 ( 
.A(n_18978),
.Y(n_19179)
);

INVx1_ASAP7_75t_L g19180 ( 
.A(n_18928),
.Y(n_19180)
);

O2A1O1Ixp33_ASAP7_75t_L g19181 ( 
.A1(n_19002),
.A2(n_8379),
.B(n_8253),
.C(n_8320),
.Y(n_19181)
);

NOR3xp33_ASAP7_75t_SL g19182 ( 
.A(n_18984),
.B(n_7130),
.C(n_7126),
.Y(n_19182)
);

NOR3xp33_ASAP7_75t_L g19183 ( 
.A(n_18918),
.B(n_5120),
.C(n_5066),
.Y(n_19183)
);

OR2x2_ASAP7_75t_L g19184 ( 
.A(n_18929),
.B(n_8873),
.Y(n_19184)
);

INVx2_ASAP7_75t_L g19185 ( 
.A(n_18949),
.Y(n_19185)
);

INVx1_ASAP7_75t_L g19186 ( 
.A(n_18988),
.Y(n_19186)
);

INVx1_ASAP7_75t_L g19187 ( 
.A(n_18982),
.Y(n_19187)
);

INVx1_ASAP7_75t_L g19188 ( 
.A(n_18960),
.Y(n_19188)
);

NOR2xp33_ASAP7_75t_L g19189 ( 
.A(n_18966),
.B(n_5897),
.Y(n_19189)
);

NOR4xp25_ASAP7_75t_SL g19190 ( 
.A(n_19009),
.B(n_8798),
.C(n_8803),
.D(n_8795),
.Y(n_19190)
);

NOR2xp33_ASAP7_75t_L g19191 ( 
.A(n_18991),
.B(n_5960),
.Y(n_19191)
);

NAND2xp5_ASAP7_75t_SL g19192 ( 
.A(n_18914),
.B(n_7367),
.Y(n_19192)
);

AOI221xp5_ASAP7_75t_L g19193 ( 
.A1(n_19040),
.A2(n_8093),
.B1(n_8110),
.B2(n_8083),
.C(n_8078),
.Y(n_19193)
);

INVx1_ASAP7_75t_L g19194 ( 
.A(n_18975),
.Y(n_19194)
);

INVx2_ASAP7_75t_L g19195 ( 
.A(n_19033),
.Y(n_19195)
);

AND3x1_ASAP7_75t_L g19196 ( 
.A(n_18964),
.B(n_19078),
.C(n_19012),
.Y(n_19196)
);

AND2x2_ASAP7_75t_L g19197 ( 
.A(n_18980),
.B(n_7120),
.Y(n_19197)
);

AOI22xp33_ASAP7_75t_L g19198 ( 
.A1(n_18997),
.A2(n_7375),
.B1(n_7377),
.B2(n_7367),
.Y(n_19198)
);

AND2x2_ASAP7_75t_L g19199 ( 
.A(n_18977),
.B(n_7120),
.Y(n_19199)
);

OR2x2_ASAP7_75t_L g19200 ( 
.A(n_19011),
.B(n_8873),
.Y(n_19200)
);

AND2x2_ASAP7_75t_L g19201 ( 
.A(n_18945),
.B(n_7120),
.Y(n_19201)
);

NAND2xp5_ASAP7_75t_L g19202 ( 
.A(n_18962),
.B(n_8078),
.Y(n_19202)
);

INVx1_ASAP7_75t_L g19203 ( 
.A(n_18934),
.Y(n_19203)
);

INVx1_ASAP7_75t_L g19204 ( 
.A(n_18938),
.Y(n_19204)
);

NAND2xp5_ASAP7_75t_L g19205 ( 
.A(n_18932),
.B(n_8083),
.Y(n_19205)
);

INVx2_ASAP7_75t_L g19206 ( 
.A(n_18940),
.Y(n_19206)
);

NAND2xp5_ASAP7_75t_L g19207 ( 
.A(n_18941),
.B(n_8083),
.Y(n_19207)
);

INVx1_ASAP7_75t_SL g19208 ( 
.A(n_19036),
.Y(n_19208)
);

XNOR2xp5_ASAP7_75t_L g19209 ( 
.A(n_19023),
.B(n_7701),
.Y(n_19209)
);

AOI322xp5_ASAP7_75t_L g19210 ( 
.A1(n_18976),
.A2(n_7632),
.A3(n_7626),
.B1(n_7036),
.B2(n_7307),
.C1(n_7254),
.C2(n_7339),
.Y(n_19210)
);

INVx1_ASAP7_75t_L g19211 ( 
.A(n_18942),
.Y(n_19211)
);

INVx1_ASAP7_75t_L g19212 ( 
.A(n_18943),
.Y(n_19212)
);

AND2x2_ASAP7_75t_L g19213 ( 
.A(n_18924),
.B(n_7120),
.Y(n_19213)
);

NAND2xp5_ASAP7_75t_L g19214 ( 
.A(n_18965),
.B(n_18967),
.Y(n_19214)
);

INVx1_ASAP7_75t_L g19215 ( 
.A(n_18972),
.Y(n_19215)
);

CKINVDCx20_ASAP7_75t_R g19216 ( 
.A(n_18936),
.Y(n_19216)
);

INVx1_ASAP7_75t_L g19217 ( 
.A(n_19043),
.Y(n_19217)
);

INVx1_ASAP7_75t_L g19218 ( 
.A(n_18913),
.Y(n_19218)
);

INVxp67_ASAP7_75t_L g19219 ( 
.A(n_18973),
.Y(n_19219)
);

INVx1_ASAP7_75t_L g19220 ( 
.A(n_18987),
.Y(n_19220)
);

INVx1_ASAP7_75t_L g19221 ( 
.A(n_19007),
.Y(n_19221)
);

AND2x2_ASAP7_75t_L g19222 ( 
.A(n_18952),
.B(n_7120),
.Y(n_19222)
);

NAND2xp5_ASAP7_75t_L g19223 ( 
.A(n_19070),
.B(n_8083),
.Y(n_19223)
);

INVx2_ASAP7_75t_SL g19224 ( 
.A(n_19148),
.Y(n_19224)
);

NOR2xp33_ASAP7_75t_L g19225 ( 
.A(n_19052),
.B(n_5960),
.Y(n_19225)
);

NAND2xp5_ASAP7_75t_L g19226 ( 
.A(n_18930),
.B(n_8093),
.Y(n_19226)
);

INVx1_ASAP7_75t_L g19227 ( 
.A(n_18933),
.Y(n_19227)
);

INVx4_ASAP7_75t_L g19228 ( 
.A(n_19045),
.Y(n_19228)
);

AND2x2_ASAP7_75t_L g19229 ( 
.A(n_18957),
.B(n_18922),
.Y(n_19229)
);

INVx2_ASAP7_75t_L g19230 ( 
.A(n_18927),
.Y(n_19230)
);

NAND2xp5_ASAP7_75t_L g19231 ( 
.A(n_18956),
.B(n_8093),
.Y(n_19231)
);

INVx2_ASAP7_75t_SL g19232 ( 
.A(n_19054),
.Y(n_19232)
);

NOR3xp33_ASAP7_75t_SL g19233 ( 
.A(n_19120),
.B(n_7130),
.C(n_7332),
.Y(n_19233)
);

INVx1_ASAP7_75t_L g19234 ( 
.A(n_19071),
.Y(n_19234)
);

INVxp67_ASAP7_75t_L g19235 ( 
.A(n_19000),
.Y(n_19235)
);

NAND2xp5_ASAP7_75t_SL g19236 ( 
.A(n_19053),
.B(n_7375),
.Y(n_19236)
);

BUFx2_ASAP7_75t_SL g19237 ( 
.A(n_18995),
.Y(n_19237)
);

INVx1_ASAP7_75t_L g19238 ( 
.A(n_19051),
.Y(n_19238)
);

INVx1_ASAP7_75t_SL g19239 ( 
.A(n_19039),
.Y(n_19239)
);

AOI32xp33_ASAP7_75t_L g19240 ( 
.A1(n_19026),
.A2(n_19047),
.A3(n_19049),
.B1(n_19140),
.B2(n_19062),
.Y(n_19240)
);

AND2x2_ASAP7_75t_L g19241 ( 
.A(n_19156),
.B(n_7150),
.Y(n_19241)
);

INVx2_ASAP7_75t_L g19242 ( 
.A(n_19102),
.Y(n_19242)
);

NOR3xp33_ASAP7_75t_SL g19243 ( 
.A(n_19004),
.B(n_7130),
.C(n_7332),
.Y(n_19243)
);

INVx1_ASAP7_75t_L g19244 ( 
.A(n_19118),
.Y(n_19244)
);

INVx1_ASAP7_75t_L g19245 ( 
.A(n_18959),
.Y(n_19245)
);

AND2x2_ASAP7_75t_L g19246 ( 
.A(n_19162),
.B(n_7150),
.Y(n_19246)
);

NAND2x1_ASAP7_75t_L g19247 ( 
.A(n_18968),
.B(n_8572),
.Y(n_19247)
);

INVx3_ASAP7_75t_SL g19248 ( 
.A(n_19068),
.Y(n_19248)
);

NOR3xp33_ASAP7_75t_SL g19249 ( 
.A(n_18951),
.B(n_7341),
.C(n_7202),
.Y(n_19249)
);

AOI21xp33_ASAP7_75t_L g19250 ( 
.A1(n_18986),
.A2(n_8320),
.B(n_8832),
.Y(n_19250)
);

INVx1_ASAP7_75t_L g19251 ( 
.A(n_18963),
.Y(n_19251)
);

AND2x2_ASAP7_75t_L g19252 ( 
.A(n_19165),
.B(n_7150),
.Y(n_19252)
);

AOI21xp5_ASAP7_75t_L g19253 ( 
.A1(n_19061),
.A2(n_19005),
.B(n_18981),
.Y(n_19253)
);

OR2x2_ASAP7_75t_L g19254 ( 
.A(n_19059),
.B(n_8873),
.Y(n_19254)
);

OR2x2_ASAP7_75t_L g19255 ( 
.A(n_18926),
.B(n_8013),
.Y(n_19255)
);

INVx2_ASAP7_75t_SL g19256 ( 
.A(n_19044),
.Y(n_19256)
);

INVx1_ASAP7_75t_L g19257 ( 
.A(n_18971),
.Y(n_19257)
);

NAND2xp5_ASAP7_75t_L g19258 ( 
.A(n_19016),
.B(n_8093),
.Y(n_19258)
);

NAND2xp5_ASAP7_75t_L g19259 ( 
.A(n_19131),
.B(n_8110),
.Y(n_19259)
);

NAND2xp5_ASAP7_75t_L g19260 ( 
.A(n_19001),
.B(n_19074),
.Y(n_19260)
);

AOI21xp33_ASAP7_75t_SL g19261 ( 
.A1(n_19046),
.A2(n_8303),
.B(n_8311),
.Y(n_19261)
);

NAND2xp5_ASAP7_75t_L g19262 ( 
.A(n_18937),
.B(n_8110),
.Y(n_19262)
);

NAND2xp5_ASAP7_75t_L g19263 ( 
.A(n_19063),
.B(n_8110),
.Y(n_19263)
);

NAND2xp33_ASAP7_75t_R g19264 ( 
.A(n_19034),
.B(n_8832),
.Y(n_19264)
);

NAND2xp5_ASAP7_75t_SL g19265 ( 
.A(n_19060),
.B(n_7375),
.Y(n_19265)
);

NAND2xp5_ASAP7_75t_L g19266 ( 
.A(n_18998),
.B(n_8111),
.Y(n_19266)
);

NOR3xp33_ASAP7_75t_SL g19267 ( 
.A(n_19069),
.B(n_7341),
.C(n_7202),
.Y(n_19267)
);

NOR3xp33_ASAP7_75t_L g19268 ( 
.A(n_19032),
.B(n_5161),
.C(n_5120),
.Y(n_19268)
);

INVx1_ASAP7_75t_L g19269 ( 
.A(n_19013),
.Y(n_19269)
);

NOR2xp33_ASAP7_75t_R g19270 ( 
.A(n_19056),
.B(n_4674),
.Y(n_19270)
);

NOR2xp33_ASAP7_75t_L g19271 ( 
.A(n_18925),
.B(n_5344),
.Y(n_19271)
);

XNOR2xp5_ASAP7_75t_L g19272 ( 
.A(n_19028),
.B(n_7701),
.Y(n_19272)
);

NAND2xp33_ASAP7_75t_R g19273 ( 
.A(n_19041),
.B(n_8832),
.Y(n_19273)
);

NAND2xp5_ASAP7_75t_L g19274 ( 
.A(n_19093),
.B(n_8111),
.Y(n_19274)
);

AND2x2_ASAP7_75t_L g19275 ( 
.A(n_18969),
.B(n_7150),
.Y(n_19275)
);

AND2x2_ASAP7_75t_L g19276 ( 
.A(n_18917),
.B(n_7150),
.Y(n_19276)
);

NOR2xp33_ASAP7_75t_L g19277 ( 
.A(n_19138),
.B(n_5344),
.Y(n_19277)
);

CKINVDCx5p33_ASAP7_75t_R g19278 ( 
.A(n_19082),
.Y(n_19278)
);

NAND2xp5_ASAP7_75t_SL g19279 ( 
.A(n_19006),
.B(n_7375),
.Y(n_19279)
);

CKINVDCx20_ASAP7_75t_R g19280 ( 
.A(n_19038),
.Y(n_19280)
);

INVx1_ASAP7_75t_L g19281 ( 
.A(n_19143),
.Y(n_19281)
);

NAND2xp5_ASAP7_75t_L g19282 ( 
.A(n_19091),
.B(n_8111),
.Y(n_19282)
);

INVx1_ASAP7_75t_L g19283 ( 
.A(n_19119),
.Y(n_19283)
);

AND2x2_ASAP7_75t_L g19284 ( 
.A(n_18950),
.B(n_7150),
.Y(n_19284)
);

INVxp67_ASAP7_75t_L g19285 ( 
.A(n_19042),
.Y(n_19285)
);

OAI22xp5_ASAP7_75t_L g19286 ( 
.A1(n_19098),
.A2(n_8124),
.B1(n_8126),
.B2(n_8111),
.Y(n_19286)
);

NOR4xp25_ASAP7_75t_SL g19287 ( 
.A(n_19149),
.B(n_8803),
.C(n_8820),
.D(n_8798),
.Y(n_19287)
);

INVx1_ASAP7_75t_L g19288 ( 
.A(n_19014),
.Y(n_19288)
);

OR2x2_ASAP7_75t_L g19289 ( 
.A(n_19020),
.B(n_8013),
.Y(n_19289)
);

INVx1_ASAP7_75t_L g19290 ( 
.A(n_19107),
.Y(n_19290)
);

NAND2xp5_ASAP7_75t_L g19291 ( 
.A(n_19086),
.B(n_8124),
.Y(n_19291)
);

INVx1_ASAP7_75t_L g19292 ( 
.A(n_19124),
.Y(n_19292)
);

INVx1_ASAP7_75t_L g19293 ( 
.A(n_18979),
.Y(n_19293)
);

INVxp67_ASAP7_75t_L g19294 ( 
.A(n_18921),
.Y(n_19294)
);

INVx1_ASAP7_75t_L g19295 ( 
.A(n_19021),
.Y(n_19295)
);

NAND2xp5_ASAP7_75t_L g19296 ( 
.A(n_19088),
.B(n_8124),
.Y(n_19296)
);

CKINVDCx5p33_ASAP7_75t_R g19297 ( 
.A(n_19058),
.Y(n_19297)
);

INVx1_ASAP7_75t_L g19298 ( 
.A(n_19152),
.Y(n_19298)
);

AND2x2_ASAP7_75t_L g19299 ( 
.A(n_19151),
.B(n_19146),
.Y(n_19299)
);

INVx1_ASAP7_75t_L g19300 ( 
.A(n_19154),
.Y(n_19300)
);

INVx1_ASAP7_75t_L g19301 ( 
.A(n_19157),
.Y(n_19301)
);

INVx1_ASAP7_75t_L g19302 ( 
.A(n_19159),
.Y(n_19302)
);

XNOR2x1_ASAP7_75t_L g19303 ( 
.A(n_19116),
.B(n_8494),
.Y(n_19303)
);

INVx1_ASAP7_75t_L g19304 ( 
.A(n_19164),
.Y(n_19304)
);

INVx1_ASAP7_75t_L g19305 ( 
.A(n_19123),
.Y(n_19305)
);

AND2x2_ASAP7_75t_L g19306 ( 
.A(n_18993),
.B(n_19076),
.Y(n_19306)
);

INVx2_ASAP7_75t_L g19307 ( 
.A(n_18953),
.Y(n_19307)
);

INVx1_ASAP7_75t_L g19308 ( 
.A(n_19072),
.Y(n_19308)
);

BUFx2_ASAP7_75t_L g19309 ( 
.A(n_18947),
.Y(n_19309)
);

INVx2_ASAP7_75t_L g19310 ( 
.A(n_18985),
.Y(n_19310)
);

AOI322xp5_ASAP7_75t_L g19311 ( 
.A1(n_19150),
.A2(n_7632),
.A3(n_7626),
.B1(n_7356),
.B2(n_7464),
.C1(n_7234),
.C2(n_7475),
.Y(n_19311)
);

XNOR2xp5_ASAP7_75t_L g19312 ( 
.A(n_19100),
.B(n_7701),
.Y(n_19312)
);

AND2x2_ASAP7_75t_L g19313 ( 
.A(n_19003),
.B(n_7186),
.Y(n_19313)
);

NOR2x1_ASAP7_75t_L g19314 ( 
.A(n_19142),
.B(n_7436),
.Y(n_19314)
);

OR2x2_ASAP7_75t_L g19315 ( 
.A(n_18974),
.B(n_8013),
.Y(n_19315)
);

CKINVDCx5p33_ASAP7_75t_R g19316 ( 
.A(n_19073),
.Y(n_19316)
);

INVx1_ASAP7_75t_L g19317 ( 
.A(n_18989),
.Y(n_19317)
);

INVx1_ASAP7_75t_L g19318 ( 
.A(n_18990),
.Y(n_19318)
);

INVx1_ASAP7_75t_L g19319 ( 
.A(n_18994),
.Y(n_19319)
);

INVx1_ASAP7_75t_L g19320 ( 
.A(n_19092),
.Y(n_19320)
);

AND2x2_ASAP7_75t_L g19321 ( 
.A(n_19015),
.B(n_19019),
.Y(n_19321)
);

CKINVDCx20_ASAP7_75t_R g19322 ( 
.A(n_19035),
.Y(n_19322)
);

NAND2xp5_ASAP7_75t_L g19323 ( 
.A(n_19114),
.B(n_8124),
.Y(n_19323)
);

INVx3_ASAP7_75t_L g19324 ( 
.A(n_19085),
.Y(n_19324)
);

INVx1_ASAP7_75t_L g19325 ( 
.A(n_19097),
.Y(n_19325)
);

NOR2xp33_ASAP7_75t_L g19326 ( 
.A(n_18939),
.B(n_5344),
.Y(n_19326)
);

NAND2xp5_ASAP7_75t_L g19327 ( 
.A(n_19077),
.B(n_8126),
.Y(n_19327)
);

AOI22xp5_ASAP7_75t_L g19328 ( 
.A1(n_19137),
.A2(n_7377),
.B1(n_7378),
.B2(n_7375),
.Y(n_19328)
);

NOR2x1_ASAP7_75t_L g19329 ( 
.A(n_19103),
.B(n_19089),
.Y(n_19329)
);

OAI322xp33_ASAP7_75t_L g19330 ( 
.A1(n_18958),
.A2(n_8178),
.A3(n_8129),
.B1(n_8196),
.B2(n_8232),
.C1(n_8149),
.C2(n_8126),
.Y(n_19330)
);

INVx1_ASAP7_75t_L g19331 ( 
.A(n_18946),
.Y(n_19331)
);

INVx1_ASAP7_75t_L g19332 ( 
.A(n_18954),
.Y(n_19332)
);

NOR4xp25_ASAP7_75t_SL g19333 ( 
.A(n_19115),
.B(n_8823),
.C(n_8827),
.D(n_8820),
.Y(n_19333)
);

OAI22xp5_ASAP7_75t_L g19334 ( 
.A1(n_19155),
.A2(n_8129),
.B1(n_8149),
.B2(n_8126),
.Y(n_19334)
);

INVx2_ASAP7_75t_L g19335 ( 
.A(n_19031),
.Y(n_19335)
);

INVx2_ASAP7_75t_L g19336 ( 
.A(n_19022),
.Y(n_19336)
);

INVx1_ASAP7_75t_L g19337 ( 
.A(n_19106),
.Y(n_19337)
);

NAND2xp5_ASAP7_75t_SL g19338 ( 
.A(n_19067),
.B(n_19153),
.Y(n_19338)
);

AOI211xp5_ASAP7_75t_L g19339 ( 
.A1(n_18931),
.A2(n_8303),
.B(n_8494),
.C(n_8433),
.Y(n_19339)
);

AND2x2_ASAP7_75t_L g19340 ( 
.A(n_19025),
.B(n_19027),
.Y(n_19340)
);

AND2x2_ASAP7_75t_L g19341 ( 
.A(n_19010),
.B(n_18970),
.Y(n_19341)
);

INVx1_ASAP7_75t_L g19342 ( 
.A(n_19109),
.Y(n_19342)
);

INVx1_ASAP7_75t_L g19343 ( 
.A(n_19112),
.Y(n_19343)
);

AOI311xp33_ASAP7_75t_L g19344 ( 
.A1(n_18915),
.A2(n_8827),
.A3(n_8843),
.B(n_8830),
.C(n_8823),
.Y(n_19344)
);

INVx1_ASAP7_75t_L g19345 ( 
.A(n_18948),
.Y(n_19345)
);

AOI211xp5_ASAP7_75t_L g19346 ( 
.A1(n_18923),
.A2(n_8303),
.B(n_8494),
.C(n_8969),
.Y(n_19346)
);

NOR3xp33_ASAP7_75t_SL g19347 ( 
.A(n_19080),
.B(n_18912),
.C(n_19104),
.Y(n_19347)
);

NOR2x1_ASAP7_75t_L g19348 ( 
.A(n_18999),
.B(n_7436),
.Y(n_19348)
);

AOI22xp33_ASAP7_75t_L g19349 ( 
.A1(n_19110),
.A2(n_7377),
.B1(n_7378),
.B2(n_7375),
.Y(n_19349)
);

NOR4xp25_ASAP7_75t_SL g19350 ( 
.A(n_18920),
.B(n_19130),
.C(n_19101),
.D(n_19128),
.Y(n_19350)
);

NAND2xp33_ASAP7_75t_L g19351 ( 
.A(n_19113),
.B(n_7377),
.Y(n_19351)
);

INVx1_ASAP7_75t_L g19352 ( 
.A(n_19048),
.Y(n_19352)
);

AND2x2_ASAP7_75t_L g19353 ( 
.A(n_19057),
.B(n_7186),
.Y(n_19353)
);

INVx1_ASAP7_75t_L g19354 ( 
.A(n_19083),
.Y(n_19354)
);

AND2x2_ASAP7_75t_L g19355 ( 
.A(n_19127),
.B(n_7186),
.Y(n_19355)
);

NAND2xp5_ASAP7_75t_L g19356 ( 
.A(n_19147),
.B(n_8129),
.Y(n_19356)
);

INVx1_ASAP7_75t_SL g19357 ( 
.A(n_19087),
.Y(n_19357)
);

INVxp67_ASAP7_75t_L g19358 ( 
.A(n_19081),
.Y(n_19358)
);

OR2x2_ASAP7_75t_L g19359 ( 
.A(n_19117),
.B(n_8013),
.Y(n_19359)
);

INVx1_ASAP7_75t_L g19360 ( 
.A(n_19111),
.Y(n_19360)
);

INVx1_ASAP7_75t_L g19361 ( 
.A(n_19064),
.Y(n_19361)
);

INVx1_ASAP7_75t_L g19362 ( 
.A(n_19090),
.Y(n_19362)
);

NAND2xp5_ASAP7_75t_L g19363 ( 
.A(n_19084),
.B(n_19144),
.Y(n_19363)
);

NAND2xp5_ASAP7_75t_L g19364 ( 
.A(n_19145),
.B(n_8129),
.Y(n_19364)
);

NAND2xp5_ASAP7_75t_L g19365 ( 
.A(n_19139),
.B(n_8149),
.Y(n_19365)
);

INVx4_ASAP7_75t_L g19366 ( 
.A(n_19121),
.Y(n_19366)
);

NAND2xp5_ASAP7_75t_L g19367 ( 
.A(n_19099),
.B(n_8149),
.Y(n_19367)
);

INVx2_ASAP7_75t_L g19368 ( 
.A(n_19018),
.Y(n_19368)
);

INVxp67_ASAP7_75t_L g19369 ( 
.A(n_19108),
.Y(n_19369)
);

INVx2_ASAP7_75t_L g19370 ( 
.A(n_19132),
.Y(n_19370)
);

CKINVDCx5p33_ASAP7_75t_R g19371 ( 
.A(n_19029),
.Y(n_19371)
);

XOR2x2_ASAP7_75t_L g19372 ( 
.A(n_19050),
.B(n_8552),
.Y(n_19372)
);

NAND2xp5_ASAP7_75t_L g19373 ( 
.A(n_19133),
.B(n_8178),
.Y(n_19373)
);

NAND2xp5_ASAP7_75t_L g19374 ( 
.A(n_19141),
.B(n_8178),
.Y(n_19374)
);

INVxp67_ASAP7_75t_L g19375 ( 
.A(n_18944),
.Y(n_19375)
);

INVx2_ASAP7_75t_L g19376 ( 
.A(n_19134),
.Y(n_19376)
);

NOR2xp33_ASAP7_75t_L g19377 ( 
.A(n_19122),
.B(n_5344),
.Y(n_19377)
);

NAND2x1_ASAP7_75t_L g19378 ( 
.A(n_19129),
.B(n_8588),
.Y(n_19378)
);

AND2x2_ASAP7_75t_L g19379 ( 
.A(n_18916),
.B(n_7186),
.Y(n_19379)
);

OR2x2_ASAP7_75t_L g19380 ( 
.A(n_19096),
.B(n_8013),
.Y(n_19380)
);

NAND2xp5_ASAP7_75t_L g19381 ( 
.A(n_19055),
.B(n_8178),
.Y(n_19381)
);

OR2x2_ASAP7_75t_L g19382 ( 
.A(n_19066),
.B(n_19126),
.Y(n_19382)
);

OAI21xp33_ASAP7_75t_SL g19383 ( 
.A1(n_19163),
.A2(n_8313),
.B(n_8311),
.Y(n_19383)
);

INVx1_ASAP7_75t_L g19384 ( 
.A(n_19094),
.Y(n_19384)
);

NAND2xp5_ASAP7_75t_L g19385 ( 
.A(n_19075),
.B(n_8196),
.Y(n_19385)
);

AOI31xp33_ASAP7_75t_L g19386 ( 
.A1(n_19179),
.A2(n_19135),
.A3(n_19079),
.B(n_19024),
.Y(n_19386)
);

AOI21xp5_ASAP7_75t_L g19387 ( 
.A1(n_19338),
.A2(n_18996),
.B(n_19037),
.Y(n_19387)
);

NAND5xp2_ASAP7_75t_SL g19388 ( 
.A(n_19297),
.B(n_19125),
.C(n_19136),
.D(n_19105),
.E(n_18961),
.Y(n_19388)
);

AOI22x1_ASAP7_75t_SL g19389 ( 
.A1(n_19280),
.A2(n_19017),
.B1(n_19030),
.B2(n_19121),
.Y(n_19389)
);

AOI21xp5_ASAP7_75t_L g19390 ( 
.A1(n_19214),
.A2(n_19158),
.B(n_19095),
.Y(n_19390)
);

INVx2_ASAP7_75t_SL g19391 ( 
.A(n_19314),
.Y(n_19391)
);

NOR2x1_ASAP7_75t_L g19392 ( 
.A(n_19228),
.B(n_19095),
.Y(n_19392)
);

NOR3x1_ASAP7_75t_L g19393 ( 
.A(n_19256),
.B(n_19065),
.C(n_8466),
.Y(n_19393)
);

NAND2xp5_ASAP7_75t_L g19394 ( 
.A(n_19228),
.B(n_8196),
.Y(n_19394)
);

AND2x2_ASAP7_75t_L g19395 ( 
.A(n_19199),
.B(n_7186),
.Y(n_19395)
);

INVx1_ASAP7_75t_L g19396 ( 
.A(n_19272),
.Y(n_19396)
);

INVx1_ASAP7_75t_L g19397 ( 
.A(n_19187),
.Y(n_19397)
);

NAND2xp5_ASAP7_75t_L g19398 ( 
.A(n_19217),
.B(n_8196),
.Y(n_19398)
);

AOI22xp5_ASAP7_75t_L g19399 ( 
.A1(n_19216),
.A2(n_7378),
.B1(n_7438),
.B2(n_7377),
.Y(n_19399)
);

NAND3xp33_ASAP7_75t_L g19400 ( 
.A(n_19240),
.B(n_4890),
.C(n_4856),
.Y(n_19400)
);

OAI211xp5_ASAP7_75t_SL g19401 ( 
.A1(n_19219),
.A2(n_19369),
.B(n_19292),
.C(n_19253),
.Y(n_19401)
);

OAI21xp5_ASAP7_75t_L g19402 ( 
.A1(n_19220),
.A2(n_8975),
.B(n_8972),
.Y(n_19402)
);

NAND2xp5_ASAP7_75t_L g19403 ( 
.A(n_19180),
.B(n_8232),
.Y(n_19403)
);

NAND2xp5_ASAP7_75t_L g19404 ( 
.A(n_19276),
.B(n_8232),
.Y(n_19404)
);

NAND2xp5_ASAP7_75t_L g19405 ( 
.A(n_19244),
.B(n_8232),
.Y(n_19405)
);

INVx1_ASAP7_75t_L g19406 ( 
.A(n_19242),
.Y(n_19406)
);

XNOR2x1_ASAP7_75t_SL g19407 ( 
.A(n_19232),
.B(n_5106),
.Y(n_19407)
);

NAND2xp5_ASAP7_75t_L g19408 ( 
.A(n_19171),
.B(n_19208),
.Y(n_19408)
);

AOI22xp5_ASAP7_75t_L g19409 ( 
.A1(n_19239),
.A2(n_7378),
.B1(n_7438),
.B2(n_7377),
.Y(n_19409)
);

NAND2xp5_ASAP7_75t_L g19410 ( 
.A(n_19168),
.B(n_8237),
.Y(n_19410)
);

NAND2xp5_ASAP7_75t_L g19411 ( 
.A(n_19172),
.B(n_8237),
.Y(n_19411)
);

NOR3xp33_ASAP7_75t_L g19412 ( 
.A(n_19188),
.B(n_5195),
.C(n_5161),
.Y(n_19412)
);

NAND2xp5_ASAP7_75t_SL g19413 ( 
.A(n_19206),
.B(n_7377),
.Y(n_19413)
);

AOI22xp5_ASAP7_75t_L g19414 ( 
.A1(n_19221),
.A2(n_7378),
.B1(n_7438),
.B2(n_7377),
.Y(n_19414)
);

OAI21xp33_ASAP7_75t_L g19415 ( 
.A1(n_19191),
.A2(n_7494),
.B(n_7440),
.Y(n_19415)
);

AND2x2_ASAP7_75t_L g19416 ( 
.A(n_19201),
.B(n_7186),
.Y(n_19416)
);

INVx2_ASAP7_75t_L g19417 ( 
.A(n_19372),
.Y(n_19417)
);

BUFx6f_ASAP7_75t_L g19418 ( 
.A(n_19248),
.Y(n_19418)
);

INVx1_ASAP7_75t_L g19419 ( 
.A(n_19312),
.Y(n_19419)
);

AOI211x1_ASAP7_75t_L g19420 ( 
.A1(n_19192),
.A2(n_9129),
.B(n_9160),
.C(n_9087),
.Y(n_19420)
);

NAND4xp75_ASAP7_75t_L g19421 ( 
.A(n_19196),
.B(n_19234),
.C(n_19238),
.D(n_19194),
.Y(n_19421)
);

AOI22xp5_ASAP7_75t_L g19422 ( 
.A1(n_19322),
.A2(n_7378),
.B1(n_7438),
.B2(n_7377),
.Y(n_19422)
);

NOR2x1_ASAP7_75t_L g19423 ( 
.A(n_19366),
.B(n_19203),
.Y(n_19423)
);

NOR2xp33_ASAP7_75t_L g19424 ( 
.A(n_19204),
.B(n_5344),
.Y(n_19424)
);

NAND2xp5_ASAP7_75t_L g19425 ( 
.A(n_19197),
.B(n_8237),
.Y(n_19425)
);

NOR2xp67_ASAP7_75t_SL g19426 ( 
.A(n_19237),
.B(n_5382),
.Y(n_19426)
);

NAND2xp5_ASAP7_75t_SL g19427 ( 
.A(n_19185),
.B(n_7377),
.Y(n_19427)
);

NAND2xp5_ASAP7_75t_L g19428 ( 
.A(n_19211),
.B(n_8237),
.Y(n_19428)
);

INVx1_ASAP7_75t_L g19429 ( 
.A(n_19213),
.Y(n_19429)
);

NAND2xp5_ASAP7_75t_L g19430 ( 
.A(n_19212),
.B(n_8240),
.Y(n_19430)
);

NAND2xp5_ASAP7_75t_L g19431 ( 
.A(n_19215),
.B(n_8240),
.Y(n_19431)
);

AO22x1_ASAP7_75t_L g19432 ( 
.A1(n_19281),
.A2(n_4890),
.B1(n_5287),
.B2(n_4856),
.Y(n_19432)
);

AOI22xp5_ASAP7_75t_L g19433 ( 
.A1(n_19293),
.A2(n_7438),
.B1(n_7444),
.B2(n_7378),
.Y(n_19433)
);

INVx1_ASAP7_75t_SL g19434 ( 
.A(n_19223),
.Y(n_19434)
);

INVx1_ASAP7_75t_L g19435 ( 
.A(n_19205),
.Y(n_19435)
);

AO22x2_ASAP7_75t_L g19436 ( 
.A1(n_19224),
.A2(n_8242),
.B1(n_8254),
.B2(n_8240),
.Y(n_19436)
);

INVx1_ASAP7_75t_L g19437 ( 
.A(n_19170),
.Y(n_19437)
);

OAI21xp5_ASAP7_75t_SL g19438 ( 
.A1(n_19218),
.A2(n_7633),
.B(n_7701),
.Y(n_19438)
);

OAI22xp5_ASAP7_75t_L g19439 ( 
.A1(n_19198),
.A2(n_19349),
.B1(n_19169),
.B2(n_19316),
.Y(n_19439)
);

AOI211x1_ASAP7_75t_L g19440 ( 
.A1(n_19236),
.A2(n_19265),
.B(n_19259),
.C(n_19279),
.Y(n_19440)
);

NAND2xp5_ASAP7_75t_L g19441 ( 
.A(n_19209),
.B(n_8240),
.Y(n_19441)
);

AND2x2_ASAP7_75t_L g19442 ( 
.A(n_19225),
.B(n_7198),
.Y(n_19442)
);

AOI21xp5_ASAP7_75t_L g19443 ( 
.A1(n_19363),
.A2(n_8975),
.B(n_8972),
.Y(n_19443)
);

AOI22xp5_ASAP7_75t_L g19444 ( 
.A1(n_19189),
.A2(n_7438),
.B1(n_7444),
.B2(n_7378),
.Y(n_19444)
);

OA22x2_ASAP7_75t_L g19445 ( 
.A1(n_19290),
.A2(n_9230),
.B1(n_8324),
.B2(n_8254),
.Y(n_19445)
);

AOI22x1_ASAP7_75t_L g19446 ( 
.A1(n_19366),
.A2(n_5414),
.B1(n_5416),
.B2(n_5382),
.Y(n_19446)
);

INVx1_ASAP7_75t_L g19447 ( 
.A(n_19229),
.Y(n_19447)
);

AOI221xp5_ASAP7_75t_L g19448 ( 
.A1(n_19283),
.A2(n_8264),
.B1(n_8270),
.B2(n_8254),
.C(n_8242),
.Y(n_19448)
);

NOR3xp33_ASAP7_75t_SL g19449 ( 
.A(n_19278),
.B(n_7341),
.C(n_7202),
.Y(n_19449)
);

AO22x2_ASAP7_75t_L g19450 ( 
.A1(n_19336),
.A2(n_8254),
.B1(n_8264),
.B2(n_8242),
.Y(n_19450)
);

NOR2xp33_ASAP7_75t_L g19451 ( 
.A(n_19235),
.B(n_5344),
.Y(n_19451)
);

NOR3xp33_ASAP7_75t_L g19452 ( 
.A(n_19260),
.B(n_5195),
.C(n_5161),
.Y(n_19452)
);

OA22x2_ASAP7_75t_L g19453 ( 
.A1(n_19376),
.A2(n_9230),
.B1(n_8264),
.B2(n_8270),
.Y(n_19453)
);

AOI22xp33_ASAP7_75t_L g19454 ( 
.A1(n_19277),
.A2(n_7438),
.B1(n_7444),
.B2(n_7378),
.Y(n_19454)
);

AOI211xp5_ASAP7_75t_L g19455 ( 
.A1(n_19186),
.A2(n_8975),
.B(n_8972),
.C(n_8313),
.Y(n_19455)
);

AOI21xp5_ASAP7_75t_L g19456 ( 
.A1(n_19351),
.A2(n_8313),
.B(n_8311),
.Y(n_19456)
);

AOI211x1_ASAP7_75t_L g19457 ( 
.A1(n_19263),
.A2(n_9129),
.B(n_9254),
.C(n_9160),
.Y(n_19457)
);

AOI22xp5_ASAP7_75t_L g19458 ( 
.A1(n_19299),
.A2(n_7438),
.B1(n_7444),
.B2(n_7378),
.Y(n_19458)
);

AOI311xp33_ASAP7_75t_L g19459 ( 
.A1(n_19308),
.A2(n_8827),
.A3(n_8843),
.B(n_8830),
.C(n_8823),
.Y(n_19459)
);

OAI22xp5_ASAP7_75t_L g19460 ( 
.A1(n_19328),
.A2(n_8264),
.B1(n_8270),
.B2(n_8242),
.Y(n_19460)
);

OA22x2_ASAP7_75t_L g19461 ( 
.A1(n_19371),
.A2(n_9230),
.B1(n_8273),
.B2(n_8276),
.Y(n_19461)
);

INVx1_ASAP7_75t_L g19462 ( 
.A(n_19321),
.Y(n_19462)
);

NAND2xp5_ASAP7_75t_L g19463 ( 
.A(n_19340),
.B(n_8270),
.Y(n_19463)
);

OAI21xp33_ASAP7_75t_L g19464 ( 
.A1(n_19270),
.A2(n_19311),
.B(n_19271),
.Y(n_19464)
);

AOI22xp5_ASAP7_75t_L g19465 ( 
.A1(n_19326),
.A2(n_7444),
.B1(n_7457),
.B2(n_7438),
.Y(n_19465)
);

INVx1_ASAP7_75t_L g19466 ( 
.A(n_19341),
.Y(n_19466)
);

AOI21xp5_ASAP7_75t_L g19467 ( 
.A1(n_19202),
.A2(n_8313),
.B(n_8311),
.Y(n_19467)
);

INVx1_ASAP7_75t_L g19468 ( 
.A(n_19207),
.Y(n_19468)
);

INVx1_ASAP7_75t_SL g19469 ( 
.A(n_19306),
.Y(n_19469)
);

NAND2xp5_ASAP7_75t_L g19470 ( 
.A(n_19230),
.B(n_8273),
.Y(n_19470)
);

CKINVDCx20_ASAP7_75t_R g19471 ( 
.A(n_19227),
.Y(n_19471)
);

NAND2xp5_ASAP7_75t_L g19472 ( 
.A(n_19370),
.B(n_19324),
.Y(n_19472)
);

INVx1_ASAP7_75t_L g19473 ( 
.A(n_19352),
.Y(n_19473)
);

INVx1_ASAP7_75t_L g19474 ( 
.A(n_19348),
.Y(n_19474)
);

AOI211xp5_ASAP7_75t_L g19475 ( 
.A1(n_19325),
.A2(n_8461),
.B(n_8466),
.C(n_8863),
.Y(n_19475)
);

AOI211xp5_ASAP7_75t_L g19476 ( 
.A1(n_19305),
.A2(n_8461),
.B(n_8466),
.C(n_8863),
.Y(n_19476)
);

NAND2xp5_ASAP7_75t_SL g19477 ( 
.A(n_19175),
.B(n_7438),
.Y(n_19477)
);

NAND2xp5_ASAP7_75t_L g19478 ( 
.A(n_19324),
.B(n_8273),
.Y(n_19478)
);

INVx1_ASAP7_75t_L g19479 ( 
.A(n_19195),
.Y(n_19479)
);

OR2x2_ASAP7_75t_L g19480 ( 
.A(n_19200),
.B(n_8013),
.Y(n_19480)
);

AOI211xp5_ASAP7_75t_L g19481 ( 
.A1(n_19384),
.A2(n_8461),
.B(n_8866),
.C(n_8863),
.Y(n_19481)
);

AOI211x1_ASAP7_75t_L g19482 ( 
.A1(n_19365),
.A2(n_9129),
.B(n_9254),
.C(n_9160),
.Y(n_19482)
);

NAND2xp5_ASAP7_75t_L g19483 ( 
.A(n_19357),
.B(n_8273),
.Y(n_19483)
);

NAND2xp5_ASAP7_75t_L g19484 ( 
.A(n_19222),
.B(n_8276),
.Y(n_19484)
);

BUFx6f_ASAP7_75t_L g19485 ( 
.A(n_19337),
.Y(n_19485)
);

NAND2xp5_ASAP7_75t_SL g19486 ( 
.A(n_19368),
.B(n_7444),
.Y(n_19486)
);

AOI21xp5_ASAP7_75t_L g19487 ( 
.A1(n_19329),
.A2(n_8361),
.B(n_8280),
.Y(n_19487)
);

INVxp67_ASAP7_75t_L g19488 ( 
.A(n_19382),
.Y(n_19488)
);

INVxp67_ASAP7_75t_L g19489 ( 
.A(n_19295),
.Y(n_19489)
);

INVx1_ASAP7_75t_SL g19490 ( 
.A(n_19335),
.Y(n_19490)
);

NAND2xp5_ASAP7_75t_L g19491 ( 
.A(n_19182),
.B(n_8276),
.Y(n_19491)
);

NOR2xp33_ASAP7_75t_L g19492 ( 
.A(n_19294),
.B(n_19285),
.Y(n_19492)
);

OAI21x1_ASAP7_75t_L g19493 ( 
.A1(n_19307),
.A2(n_9230),
.B(n_8459),
.Y(n_19493)
);

INVx1_ASAP7_75t_L g19494 ( 
.A(n_19178),
.Y(n_19494)
);

AOI21xp5_ASAP7_75t_L g19495 ( 
.A1(n_19320),
.A2(n_8361),
.B(n_8280),
.Y(n_19495)
);

OAI21x1_ASAP7_75t_SL g19496 ( 
.A1(n_19310),
.A2(n_9297),
.B(n_9254),
.Y(n_19496)
);

AOI21xp5_ASAP7_75t_L g19497 ( 
.A1(n_19342),
.A2(n_8361),
.B(n_8280),
.Y(n_19497)
);

NOR3x1_ASAP7_75t_L g19498 ( 
.A(n_19309),
.B(n_8459),
.C(n_8863),
.Y(n_19498)
);

NOR4xp25_ASAP7_75t_L g19499 ( 
.A(n_19343),
.B(n_8843),
.C(n_8877),
.D(n_8830),
.Y(n_19499)
);

NAND2xp5_ASAP7_75t_L g19500 ( 
.A(n_19241),
.B(n_8276),
.Y(n_19500)
);

INVx1_ASAP7_75t_L g19501 ( 
.A(n_19298),
.Y(n_19501)
);

NAND2xp5_ASAP7_75t_SL g19502 ( 
.A(n_19361),
.B(n_7444),
.Y(n_19502)
);

OAI21xp33_ASAP7_75t_L g19503 ( 
.A1(n_19377),
.A2(n_7528),
.B(n_7440),
.Y(n_19503)
);

NOR2xp33_ASAP7_75t_L g19504 ( 
.A(n_19358),
.B(n_5344),
.Y(n_19504)
);

AOI22xp5_ASAP7_75t_L g19505 ( 
.A1(n_19173),
.A2(n_7457),
.B1(n_7460),
.B2(n_7444),
.Y(n_19505)
);

INVx1_ASAP7_75t_L g19506 ( 
.A(n_19300),
.Y(n_19506)
);

OAI21xp33_ASAP7_75t_L g19507 ( 
.A1(n_19233),
.A2(n_7594),
.B(n_7542),
.Y(n_19507)
);

OAI21xp5_ASAP7_75t_L g19508 ( 
.A1(n_19375),
.A2(n_7907),
.B(n_8866),
.Y(n_19508)
);

NOR2x1_ASAP7_75t_L g19509 ( 
.A(n_19360),
.B(n_7542),
.Y(n_19509)
);

NAND2xp5_ASAP7_75t_SL g19510 ( 
.A(n_19301),
.B(n_19302),
.Y(n_19510)
);

NOR3xp33_ASAP7_75t_L g19511 ( 
.A(n_19304),
.B(n_5195),
.C(n_5161),
.Y(n_19511)
);

INVx1_ASAP7_75t_L g19512 ( 
.A(n_19317),
.Y(n_19512)
);

NAND2xp5_ASAP7_75t_L g19513 ( 
.A(n_19246),
.B(n_19252),
.Y(n_19513)
);

AOI211xp5_ASAP7_75t_L g19514 ( 
.A1(n_19354),
.A2(n_8866),
.B(n_8459),
.C(n_7457),
.Y(n_19514)
);

NOR3xp33_ASAP7_75t_L g19515 ( 
.A(n_19245),
.B(n_5195),
.C(n_5161),
.Y(n_19515)
);

AND2x2_ASAP7_75t_L g19516 ( 
.A(n_19275),
.B(n_19355),
.Y(n_19516)
);

AO22x2_ASAP7_75t_L g19517 ( 
.A1(n_19251),
.A2(n_8289),
.B1(n_8314),
.B2(n_8280),
.Y(n_19517)
);

OAI222xp33_ASAP7_75t_L g19518 ( 
.A1(n_19359),
.A2(n_9297),
.B1(n_7795),
.B2(n_7867),
.C1(n_7903),
.C2(n_7857),
.Y(n_19518)
);

NOR3xp33_ASAP7_75t_L g19519 ( 
.A(n_19257),
.B(n_19269),
.C(n_19288),
.Y(n_19519)
);

NAND2xp5_ASAP7_75t_L g19520 ( 
.A(n_19318),
.B(n_19319),
.Y(n_19520)
);

NAND2xp5_ASAP7_75t_L g19521 ( 
.A(n_19284),
.B(n_8289),
.Y(n_19521)
);

NAND2xp5_ASAP7_75t_L g19522 ( 
.A(n_19362),
.B(n_8289),
.Y(n_19522)
);

AOI21xp5_ASAP7_75t_L g19523 ( 
.A1(n_19350),
.A2(n_8314),
.B(n_8289),
.Y(n_19523)
);

INVx1_ASAP7_75t_L g19524 ( 
.A(n_19274),
.Y(n_19524)
);

AOI22xp5_ASAP7_75t_L g19525 ( 
.A1(n_19183),
.A2(n_7457),
.B1(n_7460),
.B2(n_7444),
.Y(n_19525)
);

NAND2xp5_ASAP7_75t_L g19526 ( 
.A(n_19243),
.B(n_8314),
.Y(n_19526)
);

NAND2xp5_ASAP7_75t_L g19527 ( 
.A(n_19267),
.B(n_8314),
.Y(n_19527)
);

AO21x1_ASAP7_75t_L g19528 ( 
.A1(n_19345),
.A2(n_8885),
.B(n_8877),
.Y(n_19528)
);

AOI211xp5_ASAP7_75t_L g19529 ( 
.A1(n_19332),
.A2(n_8866),
.B(n_7457),
.C(n_7460),
.Y(n_19529)
);

NAND2xp5_ASAP7_75t_SL g19530 ( 
.A(n_19347),
.B(n_7444),
.Y(n_19530)
);

NOR2xp33_ASAP7_75t_L g19531 ( 
.A(n_19331),
.B(n_5524),
.Y(n_19531)
);

AOI21xp5_ASAP7_75t_L g19532 ( 
.A1(n_19296),
.A2(n_8319),
.B(n_8317),
.Y(n_19532)
);

OAI21xp5_ASAP7_75t_SL g19533 ( 
.A1(n_19268),
.A2(n_7633),
.B(n_9297),
.Y(n_19533)
);

NOR3x1_ASAP7_75t_L g19534 ( 
.A(n_19282),
.B(n_8287),
.C(n_8286),
.Y(n_19534)
);

OAI22xp33_ASAP7_75t_L g19535 ( 
.A1(n_19254),
.A2(n_7460),
.B1(n_7519),
.B2(n_7457),
.Y(n_19535)
);

NAND2xp5_ASAP7_75t_L g19536 ( 
.A(n_19313),
.B(n_8317),
.Y(n_19536)
);

AOI221xp5_ASAP7_75t_L g19537 ( 
.A1(n_19367),
.A2(n_8334),
.B1(n_8340),
.B2(n_8319),
.C(n_8317),
.Y(n_19537)
);

OAI21xp33_ASAP7_75t_L g19538 ( 
.A1(n_19303),
.A2(n_7594),
.B(n_7542),
.Y(n_19538)
);

AOI211x1_ASAP7_75t_SL g19539 ( 
.A1(n_19323),
.A2(n_8319),
.B(n_8334),
.C(n_8317),
.Y(n_19539)
);

AOI22xp33_ASAP7_75t_SL g19540 ( 
.A1(n_19379),
.A2(n_7460),
.B1(n_7519),
.B2(n_7457),
.Y(n_19540)
);

AO22x2_ASAP7_75t_L g19541 ( 
.A1(n_19289),
.A2(n_8334),
.B1(n_8340),
.B2(n_8319),
.Y(n_19541)
);

NOR2xp33_ASAP7_75t_SL g19542 ( 
.A(n_19184),
.B(n_5161),
.Y(n_19542)
);

NOR3xp33_ASAP7_75t_L g19543 ( 
.A(n_19291),
.B(n_19226),
.C(n_19231),
.Y(n_19543)
);

XOR2x2_ASAP7_75t_L g19544 ( 
.A(n_19353),
.B(n_8552),
.Y(n_19544)
);

NOR2xp67_ASAP7_75t_L g19545 ( 
.A(n_19266),
.B(n_5195),
.Y(n_19545)
);

AO22x2_ASAP7_75t_L g19546 ( 
.A1(n_19287),
.A2(n_8340),
.B1(n_8355),
.B2(n_8334),
.Y(n_19546)
);

AOI21xp5_ASAP7_75t_L g19547 ( 
.A1(n_19174),
.A2(n_8355),
.B(n_8340),
.Y(n_19547)
);

OAI21xp33_ASAP7_75t_L g19548 ( 
.A1(n_19327),
.A2(n_7594),
.B(n_7542),
.Y(n_19548)
);

INVx1_ASAP7_75t_L g19549 ( 
.A(n_19262),
.Y(n_19549)
);

NOR2xp33_ASAP7_75t_L g19550 ( 
.A(n_19255),
.B(n_5524),
.Y(n_19550)
);

AOI21xp5_ASAP7_75t_L g19551 ( 
.A1(n_19364),
.A2(n_8388),
.B(n_8355),
.Y(n_19551)
);

NOR2xp33_ASAP7_75t_L g19552 ( 
.A(n_19356),
.B(n_5524),
.Y(n_19552)
);

NAND2xp5_ASAP7_75t_SL g19553 ( 
.A(n_19380),
.B(n_7457),
.Y(n_19553)
);

NAND2xp5_ASAP7_75t_L g19554 ( 
.A(n_19249),
.B(n_8355),
.Y(n_19554)
);

NAND3xp33_ASAP7_75t_L g19555 ( 
.A(n_19373),
.B(n_4890),
.C(n_4856),
.Y(n_19555)
);

OAI21xp33_ASAP7_75t_SL g19556 ( 
.A1(n_19210),
.A2(n_8214),
.B(n_8441),
.Y(n_19556)
);

AOI211x1_ASAP7_75t_L g19557 ( 
.A1(n_19385),
.A2(n_19374),
.B(n_19258),
.C(n_19381),
.Y(n_19557)
);

XNOR2x1_ASAP7_75t_SL g19558 ( 
.A(n_19190),
.B(n_5106),
.Y(n_19558)
);

NOR3x1_ASAP7_75t_L g19559 ( 
.A(n_19315),
.B(n_8287),
.C(n_8286),
.Y(n_19559)
);

NAND2xp5_ASAP7_75t_L g19560 ( 
.A(n_19176),
.B(n_8388),
.Y(n_19560)
);

AOI21xp5_ASAP7_75t_L g19561 ( 
.A1(n_19378),
.A2(n_8396),
.B(n_8388),
.Y(n_19561)
);

AOI221xp5_ASAP7_75t_L g19562 ( 
.A1(n_19286),
.A2(n_8413),
.B1(n_8421),
.B2(n_8396),
.C(n_8388),
.Y(n_19562)
);

AOI21xp5_ASAP7_75t_L g19563 ( 
.A1(n_19333),
.A2(n_8413),
.B(n_8396),
.Y(n_19563)
);

AOI221xp5_ASAP7_75t_L g19564 ( 
.A1(n_19250),
.A2(n_8421),
.B1(n_8475),
.B2(n_8413),
.C(n_8396),
.Y(n_19564)
);

AOI211x1_ASAP7_75t_L g19565 ( 
.A1(n_19344),
.A2(n_8552),
.B(n_8885),
.C(n_8877),
.Y(n_19565)
);

AOI21xp5_ASAP7_75t_L g19566 ( 
.A1(n_19247),
.A2(n_8421),
.B(n_8413),
.Y(n_19566)
);

AND4x1_ASAP7_75t_L g19567 ( 
.A(n_19181),
.B(n_7812),
.C(n_7831),
.D(n_7900),
.Y(n_19567)
);

AOI21xp5_ASAP7_75t_L g19568 ( 
.A1(n_19383),
.A2(n_8475),
.B(n_8421),
.Y(n_19568)
);

NAND2xp5_ASAP7_75t_L g19569 ( 
.A(n_19193),
.B(n_8475),
.Y(n_19569)
);

INVx1_ASAP7_75t_L g19570 ( 
.A(n_19330),
.Y(n_19570)
);

AOI211x1_ASAP7_75t_L g19571 ( 
.A1(n_19334),
.A2(n_8905),
.B(n_8912),
.C(n_8885),
.Y(n_19571)
);

AOI211xp5_ASAP7_75t_L g19572 ( 
.A1(n_19261),
.A2(n_7460),
.B(n_7519),
.C(n_7457),
.Y(n_19572)
);

NOR2x1_ASAP7_75t_L g19573 ( 
.A(n_19264),
.B(n_7594),
.Y(n_19573)
);

OA22x2_ASAP7_75t_L g19574 ( 
.A1(n_19273),
.A2(n_8485),
.B1(n_8486),
.B2(n_8475),
.Y(n_19574)
);

NAND2xp5_ASAP7_75t_L g19575 ( 
.A(n_19339),
.B(n_8485),
.Y(n_19575)
);

NOR3x1_ASAP7_75t_L g19576 ( 
.A(n_19177),
.B(n_8287),
.C(n_8286),
.Y(n_19576)
);

OA22x2_ASAP7_75t_L g19577 ( 
.A1(n_19346),
.A2(n_8486),
.B1(n_8507),
.B2(n_8485),
.Y(n_19577)
);

AOI21xp5_ASAP7_75t_L g19578 ( 
.A1(n_19338),
.A2(n_8486),
.B(n_8485),
.Y(n_19578)
);

AOI22xp5_ASAP7_75t_L g19579 ( 
.A1(n_19280),
.A2(n_7460),
.B1(n_7519),
.B2(n_7457),
.Y(n_19579)
);

NOR2xp33_ASAP7_75t_L g19580 ( 
.A(n_19228),
.B(n_5524),
.Y(n_19580)
);

INVx1_ASAP7_75t_L g19581 ( 
.A(n_19407),
.Y(n_19581)
);

AOI211xp5_ASAP7_75t_L g19582 ( 
.A1(n_19401),
.A2(n_5414),
.B(n_5416),
.C(n_5382),
.Y(n_19582)
);

XNOR2xp5_ASAP7_75t_L g19583 ( 
.A(n_19471),
.B(n_7706),
.Y(n_19583)
);

O2A1O1Ixp33_ASAP7_75t_L g19584 ( 
.A1(n_19391),
.A2(n_19472),
.B(n_19474),
.C(n_19462),
.Y(n_19584)
);

AOI21xp5_ASAP7_75t_L g19585 ( 
.A1(n_19387),
.A2(n_8507),
.B(n_8486),
.Y(n_19585)
);

AOI21xp33_ASAP7_75t_L g19586 ( 
.A1(n_19490),
.A2(n_4890),
.B(n_4856),
.Y(n_19586)
);

OAI22xp5_ASAP7_75t_L g19587 ( 
.A1(n_19400),
.A2(n_8507),
.B1(n_8569),
.B2(n_8511),
.Y(n_19587)
);

AOI22xp5_ASAP7_75t_L g19588 ( 
.A1(n_19466),
.A2(n_8802),
.B1(n_7519),
.B2(n_7531),
.Y(n_19588)
);

O2A1O1Ixp33_ASAP7_75t_L g19589 ( 
.A1(n_19510),
.A2(n_5166),
.B(n_5219),
.C(n_5122),
.Y(n_19589)
);

INVx2_ASAP7_75t_SL g19590 ( 
.A(n_19418),
.Y(n_19590)
);

AOI21xp33_ASAP7_75t_L g19591 ( 
.A1(n_19423),
.A2(n_4890),
.B(n_4856),
.Y(n_19591)
);

NAND2xp5_ASAP7_75t_L g19592 ( 
.A(n_19418),
.B(n_8507),
.Y(n_19592)
);

OAI21xp5_ASAP7_75t_SL g19593 ( 
.A1(n_19469),
.A2(n_5416),
.B(n_5414),
.Y(n_19593)
);

OAI211xp5_ASAP7_75t_L g19594 ( 
.A1(n_19397),
.A2(n_8832),
.B(n_5301),
.C(n_5483),
.Y(n_19594)
);

INVx1_ASAP7_75t_L g19595 ( 
.A(n_19418),
.Y(n_19595)
);

AOI221xp5_ASAP7_75t_L g19596 ( 
.A1(n_19386),
.A2(n_19388),
.B1(n_19439),
.B2(n_19530),
.C(n_19535),
.Y(n_19596)
);

INVx1_ASAP7_75t_SL g19597 ( 
.A(n_19389),
.Y(n_19597)
);

AOI221xp5_ASAP7_75t_L g19598 ( 
.A1(n_19406),
.A2(n_8573),
.B1(n_8576),
.B2(n_8569),
.C(n_8511),
.Y(n_19598)
);

NAND2xp5_ASAP7_75t_L g19599 ( 
.A(n_19485),
.B(n_8511),
.Y(n_19599)
);

INVx1_ASAP7_75t_L g19600 ( 
.A(n_19485),
.Y(n_19600)
);

AOI22xp5_ASAP7_75t_L g19601 ( 
.A1(n_19447),
.A2(n_8802),
.B1(n_7519),
.B2(n_7531),
.Y(n_19601)
);

XNOR2x1_ASAP7_75t_L g19602 ( 
.A(n_19421),
.B(n_19396),
.Y(n_19602)
);

AOI21xp33_ASAP7_75t_SL g19603 ( 
.A1(n_19479),
.A2(n_5166),
.B(n_5122),
.Y(n_19603)
);

INVx2_ASAP7_75t_L g19604 ( 
.A(n_19485),
.Y(n_19604)
);

HB1xp67_ASAP7_75t_L g19605 ( 
.A(n_19392),
.Y(n_19605)
);

AOI21xp33_ASAP7_75t_SL g19606 ( 
.A1(n_19570),
.A2(n_5231),
.B(n_5219),
.Y(n_19606)
);

OAI221xp5_ASAP7_75t_L g19607 ( 
.A1(n_19538),
.A2(n_7612),
.B1(n_7743),
.B2(n_7742),
.C(n_7707),
.Y(n_19607)
);

AOI21xp5_ASAP7_75t_L g19608 ( 
.A1(n_19390),
.A2(n_8569),
.B(n_8511),
.Y(n_19608)
);

AOI31xp33_ASAP7_75t_L g19609 ( 
.A1(n_19408),
.A2(n_5231),
.A3(n_5240),
.B(n_5219),
.Y(n_19609)
);

INVx1_ASAP7_75t_L g19610 ( 
.A(n_19516),
.Y(n_19610)
);

AOI221xp5_ASAP7_75t_L g19611 ( 
.A1(n_19464),
.A2(n_8576),
.B1(n_8577),
.B2(n_8573),
.C(n_8569),
.Y(n_19611)
);

AOI21xp33_ASAP7_75t_L g19612 ( 
.A1(n_19473),
.A2(n_4890),
.B(n_4856),
.Y(n_19612)
);

AOI222xp33_ASAP7_75t_L g19613 ( 
.A1(n_19556),
.A2(n_8209),
.B1(n_8205),
.B2(n_8918),
.C1(n_8912),
.C2(n_8905),
.Y(n_19613)
);

NAND2xp5_ASAP7_75t_L g19614 ( 
.A(n_19509),
.B(n_8573),
.Y(n_19614)
);

OAI22xp33_ASAP7_75t_L g19615 ( 
.A1(n_19404),
.A2(n_7519),
.B1(n_7531),
.B2(n_7460),
.Y(n_19615)
);

OAI22xp5_ASAP7_75t_L g19616 ( 
.A1(n_19454),
.A2(n_8573),
.B1(n_8577),
.B2(n_8576),
.Y(n_19616)
);

AOI211xp5_ASAP7_75t_L g19617 ( 
.A1(n_19492),
.A2(n_5416),
.B(n_5424),
.C(n_5414),
.Y(n_19617)
);

INVx1_ASAP7_75t_L g19618 ( 
.A(n_19513),
.Y(n_19618)
);

INVx2_ASAP7_75t_L g19619 ( 
.A(n_19541),
.Y(n_19619)
);

OAI22xp33_ASAP7_75t_L g19620 ( 
.A1(n_19434),
.A2(n_7519),
.B1(n_7531),
.B2(n_7460),
.Y(n_19620)
);

AOI21xp33_ASAP7_75t_L g19621 ( 
.A1(n_19488),
.A2(n_5671),
.B(n_5287),
.Y(n_19621)
);

INVx1_ASAP7_75t_L g19622 ( 
.A(n_19558),
.Y(n_19622)
);

OAI211xp5_ASAP7_75t_L g19623 ( 
.A1(n_19557),
.A2(n_8832),
.B(n_5301),
.C(n_5483),
.Y(n_19623)
);

XNOR2xp5_ASAP7_75t_L g19624 ( 
.A(n_19419),
.B(n_7706),
.Y(n_19624)
);

INVxp67_ASAP7_75t_L g19625 ( 
.A(n_19429),
.Y(n_19625)
);

NAND2xp5_ASAP7_75t_SL g19626 ( 
.A(n_19573),
.B(n_7460),
.Y(n_19626)
);

OAI22xp5_ASAP7_75t_L g19627 ( 
.A1(n_19540),
.A2(n_19555),
.B1(n_19489),
.B2(n_19506),
.Y(n_19627)
);

A2O1A1Ixp33_ASAP7_75t_L g19628 ( 
.A1(n_19580),
.A2(n_8448),
.B(n_8451),
.C(n_8441),
.Y(n_19628)
);

OAI21xp33_ASAP7_75t_L g19629 ( 
.A1(n_19415),
.A2(n_7707),
.B(n_7612),
.Y(n_19629)
);

AOI22xp33_ASAP7_75t_SL g19630 ( 
.A1(n_19501),
.A2(n_7531),
.B1(n_7544),
.B2(n_7519),
.Y(n_19630)
);

AOI322xp5_ASAP7_75t_L g19631 ( 
.A1(n_19424),
.A2(n_7178),
.A3(n_7115),
.B1(n_7356),
.B2(n_7464),
.C1(n_7339),
.C2(n_7220),
.Y(n_19631)
);

NAND2xp33_ASAP7_75t_SL g19632 ( 
.A(n_19426),
.B(n_5414),
.Y(n_19632)
);

OAI22xp5_ASAP7_75t_SL g19633 ( 
.A1(n_19512),
.A2(n_6783),
.B1(n_6858),
.B2(n_6706),
.Y(n_19633)
);

O2A1O1Ixp33_ASAP7_75t_L g19634 ( 
.A1(n_19417),
.A2(n_5240),
.B(n_5310),
.C(n_5231),
.Y(n_19634)
);

AOI221xp5_ASAP7_75t_L g19635 ( 
.A1(n_19440),
.A2(n_8578),
.B1(n_8580),
.B2(n_8577),
.C(n_8576),
.Y(n_19635)
);

AOI22xp5_ASAP7_75t_L g19636 ( 
.A1(n_19519),
.A2(n_19451),
.B1(n_19504),
.B2(n_19531),
.Y(n_19636)
);

AOI221xp5_ASAP7_75t_L g19637 ( 
.A1(n_19427),
.A2(n_8580),
.B1(n_8620),
.B2(n_8578),
.C(n_8577),
.Y(n_19637)
);

OAI21xp33_ASAP7_75t_L g19638 ( 
.A1(n_19503),
.A2(n_7707),
.B(n_7612),
.Y(n_19638)
);

AOI322xp5_ASAP7_75t_L g19639 ( 
.A1(n_19550),
.A2(n_7178),
.A3(n_7115),
.B1(n_7475),
.B2(n_7566),
.C1(n_7464),
.C2(n_7220),
.Y(n_19639)
);

OAI21xp33_ASAP7_75t_L g19640 ( 
.A1(n_19548),
.A2(n_19507),
.B(n_19520),
.Y(n_19640)
);

INVx2_ASAP7_75t_L g19641 ( 
.A(n_19541),
.Y(n_19641)
);

AOI21xp5_ASAP7_75t_L g19642 ( 
.A1(n_19435),
.A2(n_19524),
.B(n_19437),
.Y(n_19642)
);

AOI21xp5_ASAP7_75t_L g19643 ( 
.A1(n_19494),
.A2(n_8580),
.B(n_8578),
.Y(n_19643)
);

OAI22xp33_ASAP7_75t_L g19644 ( 
.A1(n_19542),
.A2(n_7531),
.B1(n_7544),
.B2(n_7519),
.Y(n_19644)
);

INVx1_ASAP7_75t_L g19645 ( 
.A(n_19394),
.Y(n_19645)
);

INVx1_ASAP7_75t_SL g19646 ( 
.A(n_19405),
.Y(n_19646)
);

INVx1_ASAP7_75t_L g19647 ( 
.A(n_19403),
.Y(n_19647)
);

INVx1_ASAP7_75t_L g19648 ( 
.A(n_19410),
.Y(n_19648)
);

INVx1_ASAP7_75t_L g19649 ( 
.A(n_19411),
.Y(n_19649)
);

HB1xp67_ASAP7_75t_L g19650 ( 
.A(n_19478),
.Y(n_19650)
);

AOI22xp5_ASAP7_75t_L g19651 ( 
.A1(n_19552),
.A2(n_8802),
.B1(n_7544),
.B2(n_7599),
.Y(n_19651)
);

AOI222xp33_ASAP7_75t_L g19652 ( 
.A1(n_19413),
.A2(n_8209),
.B1(n_8205),
.B2(n_8918),
.C1(n_8912),
.C2(n_8905),
.Y(n_19652)
);

AOI211xp5_ASAP7_75t_L g19653 ( 
.A1(n_19543),
.A2(n_5416),
.B(n_5424),
.C(n_5414),
.Y(n_19653)
);

NAND3xp33_ASAP7_75t_L g19654 ( 
.A(n_19549),
.B(n_5671),
.C(n_5287),
.Y(n_19654)
);

AOI21xp33_ASAP7_75t_L g19655 ( 
.A1(n_19468),
.A2(n_5671),
.B(n_5287),
.Y(n_19655)
);

OAI21x1_ASAP7_75t_L g19656 ( 
.A1(n_19574),
.A2(n_9239),
.B(n_9097),
.Y(n_19656)
);

OAI21xp33_ASAP7_75t_L g19657 ( 
.A1(n_19470),
.A2(n_19463),
.B(n_19398),
.Y(n_19657)
);

INVxp67_ASAP7_75t_SL g19658 ( 
.A(n_19428),
.Y(n_19658)
);

AOI22xp33_ASAP7_75t_SL g19659 ( 
.A1(n_19446),
.A2(n_7544),
.B1(n_7599),
.B2(n_7531),
.Y(n_19659)
);

AOI21xp5_ASAP7_75t_L g19660 ( 
.A1(n_19486),
.A2(n_8580),
.B(n_8578),
.Y(n_19660)
);

OAI211xp5_ASAP7_75t_SL g19661 ( 
.A1(n_19430),
.A2(n_5310),
.B(n_5342),
.C(n_5240),
.Y(n_19661)
);

OAI22xp33_ASAP7_75t_L g19662 ( 
.A1(n_19414),
.A2(n_7544),
.B1(n_7599),
.B2(n_7531),
.Y(n_19662)
);

AOI21xp33_ASAP7_75t_SL g19663 ( 
.A1(n_19431),
.A2(n_5342),
.B(n_5310),
.Y(n_19663)
);

OAI21xp5_ASAP7_75t_L g19664 ( 
.A1(n_19523),
.A2(n_7907),
.B(n_7920),
.Y(n_19664)
);

OAI22xp5_ASAP7_75t_SL g19665 ( 
.A1(n_19483),
.A2(n_6858),
.B1(n_6783),
.B2(n_8588),
.Y(n_19665)
);

NAND2xp5_ASAP7_75t_L g19666 ( 
.A(n_19545),
.B(n_8620),
.Y(n_19666)
);

OAI22xp33_ASAP7_75t_SL g19667 ( 
.A1(n_19502),
.A2(n_7487),
.B1(n_7649),
.B2(n_7522),
.Y(n_19667)
);

INVx1_ASAP7_75t_L g19668 ( 
.A(n_19522),
.Y(n_19668)
);

AOI22xp33_ASAP7_75t_L g19669 ( 
.A1(n_19452),
.A2(n_7544),
.B1(n_7599),
.B2(n_7531),
.Y(n_19669)
);

AOI22xp5_ASAP7_75t_L g19670 ( 
.A1(n_19553),
.A2(n_19412),
.B1(n_19515),
.B2(n_19511),
.Y(n_19670)
);

AOI221x1_ASAP7_75t_L g19671 ( 
.A1(n_19546),
.A2(n_8936),
.B1(n_8945),
.B2(n_8920),
.C(n_8918),
.Y(n_19671)
);

OAI21xp5_ASAP7_75t_L g19672 ( 
.A1(n_19477),
.A2(n_7907),
.B(n_7920),
.Y(n_19672)
);

INVx1_ASAP7_75t_L g19673 ( 
.A(n_19528),
.Y(n_19673)
);

NAND3xp33_ASAP7_75t_L g19674 ( 
.A(n_19572),
.B(n_5671),
.C(n_5287),
.Y(n_19674)
);

OAI21xp5_ASAP7_75t_L g19675 ( 
.A1(n_19441),
.A2(n_7932),
.B(n_7920),
.Y(n_19675)
);

INVx1_ASAP7_75t_SL g19676 ( 
.A(n_19491),
.Y(n_19676)
);

NOR4xp25_ASAP7_75t_L g19677 ( 
.A(n_19560),
.B(n_8936),
.C(n_8945),
.D(n_8920),
.Y(n_19677)
);

INVx2_ASAP7_75t_SL g19678 ( 
.A(n_19577),
.Y(n_19678)
);

NAND2xp5_ASAP7_75t_L g19679 ( 
.A(n_19449),
.B(n_8620),
.Y(n_19679)
);

INVx2_ASAP7_75t_SL g19680 ( 
.A(n_19546),
.Y(n_19680)
);

OAI21xp5_ASAP7_75t_L g19681 ( 
.A1(n_19425),
.A2(n_7932),
.B(n_7920),
.Y(n_19681)
);

OAI221xp5_ASAP7_75t_L g19682 ( 
.A1(n_19575),
.A2(n_7612),
.B1(n_7743),
.B2(n_7742),
.C(n_7707),
.Y(n_19682)
);

OAI211xp5_ASAP7_75t_SL g19683 ( 
.A1(n_19527),
.A2(n_5396),
.B(n_5464),
.C(n_5342),
.Y(n_19683)
);

O2A1O1Ixp33_ASAP7_75t_L g19684 ( 
.A1(n_19480),
.A2(n_5464),
.B(n_5503),
.C(n_5396),
.Y(n_19684)
);

OAI21xp33_ASAP7_75t_L g19685 ( 
.A1(n_19438),
.A2(n_7743),
.B(n_7742),
.Y(n_19685)
);

AOI21xp33_ASAP7_75t_L g19686 ( 
.A1(n_19484),
.A2(n_5671),
.B(n_5287),
.Y(n_19686)
);

OAI21xp5_ASAP7_75t_SL g19687 ( 
.A1(n_19539),
.A2(n_19567),
.B(n_19409),
.Y(n_19687)
);

NOR2xp33_ASAP7_75t_L g19688 ( 
.A(n_19521),
.B(n_5524),
.Y(n_19688)
);

AOI21xp5_ASAP7_75t_L g19689 ( 
.A1(n_19569),
.A2(n_8640),
.B(n_8620),
.Y(n_19689)
);

INVx1_ASAP7_75t_L g19690 ( 
.A(n_19393),
.Y(n_19690)
);

AOI211x1_ASAP7_75t_L g19691 ( 
.A1(n_19578),
.A2(n_8936),
.B(n_8945),
.C(n_8920),
.Y(n_19691)
);

INVxp67_ASAP7_75t_L g19692 ( 
.A(n_19526),
.Y(n_19692)
);

AOI21xp33_ASAP7_75t_L g19693 ( 
.A1(n_19500),
.A2(n_5671),
.B(n_8640),
.Y(n_19693)
);

AOI222xp33_ASAP7_75t_L g19694 ( 
.A1(n_19544),
.A2(n_8981),
.B1(n_8995),
.B2(n_9003),
.C1(n_8996),
.C2(n_8954),
.Y(n_19694)
);

INVxp67_ASAP7_75t_L g19695 ( 
.A(n_19554),
.Y(n_19695)
);

OA22x2_ASAP7_75t_L g19696 ( 
.A1(n_19525),
.A2(n_8640),
.B1(n_8660),
.B2(n_8658),
.Y(n_19696)
);

OAI221xp5_ASAP7_75t_SL g19697 ( 
.A1(n_19533),
.A2(n_7906),
.B1(n_7890),
.B2(n_7839),
.C(n_7684),
.Y(n_19697)
);

AOI22xp5_ASAP7_75t_L g19698 ( 
.A1(n_19458),
.A2(n_8802),
.B1(n_7544),
.B2(n_7599),
.Y(n_19698)
);

INVx2_ASAP7_75t_L g19699 ( 
.A(n_19461),
.Y(n_19699)
);

NOR2xp67_ASAP7_75t_SL g19700 ( 
.A(n_19536),
.B(n_5414),
.Y(n_19700)
);

OAI321xp33_ASAP7_75t_L g19701 ( 
.A1(n_19505),
.A2(n_7625),
.A3(n_7544),
.B1(n_7711),
.B2(n_7599),
.C(n_7531),
.Y(n_19701)
);

INVx1_ASAP7_75t_SL g19702 ( 
.A(n_19442),
.Y(n_19702)
);

OAI32xp33_ASAP7_75t_L g19703 ( 
.A1(n_19395),
.A2(n_8640),
.A3(n_8663),
.B1(n_8660),
.B2(n_8658),
.Y(n_19703)
);

INVx1_ASAP7_75t_L g19704 ( 
.A(n_19565),
.Y(n_19704)
);

NOR2xp67_ASAP7_75t_L g19705 ( 
.A(n_19487),
.B(n_5195),
.Y(n_19705)
);

INVx1_ASAP7_75t_L g19706 ( 
.A(n_19576),
.Y(n_19706)
);

NOR2xp33_ASAP7_75t_R g19707 ( 
.A(n_19416),
.B(n_5414),
.Y(n_19707)
);

INVx1_ASAP7_75t_L g19708 ( 
.A(n_19453),
.Y(n_19708)
);

XOR2x2_ASAP7_75t_L g19709 ( 
.A(n_19432),
.B(n_7742),
.Y(n_19709)
);

HB1xp67_ASAP7_75t_L g19710 ( 
.A(n_19559),
.Y(n_19710)
);

INVx1_ASAP7_75t_L g19711 ( 
.A(n_19571),
.Y(n_19711)
);

INVx1_ASAP7_75t_L g19712 ( 
.A(n_19450),
.Y(n_19712)
);

OAI221xp5_ASAP7_75t_L g19713 ( 
.A1(n_19433),
.A2(n_7743),
.B1(n_7649),
.B2(n_7705),
.C(n_7522),
.Y(n_19713)
);

CKINVDCx5p33_ASAP7_75t_R g19714 ( 
.A(n_19399),
.Y(n_19714)
);

INVx2_ASAP7_75t_L g19715 ( 
.A(n_19450),
.Y(n_19715)
);

INVx1_ASAP7_75t_L g19716 ( 
.A(n_19436),
.Y(n_19716)
);

OAI211xp5_ASAP7_75t_L g19717 ( 
.A1(n_19422),
.A2(n_5483),
.B(n_5485),
.C(n_5301),
.Y(n_19717)
);

OAI21xp5_ASAP7_75t_L g19718 ( 
.A1(n_19579),
.A2(n_7932),
.B(n_8000),
.Y(n_19718)
);

XNOR2xp5_ASAP7_75t_L g19719 ( 
.A(n_19444),
.B(n_7706),
.Y(n_19719)
);

A2O1A1Ixp33_ASAP7_75t_L g19720 ( 
.A1(n_19547),
.A2(n_8448),
.B(n_8451),
.C(n_8441),
.Y(n_19720)
);

AOI21xp33_ASAP7_75t_SL g19721 ( 
.A1(n_19499),
.A2(n_5464),
.B(n_5396),
.Y(n_19721)
);

O2A1O1Ixp5_ASAP7_75t_L g19722 ( 
.A1(n_19518),
.A2(n_19561),
.B(n_19563),
.C(n_19566),
.Y(n_19722)
);

AOI22xp5_ASAP7_75t_L g19723 ( 
.A1(n_19436),
.A2(n_8802),
.B1(n_7599),
.B2(n_7625),
.Y(n_19723)
);

XNOR2x2_ASAP7_75t_L g19724 ( 
.A(n_19420),
.B(n_7932),
.Y(n_19724)
);

INVx1_ASAP7_75t_L g19725 ( 
.A(n_19534),
.Y(n_19725)
);

NAND2xp5_ASAP7_75t_L g19726 ( 
.A(n_19532),
.B(n_8658),
.Y(n_19726)
);

OAI22xp5_ASAP7_75t_L g19727 ( 
.A1(n_19465),
.A2(n_8660),
.B1(n_8663),
.B2(n_8658),
.Y(n_19727)
);

NAND3x1_ASAP7_75t_L g19728 ( 
.A(n_19568),
.B(n_8981),
.C(n_8954),
.Y(n_19728)
);

AOI21xp5_ASAP7_75t_L g19729 ( 
.A1(n_19495),
.A2(n_8663),
.B(n_8660),
.Y(n_19729)
);

OAI21xp33_ASAP7_75t_L g19730 ( 
.A1(n_19551),
.A2(n_5831),
.B(n_5804),
.Y(n_19730)
);

OAI221xp5_ASAP7_75t_L g19731 ( 
.A1(n_19459),
.A2(n_7649),
.B1(n_7705),
.B2(n_7522),
.C(n_7487),
.Y(n_19731)
);

INVxp67_ASAP7_75t_L g19732 ( 
.A(n_19496),
.Y(n_19732)
);

INVx2_ASAP7_75t_SL g19733 ( 
.A(n_19517),
.Y(n_19733)
);

INVx2_ASAP7_75t_L g19734 ( 
.A(n_19517),
.Y(n_19734)
);

AOI21xp33_ASAP7_75t_SL g19735 ( 
.A1(n_19460),
.A2(n_5634),
.B(n_5503),
.Y(n_19735)
);

NAND2xp5_ASAP7_75t_L g19736 ( 
.A(n_19497),
.B(n_8663),
.Y(n_19736)
);

OAI22xp33_ASAP7_75t_L g19737 ( 
.A1(n_19445),
.A2(n_7599),
.B1(n_7625),
.B2(n_7544),
.Y(n_19737)
);

NOR2xp67_ASAP7_75t_L g19738 ( 
.A(n_19456),
.B(n_5301),
.Y(n_19738)
);

NOR2xp67_ASAP7_75t_L g19739 ( 
.A(n_19443),
.B(n_5301),
.Y(n_19739)
);

INVx1_ASAP7_75t_L g19740 ( 
.A(n_19457),
.Y(n_19740)
);

NOR2xp33_ASAP7_75t_L g19741 ( 
.A(n_19493),
.B(n_5524),
.Y(n_19741)
);

NAND2xp5_ASAP7_75t_L g19742 ( 
.A(n_19482),
.B(n_8670),
.Y(n_19742)
);

XOR2x2_ASAP7_75t_L g19743 ( 
.A(n_19564),
.B(n_5719),
.Y(n_19743)
);

AND2x2_ASAP7_75t_L g19744 ( 
.A(n_19498),
.B(n_7198),
.Y(n_19744)
);

NAND4xp25_ASAP7_75t_SL g19745 ( 
.A(n_19584),
.B(n_19596),
.C(n_19597),
.D(n_19610),
.Y(n_19745)
);

OAI211xp5_ASAP7_75t_L g19746 ( 
.A1(n_19640),
.A2(n_19448),
.B(n_19529),
.C(n_19476),
.Y(n_19746)
);

OAI22xp33_ASAP7_75t_L g19747 ( 
.A1(n_19590),
.A2(n_19402),
.B1(n_19508),
.B2(n_19467),
.Y(n_19747)
);

AOI221xp5_ASAP7_75t_L g19748 ( 
.A1(n_19606),
.A2(n_19537),
.B1(n_19562),
.B2(n_19514),
.C(n_19475),
.Y(n_19748)
);

NAND3xp33_ASAP7_75t_L g19749 ( 
.A(n_19605),
.B(n_19455),
.C(n_19481),
.Y(n_19749)
);

NAND4xp25_ASAP7_75t_L g19750 ( 
.A(n_19595),
.B(n_19618),
.C(n_19625),
.D(n_19702),
.Y(n_19750)
);

O2A1O1Ixp33_ASAP7_75t_L g19751 ( 
.A1(n_19600),
.A2(n_5634),
.B(n_5637),
.C(n_5503),
.Y(n_19751)
);

NOR2xp33_ASAP7_75t_SL g19752 ( 
.A(n_19604),
.B(n_5301),
.Y(n_19752)
);

OAI221xp5_ASAP7_75t_L g19753 ( 
.A1(n_19687),
.A2(n_7649),
.B1(n_7705),
.B2(n_7522),
.C(n_7487),
.Y(n_19753)
);

INVxp67_ASAP7_75t_L g19754 ( 
.A(n_19710),
.Y(n_19754)
);

AOI221xp5_ASAP7_75t_L g19755 ( 
.A1(n_19627),
.A2(n_8995),
.B1(n_8996),
.B2(n_8981),
.C(n_8954),
.Y(n_19755)
);

AOI311xp33_ASAP7_75t_L g19756 ( 
.A1(n_19690),
.A2(n_8996),
.A3(n_9028),
.B(n_9003),
.C(n_8995),
.Y(n_19756)
);

AOI221xp5_ASAP7_75t_L g19757 ( 
.A1(n_19704),
.A2(n_9036),
.B1(n_9045),
.B2(n_9028),
.C(n_9003),
.Y(n_19757)
);

AOI211xp5_ASAP7_75t_L g19758 ( 
.A1(n_19706),
.A2(n_5424),
.B(n_5440),
.C(n_5416),
.Y(n_19758)
);

INVx1_ASAP7_75t_SL g19759 ( 
.A(n_19602),
.Y(n_19759)
);

AOI211xp5_ASAP7_75t_L g19760 ( 
.A1(n_19642),
.A2(n_5424),
.B(n_5440),
.C(n_5416),
.Y(n_19760)
);

INVx1_ASAP7_75t_L g19761 ( 
.A(n_19624),
.Y(n_19761)
);

OAI221xp5_ASAP7_75t_L g19762 ( 
.A1(n_19622),
.A2(n_7649),
.B1(n_7705),
.B2(n_7522),
.C(n_7487),
.Y(n_19762)
);

AOI22xp5_ASAP7_75t_L g19763 ( 
.A1(n_19583),
.A2(n_8802),
.B1(n_8019),
.B2(n_7599),
.Y(n_19763)
);

AOI22xp5_ASAP7_75t_L g19764 ( 
.A1(n_19714),
.A2(n_8019),
.B1(n_7599),
.B2(n_7625),
.Y(n_19764)
);

AOI211xp5_ASAP7_75t_L g19765 ( 
.A1(n_19708),
.A2(n_5424),
.B(n_5440),
.C(n_5416),
.Y(n_19765)
);

AOI22xp5_ASAP7_75t_L g19766 ( 
.A1(n_19633),
.A2(n_8019),
.B1(n_7625),
.B2(n_7711),
.Y(n_19766)
);

AND4x2_ASAP7_75t_L g19767 ( 
.A(n_19608),
.B(n_7095),
.C(n_8013),
.D(n_8704),
.Y(n_19767)
);

INVx1_ASAP7_75t_L g19768 ( 
.A(n_19592),
.Y(n_19768)
);

AOI211xp5_ASAP7_75t_L g19769 ( 
.A1(n_19725),
.A2(n_19581),
.B(n_19676),
.C(n_19657),
.Y(n_19769)
);

INVx1_ASAP7_75t_L g19770 ( 
.A(n_19599),
.Y(n_19770)
);

INVx2_ASAP7_75t_SL g19771 ( 
.A(n_19626),
.Y(n_19771)
);

A2O1A1Ixp33_ASAP7_75t_L g19772 ( 
.A1(n_19722),
.A2(n_9036),
.B(n_9045),
.C(n_9028),
.Y(n_19772)
);

OAI22xp33_ASAP7_75t_L g19773 ( 
.A1(n_19699),
.A2(n_7625),
.B1(n_7711),
.B2(n_7544),
.Y(n_19773)
);

INVx2_ASAP7_75t_L g19774 ( 
.A(n_19709),
.Y(n_19774)
);

AOI222xp33_ASAP7_75t_L g19775 ( 
.A1(n_19740),
.A2(n_9045),
.B1(n_9046),
.B2(n_9070),
.C1(n_9066),
.C2(n_9036),
.Y(n_19775)
);

INVx1_ASAP7_75t_L g19776 ( 
.A(n_19680),
.Y(n_19776)
);

INVx1_ASAP7_75t_L g19777 ( 
.A(n_19619),
.Y(n_19777)
);

AOI22xp5_ASAP7_75t_L g19778 ( 
.A1(n_19654),
.A2(n_8019),
.B1(n_7711),
.B2(n_7719),
.Y(n_19778)
);

AOI21xp33_ASAP7_75t_L g19779 ( 
.A1(n_19646),
.A2(n_8673),
.B(n_8670),
.Y(n_19779)
);

XNOR2xp5_ASAP7_75t_L g19780 ( 
.A(n_19636),
.B(n_5719),
.Y(n_19780)
);

NOR2x1_ASAP7_75t_L g19781 ( 
.A(n_19673),
.B(n_5719),
.Y(n_19781)
);

AOI221xp5_ASAP7_75t_L g19782 ( 
.A1(n_19591),
.A2(n_9070),
.B1(n_9073),
.B2(n_9066),
.C(n_9046),
.Y(n_19782)
);

NOR2xp33_ASAP7_75t_L g19783 ( 
.A(n_19692),
.B(n_5524),
.Y(n_19783)
);

OAI211xp5_ASAP7_75t_L g19784 ( 
.A1(n_19695),
.A2(n_5485),
.B(n_5492),
.C(n_5483),
.Y(n_19784)
);

O2A1O1Ixp5_ASAP7_75t_L g19785 ( 
.A1(n_19641),
.A2(n_8670),
.B(n_8678),
.C(n_8673),
.Y(n_19785)
);

AOI221xp5_ASAP7_75t_L g19786 ( 
.A1(n_19678),
.A2(n_9070),
.B1(n_9073),
.B2(n_9066),
.C(n_9046),
.Y(n_19786)
);

NAND2xp5_ASAP7_75t_L g19787 ( 
.A(n_19744),
.B(n_8670),
.Y(n_19787)
);

OAI321xp33_ASAP7_75t_L g19788 ( 
.A1(n_19711),
.A2(n_7725),
.A3(n_7711),
.B1(n_7736),
.B2(n_7719),
.C(n_7625),
.Y(n_19788)
);

NOR2xp33_ASAP7_75t_L g19789 ( 
.A(n_19650),
.B(n_5601),
.Y(n_19789)
);

NAND4xp25_ASAP7_75t_L g19790 ( 
.A(n_19670),
.B(n_5726),
.C(n_5736),
.D(n_5719),
.Y(n_19790)
);

AOI221xp5_ASAP7_75t_L g19791 ( 
.A1(n_19737),
.A2(n_9085),
.B1(n_9090),
.B2(n_9079),
.C(n_9073),
.Y(n_19791)
);

BUFx2_ASAP7_75t_L g19792 ( 
.A(n_19707),
.Y(n_19792)
);

AOI211xp5_ASAP7_75t_L g19793 ( 
.A1(n_19647),
.A2(n_5424),
.B(n_5440),
.C(n_5416),
.Y(n_19793)
);

INVx2_ASAP7_75t_SL g19794 ( 
.A(n_19743),
.Y(n_19794)
);

NAND4xp25_ASAP7_75t_L g19795 ( 
.A(n_19582),
.B(n_5736),
.C(n_5726),
.D(n_5485),
.Y(n_19795)
);

AOI22xp5_ASAP7_75t_L g19796 ( 
.A1(n_19685),
.A2(n_8019),
.B1(n_7711),
.B2(n_7719),
.Y(n_19796)
);

AOI21xp5_ASAP7_75t_L g19797 ( 
.A1(n_19732),
.A2(n_8678),
.B(n_8673),
.Y(n_19797)
);

INVx1_ASAP7_75t_L g19798 ( 
.A(n_19716),
.Y(n_19798)
);

NOR3xp33_ASAP7_75t_L g19799 ( 
.A(n_19658),
.B(n_5485),
.C(n_5483),
.Y(n_19799)
);

O2A1O1Ixp33_ASAP7_75t_L g19800 ( 
.A1(n_19733),
.A2(n_5637),
.B(n_5644),
.C(n_5634),
.Y(n_19800)
);

AOI211xp5_ASAP7_75t_L g19801 ( 
.A1(n_19648),
.A2(n_5440),
.B(n_5445),
.C(n_5424),
.Y(n_19801)
);

AOI211xp5_ASAP7_75t_L g19802 ( 
.A1(n_19649),
.A2(n_5440),
.B(n_5445),
.C(n_5424),
.Y(n_19802)
);

AOI211xp5_ASAP7_75t_SL g19803 ( 
.A1(n_19668),
.A2(n_5725),
.B(n_5589),
.C(n_5393),
.Y(n_19803)
);

O2A1O1Ixp33_ASAP7_75t_L g19804 ( 
.A1(n_19645),
.A2(n_5644),
.B(n_5687),
.C(n_5637),
.Y(n_19804)
);

AOI22xp33_ASAP7_75t_L g19805 ( 
.A1(n_19674),
.A2(n_7711),
.B1(n_7719),
.B2(n_7625),
.Y(n_19805)
);

NAND3xp33_ASAP7_75t_L g19806 ( 
.A(n_19712),
.B(n_5886),
.C(n_5440),
.Y(n_19806)
);

NOR4xp25_ASAP7_75t_L g19807 ( 
.A(n_19715),
.B(n_19734),
.C(n_19614),
.D(n_19684),
.Y(n_19807)
);

AOI221x1_ASAP7_75t_L g19808 ( 
.A1(n_19632),
.A2(n_19667),
.B1(n_19721),
.B2(n_19612),
.C(n_19586),
.Y(n_19808)
);

NOR4xp75_ASAP7_75t_L g19809 ( 
.A(n_19728),
.B(n_5687),
.C(n_5720),
.D(n_5644),
.Y(n_19809)
);

XOR2xp5_ASAP7_75t_L g19810 ( 
.A(n_19719),
.B(n_19696),
.Y(n_19810)
);

AOI211xp5_ASAP7_75t_L g19811 ( 
.A1(n_19621),
.A2(n_5440),
.B(n_5445),
.C(n_5424),
.Y(n_19811)
);

AOI221xp5_ASAP7_75t_L g19812 ( 
.A1(n_19693),
.A2(n_9090),
.B1(n_9091),
.B2(n_9085),
.C(n_9079),
.Y(n_19812)
);

AOI222xp33_ASAP7_75t_L g19813 ( 
.A1(n_19705),
.A2(n_9085),
.B1(n_9090),
.B2(n_9104),
.C1(n_9091),
.C2(n_9079),
.Y(n_19813)
);

NAND3xp33_ASAP7_75t_SL g19814 ( 
.A(n_19613),
.B(n_5485),
.C(n_5483),
.Y(n_19814)
);

OAI211xp5_ASAP7_75t_L g19815 ( 
.A1(n_19593),
.A2(n_5492),
.B(n_5513),
.C(n_5485),
.Y(n_19815)
);

AOI211xp5_ASAP7_75t_SL g19816 ( 
.A1(n_19739),
.A2(n_5725),
.B(n_5589),
.C(n_5393),
.Y(n_19816)
);

INVx1_ASAP7_75t_L g19817 ( 
.A(n_19738),
.Y(n_19817)
);

OAI21xp33_ASAP7_75t_L g19818 ( 
.A1(n_19629),
.A2(n_5831),
.B(n_5804),
.Y(n_19818)
);

O2A1O1Ixp33_ASAP7_75t_L g19819 ( 
.A1(n_19666),
.A2(n_5720),
.B(n_5687),
.C(n_5726),
.Y(n_19819)
);

INVxp67_ASAP7_75t_L g19820 ( 
.A(n_19688),
.Y(n_19820)
);

OR2x2_ASAP7_75t_L g19821 ( 
.A(n_19679),
.B(n_8704),
.Y(n_19821)
);

NAND2xp5_ASAP7_75t_L g19822 ( 
.A(n_19741),
.B(n_8673),
.Y(n_19822)
);

AOI211xp5_ASAP7_75t_L g19823 ( 
.A1(n_19655),
.A2(n_5445),
.B(n_5446),
.C(n_5440),
.Y(n_19823)
);

NAND4xp25_ASAP7_75t_L g19824 ( 
.A(n_19694),
.B(n_5736),
.C(n_5726),
.D(n_5513),
.Y(n_19824)
);

AOI32xp33_ASAP7_75t_L g19825 ( 
.A1(n_19683),
.A2(n_19730),
.A3(n_19644),
.B1(n_19620),
.B2(n_19662),
.Y(n_19825)
);

AOI221xp5_ASAP7_75t_SL g19826 ( 
.A1(n_19735),
.A2(n_9106),
.B1(n_9107),
.B2(n_9104),
.C(n_9091),
.Y(n_19826)
);

AOI221xp5_ASAP7_75t_L g19827 ( 
.A1(n_19700),
.A2(n_9107),
.B1(n_9108),
.B2(n_9106),
.C(n_9104),
.Y(n_19827)
);

HB1xp67_ASAP7_75t_L g19828 ( 
.A(n_19736),
.Y(n_19828)
);

AOI22xp5_ASAP7_75t_L g19829 ( 
.A1(n_19638),
.A2(n_8019),
.B1(n_7711),
.B2(n_7725),
.Y(n_19829)
);

AOI221xp5_ASAP7_75t_L g19830 ( 
.A1(n_19603),
.A2(n_9108),
.B1(n_9120),
.B2(n_9107),
.C(n_9106),
.Y(n_19830)
);

OAI21xp5_ASAP7_75t_SL g19831 ( 
.A1(n_19589),
.A2(n_5446),
.B(n_5445),
.Y(n_19831)
);

AOI222xp33_ASAP7_75t_L g19832 ( 
.A1(n_19664),
.A2(n_9120),
.B1(n_9124),
.B2(n_9136),
.C1(n_9128),
.C2(n_9108),
.Y(n_19832)
);

OAI21xp5_ASAP7_75t_L g19833 ( 
.A1(n_19585),
.A2(n_8531),
.B(n_8291),
.Y(n_19833)
);

INVx1_ASAP7_75t_L g19834 ( 
.A(n_19726),
.Y(n_19834)
);

OAI221xp5_ASAP7_75t_L g19835 ( 
.A1(n_19659),
.A2(n_7649),
.B1(n_7705),
.B2(n_7522),
.C(n_7487),
.Y(n_19835)
);

INVx1_ASAP7_75t_SL g19836 ( 
.A(n_19742),
.Y(n_19836)
);

NAND2xp5_ASAP7_75t_L g19837 ( 
.A(n_19677),
.B(n_8679),
.Y(n_19837)
);

NAND3x1_ASAP7_75t_L g19838 ( 
.A(n_19643),
.B(n_9124),
.C(n_9120),
.Y(n_19838)
);

INVx1_ASAP7_75t_L g19839 ( 
.A(n_19691),
.Y(n_19839)
);

AOI211x1_ASAP7_75t_SL g19840 ( 
.A1(n_19661),
.A2(n_8679),
.B(n_8701),
.C(n_8678),
.Y(n_19840)
);

AOI221xp5_ASAP7_75t_L g19841 ( 
.A1(n_19663),
.A2(n_9136),
.B1(n_9137),
.B2(n_9128),
.C(n_9124),
.Y(n_19841)
);

INVx1_ASAP7_75t_L g19842 ( 
.A(n_19671),
.Y(n_19842)
);

AOI211xp5_ASAP7_75t_L g19843 ( 
.A1(n_19697),
.A2(n_5446),
.B(n_5447),
.C(n_5445),
.Y(n_19843)
);

AOI211xp5_ASAP7_75t_L g19844 ( 
.A1(n_19717),
.A2(n_5446),
.B(n_5447),
.C(n_5445),
.Y(n_19844)
);

INVx2_ASAP7_75t_L g19845 ( 
.A(n_19724),
.Y(n_19845)
);

AOI211xp5_ASAP7_75t_SL g19846 ( 
.A1(n_19609),
.A2(n_5725),
.B(n_5589),
.C(n_5393),
.Y(n_19846)
);

A2O1A1Ixp33_ASAP7_75t_L g19847 ( 
.A1(n_19634),
.A2(n_9136),
.B(n_9137),
.C(n_9128),
.Y(n_19847)
);

AOI21xp5_ASAP7_75t_L g19848 ( 
.A1(n_19713),
.A2(n_8679),
.B(n_8678),
.Y(n_19848)
);

NOR3xp33_ASAP7_75t_L g19849 ( 
.A(n_19682),
.B(n_5513),
.C(n_5492),
.Y(n_19849)
);

NAND4xp75_ASAP7_75t_L g19850 ( 
.A(n_19686),
.B(n_8588),
.C(n_5720),
.D(n_9051),
.Y(n_19850)
);

A2O1A1Ixp33_ASAP7_75t_L g19851 ( 
.A1(n_19617),
.A2(n_9141),
.B(n_9143),
.C(n_9137),
.Y(n_19851)
);

AOI21xp5_ASAP7_75t_L g19852 ( 
.A1(n_19701),
.A2(n_8701),
.B(n_8679),
.Y(n_19852)
);

OAI221xp5_ASAP7_75t_L g19853 ( 
.A1(n_19630),
.A2(n_7649),
.B1(n_7705),
.B2(n_7522),
.C(n_7487),
.Y(n_19853)
);

O2A1O1Ixp33_ASAP7_75t_L g19854 ( 
.A1(n_19615),
.A2(n_19653),
.B(n_19607),
.C(n_19720),
.Y(n_19854)
);

OAI21xp33_ASAP7_75t_SL g19855 ( 
.A1(n_19669),
.A2(n_19639),
.B(n_19631),
.Y(n_19855)
);

OAI221xp5_ASAP7_75t_L g19856 ( 
.A1(n_19731),
.A2(n_7649),
.B1(n_7705),
.B2(n_7522),
.C(n_7487),
.Y(n_19856)
);

OAI21xp5_ASAP7_75t_SL g19857 ( 
.A1(n_19698),
.A2(n_5446),
.B(n_5445),
.Y(n_19857)
);

AOI211x1_ASAP7_75t_L g19858 ( 
.A1(n_19689),
.A2(n_9143),
.B(n_9147),
.C(n_9141),
.Y(n_19858)
);

OAI31xp33_ASAP7_75t_L g19859 ( 
.A1(n_19623),
.A2(n_6961),
.A3(n_6979),
.B(n_6963),
.Y(n_19859)
);

AOI32xp33_ASAP7_75t_L g19860 ( 
.A1(n_19611),
.A2(n_8452),
.A3(n_8451),
.B1(n_8448),
.B2(n_8290),
.Y(n_19860)
);

NAND2xp5_ASAP7_75t_SL g19861 ( 
.A(n_19651),
.B(n_7725),
.Y(n_19861)
);

INVx1_ASAP7_75t_L g19862 ( 
.A(n_19703),
.Y(n_19862)
);

NAND4xp25_ASAP7_75t_L g19863 ( 
.A(n_19660),
.B(n_5736),
.C(n_5513),
.D(n_5515),
.Y(n_19863)
);

AOI222xp33_ASAP7_75t_L g19864 ( 
.A1(n_19665),
.A2(n_9143),
.B1(n_9147),
.B2(n_9175),
.C1(n_9150),
.C2(n_9141),
.Y(n_19864)
);

AOI22xp5_ASAP7_75t_L g19865 ( 
.A1(n_19587),
.A2(n_8019),
.B1(n_7711),
.B2(n_7719),
.Y(n_19865)
);

AOI221xp5_ASAP7_75t_L g19866 ( 
.A1(n_19729),
.A2(n_9175),
.B1(n_9176),
.B2(n_9150),
.C(n_9147),
.Y(n_19866)
);

AOI221x1_ASAP7_75t_SL g19867 ( 
.A1(n_19727),
.A2(n_9176),
.B1(n_9201),
.B2(n_9175),
.C(n_9150),
.Y(n_19867)
);

INVx1_ASAP7_75t_L g19868 ( 
.A(n_19723),
.Y(n_19868)
);

NAND4xp25_ASAP7_75t_L g19869 ( 
.A(n_19652),
.B(n_5513),
.C(n_5515),
.D(n_5492),
.Y(n_19869)
);

HB1xp67_ASAP7_75t_L g19870 ( 
.A(n_19656),
.Y(n_19870)
);

AOI221xp5_ASAP7_75t_L g19871 ( 
.A1(n_19675),
.A2(n_9211),
.B1(n_9217),
.B2(n_9201),
.C(n_9176),
.Y(n_19871)
);

AOI211xp5_ASAP7_75t_L g19872 ( 
.A1(n_19594),
.A2(n_5446),
.B(n_5447),
.C(n_5445),
.Y(n_19872)
);

O2A1O1Ixp5_ASAP7_75t_L g19873 ( 
.A1(n_19672),
.A2(n_8701),
.B(n_8726),
.C(n_8707),
.Y(n_19873)
);

INVx1_ASAP7_75t_SL g19874 ( 
.A(n_19588),
.Y(n_19874)
);

NAND2xp5_ASAP7_75t_L g19875 ( 
.A(n_19681),
.B(n_8701),
.Y(n_19875)
);

OAI211xp5_ASAP7_75t_L g19876 ( 
.A1(n_19635),
.A2(n_5513),
.B(n_5515),
.C(n_5492),
.Y(n_19876)
);

NAND4xp25_ASAP7_75t_L g19877 ( 
.A(n_19598),
.B(n_5515),
.C(n_5533),
.D(n_5492),
.Y(n_19877)
);

OAI211xp5_ASAP7_75t_L g19878 ( 
.A1(n_19601),
.A2(n_5533),
.B(n_5579),
.C(n_5515),
.Y(n_19878)
);

OAI211xp5_ASAP7_75t_L g19879 ( 
.A1(n_19718),
.A2(n_5533),
.B(n_5579),
.C(n_5515),
.Y(n_19879)
);

AOI211xp5_ASAP7_75t_L g19880 ( 
.A1(n_19616),
.A2(n_5447),
.B(n_5448),
.C(n_5446),
.Y(n_19880)
);

AOI22xp5_ASAP7_75t_L g19881 ( 
.A1(n_19637),
.A2(n_8019),
.B1(n_7711),
.B2(n_7725),
.Y(n_19881)
);

OAI21xp33_ASAP7_75t_L g19882 ( 
.A1(n_19628),
.A2(n_5831),
.B(n_5804),
.Y(n_19882)
);

A2O1A1Ixp33_ASAP7_75t_SL g19883 ( 
.A1(n_19610),
.A2(n_9301),
.B(n_9299),
.C(n_8726),
.Y(n_19883)
);

AOI211xp5_ASAP7_75t_L g19884 ( 
.A1(n_19584),
.A2(n_5447),
.B(n_5448),
.C(n_5446),
.Y(n_19884)
);

AOI221x1_ASAP7_75t_L g19885 ( 
.A1(n_19610),
.A2(n_9217),
.B1(n_9219),
.B2(n_9211),
.C(n_9201),
.Y(n_19885)
);

O2A1O1Ixp5_ASAP7_75t_L g19886 ( 
.A1(n_19610),
.A2(n_8707),
.B(n_8727),
.C(n_8726),
.Y(n_19886)
);

OAI321xp33_ASAP7_75t_L g19887 ( 
.A1(n_19610),
.A2(n_7736),
.A3(n_7719),
.B1(n_7803),
.B2(n_7725),
.C(n_7625),
.Y(n_19887)
);

OAI22xp5_ASAP7_75t_L g19888 ( 
.A1(n_19610),
.A2(n_8707),
.B1(n_8727),
.B2(n_8726),
.Y(n_19888)
);

XNOR2xp5_ASAP7_75t_L g19889 ( 
.A(n_19602),
.B(n_7738),
.Y(n_19889)
);

CKINVDCx16_ASAP7_75t_R g19890 ( 
.A(n_19610),
.Y(n_19890)
);

OAI21xp5_ASAP7_75t_L g19891 ( 
.A1(n_19584),
.A2(n_8531),
.B(n_8291),
.Y(n_19891)
);

AOI22xp5_ASAP7_75t_L g19892 ( 
.A1(n_19745),
.A2(n_8019),
.B1(n_7719),
.B2(n_7725),
.Y(n_19892)
);

NAND3xp33_ASAP7_75t_SL g19893 ( 
.A(n_19759),
.B(n_5579),
.C(n_5533),
.Y(n_19893)
);

NOR2xp33_ASAP7_75t_L g19894 ( 
.A(n_19890),
.B(n_5601),
.Y(n_19894)
);

OR2x2_ASAP7_75t_L g19895 ( 
.A(n_19750),
.B(n_8704),
.Y(n_19895)
);

INVx1_ASAP7_75t_L g19896 ( 
.A(n_19889),
.Y(n_19896)
);

NOR3xp33_ASAP7_75t_L g19897 ( 
.A(n_19754),
.B(n_5579),
.C(n_5533),
.Y(n_19897)
);

NAND2x1p5_ASAP7_75t_L g19898 ( 
.A(n_19781),
.B(n_19792),
.Y(n_19898)
);

AOI21xp5_ASAP7_75t_L g19899 ( 
.A1(n_19870),
.A2(n_9301),
.B(n_8727),
.Y(n_19899)
);

OAI322xp33_ASAP7_75t_L g19900 ( 
.A1(n_19776),
.A2(n_9227),
.A3(n_9217),
.B1(n_9228),
.B2(n_9242),
.C1(n_9219),
.C2(n_9211),
.Y(n_19900)
);

INVx2_ASAP7_75t_L g19901 ( 
.A(n_19798),
.Y(n_19901)
);

AND2x4_ASAP7_75t_L g19902 ( 
.A(n_19808),
.B(n_8707),
.Y(n_19902)
);

NAND2xp5_ASAP7_75t_SL g19903 ( 
.A(n_19769),
.B(n_7625),
.Y(n_19903)
);

NOR3xp33_ASAP7_75t_L g19904 ( 
.A(n_19777),
.B(n_5579),
.C(n_5533),
.Y(n_19904)
);

INVx1_ASAP7_75t_L g19905 ( 
.A(n_19780),
.Y(n_19905)
);

NAND4xp75_ASAP7_75t_L g19906 ( 
.A(n_19794),
.B(n_8588),
.C(n_9058),
.D(n_9051),
.Y(n_19906)
);

AND2x2_ASAP7_75t_L g19907 ( 
.A(n_19789),
.B(n_19761),
.Y(n_19907)
);

NAND3xp33_ASAP7_75t_L g19908 ( 
.A(n_19749),
.B(n_5886),
.C(n_5510),
.Y(n_19908)
);

INVx1_ASAP7_75t_L g19909 ( 
.A(n_19845),
.Y(n_19909)
);

HB1xp67_ASAP7_75t_L g19910 ( 
.A(n_19771),
.Y(n_19910)
);

HB1xp67_ASAP7_75t_L g19911 ( 
.A(n_19862),
.Y(n_19911)
);

INVx1_ASAP7_75t_L g19912 ( 
.A(n_19810),
.Y(n_19912)
);

NAND4xp75_ASAP7_75t_L g19913 ( 
.A(n_19768),
.B(n_8588),
.C(n_9058),
.D(n_9051),
.Y(n_19913)
);

NOR3xp33_ASAP7_75t_L g19914 ( 
.A(n_19774),
.B(n_5580),
.C(n_5579),
.Y(n_19914)
);

NAND2x1p5_ASAP7_75t_L g19915 ( 
.A(n_19817),
.B(n_19770),
.Y(n_19915)
);

NOR2x1_ASAP7_75t_L g19916 ( 
.A(n_19842),
.B(n_5580),
.Y(n_19916)
);

INVx2_ASAP7_75t_SL g19917 ( 
.A(n_19828),
.Y(n_19917)
);

NOR2x1_ASAP7_75t_L g19918 ( 
.A(n_19834),
.B(n_5580),
.Y(n_19918)
);

NOR4xp75_ASAP7_75t_L g19919 ( 
.A(n_19818),
.B(n_7343),
.C(n_7357),
.D(n_7349),
.Y(n_19919)
);

NAND3xp33_ASAP7_75t_L g19920 ( 
.A(n_19820),
.B(n_5886),
.C(n_5510),
.Y(n_19920)
);

NOR2x1_ASAP7_75t_L g19921 ( 
.A(n_19839),
.B(n_19836),
.Y(n_19921)
);

INVx1_ASAP7_75t_L g19922 ( 
.A(n_19783),
.Y(n_19922)
);

NOR3xp33_ASAP7_75t_L g19923 ( 
.A(n_19746),
.B(n_5660),
.C(n_5580),
.Y(n_19923)
);

NOR2x1_ASAP7_75t_L g19924 ( 
.A(n_19868),
.B(n_5580),
.Y(n_19924)
);

NAND2xp33_ASAP7_75t_L g19925 ( 
.A(n_19874),
.B(n_5446),
.Y(n_19925)
);

NAND3xp33_ASAP7_75t_L g19926 ( 
.A(n_19807),
.B(n_5717),
.C(n_5463),
.Y(n_19926)
);

NAND2xp5_ASAP7_75t_L g19927 ( 
.A(n_19752),
.B(n_8727),
.Y(n_19927)
);

AOI22xp5_ASAP7_75t_L g19928 ( 
.A1(n_19855),
.A2(n_8019),
.B1(n_7725),
.B2(n_7736),
.Y(n_19928)
);

NOR3xp33_ASAP7_75t_L g19929 ( 
.A(n_19747),
.B(n_5660),
.C(n_5580),
.Y(n_19929)
);

INVx1_ASAP7_75t_L g19930 ( 
.A(n_19772),
.Y(n_19930)
);

NAND4xp25_ASAP7_75t_L g19931 ( 
.A(n_19854),
.B(n_5660),
.C(n_4577),
.D(n_4583),
.Y(n_19931)
);

AOI22xp5_ASAP7_75t_L g19932 ( 
.A1(n_19849),
.A2(n_8019),
.B1(n_7725),
.B2(n_7736),
.Y(n_19932)
);

NAND2xp5_ASAP7_75t_SL g19933 ( 
.A(n_19825),
.B(n_7719),
.Y(n_19933)
);

NOR3xp33_ASAP7_75t_L g19934 ( 
.A(n_19748),
.B(n_5660),
.C(n_5806),
.Y(n_19934)
);

NOR2x1_ASAP7_75t_L g19935 ( 
.A(n_19806),
.B(n_5660),
.Y(n_19935)
);

NAND3xp33_ASAP7_75t_SL g19936 ( 
.A(n_19884),
.B(n_5660),
.C(n_5806),
.Y(n_19936)
);

NAND3xp33_ASAP7_75t_L g19937 ( 
.A(n_19765),
.B(n_5605),
.C(n_5463),
.Y(n_19937)
);

NAND4xp75_ASAP7_75t_L g19938 ( 
.A(n_19859),
.B(n_8588),
.C(n_9058),
.D(n_9051),
.Y(n_19938)
);

NAND3xp33_ASAP7_75t_L g19939 ( 
.A(n_19843),
.B(n_19758),
.C(n_19816),
.Y(n_19939)
);

NOR3xp33_ASAP7_75t_L g19940 ( 
.A(n_19787),
.B(n_5812),
.C(n_5806),
.Y(n_19940)
);

NOR2x1_ASAP7_75t_L g19941 ( 
.A(n_19814),
.B(n_5447),
.Y(n_19941)
);

NOR3xp33_ASAP7_75t_SL g19942 ( 
.A(n_19824),
.B(n_7193),
.C(n_7547),
.Y(n_19942)
);

NAND2xp5_ASAP7_75t_L g19943 ( 
.A(n_19822),
.B(n_8741),
.Y(n_19943)
);

NOR3xp33_ASAP7_75t_L g19944 ( 
.A(n_19799),
.B(n_5822),
.C(n_5812),
.Y(n_19944)
);

AO22x2_ASAP7_75t_L g19945 ( 
.A1(n_19858),
.A2(n_8746),
.B1(n_8773),
.B2(n_8741),
.Y(n_19945)
);

NAND3xp33_ASAP7_75t_L g19946 ( 
.A(n_19823),
.B(n_5605),
.C(n_5463),
.Y(n_19946)
);

NAND4xp75_ASAP7_75t_L g19947 ( 
.A(n_19861),
.B(n_19755),
.C(n_19891),
.D(n_19791),
.Y(n_19947)
);

NAND3xp33_ASAP7_75t_L g19948 ( 
.A(n_19811),
.B(n_5605),
.C(n_5463),
.Y(n_19948)
);

NAND4xp25_ASAP7_75t_L g19949 ( 
.A(n_19756),
.B(n_4577),
.C(n_4583),
.D(n_4569),
.Y(n_19949)
);

NAND3xp33_ASAP7_75t_SL g19950 ( 
.A(n_19760),
.B(n_5816),
.C(n_5812),
.Y(n_19950)
);

NOR2x1_ASAP7_75t_L g19951 ( 
.A(n_19837),
.B(n_5447),
.Y(n_19951)
);

NOR2x1_ASAP7_75t_L g19952 ( 
.A(n_19869),
.B(n_5447),
.Y(n_19952)
);

NAND3xp33_ASAP7_75t_L g19953 ( 
.A(n_19844),
.B(n_5605),
.C(n_5463),
.Y(n_19953)
);

NOR3xp33_ASAP7_75t_L g19954 ( 
.A(n_19882),
.B(n_5822),
.C(n_5812),
.Y(n_19954)
);

NAND4xp75_ASAP7_75t_L g19955 ( 
.A(n_19785),
.B(n_9058),
.C(n_9059),
.D(n_9051),
.Y(n_19955)
);

INVx1_ASAP7_75t_L g19956 ( 
.A(n_19809),
.Y(n_19956)
);

INVxp67_ASAP7_75t_L g19957 ( 
.A(n_19821),
.Y(n_19957)
);

NAND4xp75_ASAP7_75t_L g19958 ( 
.A(n_19875),
.B(n_9058),
.C(n_9059),
.D(n_9051),
.Y(n_19958)
);

NOR2x1_ASAP7_75t_L g19959 ( 
.A(n_19795),
.B(n_19863),
.Y(n_19959)
);

AOI22xp5_ASAP7_75t_L g19960 ( 
.A1(n_19773),
.A2(n_7725),
.B1(n_7736),
.B2(n_7719),
.Y(n_19960)
);

OAI22xp5_ASAP7_75t_L g19961 ( 
.A1(n_19856),
.A2(n_19805),
.B1(n_19865),
.B2(n_19753),
.Y(n_19961)
);

NOR2xp33_ASAP7_75t_L g19962 ( 
.A(n_19877),
.B(n_5601),
.Y(n_19962)
);

AOI22xp5_ASAP7_75t_L g19963 ( 
.A1(n_19790),
.A2(n_7725),
.B1(n_7736),
.B2(n_7719),
.Y(n_19963)
);

NOR3xp33_ASAP7_75t_L g19964 ( 
.A(n_19879),
.B(n_19876),
.C(n_19857),
.Y(n_19964)
);

NOR2x1_ASAP7_75t_L g19965 ( 
.A(n_19831),
.B(n_5447),
.Y(n_19965)
);

NAND4xp25_ASAP7_75t_L g19966 ( 
.A(n_19872),
.B(n_19846),
.C(n_19812),
.D(n_19840),
.Y(n_19966)
);

INVx1_ASAP7_75t_L g19967 ( 
.A(n_19838),
.Y(n_19967)
);

NAND3xp33_ASAP7_75t_L g19968 ( 
.A(n_19880),
.B(n_5707),
.C(n_5449),
.Y(n_19968)
);

NOR2xp67_ASAP7_75t_L g19969 ( 
.A(n_19815),
.B(n_5448),
.Y(n_19969)
);

NAND2xp5_ASAP7_75t_L g19970 ( 
.A(n_19800),
.B(n_8741),
.Y(n_19970)
);

INVx1_ASAP7_75t_L g19971 ( 
.A(n_19878),
.Y(n_19971)
);

NOR3xp33_ASAP7_75t_L g19972 ( 
.A(n_19819),
.B(n_5816),
.C(n_5812),
.Y(n_19972)
);

NOR3xp33_ASAP7_75t_L g19973 ( 
.A(n_19784),
.B(n_5822),
.C(n_5816),
.Y(n_19973)
);

NAND2xp33_ASAP7_75t_L g19974 ( 
.A(n_19847),
.B(n_5448),
.Y(n_19974)
);

NAND2xp5_ASAP7_75t_L g19975 ( 
.A(n_19813),
.B(n_8741),
.Y(n_19975)
);

NAND3xp33_ASAP7_75t_SL g19976 ( 
.A(n_19786),
.B(n_19751),
.C(n_19802),
.Y(n_19976)
);

OA22x2_ASAP7_75t_L g19977 ( 
.A1(n_19881),
.A2(n_8746),
.B1(n_8775),
.B2(n_8773),
.Y(n_19977)
);

NOR3xp33_ASAP7_75t_SL g19978 ( 
.A(n_19788),
.B(n_7193),
.C(n_7089),
.Y(n_19978)
);

INVx1_ASAP7_75t_L g19979 ( 
.A(n_19886),
.Y(n_19979)
);

NOR3xp33_ASAP7_75t_L g19980 ( 
.A(n_19762),
.B(n_5822),
.C(n_5816),
.Y(n_19980)
);

NOR3xp33_ASAP7_75t_L g19981 ( 
.A(n_19782),
.B(n_5822),
.C(n_5816),
.Y(n_19981)
);

AOI22xp5_ASAP7_75t_L g19982 ( 
.A1(n_19778),
.A2(n_19793),
.B1(n_19801),
.B2(n_19766),
.Y(n_19982)
);

NOR3xp33_ASAP7_75t_L g19983 ( 
.A(n_19804),
.B(n_19873),
.C(n_19797),
.Y(n_19983)
);

NAND2x1p5_ASAP7_75t_L g19984 ( 
.A(n_19796),
.B(n_5448),
.Y(n_19984)
);

NOR2x1p5_ASAP7_75t_L g19985 ( 
.A(n_19850),
.B(n_5448),
.Y(n_19985)
);

NAND4xp75_ASAP7_75t_L g19986 ( 
.A(n_19826),
.B(n_9059),
.C(n_9058),
.D(n_4580),
.Y(n_19986)
);

NOR2x1_ASAP7_75t_L g19987 ( 
.A(n_19851),
.B(n_5448),
.Y(n_19987)
);

INVx1_ASAP7_75t_L g19988 ( 
.A(n_19867),
.Y(n_19988)
);

NAND2xp5_ASAP7_75t_L g19989 ( 
.A(n_19803),
.B(n_8746),
.Y(n_19989)
);

NAND3xp33_ASAP7_75t_L g19990 ( 
.A(n_19864),
.B(n_5540),
.C(n_5469),
.Y(n_19990)
);

INVx1_ASAP7_75t_L g19991 ( 
.A(n_19832),
.Y(n_19991)
);

INVx1_ASAP7_75t_L g19992 ( 
.A(n_19888),
.Y(n_19992)
);

NAND2xp5_ASAP7_75t_L g19993 ( 
.A(n_19841),
.B(n_8746),
.Y(n_19993)
);

NAND4xp25_ASAP7_75t_L g19994 ( 
.A(n_19883),
.B(n_19830),
.C(n_19779),
.D(n_19827),
.Y(n_19994)
);

NOR3xp33_ASAP7_75t_L g19995 ( 
.A(n_19887),
.B(n_5920),
.C(n_5904),
.Y(n_19995)
);

AND2x4_ASAP7_75t_L g19996 ( 
.A(n_19848),
.B(n_8773),
.Y(n_19996)
);

NOR3xp33_ASAP7_75t_L g19997 ( 
.A(n_19835),
.B(n_5920),
.C(n_5904),
.Y(n_19997)
);

NAND2xp5_ASAP7_75t_L g19998 ( 
.A(n_19871),
.B(n_8773),
.Y(n_19998)
);

NOR2xp33_ASAP7_75t_L g19999 ( 
.A(n_19853),
.B(n_5601),
.Y(n_19999)
);

NAND4xp75_ASAP7_75t_L g20000 ( 
.A(n_19885),
.B(n_9059),
.C(n_4631),
.D(n_4572),
.Y(n_20000)
);

INVx1_ASAP7_75t_L g20001 ( 
.A(n_19866),
.Y(n_20001)
);

AND2x2_ASAP7_75t_L g20002 ( 
.A(n_19829),
.B(n_6996),
.Y(n_20002)
);

NOR3x1_ASAP7_75t_L g20003 ( 
.A(n_19833),
.B(n_8531),
.C(n_8532),
.Y(n_20003)
);

INVx1_ASAP7_75t_L g20004 ( 
.A(n_19852),
.Y(n_20004)
);

AOI22xp5_ASAP7_75t_L g20005 ( 
.A1(n_19764),
.A2(n_7803),
.B1(n_7736),
.B2(n_6960),
.Y(n_20005)
);

BUFx2_ASAP7_75t_L g20006 ( 
.A(n_19757),
.Y(n_20006)
);

NOR3x1_ASAP7_75t_L g20007 ( 
.A(n_19767),
.B(n_8531),
.C(n_8532),
.Y(n_20007)
);

NOR2x1_ASAP7_75t_L g20008 ( 
.A(n_19775),
.B(n_5448),
.Y(n_20008)
);

NOR2xp33_ASAP7_75t_L g20009 ( 
.A(n_19763),
.B(n_5601),
.Y(n_20009)
);

INVx1_ASAP7_75t_L g20010 ( 
.A(n_19860),
.Y(n_20010)
);

AND2x2_ASAP7_75t_L g20011 ( 
.A(n_19890),
.B(n_6996),
.Y(n_20011)
);

INVx2_ASAP7_75t_SL g20012 ( 
.A(n_19889),
.Y(n_20012)
);

NAND2xp5_ASAP7_75t_L g20013 ( 
.A(n_19890),
.B(n_8775),
.Y(n_20013)
);

INVx1_ASAP7_75t_L g20014 ( 
.A(n_19889),
.Y(n_20014)
);

INVx1_ASAP7_75t_L g20015 ( 
.A(n_19889),
.Y(n_20015)
);

INVx1_ASAP7_75t_L g20016 ( 
.A(n_19889),
.Y(n_20016)
);

NAND3xp33_ASAP7_75t_SL g20017 ( 
.A(n_19759),
.B(n_5920),
.C(n_5904),
.Y(n_20017)
);

INVx1_ASAP7_75t_SL g20018 ( 
.A(n_19759),
.Y(n_20018)
);

OAI22xp5_ASAP7_75t_L g20019 ( 
.A1(n_19890),
.A2(n_8807),
.B1(n_8816),
.B2(n_8775),
.Y(n_20019)
);

INVx1_ASAP7_75t_L g20020 ( 
.A(n_19889),
.Y(n_20020)
);

AOI21xp5_ASAP7_75t_L g20021 ( 
.A1(n_19745),
.A2(n_9301),
.B(n_9299),
.Y(n_20021)
);

A2O1A1Ixp33_ASAP7_75t_SL g20022 ( 
.A1(n_19745),
.A2(n_8807),
.B(n_8816),
.C(n_8775),
.Y(n_20022)
);

NOR2x1_ASAP7_75t_L g20023 ( 
.A(n_19750),
.B(n_5448),
.Y(n_20023)
);

OAI22xp5_ASAP7_75t_L g20024 ( 
.A1(n_19890),
.A2(n_8816),
.B1(n_8828),
.B2(n_8807),
.Y(n_20024)
);

AOI21xp5_ASAP7_75t_SL g20025 ( 
.A1(n_19967),
.A2(n_5453),
.B(n_5449),
.Y(n_20025)
);

NAND5xp2_ASAP7_75t_L g20026 ( 
.A(n_19912),
.B(n_7095),
.C(n_7901),
.D(n_7900),
.E(n_7839),
.Y(n_20026)
);

AOI22xp5_ASAP7_75t_L g20027 ( 
.A1(n_20018),
.A2(n_8816),
.B1(n_8828),
.B2(n_8807),
.Y(n_20027)
);

INVx1_ASAP7_75t_L g20028 ( 
.A(n_19911),
.Y(n_20028)
);

NAND3xp33_ASAP7_75t_SL g20029 ( 
.A(n_19901),
.B(n_5920),
.C(n_5904),
.Y(n_20029)
);

NOR3xp33_ASAP7_75t_SL g20030 ( 
.A(n_19909),
.B(n_7193),
.C(n_7089),
.Y(n_20030)
);

NAND4xp25_ASAP7_75t_L g20031 ( 
.A(n_19896),
.B(n_4577),
.C(n_4583),
.D(n_4569),
.Y(n_20031)
);

INVx1_ASAP7_75t_L g20032 ( 
.A(n_19910),
.Y(n_20032)
);

NOR2x1p5_ASAP7_75t_L g20033 ( 
.A(n_20014),
.B(n_5449),
.Y(n_20033)
);

INVx2_ASAP7_75t_L g20034 ( 
.A(n_19895),
.Y(n_20034)
);

NOR2xp33_ASAP7_75t_L g20035 ( 
.A(n_19933),
.B(n_5601),
.Y(n_20035)
);

OR5x1_ASAP7_75t_L g20036 ( 
.A(n_19966),
.B(n_7095),
.C(n_8716),
.D(n_8704),
.E(n_8013),
.Y(n_20036)
);

AOI221x1_ASAP7_75t_L g20037 ( 
.A1(n_20004),
.A2(n_9228),
.B1(n_9242),
.B2(n_9227),
.C(n_9219),
.Y(n_20037)
);

O2A1O1Ixp33_ASAP7_75t_L g20038 ( 
.A1(n_19917),
.A2(n_4572),
.B(n_7409),
.C(n_7406),
.Y(n_20038)
);

INVx1_ASAP7_75t_L g20039 ( 
.A(n_20013),
.Y(n_20039)
);

NAND3xp33_ASAP7_75t_SL g20040 ( 
.A(n_19898),
.B(n_5920),
.C(n_5904),
.Y(n_20040)
);

O2A1O1Ixp33_ASAP7_75t_L g20041 ( 
.A1(n_20012),
.A2(n_7409),
.B(n_7412),
.C(n_7406),
.Y(n_20041)
);

OAI311xp33_ASAP7_75t_L g20042 ( 
.A1(n_19928),
.A2(n_7901),
.A3(n_7906),
.B1(n_7890),
.C1(n_7839),
.Y(n_20042)
);

NAND4xp25_ASAP7_75t_SL g20043 ( 
.A(n_20021),
.B(n_7906),
.C(n_7890),
.D(n_9227),
.Y(n_20043)
);

NOR2xp67_ASAP7_75t_L g20044 ( 
.A(n_20015),
.B(n_5449),
.Y(n_20044)
);

NOR5xp2_ASAP7_75t_L g20045 ( 
.A(n_19957),
.B(n_7708),
.C(n_7712),
.D(n_7779),
.E(n_7752),
.Y(n_20045)
);

OAI21xp33_ASAP7_75t_L g20046 ( 
.A1(n_19894),
.A2(n_5930),
.B(n_5892),
.Y(n_20046)
);

NAND3xp33_ASAP7_75t_L g20047 ( 
.A(n_19921),
.B(n_5453),
.C(n_5449),
.Y(n_20047)
);

OAI211xp5_ASAP7_75t_L g20048 ( 
.A1(n_20016),
.A2(n_5453),
.B(n_5458),
.C(n_5449),
.Y(n_20048)
);

A2O1A1Ixp33_ASAP7_75t_L g20049 ( 
.A1(n_19902),
.A2(n_9301),
.B(n_9299),
.C(n_8839),
.Y(n_20049)
);

NOR3xp33_ASAP7_75t_L g20050 ( 
.A(n_20020),
.B(n_5937),
.C(n_5934),
.Y(n_20050)
);

NAND4xp25_ASAP7_75t_L g20051 ( 
.A(n_20022),
.B(n_4569),
.C(n_4583),
.D(n_4577),
.Y(n_20051)
);

NAND4xp75_ASAP7_75t_L g20052 ( 
.A(n_19907),
.B(n_9059),
.C(n_9242),
.D(n_9228),
.Y(n_20052)
);

NAND2xp5_ASAP7_75t_L g20053 ( 
.A(n_20011),
.B(n_8828),
.Y(n_20053)
);

OAI211xp5_ASAP7_75t_L g20054 ( 
.A1(n_19988),
.A2(n_5453),
.B(n_5458),
.C(n_5449),
.Y(n_20054)
);

AOI221x1_ASAP7_75t_L g20055 ( 
.A1(n_19905),
.A2(n_9252),
.B1(n_8840),
.B2(n_8864),
.C(n_8839),
.Y(n_20055)
);

AOI221xp5_ASAP7_75t_L g20056 ( 
.A1(n_19961),
.A2(n_9252),
.B1(n_8828),
.B2(n_8864),
.C(n_8840),
.Y(n_20056)
);

OAI21xp5_ASAP7_75t_SL g20057 ( 
.A1(n_19915),
.A2(n_5453),
.B(n_5449),
.Y(n_20057)
);

NAND4xp25_ASAP7_75t_L g20058 ( 
.A(n_20023),
.B(n_4584),
.C(n_4607),
.D(n_4569),
.Y(n_20058)
);

OAI22xp5_ASAP7_75t_L g20059 ( 
.A1(n_19926),
.A2(n_8840),
.B1(n_8864),
.B2(n_8839),
.Y(n_20059)
);

NOR3xp33_ASAP7_75t_L g20060 ( 
.A(n_19922),
.B(n_5937),
.C(n_5934),
.Y(n_20060)
);

AOI211x1_ASAP7_75t_L g20061 ( 
.A1(n_19908),
.A2(n_9252),
.B(n_7349),
.C(n_7357),
.Y(n_20061)
);

OAI211xp5_ASAP7_75t_SL g20062 ( 
.A1(n_19991),
.A2(n_8840),
.B(n_8864),
.C(n_8839),
.Y(n_20062)
);

NOR2xp33_ASAP7_75t_L g20063 ( 
.A(n_19903),
.B(n_5601),
.Y(n_20063)
);

AOI21xp5_ASAP7_75t_L g20064 ( 
.A1(n_20010),
.A2(n_8882),
.B(n_8872),
.Y(n_20064)
);

AOI322xp5_ASAP7_75t_L g20065 ( 
.A1(n_19902),
.A2(n_9299),
.A3(n_8882),
.B1(n_8896),
.B2(n_8925),
.C1(n_8955),
.C2(n_8949),
.Y(n_20065)
);

NAND4xp25_ASAP7_75t_L g20066 ( 
.A(n_19916),
.B(n_4584),
.C(n_4607),
.D(n_6171),
.Y(n_20066)
);

AND5x1_ASAP7_75t_L g20067 ( 
.A(n_19982),
.B(n_7095),
.C(n_8716),
.D(n_8704),
.E(n_8013),
.Y(n_20067)
);

NAND2xp5_ASAP7_75t_L g20068 ( 
.A(n_19999),
.B(n_8872),
.Y(n_20068)
);

NAND3xp33_ASAP7_75t_SL g20069 ( 
.A(n_20001),
.B(n_5937),
.C(n_5934),
.Y(n_20069)
);

AOI211xp5_ASAP7_75t_L g20070 ( 
.A1(n_19971),
.A2(n_5453),
.B(n_5458),
.C(n_5449),
.Y(n_20070)
);

NAND3xp33_ASAP7_75t_L g20071 ( 
.A(n_19930),
.B(n_5458),
.C(n_5453),
.Y(n_20071)
);

NAND3xp33_ASAP7_75t_SL g20072 ( 
.A(n_20006),
.B(n_5937),
.C(n_5934),
.Y(n_20072)
);

OAI221xp5_ASAP7_75t_L g20073 ( 
.A1(n_19956),
.A2(n_5463),
.B1(n_5469),
.B2(n_5458),
.C(n_5453),
.Y(n_20073)
);

NAND3xp33_ASAP7_75t_SL g20074 ( 
.A(n_19992),
.B(n_5937),
.C(n_5934),
.Y(n_20074)
);

NAND2xp5_ASAP7_75t_SL g20075 ( 
.A(n_19959),
.B(n_7736),
.Y(n_20075)
);

NAND3xp33_ASAP7_75t_SL g20076 ( 
.A(n_19979),
.B(n_5994),
.C(n_5964),
.Y(n_20076)
);

NOR2x1_ASAP7_75t_L g20077 ( 
.A(n_19924),
.B(n_5453),
.Y(n_20077)
);

AOI221xp5_ASAP7_75t_L g20078 ( 
.A1(n_19964),
.A2(n_8872),
.B1(n_8925),
.B2(n_8896),
.C(n_8882),
.Y(n_20078)
);

NAND4xp25_ASAP7_75t_SL g20079 ( 
.A(n_19929),
.B(n_8882),
.C(n_8896),
.D(n_8872),
.Y(n_20079)
);

AOI221xp5_ASAP7_75t_L g20080 ( 
.A1(n_19976),
.A2(n_8896),
.B1(n_8955),
.B2(n_8949),
.C(n_8925),
.Y(n_20080)
);

OAI211xp5_ASAP7_75t_L g20081 ( 
.A1(n_19994),
.A2(n_5463),
.B(n_5469),
.C(n_5458),
.Y(n_20081)
);

NAND3xp33_ASAP7_75t_SL g20082 ( 
.A(n_19983),
.B(n_5994),
.C(n_5964),
.Y(n_20082)
);

NAND4xp25_ASAP7_75t_L g20083 ( 
.A(n_19939),
.B(n_4584),
.C(n_4607),
.D(n_6171),
.Y(n_20083)
);

NOR4xp25_ASAP7_75t_L g20084 ( 
.A(n_19925),
.B(n_8949),
.C(n_8955),
.D(n_8925),
.Y(n_20084)
);

OAI211xp5_ASAP7_75t_L g20085 ( 
.A1(n_19935),
.A2(n_5463),
.B(n_5469),
.C(n_5458),
.Y(n_20085)
);

AOI211xp5_ASAP7_75t_L g20086 ( 
.A1(n_19923),
.A2(n_5463),
.B(n_5469),
.C(n_5458),
.Y(n_20086)
);

NOR3xp33_ASAP7_75t_L g20087 ( 
.A(n_19947),
.B(n_5994),
.C(n_5964),
.Y(n_20087)
);

NAND2xp5_ASAP7_75t_L g20088 ( 
.A(n_19918),
.B(n_8949),
.Y(n_20088)
);

OAI221xp5_ASAP7_75t_L g20089 ( 
.A1(n_19892),
.A2(n_5484),
.B1(n_5500),
.B2(n_5469),
.C(n_5458),
.Y(n_20089)
);

NAND4xp75_ASAP7_75t_L g20090 ( 
.A(n_19951),
.B(n_9059),
.C(n_8959),
.D(n_8977),
.Y(n_20090)
);

AOI21xp5_ASAP7_75t_L g20091 ( 
.A1(n_19974),
.A2(n_8959),
.B(n_8955),
.Y(n_20091)
);

NOR4xp25_ASAP7_75t_L g20092 ( 
.A(n_19893),
.B(n_8977),
.C(n_8992),
.D(n_8959),
.Y(n_20092)
);

AOI21xp5_ASAP7_75t_L g20093 ( 
.A1(n_19934),
.A2(n_8977),
.B(n_8959),
.Y(n_20093)
);

NAND2xp5_ASAP7_75t_L g20094 ( 
.A(n_19962),
.B(n_8977),
.Y(n_20094)
);

NAND4xp25_ASAP7_75t_L g20095 ( 
.A(n_19931),
.B(n_19914),
.C(n_19897),
.D(n_19904),
.Y(n_20095)
);

NAND4xp25_ASAP7_75t_L g20096 ( 
.A(n_19920),
.B(n_4584),
.C(n_4607),
.D(n_6872),
.Y(n_20096)
);

NAND3xp33_ASAP7_75t_L g20097 ( 
.A(n_19942),
.B(n_5484),
.C(n_5469),
.Y(n_20097)
);

AOI221xp5_ASAP7_75t_L g20098 ( 
.A1(n_20017),
.A2(n_8992),
.B1(n_9049),
.B2(n_9043),
.C(n_9030),
.Y(n_20098)
);

OAI221xp5_ASAP7_75t_L g20099 ( 
.A1(n_19941),
.A2(n_19969),
.B1(n_19952),
.B2(n_19954),
.C(n_19984),
.Y(n_20099)
);

NOR2x1p5_ASAP7_75t_L g20100 ( 
.A(n_19936),
.B(n_5469),
.Y(n_20100)
);

INVx1_ASAP7_75t_L g20101 ( 
.A(n_19987),
.Y(n_20101)
);

NOR4xp25_ASAP7_75t_L g20102 ( 
.A(n_19950),
.B(n_9030),
.C(n_9043),
.D(n_8992),
.Y(n_20102)
);

NAND5xp2_ASAP7_75t_L g20103 ( 
.A(n_19997),
.B(n_7095),
.C(n_5646),
.D(n_6324),
.E(n_6890),
.Y(n_20103)
);

AOI221xp5_ASAP7_75t_L g20104 ( 
.A1(n_19944),
.A2(n_20009),
.B1(n_19981),
.B2(n_19980),
.C(n_19953),
.Y(n_20104)
);

NAND2xp5_ASAP7_75t_L g20105 ( 
.A(n_19985),
.B(n_8992),
.Y(n_20105)
);

OAI211xp5_ASAP7_75t_SL g20106 ( 
.A1(n_19943),
.A2(n_19975),
.B(n_19932),
.C(n_19965),
.Y(n_20106)
);

NOR3xp33_ASAP7_75t_L g20107 ( 
.A(n_19949),
.B(n_5994),
.C(n_5964),
.Y(n_20107)
);

OAI211xp5_ASAP7_75t_SL g20108 ( 
.A1(n_19993),
.A2(n_9043),
.B(n_9049),
.C(n_9030),
.Y(n_20108)
);

NAND3xp33_ASAP7_75t_L g20109 ( 
.A(n_19946),
.B(n_5484),
.C(n_5469),
.Y(n_20109)
);

NOR2x1_ASAP7_75t_L g20110 ( 
.A(n_20008),
.B(n_5484),
.Y(n_20110)
);

AND2x4_ASAP7_75t_L g20111 ( 
.A(n_19948),
.B(n_9030),
.Y(n_20111)
);

NAND3xp33_ASAP7_75t_L g20112 ( 
.A(n_19972),
.B(n_5500),
.C(n_5484),
.Y(n_20112)
);

NAND4xp25_ASAP7_75t_L g20113 ( 
.A(n_20002),
.B(n_19940),
.C(n_19968),
.D(n_19937),
.Y(n_20113)
);

NAND2xp5_ASAP7_75t_L g20114 ( 
.A(n_19996),
.B(n_9043),
.Y(n_20114)
);

NOR2xp67_ASAP7_75t_L g20115 ( 
.A(n_19927),
.B(n_5484),
.Y(n_20115)
);

NAND2xp5_ASAP7_75t_SL g20116 ( 
.A(n_19963),
.B(n_7736),
.Y(n_20116)
);

AOI221xp5_ASAP7_75t_L g20117 ( 
.A1(n_19996),
.A2(n_9049),
.B1(n_9098),
.B2(n_9068),
.C(n_9062),
.Y(n_20117)
);

NAND5xp2_ASAP7_75t_L g20118 ( 
.A(n_19973),
.B(n_7095),
.C(n_6890),
.D(n_6873),
.E(n_6858),
.Y(n_20118)
);

OAI211xp5_ASAP7_75t_SL g20119 ( 
.A1(n_19998),
.A2(n_9062),
.B(n_9068),
.C(n_9049),
.Y(n_20119)
);

AOI211xp5_ASAP7_75t_L g20120 ( 
.A1(n_19970),
.A2(n_5500),
.B(n_5510),
.C(n_5484),
.Y(n_20120)
);

NAND2xp5_ASAP7_75t_L g20121 ( 
.A(n_19977),
.B(n_9062),
.Y(n_20121)
);

NAND2xp5_ASAP7_75t_L g20122 ( 
.A(n_19945),
.B(n_9062),
.Y(n_20122)
);

OAI211xp5_ASAP7_75t_SL g20123 ( 
.A1(n_19978),
.A2(n_9098),
.B(n_9102),
.C(n_9068),
.Y(n_20123)
);

NAND2xp5_ASAP7_75t_SL g20124 ( 
.A(n_19899),
.B(n_7736),
.Y(n_20124)
);

OAI221xp5_ASAP7_75t_L g20125 ( 
.A1(n_19989),
.A2(n_5510),
.B1(n_5540),
.B2(n_5500),
.C(n_5484),
.Y(n_20125)
);

A2O1A1Ixp33_ASAP7_75t_L g20126 ( 
.A1(n_19990),
.A2(n_9098),
.B(n_9102),
.C(n_9068),
.Y(n_20126)
);

NAND5xp2_ASAP7_75t_L g20127 ( 
.A(n_19995),
.B(n_7095),
.C(n_6890),
.D(n_6858),
.E(n_7274),
.Y(n_20127)
);

NAND5xp2_ASAP7_75t_L g20128 ( 
.A(n_20005),
.B(n_19960),
.C(n_19945),
.D(n_19919),
.E(n_20007),
.Y(n_20128)
);

CKINVDCx20_ASAP7_75t_R g20129 ( 
.A(n_20019),
.Y(n_20129)
);

NOR3xp33_ASAP7_75t_L g20130 ( 
.A(n_20024),
.B(n_19938),
.C(n_19986),
.Y(n_20130)
);

NOR2x1_ASAP7_75t_L g20131 ( 
.A(n_20000),
.B(n_5484),
.Y(n_20131)
);

NAND5xp2_ASAP7_75t_L g20132 ( 
.A(n_19955),
.B(n_7095),
.C(n_6890),
.D(n_7277),
.E(n_7274),
.Y(n_20132)
);

OAI211xp5_ASAP7_75t_L g20133 ( 
.A1(n_19900),
.A2(n_5510),
.B(n_5540),
.C(n_5500),
.Y(n_20133)
);

NAND5xp2_ASAP7_75t_L g20134 ( 
.A(n_20003),
.B(n_6890),
.C(n_7277),
.D(n_7286),
.E(n_7274),
.Y(n_20134)
);

NOR2xp33_ASAP7_75t_L g20135 ( 
.A(n_19958),
.B(n_5500),
.Y(n_20135)
);

AOI22xp5_ASAP7_75t_L g20136 ( 
.A1(n_20028),
.A2(n_19906),
.B1(n_19913),
.B2(n_7803),
.Y(n_20136)
);

INVx1_ASAP7_75t_L g20137 ( 
.A(n_20032),
.Y(n_20137)
);

INVx2_ASAP7_75t_L g20138 ( 
.A(n_20033),
.Y(n_20138)
);

INVx1_ASAP7_75t_L g20139 ( 
.A(n_20101),
.Y(n_20139)
);

BUFx2_ASAP7_75t_L g20140 ( 
.A(n_20129),
.Y(n_20140)
);

AOI221xp5_ASAP7_75t_L g20141 ( 
.A1(n_20130),
.A2(n_9237),
.B1(n_9112),
.B2(n_9102),
.C(n_9103),
.Y(n_20141)
);

NAND4xp25_ASAP7_75t_L g20142 ( 
.A(n_20034),
.B(n_20128),
.C(n_20106),
.D(n_20104),
.Y(n_20142)
);

NOR2xp67_ASAP7_75t_L g20143 ( 
.A(n_20099),
.B(n_20039),
.Y(n_20143)
);

HB1xp67_ASAP7_75t_L g20144 ( 
.A(n_20044),
.Y(n_20144)
);

INVx1_ASAP7_75t_L g20145 ( 
.A(n_20110),
.Y(n_20145)
);

NAND4xp75_ASAP7_75t_L g20146 ( 
.A(n_20075),
.B(n_9102),
.C(n_9103),
.D(n_9098),
.Y(n_20146)
);

HB1xp67_ASAP7_75t_L g20147 ( 
.A(n_20077),
.Y(n_20147)
);

AND2x2_ASAP7_75t_L g20148 ( 
.A(n_20035),
.B(n_6961),
.Y(n_20148)
);

NOR2x1_ASAP7_75t_L g20149 ( 
.A(n_20047),
.B(n_5500),
.Y(n_20149)
);

INVx1_ASAP7_75t_SL g20150 ( 
.A(n_20094),
.Y(n_20150)
);

XOR2xp5_ASAP7_75t_L g20151 ( 
.A(n_20113),
.B(n_5500),
.Y(n_20151)
);

OR2x2_ASAP7_75t_L g20152 ( 
.A(n_20134),
.B(n_20058),
.Y(n_20152)
);

AOI22xp5_ASAP7_75t_L g20153 ( 
.A1(n_20087),
.A2(n_7803),
.B1(n_6960),
.B2(n_7014),
.Y(n_20153)
);

INVx1_ASAP7_75t_L g20154 ( 
.A(n_20095),
.Y(n_20154)
);

NAND2xp5_ASAP7_75t_L g20155 ( 
.A(n_20115),
.B(n_9103),
.Y(n_20155)
);

INVx1_ASAP7_75t_L g20156 ( 
.A(n_20100),
.Y(n_20156)
);

NOR2x1_ASAP7_75t_L g20157 ( 
.A(n_20025),
.B(n_5500),
.Y(n_20157)
);

INVx5_ASAP7_75t_L g20158 ( 
.A(n_20111),
.Y(n_20158)
);

INVx1_ASAP7_75t_SL g20159 ( 
.A(n_20068),
.Y(n_20159)
);

INVx1_ASAP7_75t_L g20160 ( 
.A(n_20116),
.Y(n_20160)
);

XOR2x2_ASAP7_75t_L g20161 ( 
.A(n_20071),
.B(n_6171),
.Y(n_20161)
);

NOR2xp33_ASAP7_75t_L g20162 ( 
.A(n_20063),
.B(n_5510),
.Y(n_20162)
);

INVx1_ASAP7_75t_L g20163 ( 
.A(n_20105),
.Y(n_20163)
);

INVx1_ASAP7_75t_L g20164 ( 
.A(n_20135),
.Y(n_20164)
);

NOR2x1_ASAP7_75t_L g20165 ( 
.A(n_20051),
.B(n_5510),
.Y(n_20165)
);

INVx1_ASAP7_75t_L g20166 ( 
.A(n_20124),
.Y(n_20166)
);

NOR2x1_ASAP7_75t_L g20167 ( 
.A(n_20085),
.B(n_5510),
.Y(n_20167)
);

NAND3xp33_ASAP7_75t_L g20168 ( 
.A(n_20050),
.B(n_5540),
.C(n_5510),
.Y(n_20168)
);

AND2x2_ASAP7_75t_SL g20169 ( 
.A(n_20060),
.B(n_5550),
.Y(n_20169)
);

NOR2x1_ASAP7_75t_L g20170 ( 
.A(n_20123),
.B(n_5540),
.Y(n_20170)
);

NAND4xp75_ASAP7_75t_L g20171 ( 
.A(n_20131),
.B(n_9112),
.C(n_9125),
.D(n_9103),
.Y(n_20171)
);

NAND4xp75_ASAP7_75t_L g20172 ( 
.A(n_20064),
.B(n_9125),
.C(n_9127),
.D(n_9112),
.Y(n_20172)
);

AND3x4_ASAP7_75t_L g20173 ( 
.A(n_20030),
.B(n_6963),
.C(n_6961),
.Y(n_20173)
);

NOR2x1p5_ASAP7_75t_L g20174 ( 
.A(n_20072),
.B(n_5540),
.Y(n_20174)
);

OAI22xp5_ASAP7_75t_L g20175 ( 
.A1(n_20097),
.A2(n_9125),
.B1(n_9127),
.B2(n_9112),
.Y(n_20175)
);

INVx1_ASAP7_75t_L g20176 ( 
.A(n_20122),
.Y(n_20176)
);

OR2x2_ASAP7_75t_L g20177 ( 
.A(n_20066),
.B(n_8704),
.Y(n_20177)
);

NOR2x1_ASAP7_75t_L g20178 ( 
.A(n_20076),
.B(n_5540),
.Y(n_20178)
);

INVx1_ASAP7_75t_L g20179 ( 
.A(n_20088),
.Y(n_20179)
);

OAI22xp5_ASAP7_75t_L g20180 ( 
.A1(n_20112),
.A2(n_9127),
.B1(n_9139),
.B2(n_9125),
.Y(n_20180)
);

INVx1_ASAP7_75t_L g20181 ( 
.A(n_20121),
.Y(n_20181)
);

OAI221xp5_ASAP7_75t_L g20182 ( 
.A1(n_20081),
.A2(n_5553),
.B1(n_5587),
.B2(n_5550),
.C(n_5540),
.Y(n_20182)
);

NOR3xp33_ASAP7_75t_L g20183 ( 
.A(n_20082),
.B(n_5994),
.C(n_5964),
.Y(n_20183)
);

XOR2xp5_ASAP7_75t_L g20184 ( 
.A(n_20096),
.B(n_5540),
.Y(n_20184)
);

NAND2x1p5_ASAP7_75t_L g20185 ( 
.A(n_20111),
.B(n_5550),
.Y(n_20185)
);

NAND2xp5_ASAP7_75t_L g20186 ( 
.A(n_20086),
.B(n_9127),
.Y(n_20186)
);

NOR2x1_ASAP7_75t_L g20187 ( 
.A(n_20062),
.B(n_5550),
.Y(n_20187)
);

INVxp33_ASAP7_75t_SL g20188 ( 
.A(n_20053),
.Y(n_20188)
);

AO22x2_ASAP7_75t_L g20189 ( 
.A1(n_20054),
.A2(n_9153),
.B1(n_9154),
.B2(n_9139),
.Y(n_20189)
);

NAND2xp5_ASAP7_75t_L g20190 ( 
.A(n_20102),
.B(n_9139),
.Y(n_20190)
);

INVx1_ASAP7_75t_L g20191 ( 
.A(n_20114),
.Y(n_20191)
);

AND2x4_ASAP7_75t_L g20192 ( 
.A(n_20107),
.B(n_6961),
.Y(n_20192)
);

NAND2xp5_ASAP7_75t_L g20193 ( 
.A(n_20120),
.B(n_9139),
.Y(n_20193)
);

INVx1_ASAP7_75t_L g20194 ( 
.A(n_20133),
.Y(n_20194)
);

NAND2xp5_ASAP7_75t_L g20195 ( 
.A(n_20092),
.B(n_20061),
.Y(n_20195)
);

AND3x4_ASAP7_75t_L g20196 ( 
.A(n_20084),
.B(n_6979),
.C(n_6963),
.Y(n_20196)
);

INVx1_ASAP7_75t_L g20197 ( 
.A(n_20069),
.Y(n_20197)
);

INVx1_ASAP7_75t_L g20198 ( 
.A(n_20040),
.Y(n_20198)
);

NAND2xp5_ASAP7_75t_L g20199 ( 
.A(n_20046),
.B(n_9153),
.Y(n_20199)
);

NOR2x1_ASAP7_75t_L g20200 ( 
.A(n_20029),
.B(n_5550),
.Y(n_20200)
);

NAND4xp75_ASAP7_75t_L g20201 ( 
.A(n_20037),
.B(n_9154),
.C(n_9159),
.D(n_9153),
.Y(n_20201)
);

NOR2x1_ASAP7_75t_L g20202 ( 
.A(n_20074),
.B(n_5550),
.Y(n_20202)
);

HB1xp67_ASAP7_75t_L g20203 ( 
.A(n_20079),
.Y(n_20203)
);

NAND4xp75_ASAP7_75t_L g20204 ( 
.A(n_20055),
.B(n_9154),
.C(n_9159),
.D(n_9153),
.Y(n_20204)
);

OAI22xp5_ASAP7_75t_L g20205 ( 
.A1(n_20109),
.A2(n_9159),
.B1(n_9182),
.B2(n_9154),
.Y(n_20205)
);

NOR2x1_ASAP7_75t_L g20206 ( 
.A(n_20057),
.B(n_5550),
.Y(n_20206)
);

NAND4xp75_ASAP7_75t_L g20207 ( 
.A(n_20027),
.B(n_9182),
.C(n_9184),
.D(n_9159),
.Y(n_20207)
);

INVx2_ASAP7_75t_SL g20208 ( 
.A(n_20045),
.Y(n_20208)
);

NAND2xp5_ASAP7_75t_L g20209 ( 
.A(n_20070),
.B(n_9182),
.Y(n_20209)
);

OAI22xp5_ASAP7_75t_L g20210 ( 
.A1(n_20089),
.A2(n_20073),
.B1(n_20048),
.B2(n_20126),
.Y(n_20210)
);

AO22x2_ASAP7_75t_L g20211 ( 
.A1(n_20090),
.A2(n_9184),
.B1(n_9188),
.B2(n_9182),
.Y(n_20211)
);

AND2x2_ASAP7_75t_L g20212 ( 
.A(n_20049),
.B(n_6963),
.Y(n_20212)
);

INVx3_ASAP7_75t_L g20213 ( 
.A(n_20119),
.Y(n_20213)
);

NOR2xp33_ASAP7_75t_L g20214 ( 
.A(n_20031),
.B(n_5550),
.Y(n_20214)
);

INVx1_ASAP7_75t_L g20215 ( 
.A(n_20108),
.Y(n_20215)
);

NAND4xp75_ASAP7_75t_L g20216 ( 
.A(n_20056),
.B(n_9188),
.C(n_9193),
.D(n_9184),
.Y(n_20216)
);

AND2x2_ASAP7_75t_L g20217 ( 
.A(n_20038),
.B(n_6979),
.Y(n_20217)
);

AO22x2_ASAP7_75t_L g20218 ( 
.A1(n_20091),
.A2(n_9188),
.B1(n_9193),
.B2(n_9184),
.Y(n_20218)
);

AND2x4_ASAP7_75t_L g20219 ( 
.A(n_20093),
.B(n_6979),
.Y(n_20219)
);

INVx1_ASAP7_75t_L g20220 ( 
.A(n_20083),
.Y(n_20220)
);

NOR2x1_ASAP7_75t_L g20221 ( 
.A(n_20043),
.B(n_5550),
.Y(n_20221)
);

AOI221xp5_ASAP7_75t_L g20222 ( 
.A1(n_20042),
.A2(n_9188),
.B1(n_9193),
.B2(n_9207),
.C(n_9194),
.Y(n_20222)
);

XNOR2x1_ASAP7_75t_L g20223 ( 
.A(n_20052),
.B(n_5553),
.Y(n_20223)
);

AOI22xp5_ASAP7_75t_L g20224 ( 
.A1(n_20125),
.A2(n_7803),
.B1(n_6960),
.B2(n_7014),
.Y(n_20224)
);

BUFx2_ASAP7_75t_L g20225 ( 
.A(n_20098),
.Y(n_20225)
);

NOR2xp67_ASAP7_75t_L g20226 ( 
.A(n_20132),
.B(n_5553),
.Y(n_20226)
);

NAND2x1p5_ASAP7_75t_SL g20227 ( 
.A(n_20127),
.B(n_5731),
.Y(n_20227)
);

INVx2_ASAP7_75t_SL g20228 ( 
.A(n_20059),
.Y(n_20228)
);

INVx2_ASAP7_75t_L g20229 ( 
.A(n_20036),
.Y(n_20229)
);

NOR2x1_ASAP7_75t_L g20230 ( 
.A(n_20026),
.B(n_20103),
.Y(n_20230)
);

OR2x2_ASAP7_75t_L g20231 ( 
.A(n_20118),
.B(n_8704),
.Y(n_20231)
);

AOI22xp5_ASAP7_75t_L g20232 ( 
.A1(n_20078),
.A2(n_7803),
.B1(n_6960),
.B2(n_7014),
.Y(n_20232)
);

NAND3xp33_ASAP7_75t_SL g20233 ( 
.A(n_20137),
.B(n_20080),
.C(n_20041),
.Y(n_20233)
);

INVx2_ASAP7_75t_L g20234 ( 
.A(n_20140),
.Y(n_20234)
);

NOR2xp67_ASAP7_75t_L g20235 ( 
.A(n_20208),
.B(n_20065),
.Y(n_20235)
);

NAND4xp25_ASAP7_75t_SL g20236 ( 
.A(n_20139),
.B(n_20117),
.C(n_20067),
.D(n_9194),
.Y(n_20236)
);

NAND3xp33_ASAP7_75t_L g20237 ( 
.A(n_20142),
.B(n_5587),
.C(n_5553),
.Y(n_20237)
);

AOI21xp5_ASAP7_75t_L g20238 ( 
.A1(n_20143),
.A2(n_9207),
.B(n_9193),
.Y(n_20238)
);

NOR4xp25_ASAP7_75t_L g20239 ( 
.A(n_20164),
.B(n_9207),
.C(n_9237),
.D(n_9194),
.Y(n_20239)
);

AND3x4_ASAP7_75t_L g20240 ( 
.A(n_20230),
.B(n_7031),
.C(n_7010),
.Y(n_20240)
);

NOR4xp25_ASAP7_75t_L g20241 ( 
.A(n_20154),
.B(n_20181),
.C(n_20150),
.D(n_20156),
.Y(n_20241)
);

NOR3xp33_ASAP7_75t_SL g20242 ( 
.A(n_20179),
.B(n_7089),
.C(n_7085),
.Y(n_20242)
);

AOI211xp5_ASAP7_75t_SL g20243 ( 
.A1(n_20163),
.A2(n_20191),
.B(n_20144),
.C(n_20147),
.Y(n_20243)
);

NAND3xp33_ASAP7_75t_L g20244 ( 
.A(n_20203),
.B(n_5587),
.C(n_5553),
.Y(n_20244)
);

NAND2xp5_ASAP7_75t_L g20245 ( 
.A(n_20136),
.B(n_9194),
.Y(n_20245)
);

NAND4xp75_ASAP7_75t_L g20246 ( 
.A(n_20176),
.B(n_5756),
.C(n_5741),
.D(n_9207),
.Y(n_20246)
);

OR2x6_ASAP7_75t_L g20247 ( 
.A(n_20138),
.B(n_5553),
.Y(n_20247)
);

NOR3xp33_ASAP7_75t_SL g20248 ( 
.A(n_20166),
.B(n_7085),
.C(n_7208),
.Y(n_20248)
);

NOR3xp33_ASAP7_75t_L g20249 ( 
.A(n_20159),
.B(n_6114),
.C(n_6074),
.Y(n_20249)
);

NAND4xp25_ASAP7_75t_SL g20250 ( 
.A(n_20152),
.B(n_9267),
.C(n_9237),
.D(n_7566),
.Y(n_20250)
);

NAND2xp5_ASAP7_75t_L g20251 ( 
.A(n_20226),
.B(n_9237),
.Y(n_20251)
);

INVx1_ASAP7_75t_L g20252 ( 
.A(n_20151),
.Y(n_20252)
);

NAND5xp2_ASAP7_75t_L g20253 ( 
.A(n_20188),
.B(n_7798),
.C(n_7868),
.D(n_7248),
.E(n_7245),
.Y(n_20253)
);

OAI221xp5_ASAP7_75t_SL g20254 ( 
.A1(n_20229),
.A2(n_7684),
.B1(n_7676),
.B2(n_7668),
.C(n_7412),
.Y(n_20254)
);

NOR3xp33_ASAP7_75t_SL g20255 ( 
.A(n_20145),
.B(n_20160),
.C(n_20197),
.Y(n_20255)
);

NOR3xp33_ASAP7_75t_L g20256 ( 
.A(n_20228),
.B(n_6114),
.C(n_6074),
.Y(n_20256)
);

AOI31xp33_ASAP7_75t_L g20257 ( 
.A1(n_20220),
.A2(n_5756),
.A3(n_7777),
.B(n_7738),
.Y(n_20257)
);

NOR4xp25_ASAP7_75t_L g20258 ( 
.A(n_20194),
.B(n_9267),
.C(n_7566),
.D(n_7583),
.Y(n_20258)
);

NAND3xp33_ASAP7_75t_SL g20259 ( 
.A(n_20225),
.B(n_6114),
.C(n_6074),
.Y(n_20259)
);

NOR3xp33_ASAP7_75t_L g20260 ( 
.A(n_20198),
.B(n_6114),
.C(n_6074),
.Y(n_20260)
);

NAND2xp5_ASAP7_75t_L g20261 ( 
.A(n_20169),
.B(n_20213),
.Y(n_20261)
);

NAND4xp25_ASAP7_75t_L g20262 ( 
.A(n_20215),
.B(n_20195),
.C(n_20214),
.D(n_20210),
.Y(n_20262)
);

NAND4xp25_ASAP7_75t_L g20263 ( 
.A(n_20221),
.B(n_20162),
.C(n_20165),
.D(n_20148),
.Y(n_20263)
);

NOR2xp33_ASAP7_75t_L g20264 ( 
.A(n_20158),
.B(n_20192),
.Y(n_20264)
);

INVx1_ASAP7_75t_L g20265 ( 
.A(n_20158),
.Y(n_20265)
);

INVx1_ASAP7_75t_L g20266 ( 
.A(n_20158),
.Y(n_20266)
);

NOR2x2_ASAP7_75t_L g20267 ( 
.A(n_20227),
.B(n_20184),
.Y(n_20267)
);

NOR3xp33_ASAP7_75t_L g20268 ( 
.A(n_20231),
.B(n_6114),
.C(n_6074),
.Y(n_20268)
);

AND5x1_ASAP7_75t_L g20269 ( 
.A(n_20153),
.B(n_8704),
.C(n_8716),
.D(n_9151),
.E(n_9067),
.Y(n_20269)
);

OR2x2_ASAP7_75t_L g20270 ( 
.A(n_20219),
.B(n_8704),
.Y(n_20270)
);

NOR3xp33_ASAP7_75t_L g20271 ( 
.A(n_20168),
.B(n_6121),
.C(n_6118),
.Y(n_20271)
);

AND2x4_ASAP7_75t_L g20272 ( 
.A(n_20174),
.B(n_20212),
.Y(n_20272)
);

NOR3xp33_ASAP7_75t_L g20273 ( 
.A(n_20217),
.B(n_6121),
.C(n_6118),
.Y(n_20273)
);

AND2x4_ASAP7_75t_L g20274 ( 
.A(n_20157),
.B(n_9267),
.Y(n_20274)
);

NAND2xp5_ASAP7_75t_L g20275 ( 
.A(n_20223),
.B(n_9267),
.Y(n_20275)
);

AOI21xp5_ASAP7_75t_L g20276 ( 
.A1(n_20190),
.A2(n_7409),
.B(n_7406),
.Y(n_20276)
);

AND4x1_ASAP7_75t_L g20277 ( 
.A(n_20202),
.B(n_7847),
.C(n_7870),
.D(n_7852),
.Y(n_20277)
);

AOI21xp5_ASAP7_75t_L g20278 ( 
.A1(n_20155),
.A2(n_7409),
.B(n_7406),
.Y(n_20278)
);

OAI211xp5_ASAP7_75t_SL g20279 ( 
.A1(n_20178),
.A2(n_5589),
.B(n_5393),
.C(n_5756),
.Y(n_20279)
);

NOR5xp2_ASAP7_75t_L g20280 ( 
.A(n_20182),
.B(n_7708),
.C(n_7712),
.D(n_7779),
.E(n_7752),
.Y(n_20280)
);

NOR3xp33_ASAP7_75t_SL g20281 ( 
.A(n_20199),
.B(n_7085),
.C(n_7208),
.Y(n_20281)
);

NAND4xp25_ASAP7_75t_L g20282 ( 
.A(n_20200),
.B(n_20170),
.C(n_20183),
.D(n_20187),
.Y(n_20282)
);

AND2x4_ASAP7_75t_L g20283 ( 
.A(n_20206),
.B(n_5553),
.Y(n_20283)
);

INVx2_ASAP7_75t_L g20284 ( 
.A(n_20185),
.Y(n_20284)
);

AND2x2_ASAP7_75t_L g20285 ( 
.A(n_20177),
.B(n_8716),
.Y(n_20285)
);

NAND4xp75_ASAP7_75t_L g20286 ( 
.A(n_20167),
.B(n_7615),
.C(n_7631),
.D(n_7629),
.Y(n_20286)
);

NOR3xp33_ASAP7_75t_L g20287 ( 
.A(n_20186),
.B(n_6121),
.C(n_6118),
.Y(n_20287)
);

OR2x2_ASAP7_75t_L g20288 ( 
.A(n_20161),
.B(n_8716),
.Y(n_20288)
);

NAND3xp33_ASAP7_75t_SL g20289 ( 
.A(n_20196),
.B(n_6121),
.C(n_6118),
.Y(n_20289)
);

OA22x2_ASAP7_75t_L g20290 ( 
.A1(n_20173),
.A2(n_9239),
.B1(n_9246),
.B2(n_9097),
.Y(n_20290)
);

NOR3xp33_ASAP7_75t_SL g20291 ( 
.A(n_20193),
.B(n_7229),
.C(n_7208),
.Y(n_20291)
);

INVx1_ASAP7_75t_L g20292 ( 
.A(n_20211),
.Y(n_20292)
);

AND2x4_ASAP7_75t_L g20293 ( 
.A(n_20149),
.B(n_5553),
.Y(n_20293)
);

NAND3xp33_ASAP7_75t_SL g20294 ( 
.A(n_20209),
.B(n_6121),
.C(n_6118),
.Y(n_20294)
);

NOR4xp25_ASAP7_75t_L g20295 ( 
.A(n_20141),
.B(n_7583),
.C(n_7584),
.D(n_7475),
.Y(n_20295)
);

OAI22xp5_ASAP7_75t_L g20296 ( 
.A1(n_20232),
.A2(n_20224),
.B1(n_20211),
.B2(n_20171),
.Y(n_20296)
);

NAND4xp75_ASAP7_75t_L g20297 ( 
.A(n_20222),
.B(n_20189),
.C(n_20146),
.D(n_20218),
.Y(n_20297)
);

NAND4xp75_ASAP7_75t_L g20298 ( 
.A(n_20189),
.B(n_7615),
.C(n_7631),
.D(n_7629),
.Y(n_20298)
);

NOR3xp33_ASAP7_75t_L g20299 ( 
.A(n_20207),
.B(n_20216),
.C(n_20172),
.Y(n_20299)
);

AOI211xp5_ASAP7_75t_L g20300 ( 
.A1(n_20175),
.A2(n_5587),
.B(n_5595),
.C(n_5553),
.Y(n_20300)
);

OA22x2_ASAP7_75t_L g20301 ( 
.A1(n_20180),
.A2(n_20205),
.B1(n_20218),
.B2(n_20201),
.Y(n_20301)
);

NOR3xp33_ASAP7_75t_L g20302 ( 
.A(n_20204),
.B(n_6140),
.C(n_6123),
.Y(n_20302)
);

NOR3xp33_ASAP7_75t_SL g20303 ( 
.A(n_20142),
.B(n_7229),
.C(n_7343),
.Y(n_20303)
);

AND2x2_ASAP7_75t_L g20304 ( 
.A(n_20137),
.B(n_8716),
.Y(n_20304)
);

NOR4xp25_ASAP7_75t_L g20305 ( 
.A(n_20142),
.B(n_7584),
.C(n_7597),
.D(n_7583),
.Y(n_20305)
);

CKINVDCx20_ASAP7_75t_R g20306 ( 
.A(n_20140),
.Y(n_20306)
);

NOR3xp33_ASAP7_75t_SL g20307 ( 
.A(n_20142),
.B(n_7229),
.C(n_7343),
.Y(n_20307)
);

NAND4xp25_ASAP7_75t_L g20308 ( 
.A(n_20142),
.B(n_6278),
.C(n_6290),
.D(n_6171),
.Y(n_20308)
);

INVx1_ASAP7_75t_L g20309 ( 
.A(n_20151),
.Y(n_20309)
);

NOR4xp25_ASAP7_75t_L g20310 ( 
.A(n_20142),
.B(n_7597),
.C(n_7602),
.D(n_7584),
.Y(n_20310)
);

CKINVDCx6p67_ASAP7_75t_R g20311 ( 
.A(n_20140),
.Y(n_20311)
);

AND2x2_ASAP7_75t_L g20312 ( 
.A(n_20137),
.B(n_8716),
.Y(n_20312)
);

OAI211xp5_ASAP7_75t_SL g20313 ( 
.A1(n_20137),
.A2(n_5234),
.B(n_5320),
.C(n_5237),
.Y(n_20313)
);

NAND3xp33_ASAP7_75t_SL g20314 ( 
.A(n_20137),
.B(n_6140),
.C(n_6123),
.Y(n_20314)
);

INVx1_ASAP7_75t_L g20315 ( 
.A(n_20151),
.Y(n_20315)
);

AND2x4_ASAP7_75t_L g20316 ( 
.A(n_20137),
.B(n_7010),
.Y(n_20316)
);

AND2x4_ASAP7_75t_L g20317 ( 
.A(n_20316),
.B(n_7010),
.Y(n_20317)
);

NOR2xp33_ASAP7_75t_L g20318 ( 
.A(n_20311),
.B(n_20234),
.Y(n_20318)
);

NAND4xp25_ASAP7_75t_L g20319 ( 
.A(n_20243),
.B(n_6290),
.C(n_6310),
.D(n_6278),
.Y(n_20319)
);

INVxp67_ASAP7_75t_SL g20320 ( 
.A(n_20265),
.Y(n_20320)
);

INVx1_ASAP7_75t_L g20321 ( 
.A(n_20266),
.Y(n_20321)
);

NAND5xp2_ASAP7_75t_L g20322 ( 
.A(n_20255),
.B(n_20264),
.C(n_20315),
.D(n_20309),
.E(n_20252),
.Y(n_20322)
);

AOI21xp5_ASAP7_75t_L g20323 ( 
.A1(n_20261),
.A2(n_5595),
.B(n_5587),
.Y(n_20323)
);

INVx1_ASAP7_75t_L g20324 ( 
.A(n_20306),
.Y(n_20324)
);

NAND4xp25_ASAP7_75t_L g20325 ( 
.A(n_20262),
.B(n_6290),
.C(n_6310),
.D(n_6278),
.Y(n_20325)
);

HB1xp67_ASAP7_75t_L g20326 ( 
.A(n_20235),
.Y(n_20326)
);

AND4x1_ASAP7_75t_L g20327 ( 
.A(n_20241),
.B(n_7852),
.C(n_7870),
.D(n_7847),
.Y(n_20327)
);

NOR3xp33_ASAP7_75t_L g20328 ( 
.A(n_20233),
.B(n_6140),
.C(n_6123),
.Y(n_20328)
);

NOR2x1p5_ASAP7_75t_L g20329 ( 
.A(n_20263),
.B(n_5587),
.Y(n_20329)
);

NAND2x1_ASAP7_75t_L g20330 ( 
.A(n_20272),
.B(n_5587),
.Y(n_20330)
);

NAND3xp33_ASAP7_75t_SL g20331 ( 
.A(n_20284),
.B(n_6140),
.C(n_6123),
.Y(n_20331)
);

OAI221xp5_ASAP7_75t_L g20332 ( 
.A1(n_20268),
.A2(n_5605),
.B1(n_5619),
.B2(n_5595),
.C(n_5587),
.Y(n_20332)
);

AOI22xp33_ASAP7_75t_L g20333 ( 
.A1(n_20237),
.A2(n_6960),
.B1(n_7014),
.B2(n_6916),
.Y(n_20333)
);

INVx1_ASAP7_75t_SL g20334 ( 
.A(n_20267),
.Y(n_20334)
);

XNOR2xp5_ASAP7_75t_L g20335 ( 
.A(n_20297),
.B(n_7738),
.Y(n_20335)
);

XOR2xp5_ASAP7_75t_L g20336 ( 
.A(n_20272),
.B(n_20282),
.Y(n_20336)
);

OAI22xp5_ASAP7_75t_L g20337 ( 
.A1(n_20247),
.A2(n_5595),
.B1(n_5605),
.B2(n_5587),
.Y(n_20337)
);

OAI211xp5_ASAP7_75t_SL g20338 ( 
.A1(n_20292),
.A2(n_5237),
.B(n_5343),
.C(n_5320),
.Y(n_20338)
);

AOI21xp5_ASAP7_75t_L g20339 ( 
.A1(n_20296),
.A2(n_5605),
.B(n_5595),
.Y(n_20339)
);

AO22x2_ASAP7_75t_L g20340 ( 
.A1(n_20299),
.A2(n_20289),
.B1(n_20240),
.B2(n_20245),
.Y(n_20340)
);

OAI211xp5_ASAP7_75t_L g20341 ( 
.A1(n_20305),
.A2(n_5605),
.B(n_5619),
.C(n_5595),
.Y(n_20341)
);

INVx5_ASAP7_75t_L g20342 ( 
.A(n_20247),
.Y(n_20342)
);

NOR2x1p5_ASAP7_75t_L g20343 ( 
.A(n_20308),
.B(n_5595),
.Y(n_20343)
);

NAND4xp25_ASAP7_75t_L g20344 ( 
.A(n_20251),
.B(n_6290),
.C(n_6310),
.D(n_6278),
.Y(n_20344)
);

AOI31xp33_ASAP7_75t_L g20345 ( 
.A1(n_20304),
.A2(n_7777),
.A3(n_7781),
.B(n_7738),
.Y(n_20345)
);

INVx2_ASAP7_75t_L g20346 ( 
.A(n_20301),
.Y(n_20346)
);

HB1xp67_ASAP7_75t_L g20347 ( 
.A(n_20236),
.Y(n_20347)
);

AOI22xp5_ASAP7_75t_L g20348 ( 
.A1(n_20312),
.A2(n_20273),
.B1(n_20260),
.B2(n_20244),
.Y(n_20348)
);

NOR3xp33_ASAP7_75t_SL g20349 ( 
.A(n_20294),
.B(n_7357),
.C(n_7349),
.Y(n_20349)
);

NAND3xp33_ASAP7_75t_L g20350 ( 
.A(n_20303),
.B(n_5605),
.C(n_5595),
.Y(n_20350)
);

NOR3xp33_ASAP7_75t_L g20351 ( 
.A(n_20275),
.B(n_6140),
.C(n_6123),
.Y(n_20351)
);

XOR2xp5_ASAP7_75t_L g20352 ( 
.A(n_20288),
.B(n_5595),
.Y(n_20352)
);

AOI211xp5_ASAP7_75t_L g20353 ( 
.A1(n_20310),
.A2(n_5641),
.B(n_5673),
.C(n_5619),
.Y(n_20353)
);

AOI22xp5_ASAP7_75t_L g20354 ( 
.A1(n_20307),
.A2(n_5641),
.B1(n_5673),
.B2(n_5619),
.Y(n_20354)
);

HB1xp67_ASAP7_75t_L g20355 ( 
.A(n_20293),
.Y(n_20355)
);

INVx1_ASAP7_75t_L g20356 ( 
.A(n_20283),
.Y(n_20356)
);

NAND4xp25_ASAP7_75t_L g20357 ( 
.A(n_20238),
.B(n_6572),
.C(n_6606),
.D(n_6310),
.Y(n_20357)
);

AOI211xp5_ASAP7_75t_SL g20358 ( 
.A1(n_20249),
.A2(n_5320),
.B(n_5343),
.C(n_5237),
.Y(n_20358)
);

NAND2xp5_ASAP7_75t_L g20359 ( 
.A(n_20242),
.B(n_8716),
.Y(n_20359)
);

NOR3xp33_ASAP7_75t_L g20360 ( 
.A(n_20259),
.B(n_20314),
.C(n_20287),
.Y(n_20360)
);

INVx2_ASAP7_75t_L g20361 ( 
.A(n_20283),
.Y(n_20361)
);

NOR4xp25_ASAP7_75t_L g20362 ( 
.A(n_20279),
.B(n_7602),
.C(n_7638),
.D(n_7597),
.Y(n_20362)
);

AND2x4_ASAP7_75t_L g20363 ( 
.A(n_20248),
.B(n_7010),
.Y(n_20363)
);

INVx1_ASAP7_75t_L g20364 ( 
.A(n_20293),
.Y(n_20364)
);

OAI211xp5_ASAP7_75t_L g20365 ( 
.A1(n_20295),
.A2(n_5641),
.B(n_5673),
.C(n_5619),
.Y(n_20365)
);

OAI222xp33_ASAP7_75t_L g20366 ( 
.A1(n_20276),
.A2(n_7867),
.B1(n_7795),
.B2(n_7903),
.C1(n_7857),
.C2(n_7722),
.Y(n_20366)
);

XNOR2xp5_ASAP7_75t_L g20367 ( 
.A(n_20300),
.B(n_7738),
.Y(n_20367)
);

NOR3xp33_ASAP7_75t_L g20368 ( 
.A(n_20256),
.B(n_6572),
.C(n_6310),
.Y(n_20368)
);

AND2x2_ASAP7_75t_L g20369 ( 
.A(n_20281),
.B(n_8716),
.Y(n_20369)
);

AND2x4_ASAP7_75t_L g20370 ( 
.A(n_20291),
.B(n_7031),
.Y(n_20370)
);

AND4x1_ASAP7_75t_L g20371 ( 
.A(n_20258),
.B(n_7852),
.C(n_7870),
.D(n_7847),
.Y(n_20371)
);

OA21x2_ASAP7_75t_L g20372 ( 
.A1(n_20274),
.A2(n_8532),
.B(n_8510),
.Y(n_20372)
);

INVx2_ASAP7_75t_L g20373 ( 
.A(n_20274),
.Y(n_20373)
);

INVx1_ASAP7_75t_L g20374 ( 
.A(n_20298),
.Y(n_20374)
);

AOI22xp33_ASAP7_75t_L g20375 ( 
.A1(n_20271),
.A2(n_6960),
.B1(n_7014),
.B2(n_6916),
.Y(n_20375)
);

INVx1_ASAP7_75t_L g20376 ( 
.A(n_20286),
.Y(n_20376)
);

NOR3xp33_ASAP7_75t_L g20377 ( 
.A(n_20250),
.B(n_6606),
.C(n_6572),
.Y(n_20377)
);

HB1xp67_ASAP7_75t_L g20378 ( 
.A(n_20246),
.Y(n_20378)
);

AOI22xp5_ASAP7_75t_L g20379 ( 
.A1(n_20285),
.A2(n_20302),
.B1(n_20278),
.B2(n_20313),
.Y(n_20379)
);

NOR3x2_ASAP7_75t_L g20380 ( 
.A(n_20280),
.B(n_5901),
.C(n_5641),
.Y(n_20380)
);

NAND4xp25_ASAP7_75t_L g20381 ( 
.A(n_20253),
.B(n_6606),
.C(n_6608),
.D(n_6572),
.Y(n_20381)
);

AOI22xp33_ASAP7_75t_L g20382 ( 
.A1(n_20270),
.A2(n_6960),
.B1(n_7018),
.B2(n_7014),
.Y(n_20382)
);

AND2x2_ASAP7_75t_L g20383 ( 
.A(n_20277),
.B(n_7031),
.Y(n_20383)
);

INVx1_ASAP7_75t_L g20384 ( 
.A(n_20257),
.Y(n_20384)
);

INVx1_ASAP7_75t_L g20385 ( 
.A(n_20239),
.Y(n_20385)
);

A2O1A1Ixp33_ASAP7_75t_L g20386 ( 
.A1(n_20318),
.A2(n_20254),
.B(n_20269),
.C(n_20290),
.Y(n_20386)
);

AOI221xp5_ASAP7_75t_L g20387 ( 
.A1(n_20320),
.A2(n_5673),
.B1(n_5678),
.B2(n_5641),
.C(n_5619),
.Y(n_20387)
);

OAI221xp5_ASAP7_75t_L g20388 ( 
.A1(n_20324),
.A2(n_5673),
.B1(n_5678),
.B2(n_5641),
.C(n_5619),
.Y(n_20388)
);

AOI22xp5_ASAP7_75t_L g20389 ( 
.A1(n_20326),
.A2(n_5641),
.B1(n_5673),
.B2(n_5619),
.Y(n_20389)
);

INVx3_ASAP7_75t_L g20390 ( 
.A(n_20346),
.Y(n_20390)
);

HB1xp67_ASAP7_75t_L g20391 ( 
.A(n_20321),
.Y(n_20391)
);

INVx1_ASAP7_75t_L g20392 ( 
.A(n_20335),
.Y(n_20392)
);

INVx2_ASAP7_75t_L g20393 ( 
.A(n_20361),
.Y(n_20393)
);

NAND2x1_ASAP7_75t_SL g20394 ( 
.A(n_20347),
.B(n_20355),
.Y(n_20394)
);

AOI31xp33_ASAP7_75t_L g20395 ( 
.A1(n_20334),
.A2(n_7777),
.A3(n_7781),
.B(n_7738),
.Y(n_20395)
);

OAI22xp33_ASAP7_75t_L g20396 ( 
.A1(n_20376),
.A2(n_5641),
.B1(n_5673),
.B2(n_5619),
.Y(n_20396)
);

NAND2xp5_ASAP7_75t_L g20397 ( 
.A(n_20329),
.B(n_5641),
.Y(n_20397)
);

AOI21xp33_ASAP7_75t_SL g20398 ( 
.A1(n_20374),
.A2(n_8287),
.B(n_8286),
.Y(n_20398)
);

INVx1_ASAP7_75t_L g20399 ( 
.A(n_20336),
.Y(n_20399)
);

INVx2_ASAP7_75t_L g20400 ( 
.A(n_20373),
.Y(n_20400)
);

NAND2xp5_ASAP7_75t_L g20401 ( 
.A(n_20384),
.B(n_5673),
.Y(n_20401)
);

NAND3xp33_ASAP7_75t_SL g20402 ( 
.A(n_20364),
.B(n_6606),
.C(n_6572),
.Y(n_20402)
);

NAND4xp25_ASAP7_75t_L g20403 ( 
.A(n_20322),
.B(n_20385),
.C(n_20348),
.D(n_20379),
.Y(n_20403)
);

AO22x2_ASAP7_75t_L g20404 ( 
.A1(n_20356),
.A2(n_6608),
.B1(n_6629),
.B2(n_6606),
.Y(n_20404)
);

XOR2xp5_ASAP7_75t_L g20405 ( 
.A(n_20340),
.B(n_5673),
.Y(n_20405)
);

OAI22xp5_ASAP7_75t_L g20406 ( 
.A1(n_20352),
.A2(n_5707),
.B1(n_5711),
.B2(n_5678),
.Y(n_20406)
);

INVx2_ASAP7_75t_L g20407 ( 
.A(n_20340),
.Y(n_20407)
);

NOR2xp33_ASAP7_75t_R g20408 ( 
.A(n_20342),
.B(n_5678),
.Y(n_20408)
);

INVx1_ASAP7_75t_L g20409 ( 
.A(n_20378),
.Y(n_20409)
);

INVxp33_ASAP7_75t_L g20410 ( 
.A(n_20360),
.Y(n_20410)
);

AOI22xp5_ASAP7_75t_L g20411 ( 
.A1(n_20328),
.A2(n_5707),
.B1(n_5711),
.B2(n_5678),
.Y(n_20411)
);

NOR2xp67_ASAP7_75t_L g20412 ( 
.A(n_20342),
.B(n_5678),
.Y(n_20412)
);

INVx1_ASAP7_75t_L g20413 ( 
.A(n_20342),
.Y(n_20413)
);

AOI22xp5_ASAP7_75t_L g20414 ( 
.A1(n_20317),
.A2(n_5707),
.B1(n_5711),
.B2(n_5678),
.Y(n_20414)
);

AOI211x1_ASAP7_75t_L g20415 ( 
.A1(n_20365),
.A2(n_7376),
.B(n_7388),
.C(n_7365),
.Y(n_20415)
);

INVx1_ASAP7_75t_L g20416 ( 
.A(n_20380),
.Y(n_20416)
);

NOR2x1_ASAP7_75t_L g20417 ( 
.A(n_20330),
.B(n_5678),
.Y(n_20417)
);

OAI21xp33_ASAP7_75t_L g20418 ( 
.A1(n_20339),
.A2(n_20381),
.B(n_20363),
.Y(n_20418)
);

NOR2x1p5_ASAP7_75t_L g20419 ( 
.A(n_20370),
.B(n_5678),
.Y(n_20419)
);

OAI221xp5_ASAP7_75t_SL g20420 ( 
.A1(n_20375),
.A2(n_7406),
.B1(n_7437),
.B2(n_7412),
.C(n_7409),
.Y(n_20420)
);

INVx2_ASAP7_75t_L g20421 ( 
.A(n_20343),
.Y(n_20421)
);

HB1xp67_ASAP7_75t_L g20422 ( 
.A(n_20383),
.Y(n_20422)
);

XNOR2xp5_ASAP7_75t_L g20423 ( 
.A(n_20353),
.B(n_7777),
.Y(n_20423)
);

INVx1_ASAP7_75t_L g20424 ( 
.A(n_20341),
.Y(n_20424)
);

NAND2xp5_ASAP7_75t_L g20425 ( 
.A(n_20377),
.B(n_5707),
.Y(n_20425)
);

AOI221xp5_ASAP7_75t_L g20426 ( 
.A1(n_20362),
.A2(n_5716),
.B1(n_5717),
.B2(n_5711),
.C(n_5707),
.Y(n_20426)
);

HB1xp67_ASAP7_75t_L g20427 ( 
.A(n_20367),
.Y(n_20427)
);

OAI22xp5_ASAP7_75t_L g20428 ( 
.A1(n_20332),
.A2(n_5711),
.B1(n_5716),
.B2(n_5707),
.Y(n_20428)
);

INVx2_ASAP7_75t_L g20429 ( 
.A(n_20369),
.Y(n_20429)
);

INVx2_ASAP7_75t_L g20430 ( 
.A(n_20359),
.Y(n_20430)
);

AOI32xp33_ASAP7_75t_L g20431 ( 
.A1(n_20368),
.A2(n_6682),
.A3(n_6742),
.B1(n_6629),
.B2(n_6608),
.Y(n_20431)
);

INVx2_ASAP7_75t_SL g20432 ( 
.A(n_20371),
.Y(n_20432)
);

OAI22xp33_ASAP7_75t_R g20433 ( 
.A1(n_20349),
.A2(n_7402),
.B1(n_7323),
.B2(n_7278),
.Y(n_20433)
);

NAND4xp25_ASAP7_75t_SL g20434 ( 
.A(n_20323),
.B(n_7638),
.C(n_7602),
.D(n_7376),
.Y(n_20434)
);

OAI22xp5_ASAP7_75t_L g20435 ( 
.A1(n_20350),
.A2(n_5711),
.B1(n_5716),
.B2(n_5707),
.Y(n_20435)
);

NAND2xp5_ASAP7_75t_SL g20436 ( 
.A(n_20351),
.B(n_5707),
.Y(n_20436)
);

INVx2_ASAP7_75t_L g20437 ( 
.A(n_20354),
.Y(n_20437)
);

NAND5xp2_ASAP7_75t_L g20438 ( 
.A(n_20358),
.B(n_7798),
.C(n_7868),
.D(n_7248),
.E(n_7245),
.Y(n_20438)
);

INVx2_ASAP7_75t_SL g20439 ( 
.A(n_20327),
.Y(n_20439)
);

HB1xp67_ASAP7_75t_L g20440 ( 
.A(n_20331),
.Y(n_20440)
);

NAND2xp5_ASAP7_75t_L g20441 ( 
.A(n_20357),
.B(n_5711),
.Y(n_20441)
);

AOI21xp5_ASAP7_75t_SL g20442 ( 
.A1(n_20337),
.A2(n_5716),
.B(n_5711),
.Y(n_20442)
);

OAI22xp5_ASAP7_75t_L g20443 ( 
.A1(n_20382),
.A2(n_5716),
.B1(n_5717),
.B2(n_5711),
.Y(n_20443)
);

NAND3xp33_ASAP7_75t_SL g20444 ( 
.A(n_20333),
.B(n_6629),
.C(n_6608),
.Y(n_20444)
);

INVx1_ASAP7_75t_L g20445 ( 
.A(n_20391),
.Y(n_20445)
);

OAI22xp5_ASAP7_75t_SL g20446 ( 
.A1(n_20399),
.A2(n_20319),
.B1(n_20325),
.B2(n_20338),
.Y(n_20446)
);

INVx1_ASAP7_75t_L g20447 ( 
.A(n_20390),
.Y(n_20447)
);

INVx1_ASAP7_75t_L g20448 ( 
.A(n_20390),
.Y(n_20448)
);

XNOR2xp5_ASAP7_75t_L g20449 ( 
.A(n_20403),
.B(n_20344),
.Y(n_20449)
);

INVx1_ASAP7_75t_L g20450 ( 
.A(n_20405),
.Y(n_20450)
);

XOR2xp5_ASAP7_75t_L g20451 ( 
.A(n_20410),
.B(n_20345),
.Y(n_20451)
);

INVx2_ASAP7_75t_SL g20452 ( 
.A(n_20394),
.Y(n_20452)
);

INVx1_ASAP7_75t_L g20453 ( 
.A(n_20413),
.Y(n_20453)
);

AOI22x1_ASAP7_75t_L g20454 ( 
.A1(n_20393),
.A2(n_20366),
.B1(n_20372),
.B2(n_5717),
.Y(n_20454)
);

INVx2_ASAP7_75t_L g20455 ( 
.A(n_20419),
.Y(n_20455)
);

INVx1_ASAP7_75t_L g20456 ( 
.A(n_20416),
.Y(n_20456)
);

NOR2xp33_ASAP7_75t_SL g20457 ( 
.A(n_20400),
.B(n_5716),
.Y(n_20457)
);

INVx1_ASAP7_75t_L g20458 ( 
.A(n_20422),
.Y(n_20458)
);

INVx1_ASAP7_75t_L g20459 ( 
.A(n_20407),
.Y(n_20459)
);

INVx1_ASAP7_75t_L g20460 ( 
.A(n_20392),
.Y(n_20460)
);

INVx1_ASAP7_75t_L g20461 ( 
.A(n_20409),
.Y(n_20461)
);

XNOR2xp5_ASAP7_75t_SL g20462 ( 
.A(n_20427),
.B(n_20372),
.Y(n_20462)
);

AOI22xp5_ASAP7_75t_L g20463 ( 
.A1(n_20401),
.A2(n_5717),
.B1(n_5716),
.B2(n_6916),
.Y(n_20463)
);

XOR2xp5_ASAP7_75t_L g20464 ( 
.A(n_20440),
.B(n_5716),
.Y(n_20464)
);

NAND2xp33_ASAP7_75t_L g20465 ( 
.A(n_20429),
.B(n_20386),
.Y(n_20465)
);

NOR2xp33_ASAP7_75t_L g20466 ( 
.A(n_20418),
.B(n_5716),
.Y(n_20466)
);

NAND2xp5_ASAP7_75t_L g20467 ( 
.A(n_20439),
.B(n_5717),
.Y(n_20467)
);

INVx1_ASAP7_75t_L g20468 ( 
.A(n_20432),
.Y(n_20468)
);

INVx2_ASAP7_75t_L g20469 ( 
.A(n_20421),
.Y(n_20469)
);

INVx1_ASAP7_75t_L g20470 ( 
.A(n_20424),
.Y(n_20470)
);

INVx1_ASAP7_75t_L g20471 ( 
.A(n_20437),
.Y(n_20471)
);

INVx1_ASAP7_75t_L g20472 ( 
.A(n_20430),
.Y(n_20472)
);

XNOR2x1_ASAP7_75t_L g20473 ( 
.A(n_20423),
.B(n_5717),
.Y(n_20473)
);

OAI22xp5_ASAP7_75t_L g20474 ( 
.A1(n_20397),
.A2(n_5717),
.B1(n_7705),
.B2(n_7487),
.Y(n_20474)
);

AOI22xp5_ASAP7_75t_L g20475 ( 
.A1(n_20412),
.A2(n_5717),
.B1(n_6960),
.B2(n_6916),
.Y(n_20475)
);

INVx1_ASAP7_75t_L g20476 ( 
.A(n_20425),
.Y(n_20476)
);

AOI22xp5_ASAP7_75t_L g20477 ( 
.A1(n_20441),
.A2(n_6960),
.B1(n_7014),
.B2(n_6916),
.Y(n_20477)
);

INVx4_ASAP7_75t_L g20478 ( 
.A(n_20408),
.Y(n_20478)
);

INVx1_ASAP7_75t_L g20479 ( 
.A(n_20417),
.Y(n_20479)
);

AOI22xp5_ASAP7_75t_L g20480 ( 
.A1(n_20444),
.A2(n_7014),
.B1(n_7018),
.B2(n_6916),
.Y(n_20480)
);

INVxp67_ASAP7_75t_SL g20481 ( 
.A(n_20436),
.Y(n_20481)
);

INVx1_ASAP7_75t_SL g20482 ( 
.A(n_20389),
.Y(n_20482)
);

INVx1_ASAP7_75t_L g20483 ( 
.A(n_20442),
.Y(n_20483)
);

INVx1_ASAP7_75t_L g20484 ( 
.A(n_20396),
.Y(n_20484)
);

XOR2xp5_ASAP7_75t_L g20485 ( 
.A(n_20402),
.B(n_5965),
.Y(n_20485)
);

INVx1_ASAP7_75t_L g20486 ( 
.A(n_20415),
.Y(n_20486)
);

INVxp67_ASAP7_75t_L g20487 ( 
.A(n_20434),
.Y(n_20487)
);

BUFx2_ASAP7_75t_L g20488 ( 
.A(n_20452),
.Y(n_20488)
);

NOR2x1p5_ASAP7_75t_L g20489 ( 
.A(n_20445),
.B(n_20438),
.Y(n_20489)
);

AOI22xp33_ASAP7_75t_SL g20490 ( 
.A1(n_20447),
.A2(n_20428),
.B1(n_20406),
.B2(n_20435),
.Y(n_20490)
);

INVxp67_ASAP7_75t_SL g20491 ( 
.A(n_20459),
.Y(n_20491)
);

INVx3_ASAP7_75t_L g20492 ( 
.A(n_20448),
.Y(n_20492)
);

HB1xp67_ASAP7_75t_L g20493 ( 
.A(n_20461),
.Y(n_20493)
);

BUFx10_ASAP7_75t_L g20494 ( 
.A(n_20453),
.Y(n_20494)
);

BUFx2_ASAP7_75t_L g20495 ( 
.A(n_20458),
.Y(n_20495)
);

INVx1_ASAP7_75t_L g20496 ( 
.A(n_20462),
.Y(n_20496)
);

BUFx6f_ASAP7_75t_L g20497 ( 
.A(n_20469),
.Y(n_20497)
);

INVx1_ASAP7_75t_SL g20498 ( 
.A(n_20468),
.Y(n_20498)
);

INVx1_ASAP7_75t_L g20499 ( 
.A(n_20471),
.Y(n_20499)
);

INVx1_ASAP7_75t_L g20500 ( 
.A(n_20456),
.Y(n_20500)
);

INVx2_ASAP7_75t_L g20501 ( 
.A(n_20454),
.Y(n_20501)
);

AOI22xp33_ASAP7_75t_L g20502 ( 
.A1(n_20470),
.A2(n_20426),
.B1(n_20433),
.B2(n_20411),
.Y(n_20502)
);

OAI31xp67_ASAP7_75t_L g20503 ( 
.A1(n_20455),
.A2(n_20431),
.A3(n_20395),
.B(n_20420),
.Y(n_20503)
);

NAND2xp5_ASAP7_75t_L g20504 ( 
.A(n_20457),
.B(n_20387),
.Y(n_20504)
);

INVx4_ASAP7_75t_L g20505 ( 
.A(n_20478),
.Y(n_20505)
);

INVx2_ASAP7_75t_L g20506 ( 
.A(n_20478),
.Y(n_20506)
);

INVx2_ASAP7_75t_SL g20507 ( 
.A(n_20460),
.Y(n_20507)
);

OAI22xp5_ASAP7_75t_SL g20508 ( 
.A1(n_20451),
.A2(n_20388),
.B1(n_20414),
.B2(n_20443),
.Y(n_20508)
);

XNOR2xp5_ASAP7_75t_L g20509 ( 
.A(n_20449),
.B(n_20404),
.Y(n_20509)
);

NOR2x1_ASAP7_75t_L g20510 ( 
.A(n_20465),
.B(n_20404),
.Y(n_20510)
);

AOI21xp5_ASAP7_75t_L g20511 ( 
.A1(n_20472),
.A2(n_20398),
.B(n_7409),
.Y(n_20511)
);

OAI22xp5_ASAP7_75t_L g20512 ( 
.A1(n_20464),
.A2(n_7014),
.B1(n_7018),
.B2(n_6916),
.Y(n_20512)
);

CKINVDCx20_ASAP7_75t_R g20513 ( 
.A(n_20446),
.Y(n_20513)
);

HB1xp67_ASAP7_75t_L g20514 ( 
.A(n_20487),
.Y(n_20514)
);

INVx1_ASAP7_75t_L g20515 ( 
.A(n_20479),
.Y(n_20515)
);

INVx1_ASAP7_75t_L g20516 ( 
.A(n_20486),
.Y(n_20516)
);

OAI211xp5_ASAP7_75t_L g20517 ( 
.A1(n_20450),
.A2(n_6608),
.B(n_6682),
.C(n_6629),
.Y(n_20517)
);

AOI211xp5_ASAP7_75t_L g20518 ( 
.A1(n_20498),
.A2(n_20499),
.B(n_20500),
.C(n_20496),
.Y(n_20518)
);

NOR2x1_ASAP7_75t_L g20519 ( 
.A(n_20510),
.B(n_20488),
.Y(n_20519)
);

INVx1_ASAP7_75t_SL g20520 ( 
.A(n_20495),
.Y(n_20520)
);

INVxp67_ASAP7_75t_SL g20521 ( 
.A(n_20493),
.Y(n_20521)
);

INVx1_ASAP7_75t_L g20522 ( 
.A(n_20491),
.Y(n_20522)
);

INVx1_ASAP7_75t_L g20523 ( 
.A(n_20494),
.Y(n_20523)
);

NOR4xp75_ASAP7_75t_L g20524 ( 
.A(n_20507),
.B(n_20467),
.C(n_20481),
.D(n_20476),
.Y(n_20524)
);

NOR4xp25_ASAP7_75t_L g20525 ( 
.A(n_20515),
.B(n_20516),
.C(n_20492),
.D(n_20506),
.Y(n_20525)
);

INVx1_ASAP7_75t_L g20526 ( 
.A(n_20497),
.Y(n_20526)
);

OAI321xp33_ASAP7_75t_L g20527 ( 
.A1(n_20497),
.A2(n_20484),
.A3(n_20483),
.B1(n_20466),
.B2(n_20480),
.C(n_20474),
.Y(n_20527)
);

AND2x2_ASAP7_75t_L g20528 ( 
.A(n_20514),
.B(n_20505),
.Y(n_20528)
);

INVxp67_ASAP7_75t_SL g20529 ( 
.A(n_20489),
.Y(n_20529)
);

NAND3xp33_ASAP7_75t_SL g20530 ( 
.A(n_20513),
.B(n_20482),
.C(n_20485),
.Y(n_20530)
);

HB1xp67_ASAP7_75t_L g20531 ( 
.A(n_20501),
.Y(n_20531)
);

AND3x4_ASAP7_75t_L g20532 ( 
.A(n_20503),
.B(n_20473),
.C(n_20477),
.Y(n_20532)
);

OR2x2_ASAP7_75t_L g20533 ( 
.A(n_20502),
.B(n_20475),
.Y(n_20533)
);

XNOR2xp5_ASAP7_75t_L g20534 ( 
.A(n_20509),
.B(n_20463),
.Y(n_20534)
);

AOI22xp5_ASAP7_75t_L g20535 ( 
.A1(n_20508),
.A2(n_7018),
.B1(n_7050),
.B2(n_6916),
.Y(n_20535)
);

OAI221xp5_ASAP7_75t_L g20536 ( 
.A1(n_20490),
.A2(n_5814),
.B1(n_5827),
.B2(n_5784),
.C(n_5780),
.Y(n_20536)
);

NAND2xp5_ASAP7_75t_L g20537 ( 
.A(n_20504),
.B(n_7798),
.Y(n_20537)
);

OAI22xp5_ASAP7_75t_SL g20538 ( 
.A1(n_20520),
.A2(n_20511),
.B1(n_20512),
.B2(n_20517),
.Y(n_20538)
);

INVx2_ASAP7_75t_L g20539 ( 
.A(n_20528),
.Y(n_20539)
);

INVx2_ASAP7_75t_L g20540 ( 
.A(n_20519),
.Y(n_20540)
);

AOI22xp5_ASAP7_75t_L g20541 ( 
.A1(n_20521),
.A2(n_5784),
.B1(n_5814),
.B2(n_5780),
.Y(n_20541)
);

AO22x2_ASAP7_75t_L g20542 ( 
.A1(n_20532),
.A2(n_7868),
.B1(n_7798),
.B2(n_6682),
.Y(n_20542)
);

XOR2x2_ASAP7_75t_L g20543 ( 
.A(n_20518),
.B(n_6629),
.Y(n_20543)
);

OAI21xp5_ASAP7_75t_L g20544 ( 
.A1(n_20525),
.A2(n_8290),
.B(n_8365),
.Y(n_20544)
);

INVx1_ASAP7_75t_L g20545 ( 
.A(n_20522),
.Y(n_20545)
);

NAND2xp5_ASAP7_75t_SL g20546 ( 
.A(n_20523),
.B(n_5780),
.Y(n_20546)
);

INVx1_ASAP7_75t_L g20547 ( 
.A(n_20531),
.Y(n_20547)
);

INVx1_ASAP7_75t_L g20548 ( 
.A(n_20526),
.Y(n_20548)
);

INVx2_ASAP7_75t_L g20549 ( 
.A(n_20533),
.Y(n_20549)
);

AO22x2_ASAP7_75t_L g20550 ( 
.A1(n_20530),
.A2(n_7868),
.B1(n_7798),
.B2(n_6742),
.Y(n_20550)
);

INVx1_ASAP7_75t_L g20551 ( 
.A(n_20529),
.Y(n_20551)
);

OAI22xp5_ASAP7_75t_SL g20552 ( 
.A1(n_20534),
.A2(n_5784),
.B1(n_5814),
.B2(n_5780),
.Y(n_20552)
);

AND2x2_ASAP7_75t_SL g20553 ( 
.A(n_20540),
.B(n_20524),
.Y(n_20553)
);

NAND5xp2_ASAP7_75t_L g20554 ( 
.A(n_20551),
.B(n_20527),
.C(n_20537),
.D(n_20535),
.E(n_20536),
.Y(n_20554)
);

OA22x2_ASAP7_75t_L g20555 ( 
.A1(n_20547),
.A2(n_8532),
.B1(n_7409),
.B2(n_7412),
.Y(n_20555)
);

NOR2xp67_ASAP7_75t_L g20556 ( 
.A(n_20539),
.B(n_6682),
.Y(n_20556)
);

NAND4xp25_ASAP7_75t_L g20557 ( 
.A(n_20548),
.B(n_6742),
.C(n_6791),
.D(n_6682),
.Y(n_20557)
);

OAI22xp5_ASAP7_75t_L g20558 ( 
.A1(n_20549),
.A2(n_5814),
.B1(n_5827),
.B2(n_5784),
.Y(n_20558)
);

AOI22xp33_ASAP7_75t_L g20559 ( 
.A1(n_20545),
.A2(n_7018),
.B1(n_7050),
.B2(n_6916),
.Y(n_20559)
);

INVx2_ASAP7_75t_L g20560 ( 
.A(n_20543),
.Y(n_20560)
);

AOI21xp33_ASAP7_75t_L g20561 ( 
.A1(n_20538),
.A2(n_5814),
.B(n_5784),
.Y(n_20561)
);

OR2x2_ASAP7_75t_L g20562 ( 
.A(n_20546),
.B(n_7406),
.Y(n_20562)
);

AOI22xp33_ASAP7_75t_SL g20563 ( 
.A1(n_20553),
.A2(n_20544),
.B1(n_20552),
.B2(n_20550),
.Y(n_20563)
);

AOI22xp33_ASAP7_75t_L g20564 ( 
.A1(n_20560),
.A2(n_20541),
.B1(n_20542),
.B2(n_7050),
.Y(n_20564)
);

INVx1_ASAP7_75t_L g20565 ( 
.A(n_20554),
.Y(n_20565)
);

XNOR2xp5_ASAP7_75t_L g20566 ( 
.A(n_20556),
.B(n_20562),
.Y(n_20566)
);

OAI21xp5_ASAP7_75t_L g20567 ( 
.A1(n_20561),
.A2(n_20558),
.B(n_20559),
.Y(n_20567)
);

INVx1_ASAP7_75t_L g20568 ( 
.A(n_20557),
.Y(n_20568)
);

INVx1_ASAP7_75t_L g20569 ( 
.A(n_20555),
.Y(n_20569)
);

AOI21xp5_ASAP7_75t_L g20570 ( 
.A1(n_20565),
.A2(n_5814),
.B(n_5784),
.Y(n_20570)
);

AOI222xp33_ASAP7_75t_SL g20571 ( 
.A1(n_20569),
.A2(n_7638),
.B1(n_5363),
.B2(n_5237),
.C1(n_5343),
.C2(n_5320),
.Y(n_20571)
);

OAI221xp5_ASAP7_75t_L g20572 ( 
.A1(n_20563),
.A2(n_5865),
.B1(n_5938),
.B2(n_5864),
.C(n_5827),
.Y(n_20572)
);

AOI21xp5_ASAP7_75t_L g20573 ( 
.A1(n_20566),
.A2(n_5864),
.B(n_5827),
.Y(n_20573)
);

NAND2xp5_ASAP7_75t_L g20574 ( 
.A(n_20568),
.B(n_5827),
.Y(n_20574)
);

XNOR2xp5_ASAP7_75t_L g20575 ( 
.A(n_20574),
.B(n_20564),
.Y(n_20575)
);

AOI22xp33_ASAP7_75t_L g20576 ( 
.A1(n_20570),
.A2(n_20567),
.B1(n_7050),
.B2(n_7065),
.Y(n_20576)
);

AOI21x1_ASAP7_75t_L g20577 ( 
.A1(n_20573),
.A2(n_7781),
.B(n_7777),
.Y(n_20577)
);

AOI22xp33_ASAP7_75t_L g20578 ( 
.A1(n_20572),
.A2(n_7050),
.B1(n_7065),
.B2(n_7018),
.Y(n_20578)
);

OR2x2_ASAP7_75t_L g20579 ( 
.A(n_20571),
.B(n_5827),
.Y(n_20579)
);

OAI21xp5_ASAP7_75t_L g20580 ( 
.A1(n_20575),
.A2(n_8370),
.B(n_8365),
.Y(n_20580)
);

OAI22xp5_ASAP7_75t_L g20581 ( 
.A1(n_20579),
.A2(n_5864),
.B1(n_5865),
.B2(n_5827),
.Y(n_20581)
);

AOI22xp5_ASAP7_75t_L g20582 ( 
.A1(n_20576),
.A2(n_20578),
.B1(n_20577),
.B2(n_5865),
.Y(n_20582)
);

AOI21xp5_ASAP7_75t_L g20583 ( 
.A1(n_20575),
.A2(n_5865),
.B(n_5864),
.Y(n_20583)
);

CKINVDCx20_ASAP7_75t_R g20584 ( 
.A(n_20582),
.Y(n_20584)
);

INVx1_ASAP7_75t_L g20585 ( 
.A(n_20583),
.Y(n_20585)
);

INVxp67_ASAP7_75t_L g20586 ( 
.A(n_20585),
.Y(n_20586)
);

NAND2xp5_ASAP7_75t_L g20587 ( 
.A(n_20584),
.B(n_20581),
.Y(n_20587)
);

OA21x2_ASAP7_75t_L g20588 ( 
.A1(n_20585),
.A2(n_20580),
.B(n_8510),
.Y(n_20588)
);

OAI221xp5_ASAP7_75t_R g20589 ( 
.A1(n_20586),
.A2(n_7600),
.B1(n_7248),
.B2(n_7245),
.C(n_8131),
.Y(n_20589)
);

AOI22xp33_ASAP7_75t_L g20590 ( 
.A1(n_20589),
.A2(n_20587),
.B1(n_20588),
.B2(n_5865),
.Y(n_20590)
);

AOI211xp5_ASAP7_75t_L g20591 ( 
.A1(n_20590),
.A2(n_5865),
.B(n_5938),
.C(n_5864),
.Y(n_20591)
);


endmodule