module real_aes_2205_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_0), .B(n_501), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_1), .A2(n_503), .B(n_504), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_2), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_3), .B(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_4), .B(n_268), .Y(n_536) );
INVx1_ASAP7_75t_L g154 ( .A(n_5), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_6), .B(n_173), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_7), .B(n_268), .Y(n_563) );
INVx1_ASAP7_75t_L g237 ( .A(n_8), .Y(n_237) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_9), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_10), .Y(n_202) );
NAND2xp33_ASAP7_75t_L g525 ( .A(n_11), .B(n_265), .Y(n_525) );
INVx2_ASAP7_75t_L g143 ( .A(n_12), .Y(n_143) );
AOI221x1_ASAP7_75t_L g569 ( .A1(n_13), .A2(n_25), .B1(n_501), .B2(n_503), .C(n_570), .Y(n_569) );
NOR3xp33_ASAP7_75t_L g107 ( .A(n_14), .B(n_108), .C(n_110), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g122 ( .A(n_14), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_15), .B(n_501), .Y(n_521) );
INVx1_ASAP7_75t_L g266 ( .A(n_16), .Y(n_266) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_17), .A2(n_218), .B(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_18), .B(n_177), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_19), .B(n_268), .Y(n_513) );
AO21x1_ASAP7_75t_L g531 ( .A1(n_20), .A2(n_501), .B(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g105 ( .A(n_21), .Y(n_105) );
INVx1_ASAP7_75t_L g263 ( .A(n_22), .Y(n_263) );
INVx1_ASAP7_75t_SL g183 ( .A(n_23), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_24), .B(n_160), .Y(n_253) );
CKINVDCx20_ASAP7_75t_R g788 ( .A(n_26), .Y(n_788) );
AOI33xp33_ASAP7_75t_L g223 ( .A1(n_27), .A2(n_54), .A3(n_149), .B1(n_158), .B2(n_224), .B3(n_225), .Y(n_223) );
NAND2x1_ASAP7_75t_L g544 ( .A(n_28), .B(n_268), .Y(n_544) );
NAND2x1_ASAP7_75t_L g562 ( .A(n_29), .B(n_265), .Y(n_562) );
INVx1_ASAP7_75t_L g194 ( .A(n_30), .Y(n_194) );
OA21x2_ASAP7_75t_L g142 ( .A1(n_31), .A2(n_86), .B(n_143), .Y(n_142) );
OR2x2_ASAP7_75t_L g174 ( .A(n_31), .B(n_86), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_32), .B(n_168), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_33), .B(n_265), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_34), .B(n_268), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_35), .B(n_265), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_36), .A2(n_503), .B(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g148 ( .A(n_37), .Y(n_148) );
AND2x2_ASAP7_75t_L g166 ( .A(n_37), .B(n_154), .Y(n_166) );
AND2x2_ASAP7_75t_L g172 ( .A(n_37), .B(n_151), .Y(n_172) );
INVxp67_ASAP7_75t_L g110 ( .A(n_38), .Y(n_110) );
OR2x6_ASAP7_75t_L g124 ( .A(n_38), .B(n_104), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_39), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_40), .B(n_501), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_41), .B(n_168), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g246 ( .A1(n_42), .A2(n_141), .B1(n_173), .B2(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_43), .B(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_44), .B(n_160), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_45), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_46), .B(n_265), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_47), .Y(n_804) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_48), .B(n_218), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_49), .B(n_160), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_50), .A2(n_503), .B(n_561), .Y(n_560) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_51), .Y(n_250) );
OAI222xp33_ASAP7_75t_L g126 ( .A1(n_52), .A2(n_127), .B1(n_784), .B2(n_785), .C1(n_788), .C2(n_789), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_52), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_53), .B(n_265), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_55), .B(n_160), .Y(n_213) );
INVx1_ASAP7_75t_L g153 ( .A(n_56), .Y(n_153) );
INVx1_ASAP7_75t_L g162 ( .A(n_56), .Y(n_162) );
AND2x2_ASAP7_75t_L g214 ( .A(n_57), .B(n_177), .Y(n_214) );
AOI221xp5_ASAP7_75t_L g235 ( .A1(n_58), .A2(n_74), .B1(n_146), .B2(n_168), .C(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_59), .B(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_60), .B(n_268), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_61), .B(n_141), .Y(n_204) );
AOI21xp5_ASAP7_75t_SL g145 ( .A1(n_62), .A2(n_146), .B(n_155), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_63), .A2(n_503), .B(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g260 ( .A(n_64), .Y(n_260) );
AO21x1_ASAP7_75t_L g533 ( .A1(n_65), .A2(n_503), .B(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_66), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g212 ( .A(n_67), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_68), .B(n_501), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_69), .A2(n_146), .B(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g555 ( .A(n_70), .B(n_178), .Y(n_555) );
INVx1_ASAP7_75t_L g151 ( .A(n_71), .Y(n_151) );
INVx1_ASAP7_75t_L g164 ( .A(n_71), .Y(n_164) );
AND2x2_ASAP7_75t_L g565 ( .A(n_72), .B(n_140), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_73), .B(n_168), .Y(n_226) );
AND2x2_ASAP7_75t_L g185 ( .A(n_75), .B(n_140), .Y(n_185) );
INVx1_ASAP7_75t_L g261 ( .A(n_76), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_77), .A2(n_146), .B(n_182), .Y(n_181) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_78), .A2(n_146), .B(n_217), .C(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g106 ( .A(n_79), .Y(n_106) );
AND2x2_ASAP7_75t_L g498 ( .A(n_80), .B(n_140), .Y(n_498) );
AND2x2_ASAP7_75t_SL g139 ( .A(n_81), .B(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_82), .B(n_501), .Y(n_515) );
OAI22xp5_ASAP7_75t_SL g799 ( .A1(n_83), .A2(n_489), .B1(n_800), .B2(n_801), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_83), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g220 ( .A1(n_84), .A2(n_146), .B1(n_221), .B2(n_222), .Y(n_220) );
AND2x2_ASAP7_75t_L g532 ( .A(n_85), .B(n_173), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_87), .B(n_265), .Y(n_514) );
AND2x2_ASAP7_75t_L g547 ( .A(n_88), .B(n_140), .Y(n_547) );
INVx1_ASAP7_75t_L g156 ( .A(n_89), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_90), .B(n_268), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_91), .A2(n_503), .B(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_92), .B(n_265), .Y(n_571) );
AND2x2_ASAP7_75t_L g227 ( .A(n_93), .B(n_140), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_94), .B(n_268), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_95), .A2(n_192), .B(n_193), .C(n_196), .Y(n_191) );
INVx1_ASAP7_75t_SL g114 ( .A(n_96), .Y(n_114) );
BUFx2_ASAP7_75t_SL g797 ( .A(n_96), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_97), .A2(n_503), .B(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_98), .B(n_160), .Y(n_159) );
AOI21xp33_ASAP7_75t_SL g99 ( .A1(n_100), .A2(n_111), .B(n_803), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_SL g805 ( .A(n_101), .Y(n_805) );
INVx2_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_SL g102 ( .A(n_103), .B(n_107), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
OA21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_126), .B(n_793), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_115), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
INVxp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g798 ( .A1(n_116), .A2(n_799), .B(n_802), .Y(n_798) );
NOR2xp33_ASAP7_75t_SL g116 ( .A(n_117), .B(n_125), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_120), .Y(n_802) );
BUFx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
OR2x6_ASAP7_75t_SL g488 ( .A(n_122), .B(n_123), .Y(n_488) );
AND2x6_ASAP7_75t_SL g783 ( .A(n_122), .B(n_124), .Y(n_783) );
OR2x2_ASAP7_75t_L g787 ( .A(n_122), .B(n_124), .Y(n_787) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
OAI22x1_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_486), .B1(n_489), .B2(n_782), .Y(n_128) );
AOI22x1_ASAP7_75t_L g789 ( .A1(n_129), .A2(n_487), .B1(n_790), .B2(n_792), .Y(n_789) );
INVx1_ASAP7_75t_SL g129 ( .A(n_130), .Y(n_129) );
AND3x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_376), .C(n_439), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_340), .Y(n_132) );
NOR3xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_281), .C(n_310), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g134 ( .A(n_135), .B(n_270), .Y(n_134) );
AOI22xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_186), .B1(n_228), .B2(n_240), .Y(n_135) );
NAND2x1_ASAP7_75t_L g425 ( .A(n_136), .B(n_271), .Y(n_425) );
INVx2_ASAP7_75t_SL g136 ( .A(n_137), .Y(n_136) );
OR2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_175), .Y(n_137) );
INVx2_ASAP7_75t_L g242 ( .A(n_138), .Y(n_242) );
INVx4_ASAP7_75t_L g286 ( .A(n_138), .Y(n_286) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_138), .Y(n_306) );
AND2x4_ASAP7_75t_L g317 ( .A(n_138), .B(n_285), .Y(n_317) );
AND2x2_ASAP7_75t_L g323 ( .A(n_138), .B(n_245), .Y(n_323) );
NOR2x1_ASAP7_75t_SL g453 ( .A(n_138), .B(n_256), .Y(n_453) );
OR2x6_ASAP7_75t_L g138 ( .A(n_139), .B(n_144), .Y(n_138) );
OAI22xp5_ASAP7_75t_L g190 ( .A1(n_140), .A2(n_191), .B1(n_197), .B2(n_198), .Y(n_190) );
INVx3_ASAP7_75t_L g198 ( .A(n_140), .Y(n_198) );
INVx4_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_141), .B(n_201), .Y(n_200) );
INVx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx4f_ASAP7_75t_L g218 ( .A(n_142), .Y(n_218) );
AND2x4_ASAP7_75t_L g173 ( .A(n_143), .B(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_SL g178 ( .A(n_143), .B(n_174), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_167), .B(n_173), .Y(n_144) );
INVxp67_ASAP7_75t_L g203 ( .A(n_146), .Y(n_203) );
AND2x4_ASAP7_75t_L g146 ( .A(n_147), .B(n_152), .Y(n_146) );
NOR2x1p5_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
INVx1_ASAP7_75t_L g225 ( .A(n_149), .Y(n_225) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
OR2x6_ASAP7_75t_L g157 ( .A(n_150), .B(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x6_ASAP7_75t_L g265 ( .A(n_151), .B(n_161), .Y(n_265) );
AND2x6_ASAP7_75t_L g503 ( .A(n_152), .B(n_172), .Y(n_503) );
AND2x2_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
INVx2_ASAP7_75t_L g158 ( .A(n_153), .Y(n_158) );
AND2x4_ASAP7_75t_L g268 ( .A(n_153), .B(n_163), .Y(n_268) );
HB1xp67_ASAP7_75t_L g170 ( .A(n_154), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_159), .C(n_165), .Y(n_155) );
O2A1O1Ixp33_ASAP7_75t_SL g182 ( .A1(n_157), .A2(n_165), .B(n_183), .C(n_184), .Y(n_182) );
INVxp67_ASAP7_75t_L g192 ( .A(n_157), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g211 ( .A1(n_157), .A2(n_165), .B(n_212), .C(n_213), .Y(n_211) );
O2A1O1Ixp33_ASAP7_75t_SL g236 ( .A1(n_157), .A2(n_165), .B(n_237), .C(n_238), .Y(n_236) );
INVx2_ASAP7_75t_L g255 ( .A(n_157), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g259 ( .A1(n_157), .A2(n_195), .B1(n_260), .B2(n_261), .Y(n_259) );
AND2x2_ASAP7_75t_L g169 ( .A(n_158), .B(n_170), .Y(n_169) );
INVxp33_ASAP7_75t_L g224 ( .A(n_158), .Y(n_224) );
INVx1_ASAP7_75t_L g195 ( .A(n_160), .Y(n_195) );
AND2x4_ASAP7_75t_L g501 ( .A(n_160), .B(n_166), .Y(n_501) );
AND2x4_ASAP7_75t_L g160 ( .A(n_161), .B(n_163), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g221 ( .A(n_165), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_165), .A2(n_253), .B(n_254), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_165), .B(n_173), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_165), .A2(n_505), .B(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_165), .A2(n_513), .B(n_514), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_165), .A2(n_524), .B(n_525), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_165), .A2(n_535), .B(n_536), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_165), .A2(n_544), .B(n_545), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_165), .A2(n_552), .B(n_553), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_165), .A2(n_562), .B(n_563), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_165), .A2(n_571), .B(n_572), .Y(n_570) );
INVx5_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_166), .Y(n_196) );
INVx1_ASAP7_75t_L g205 ( .A(n_168), .Y(n_205) );
AND2x4_ASAP7_75t_L g168 ( .A(n_169), .B(n_171), .Y(n_168) );
INVx1_ASAP7_75t_L g248 ( .A(n_169), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_171), .Y(n_249) );
BUFx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_SL g509 ( .A(n_173), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_173), .A2(n_521), .B(n_522), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_173), .B(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g289 ( .A(n_175), .Y(n_289) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_175), .Y(n_303) );
INVx1_ASAP7_75t_L g314 ( .A(n_175), .Y(n_314) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_175), .Y(n_326) );
AND2x2_ASAP7_75t_L g358 ( .A(n_175), .B(n_256), .Y(n_358) );
AND2x2_ASAP7_75t_L g390 ( .A(n_175), .B(n_274), .Y(n_390) );
INVx1_ASAP7_75t_L g397 ( .A(n_175), .Y(n_397) );
AO21x2_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_179), .B(n_185), .Y(n_175) );
AO21x2_ASAP7_75t_L g558 ( .A1(n_176), .A2(n_559), .B(n_565), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_177), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_177), .A2(n_500), .B(n_502), .Y(n_499) );
OA21x2_ASAP7_75t_L g568 ( .A1(n_177), .A2(n_569), .B(n_573), .Y(n_568) );
OA21x2_ASAP7_75t_L g608 ( .A1(n_177), .A2(n_569), .B(n_573), .Y(n_608) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
AND2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_206), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g339 ( .A(n_188), .B(n_278), .Y(n_339) );
INVx2_ASAP7_75t_L g413 ( .A(n_188), .Y(n_413) );
AND2x2_ASAP7_75t_L g436 ( .A(n_188), .B(n_206), .Y(n_436) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_189), .B(n_231), .Y(n_277) );
INVx2_ASAP7_75t_L g298 ( .A(n_189), .Y(n_298) );
AND2x4_ASAP7_75t_L g320 ( .A(n_189), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g355 ( .A(n_189), .Y(n_355) );
AND2x2_ASAP7_75t_L g432 ( .A(n_189), .B(n_234), .Y(n_432) );
OR2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_199), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
AO21x2_ASAP7_75t_L g207 ( .A1(n_198), .A2(n_208), .B(n_214), .Y(n_207) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_198), .A2(n_208), .B(n_214), .Y(n_231) );
AO21x2_ASAP7_75t_L g540 ( .A1(n_198), .A2(n_541), .B(n_547), .Y(n_540) );
AO21x2_ASAP7_75t_L g548 ( .A1(n_198), .A2(n_549), .B(n_555), .Y(n_548) );
AO21x2_ASAP7_75t_L g576 ( .A1(n_198), .A2(n_541), .B(n_547), .Y(n_576) );
AO21x2_ASAP7_75t_L g594 ( .A1(n_198), .A2(n_549), .B(n_555), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_203), .B1(n_204), .B2(n_205), .Y(n_199) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g403 ( .A(n_206), .Y(n_403) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_215), .Y(n_206) );
NOR2xp67_ASAP7_75t_L g328 ( .A(n_207), .B(n_298), .Y(n_328) );
AND2x2_ASAP7_75t_L g333 ( .A(n_207), .B(n_298), .Y(n_333) );
INVx2_ASAP7_75t_L g346 ( .A(n_207), .Y(n_346) );
NOR2x1_ASAP7_75t_L g394 ( .A(n_207), .B(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
AND2x4_ASAP7_75t_L g319 ( .A(n_215), .B(n_230), .Y(n_319) );
AND2x2_ASAP7_75t_L g334 ( .A(n_215), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g387 ( .A(n_215), .Y(n_387) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_216), .B(n_234), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_216), .B(n_231), .Y(n_391) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_219), .B(n_227), .Y(n_216) );
AO21x2_ASAP7_75t_L g280 ( .A1(n_217), .A2(n_219), .B(n_227), .Y(n_280) );
INVx2_ASAP7_75t_SL g217 ( .A(n_218), .Y(n_217) );
OA21x2_ASAP7_75t_L g234 ( .A1(n_218), .A2(n_235), .B(n_239), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_220), .B(n_226), .Y(n_219) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVxp33_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NAND2x1p5_ASAP7_75t_L g229 ( .A(n_230), .B(n_232), .Y(n_229) );
INVx3_ASAP7_75t_L g295 ( .A(n_230), .Y(n_295) );
INVx3_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_231), .Y(n_293) );
AND2x2_ASAP7_75t_L g462 ( .A(n_231), .B(n_463), .Y(n_462) );
INVx3_ASAP7_75t_L g350 ( .A(n_232), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_232), .B(n_387), .Y(n_482) );
BUFx3_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g297 ( .A(n_233), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x4_ASAP7_75t_L g278 ( .A(n_234), .B(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g321 ( .A(n_234), .Y(n_321) );
INVxp67_ASAP7_75t_L g335 ( .A(n_234), .Y(n_335) );
INVx1_ASAP7_75t_L g395 ( .A(n_234), .Y(n_395) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_234), .Y(n_463) );
INVx1_ASAP7_75t_L g447 ( .A(n_240), .Y(n_447) );
NOR2x1_ASAP7_75t_L g240 ( .A(n_241), .B(n_243), .Y(n_240) );
NOR2x1_ASAP7_75t_L g367 ( .A(n_241), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g401 ( .A(n_242), .B(n_273), .Y(n_401) );
OR2x2_ASAP7_75t_L g437 ( .A(n_243), .B(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g419 ( .A(n_244), .B(n_397), .Y(n_419) );
AND2x2_ASAP7_75t_L g471 ( .A(n_244), .B(n_306), .Y(n_471) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_256), .Y(n_244) );
AND2x4_ASAP7_75t_L g273 ( .A(n_245), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g285 ( .A(n_245), .Y(n_285) );
INVx2_ASAP7_75t_L g302 ( .A(n_245), .Y(n_302) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_245), .Y(n_480) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_251), .Y(n_245) );
NOR3xp33_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .C(n_250), .Y(n_247) );
INVx3_ASAP7_75t_L g274 ( .A(n_256), .Y(n_274) );
INVx2_ASAP7_75t_L g368 ( .A(n_256), .Y(n_368) );
AND2x4_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
OAI21xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_262), .B(n_269), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_264), .B1(n_266), .B2(n_267), .Y(n_262) );
INVxp67_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVxp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_275), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_272), .B(n_348), .Y(n_365) );
NOR2x1_ASAP7_75t_L g407 ( .A(n_272), .B(n_286), .Y(n_407) );
INVx4_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_273), .B(n_348), .Y(n_485) );
AND2x2_ASAP7_75t_L g301 ( .A(n_274), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g315 ( .A(n_274), .Y(n_315) );
AOI22xp5_ASAP7_75t_SL g363 ( .A1(n_275), .A2(n_364), .B1(n_365), .B2(n_366), .Y(n_363) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
NAND2x1p5_ASAP7_75t_L g360 ( .A(n_276), .B(n_334), .Y(n_360) );
INVx2_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g421 ( .A(n_277), .B(n_309), .Y(n_421) );
AND2x2_ASAP7_75t_L g291 ( .A(n_278), .B(n_292), .Y(n_291) );
AND2x4_ASAP7_75t_L g327 ( .A(n_278), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g423 ( .A(n_278), .B(n_413), .Y(n_423) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x4_ASAP7_75t_L g345 ( .A(n_280), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g371 ( .A(n_280), .Y(n_371) );
AND2x2_ASAP7_75t_L g461 ( .A(n_280), .B(n_298), .Y(n_461) );
OAI221xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_290), .B1(n_294), .B2(n_299), .C(n_304), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_287), .Y(n_283) );
INVx1_ASAP7_75t_L g362 ( .A(n_284), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_284), .B(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_284), .B(n_358), .Y(n_477) );
AND2x4_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
NOR2xp67_ASAP7_75t_SL g330 ( .A(n_286), .B(n_331), .Y(n_330) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_286), .Y(n_343) );
OR2x2_ASAP7_75t_L g427 ( .A(n_286), .B(n_428), .Y(n_427) );
AND2x4_ASAP7_75t_SL g479 ( .A(n_286), .B(n_480), .Y(n_479) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx3_ASAP7_75t_L g348 ( .A(n_288), .Y(n_348) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_289), .Y(n_438) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AOI221x1_ASAP7_75t_L g378 ( .A1(n_291), .A2(n_379), .B1(n_381), .B2(n_384), .C(n_388), .Y(n_378) );
AND2x2_ASAP7_75t_L g364 ( .A(n_292), .B(n_320), .Y(n_364) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
AND2x2_ASAP7_75t_L g307 ( .A(n_295), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_295), .B(n_297), .Y(n_434) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
AND2x2_ASAP7_75t_SL g305 ( .A(n_301), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_301), .B(n_314), .Y(n_331) );
INVx2_ASAP7_75t_L g338 ( .A(n_301), .Y(n_338) );
INVx1_ASAP7_75t_L g383 ( .A(n_302), .Y(n_383) );
BUFx2_ASAP7_75t_L g472 ( .A(n_303), .Y(n_472) );
NAND2xp33_ASAP7_75t_SL g304 ( .A(n_305), .B(n_307), .Y(n_304) );
OR2x6_ASAP7_75t_L g337 ( .A(n_306), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g418 ( .A(n_306), .B(n_358), .Y(n_418) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_329), .Y(n_310) );
AOI22xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_318), .B1(n_322), .B2(n_327), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_313), .B(n_316), .Y(n_312) );
AND2x2_ASAP7_75t_SL g375 ( .A(n_313), .B(n_317), .Y(n_375) );
AND2x4_ASAP7_75t_L g381 ( .A(n_313), .B(n_382), .Y(n_381) );
AND2x4_ASAP7_75t_SL g313 ( .A(n_314), .B(n_315), .Y(n_313) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_314), .Y(n_406) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_317), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_317), .B(n_348), .Y(n_380) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_317), .Y(n_464) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AND2x2_ASAP7_75t_L g411 ( .A(n_319), .B(n_412), .Y(n_411) );
INVx3_ASAP7_75t_L g372 ( .A(n_320), .Y(n_372) );
NAND2x1_ASAP7_75t_SL g416 ( .A(n_320), .B(n_371), .Y(n_416) );
AND2x2_ASAP7_75t_L g450 ( .A(n_320), .B(n_345), .Y(n_450) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_332), .B1(n_336), .B2(n_339), .Y(n_329) );
BUFx2_ASAP7_75t_L g445 ( .A(n_331), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_332), .A2(n_401), .B1(n_475), .B2(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
NAND2x1p5_ASAP7_75t_L g386 ( .A(n_333), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g353 ( .A(n_334), .B(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND3xp33_ASAP7_75t_L g469 ( .A(n_338), .B(n_470), .C(n_472), .Y(n_469) );
INVx1_ASAP7_75t_L g373 ( .A(n_339), .Y(n_373) );
AOI211x1_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_349), .B(n_351), .C(n_369), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_344), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_347), .Y(n_344) );
AND2x2_ASAP7_75t_L g431 ( .A(n_345), .B(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_345), .B(n_412), .Y(n_443) );
AND2x2_ASAP7_75t_L g475 ( .A(n_345), .B(n_413), .Y(n_475) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g456 ( .A(n_348), .Y(n_456) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g385 ( .A(n_350), .B(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_352), .B(n_363), .Y(n_351) );
AOI22xp5_ASAP7_75t_SL g352 ( .A1(n_353), .A2(n_356), .B1(n_359), .B2(n_361), .Y(n_352) );
BUFx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g393 ( .A(n_355), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g408 ( .A(n_355), .Y(n_408) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_SL g478 ( .A(n_358), .B(n_479), .Y(n_478) );
INVx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVxp67_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g414 ( .A(n_367), .B(n_397), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_373), .B(n_374), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_371), .B(n_393), .Y(n_468) );
OR2x2_ASAP7_75t_L g446 ( .A(n_372), .B(n_391), .Y(n_446) );
INVx1_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND3x1_ASAP7_75t_L g377 ( .A(n_378), .B(n_398), .C(n_422), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_381), .A2(n_411), .B1(n_414), .B2(n_415), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_382), .B(n_397), .Y(n_396) );
INVx2_ASAP7_75t_SL g455 ( .A(n_382), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_382), .B(n_456), .Y(n_459) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OAI222xp33_ASAP7_75t_L g442 ( .A1(n_386), .A2(n_443), .B1(n_444), .B2(n_445), .C1(n_446), .C2(n_447), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_391), .B1(n_392), .B2(n_396), .Y(n_388) );
INVx1_ASAP7_75t_SL g428 ( .A(n_390), .Y(n_428) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g465 ( .A(n_394), .B(n_461), .Y(n_465) );
NOR2x1_ASAP7_75t_L g398 ( .A(n_399), .B(n_409), .Y(n_398) );
AOI21xp5_ASAP7_75t_SL g399 ( .A1(n_400), .A2(n_402), .B(n_408), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_417), .Y(n_409) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_416), .B(n_430), .Y(n_429) );
OAI21xp5_ASAP7_75t_SL g417 ( .A1(n_418), .A2(n_419), .B(n_420), .Y(n_417) );
INVx1_ASAP7_75t_L g444 ( .A(n_419), .Y(n_444) );
INVx1_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_424), .B1(n_426), .B2(n_429), .C(n_433), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVxp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B(n_437), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVxp67_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
NAND3x1_ASAP7_75t_L g440 ( .A(n_441), .B(n_466), .C(n_473), .Y(n_440) );
NOR2x1_ASAP7_75t_L g441 ( .A(n_442), .B(n_448), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_457), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_450), .B(n_451), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_454), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_452), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_460), .B1(n_464), .B2(n_465), .Y(n_457) );
AND2x4_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_467), .B(n_469), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_483), .Y(n_473) );
AOI22xp5_ASAP7_75t_SL g474 ( .A1(n_475), .A2(n_476), .B1(n_478), .B2(n_481), .Y(n_474) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVxp67_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
CKINVDCx11_ASAP7_75t_R g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g801 ( .A(n_489), .Y(n_801) );
INVx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g792 ( .A(n_490), .Y(n_792) );
AND2x4_ASAP7_75t_L g490 ( .A(n_491), .B(n_691), .Y(n_490) );
NOR4xp25_ASAP7_75t_L g491 ( .A(n_492), .B(n_609), .C(n_635), .D(n_675), .Y(n_491) );
OAI211xp5_ASAP7_75t_SL g492 ( .A1(n_493), .A2(n_526), .B(n_556), .C(n_595), .Y(n_492) );
INVxp67_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_507), .Y(n_494) );
AND2x2_ASAP7_75t_L g762 ( .A(n_495), .B(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_496), .B(n_507), .Y(n_629) );
BUFx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g557 ( .A(n_497), .B(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_497), .B(n_582), .Y(n_581) );
INVx5_ASAP7_75t_L g615 ( .A(n_497), .Y(n_615) );
NOR2x1_ASAP7_75t_SL g657 ( .A(n_497), .B(n_508), .Y(n_657) );
AND2x2_ASAP7_75t_L g713 ( .A(n_497), .B(n_519), .Y(n_713) );
OR2x6_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_518), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_508), .B(n_519), .Y(n_585) );
AND2x2_ASAP7_75t_L g646 ( .A(n_508), .B(n_615), .Y(n_646) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .B(n_516), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_509), .B(n_517), .Y(n_516) );
AO21x2_ASAP7_75t_L g599 ( .A1(n_509), .A2(n_510), .B(n_516), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_515), .Y(n_510) );
AND2x2_ASAP7_75t_L g658 ( .A(n_518), .B(n_582), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_518), .B(n_663), .Y(n_662) );
OR2x2_ASAP7_75t_L g702 ( .A(n_518), .B(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g735 ( .A(n_518), .B(n_557), .Y(n_735) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g579 ( .A(n_519), .Y(n_579) );
AND2x2_ASAP7_75t_L g612 ( .A(n_519), .B(n_613), .Y(n_612) );
BUFx3_ASAP7_75t_L g647 ( .A(n_519), .Y(n_647) );
OR2x2_ASAP7_75t_L g723 ( .A(n_519), .B(n_582), .Y(n_723) );
INVx1_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_539), .Y(n_527) );
AOI211x1_ASAP7_75t_SL g652 ( .A1(n_528), .A2(n_644), .B(n_653), .C(n_655), .Y(n_652) );
AND2x2_ASAP7_75t_SL g697 ( .A(n_528), .B(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_528), .B(n_695), .Y(n_742) );
BUFx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g592 ( .A(n_529), .Y(n_592) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g567 ( .A(n_530), .Y(n_567) );
OAI21x1_ASAP7_75t_SL g530 ( .A1(n_531), .A2(n_533), .B(n_537), .Y(n_530) );
INVx1_ASAP7_75t_L g538 ( .A(n_532), .Y(n_538) );
AOI322xp5_ASAP7_75t_L g556 ( .A1(n_539), .A2(n_557), .A3(n_566), .B1(n_574), .B2(n_577), .C1(n_583), .C2(n_586), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_539), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_548), .Y(n_539) );
INVx2_ASAP7_75t_L g590 ( .A(n_540), .Y(n_590) );
INVxp67_ASAP7_75t_L g632 ( .A(n_540), .Y(n_632) );
BUFx3_ASAP7_75t_L g696 ( .A(n_540), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_546), .Y(n_541) );
INVx2_ASAP7_75t_L g605 ( .A(n_548), .Y(n_605) );
AND2x2_ASAP7_75t_L g654 ( .A(n_548), .B(n_568), .Y(n_654) );
AND2x2_ASAP7_75t_L g698 ( .A(n_548), .B(n_607), .Y(n_698) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_550), .B(n_554), .Y(n_549) );
AND2x2_ASAP7_75t_L g583 ( .A(n_557), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_557), .B(n_768), .Y(n_767) );
AND2x2_ASAP7_75t_SL g777 ( .A(n_557), .B(n_612), .Y(n_777) );
INVx4_ASAP7_75t_L g582 ( .A(n_558), .Y(n_582) );
AND2x2_ASAP7_75t_L g614 ( .A(n_558), .B(n_615), .Y(n_614) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_558), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_564), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g676 ( .A(n_566), .B(n_651), .Y(n_676) );
INVx1_ASAP7_75t_SL g715 ( .A(n_566), .Y(n_715) );
AND2x4_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
AND2x4_ASAP7_75t_L g606 ( .A(n_567), .B(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_567), .B(n_605), .Y(n_674) );
AND2x2_ASAP7_75t_L g726 ( .A(n_567), .B(n_576), .Y(n_726) );
OR2x2_ASAP7_75t_L g750 ( .A(n_567), .B(n_568), .Y(n_750) );
AND2x2_ASAP7_75t_L g574 ( .A(n_568), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g624 ( .A(n_568), .B(n_605), .Y(n_624) );
AND2x2_ASAP7_75t_SL g680 ( .A(n_568), .B(n_592), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_574), .B(n_687), .Y(n_704) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
BUFx2_ASAP7_75t_L g639 ( .A(n_576), .Y(n_639) );
AND2x4_ASAP7_75t_SL g679 ( .A(n_576), .B(n_593), .Y(n_679) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .Y(n_577) );
OR2x2_ASAP7_75t_L g627 ( .A(n_578), .B(n_581), .Y(n_627) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g596 ( .A(n_579), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g744 ( .A(n_579), .B(n_657), .Y(n_744) );
AND2x2_ASAP7_75t_L g760 ( .A(n_579), .B(n_614), .Y(n_760) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AOI311xp33_ASAP7_75t_L g730 ( .A1(n_581), .A2(n_669), .A3(n_731), .B(n_733), .C(n_740), .Y(n_730) );
AND2x4_ASAP7_75t_L g597 ( .A(n_582), .B(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g601 ( .A(n_582), .Y(n_601) );
NAND2x1p5_ASAP7_75t_L g671 ( .A(n_582), .B(n_615), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_582), .B(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g714 ( .A(n_582), .B(n_701), .Y(n_714) );
AND2x2_ASAP7_75t_L g600 ( .A(n_584), .B(n_601), .Y(n_600) );
INVxp67_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
INVxp67_ASAP7_75t_SL g618 ( .A(n_585), .Y(n_618) );
OR2x2_ASAP7_75t_L g707 ( .A(n_585), .B(n_671), .Y(n_707) );
INVx1_ASAP7_75t_L g763 ( .A(n_585), .Y(n_763) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_591), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g672 ( .A(n_589), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g686 ( .A(n_589), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g761 ( .A(n_589), .B(n_634), .Y(n_761) );
BUFx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g604 ( .A(n_590), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g623 ( .A(n_590), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g685 ( .A(n_591), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_591), .A2(n_741), .B1(n_742), .B2(n_743), .Y(n_740) );
OR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
AND2x2_ASAP7_75t_L g634 ( .A(n_592), .B(n_605), .Y(n_634) );
AND2x4_ASAP7_75t_L g687 ( .A(n_592), .B(n_594), .Y(n_687) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
OAI21xp33_ASAP7_75t_SL g595 ( .A1(n_596), .A2(n_600), .B(n_602), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_596), .A2(n_682), .B1(n_686), .B2(n_688), .Y(n_681) );
AND2x2_ASAP7_75t_SL g641 ( .A(n_597), .B(n_615), .Y(n_641) );
INVx2_ASAP7_75t_L g703 ( .A(n_597), .Y(n_703) );
AND2x2_ASAP7_75t_L g717 ( .A(n_597), .B(n_713), .Y(n_717) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g613 ( .A(n_599), .Y(n_613) );
INVx1_ASAP7_75t_L g666 ( .A(n_599), .Y(n_666) );
INVx1_ASAP7_75t_L g617 ( .A(n_601), .Y(n_617) );
AND3x2_ASAP7_75t_L g645 ( .A(n_601), .B(n_646), .C(n_647), .Y(n_645) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
INVx1_ASAP7_75t_L g709 ( .A(n_604), .Y(n_709) );
AND2x2_ASAP7_75t_L g637 ( .A(n_606), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g708 ( .A(n_606), .B(n_709), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_606), .A2(n_720), .B1(n_724), .B2(n_727), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_606), .B(n_754), .Y(n_758) );
BUFx2_ASAP7_75t_L g649 ( .A(n_607), .Y(n_649) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g620 ( .A(n_608), .Y(n_620) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_608), .Y(n_739) );
OAI221xp5_ASAP7_75t_SL g609 ( .A1(n_610), .A2(n_619), .B1(n_621), .B2(n_622), .C(n_625), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_616), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
INVx1_ASAP7_75t_L g701 ( .A(n_613), .Y(n_701) );
INVx2_ASAP7_75t_SL g690 ( .A(n_614), .Y(n_690) );
AND2x2_ASAP7_75t_L g772 ( .A(n_614), .B(n_639), .Y(n_772) );
INVx4_ASAP7_75t_L g663 ( .A(n_615), .Y(n_663) );
INVx1_ASAP7_75t_L g621 ( .A(n_616), .Y(n_621) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
AND2x4_ASAP7_75t_L g732 ( .A(n_620), .B(n_687), .Y(n_732) );
INVx1_ASAP7_75t_SL g771 ( .A(n_620), .Y(n_771) );
AND2x2_ASAP7_75t_L g776 ( .A(n_620), .B(n_679), .Y(n_776) );
INVx1_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g718 ( .A(n_624), .Y(n_718) );
OAI21xp5_ASAP7_75t_SL g625 ( .A1(n_626), .A2(n_628), .B(n_630), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx1_ASAP7_75t_L g651 ( .A(n_632), .Y(n_651) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g648 ( .A(n_634), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g738 ( .A(n_634), .B(n_739), .Y(n_738) );
OAI211xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_640), .B(n_642), .C(n_659), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g731 ( .A(n_638), .B(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_639), .B(n_654), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_639), .B(n_749), .Y(n_748) );
AND2x2_ASAP7_75t_L g764 ( .A(n_639), .B(n_687), .Y(n_764) );
OAI221xp5_ASAP7_75t_SL g675 ( .A1(n_640), .A2(n_664), .B1(n_676), .B2(n_677), .C(n_681), .Y(n_675) );
INVx3_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g746 ( .A(n_641), .B(n_647), .Y(n_746) );
OAI32xp33_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_648), .A3(n_650), .B1(n_652), .B2(n_656), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVxp67_ASAP7_75t_SL g736 ( .A(n_646), .Y(n_736) );
INVx2_ASAP7_75t_L g669 ( .A(n_647), .Y(n_669) );
O2A1O1Ixp33_ASAP7_75t_L g778 ( .A1(n_647), .A2(n_699), .B(n_779), .C(n_780), .Y(n_778) );
INVx1_ASAP7_75t_L g684 ( .A(n_649), .Y(n_684) );
OR2x2_ASAP7_75t_L g780 ( .A(n_649), .B(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_653), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g741 ( .A(n_656), .Y(n_741) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
INVx1_ASAP7_75t_L g722 ( .A(n_657), .Y(n_722) );
OAI21xp33_ASAP7_75t_SL g659 ( .A1(n_660), .A2(n_668), .B(n_672), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OR2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .Y(n_661) );
OR2x2_ASAP7_75t_L g699 ( .A(n_662), .B(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_663), .B(n_666), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_667), .Y(n_664) );
AOI221xp5_ASAP7_75t_L g765 ( .A1(n_665), .A2(n_697), .B1(n_766), .B2(n_769), .C(n_773), .Y(n_765) );
INVx2_ASAP7_75t_L g768 ( .A(n_665), .Y(n_768) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
OR2x2_ASAP7_75t_L g689 ( .A(n_669), .B(n_690), .Y(n_689) );
AND2x4_ASAP7_75t_L g756 ( .A(n_669), .B(n_714), .Y(n_756) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVxp67_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
INVx1_ASAP7_75t_L g754 ( .A(n_679), .Y(n_754) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_687), .B(n_717), .Y(n_774) );
INVx2_ASAP7_75t_L g781 ( .A(n_687), .Y(n_781) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OAI221xp5_ASAP7_75t_L g751 ( .A1(n_689), .A2(n_752), .B1(n_755), .B2(n_757), .C(n_759), .Y(n_751) );
AND5x1_ASAP7_75t_L g691 ( .A(n_692), .B(n_730), .C(n_745), .D(n_765), .E(n_775), .Y(n_691) );
NOR2xp33_ASAP7_75t_SL g692 ( .A(n_693), .B(n_710), .Y(n_692) );
OAI221xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_699), .B1(n_702), .B2(n_704), .C(n_705), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_695), .B(n_697), .Y(n_694) );
INVx1_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_708), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OAI221xp5_ASAP7_75t_SL g710 ( .A1(n_711), .A2(n_715), .B1(n_716), .B2(n_718), .C(n_719), .Y(n_710) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
AND2x4_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_715), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
OR2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
OR2x2_ASAP7_75t_L g728 ( .A(n_723), .B(n_729), .Y(n_728) );
CKINVDCx16_ASAP7_75t_R g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
AOI21xp33_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_736), .B(n_737), .Y(n_733) );
INVx1_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AOI21xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_747), .B(n_751), .Y(n_745) );
INVx1_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVxp67_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVxp67_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
AOI22xp5_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_761), .B1(n_762), .B2(n_764), .Y(n_759) );
O2A1O1Ixp33_ASAP7_75t_L g775 ( .A1(n_761), .A2(n_776), .B(n_777), .C(n_778), .Y(n_775) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
INVx1_ASAP7_75t_L g779 ( .A(n_772), .Y(n_779) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
CKINVDCx11_ASAP7_75t_R g782 ( .A(n_783), .Y(n_782) );
CKINVDCx5p33_ASAP7_75t_R g791 ( .A(n_783), .Y(n_791) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx3_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx3_ASAP7_75t_SL g790 ( .A(n_791), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_794), .B(n_798), .Y(n_793) );
CKINVDCx5p33_ASAP7_75t_R g794 ( .A(n_795), .Y(n_794) );
CKINVDCx11_ASAP7_75t_R g795 ( .A(n_796), .Y(n_795) );
CKINVDCx8_ASAP7_75t_R g796 ( .A(n_797), .Y(n_796) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
endmodule