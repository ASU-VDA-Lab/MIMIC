module fake_jpeg_30695_n_133 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_133);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

BUFx10_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_25),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_4),
.B(n_30),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_59),
.B(n_53),
.Y(n_75)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_60),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_64),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_51),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_51),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_63),
.B(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_66),
.B(n_71),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_74),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_57),
.B(n_56),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_64),
.A2(n_43),
.B1(n_53),
.B2(n_54),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_72),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_76),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_58),
.B(n_55),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_44),
.Y(n_84)
);

NOR2x1_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_47),
.Y(n_78)
);

NOR2xp67_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_61),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_23),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_65),
.C(n_5),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_88),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_45),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_89),
.Y(n_94)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_46),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_0),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_2),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_92),
.A2(n_72),
.B(n_4),
.Y(n_97)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_13),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_106),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_110),
.B1(n_98),
.B2(n_95),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_26),
.C(n_27),
.Y(n_120)
);

A2O1A1O1Ixp25_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_22),
.B(n_38),
.C(n_37),
.D(n_9),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_107),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_3),
.B(n_5),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_105),
.B(n_21),
.Y(n_117)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_24),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_103),
.B(n_109),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_6),
.B(n_10),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_14),
.Y(n_107)
);

OAI32xp33_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_16),
.A3(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_108)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_83),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_20),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_118),
.Y(n_125)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_119),
.B(n_120),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_98),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_124),
.C(n_94),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_106),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_SL g126 ( 
.A1(n_125),
.A2(n_118),
.B(n_114),
.C(n_116),
.Y(n_126)
);

AOI21x1_ASAP7_75t_L g128 ( 
.A1(n_126),
.A2(n_127),
.B(n_122),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_112),
.B1(n_121),
.B2(n_31),
.Y(n_129)
);

MAJx2_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_28),
.C(n_29),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_130),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_36),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_132),
.B(n_41),
.Y(n_133)
);


endmodule