module fake_netlist_6_3077_n_1759 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1759);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1759;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_32),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_3),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_79),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_141),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_122),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_101),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_56),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_10),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_102),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

BUFx2_ASAP7_75t_SL g166 ( 
.A(n_53),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_139),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_23),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_57),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_107),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_67),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_7),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_26),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_129),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_138),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_144),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_92),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_135),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_84),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_119),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_111),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_36),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_31),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_58),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_120),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_42),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_8),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_36),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_91),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_4),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_3),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_94),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_128),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_42),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_95),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_54),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_41),
.Y(n_198)
);

BUFx10_ASAP7_75t_L g199 ( 
.A(n_105),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_68),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_41),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_99),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_48),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_6),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_9),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_18),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_27),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_106),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_145),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_69),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_45),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_35),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_131),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_24),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_52),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_38),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_112),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_150),
.Y(n_218)
);

INVxp33_ASAP7_75t_L g219 ( 
.A(n_132),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_146),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_28),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_89),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_77),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_40),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_108),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_39),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_50),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_5),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_59),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_86),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_9),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_4),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_83),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_62),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_30),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_88),
.Y(n_236)
);

INVxp33_ASAP7_75t_L g237 ( 
.A(n_44),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_74),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_34),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_64),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_47),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_65),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_104),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_126),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_18),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_96),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_90),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_87),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_117),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_39),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_25),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_140),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_20),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_14),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_149),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_49),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_124),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_76),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_10),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_27),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_97),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_148),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_130),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_100),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_93),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_82),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_66),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_29),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_8),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_143),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_142),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_30),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_152),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_20),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_110),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_13),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_98),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_116),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_7),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_78),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_15),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_72),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_85),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_23),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_121),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_61),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_34),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_55),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_11),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_17),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_37),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_81),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_109),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_21),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_80),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_28),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_22),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_12),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_13),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_125),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_47),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_6),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_17),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_294),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_294),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_294),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_183),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_294),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_294),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_172),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_270),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_193),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_189),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_164),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_194),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_172),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_196),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_198),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_161),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_198),
.Y(n_320)
);

INVxp33_ASAP7_75t_SL g321 ( 
.A(n_153),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_248),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_197),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_284),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_284),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_200),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_202),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_163),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_303),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_303),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_191),
.Y(n_331)
);

INVxp33_ASAP7_75t_L g332 ( 
.A(n_237),
.Y(n_332)
);

INVxp33_ASAP7_75t_SL g333 ( 
.A(n_153),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_174),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_248),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_203),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_207),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_226),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_228),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_208),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_213),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_231),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_251),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_296),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_265),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_265),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_253),
.Y(n_347)
);

INVxp33_ASAP7_75t_SL g348 ( 
.A(n_168),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_269),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_215),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_272),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_279),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_290),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_220),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_291),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_227),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_155),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_164),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_155),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_229),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_168),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_234),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_232),
.Y(n_363)
);

INVxp33_ASAP7_75t_SL g364 ( 
.A(n_173),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_219),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_238),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_240),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_232),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_165),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_165),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_173),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_233),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_164),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_247),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_154),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_233),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_236),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_375),
.B(n_210),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_304),
.B(n_236),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_322),
.B(n_156),
.Y(n_380)
);

OA21x2_ASAP7_75t_L g381 ( 
.A1(n_314),
.A2(n_170),
.B(n_159),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_304),
.B(n_305),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_305),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_306),
.B(n_178),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_314),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_314),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_358),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_319),
.A2(n_162),
.B1(n_260),
.B2(n_299),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_306),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_358),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_308),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_358),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_344),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_373),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_373),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_335),
.B(n_182),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_328),
.A2(n_274),
.B1(n_289),
.B2(n_298),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_346),
.B(n_167),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_345),
.B(n_186),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_373),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_312),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_308),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_332),
.A2(n_302),
.B1(n_301),
.B2(n_298),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_309),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_345),
.B(n_190),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_309),
.B(n_157),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_369),
.B(n_370),
.Y(n_407)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_315),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_317),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_369),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_345),
.B(n_217),
.Y(n_411)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_323),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_370),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_372),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_372),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_376),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_377),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_377),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_376),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_365),
.B(n_218),
.Y(n_420)
);

OA21x2_ASAP7_75t_L g421 ( 
.A1(n_310),
.A2(n_244),
.B(n_300),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_310),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_357),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_326),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_334),
.Y(n_425)
);

OAI21x1_ASAP7_75t_L g426 ( 
.A1(n_316),
.A2(n_223),
.B(n_222),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_316),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_357),
.B(n_157),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_341),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_318),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_331),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_361),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_318),
.B(n_225),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_359),
.B(n_158),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_331),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_338),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_338),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_339),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_320),
.B(n_243),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_327),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_320),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_339),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_336),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_342),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_342),
.Y(n_445)
);

CKINVDCx8_ASAP7_75t_R g446 ( 
.A(n_361),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_382),
.Y(n_447)
);

AO21x2_ASAP7_75t_L g448 ( 
.A1(n_426),
.A2(n_249),
.B(n_246),
.Y(n_448)
);

INVx8_ASAP7_75t_L g449 ( 
.A(n_378),
.Y(n_449)
);

INVx6_ASAP7_75t_L g450 ( 
.A(n_384),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_382),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_384),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_378),
.B(n_340),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_398),
.A2(n_311),
.B1(n_420),
.B2(n_401),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_423),
.Y(n_455)
);

INVx4_ASAP7_75t_SL g456 ( 
.A(n_386),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_382),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_382),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_393),
.Y(n_459)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_402),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_382),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_398),
.B(n_371),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_378),
.B(n_350),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_386),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_386),
.Y(n_465)
);

OAI22xp33_ASAP7_75t_L g466 ( 
.A1(n_446),
.A2(n_224),
.B1(n_192),
.B2(n_195),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_383),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_432),
.B(n_354),
.Y(n_468)
);

INVx4_ASAP7_75t_SL g469 ( 
.A(n_386),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_408),
.B(n_356),
.Y(n_470)
);

AND2x6_ASAP7_75t_L g471 ( 
.A(n_380),
.B(n_164),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_420),
.B(n_380),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_402),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_384),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_425),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_383),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_399),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_389),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_389),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_408),
.B(n_360),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_386),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_391),
.Y(n_482)
);

INVx5_ASAP7_75t_L g483 ( 
.A(n_386),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_386),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_408),
.B(n_362),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_390),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_391),
.Y(n_487)
);

INVx4_ASAP7_75t_L g488 ( 
.A(n_402),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_404),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_384),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_412),
.B(n_366),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_384),
.Y(n_492)
);

INVx5_ASAP7_75t_L g493 ( 
.A(n_390),
.Y(n_493)
);

NAND2xp33_ASAP7_75t_L g494 ( 
.A(n_420),
.B(n_164),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_412),
.B(n_367),
.Y(n_495)
);

AOI22xp33_ASAP7_75t_L g496 ( 
.A1(n_380),
.A2(n_333),
.B1(n_348),
.B2(n_364),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_404),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_396),
.B(n_374),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_422),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_429),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_390),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_412),
.B(n_321),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_379),
.Y(n_503)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_432),
.B(n_393),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_396),
.A2(n_166),
.B1(n_337),
.B2(n_307),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_440),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_422),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_379),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_379),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_412),
.B(n_313),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_399),
.B(n_405),
.Y(n_511)
);

OAI22xp33_ASAP7_75t_L g512 ( 
.A1(n_446),
.A2(n_211),
.B1(n_216),
.B2(n_214),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_396),
.B(n_177),
.Y(n_513)
);

INVx2_ASAP7_75t_SL g514 ( 
.A(n_399),
.Y(n_514)
);

INVx11_ASAP7_75t_L g515 ( 
.A(n_446),
.Y(n_515)
);

AO22x2_ASAP7_75t_L g516 ( 
.A1(n_403),
.A2(n_286),
.B1(n_252),
.B2(n_258),
.Y(n_516)
);

BUFx10_ASAP7_75t_L g517 ( 
.A(n_424),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_422),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_379),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_379),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_422),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_407),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_422),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_422),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_405),
.B(n_209),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_405),
.B(n_411),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_390),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_411),
.A2(n_353),
.B1(n_343),
.B2(n_349),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_443),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_407),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_422),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_407),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_409),
.B(n_199),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_411),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_403),
.B(n_199),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_390),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_427),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_433),
.B(n_343),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_406),
.B(n_277),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_402),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_406),
.B(n_256),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_427),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_407),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_402),
.Y(n_544)
);

BUFx10_ASAP7_75t_L g545 ( 
.A(n_433),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_407),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_427),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_431),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_427),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_431),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_427),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_435),
.Y(n_552)
);

NAND3xp33_ASAP7_75t_L g553 ( 
.A(n_428),
.B(n_201),
.C(n_204),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_388),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_433),
.B(n_257),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_427),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_433),
.B(n_439),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_427),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_441),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_435),
.Y(n_560)
);

INVx1_ASAP7_75t_SL g561 ( 
.A(n_388),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_428),
.B(n_199),
.Y(n_562)
);

AND2x6_ASAP7_75t_L g563 ( 
.A(n_433),
.B(n_261),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_441),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_441),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_423),
.B(n_324),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_434),
.B(n_368),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_423),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_434),
.B(n_359),
.Y(n_569)
);

CKINVDCx6p67_ASAP7_75t_R g570 ( 
.A(n_439),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_410),
.B(n_324),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_390),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_402),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_439),
.B(n_262),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_436),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_441),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_439),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_439),
.B(n_158),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_390),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_410),
.B(n_325),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_421),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_436),
.Y(n_582)
);

NOR2x1p5_ASAP7_75t_L g583 ( 
.A(n_437),
.B(n_184),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_441),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_421),
.A2(n_349),
.B1(n_347),
.B2(n_355),
.Y(n_585)
);

INVxp67_ASAP7_75t_L g586 ( 
.A(n_397),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_437),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_438),
.B(n_160),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_421),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_441),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_417),
.B(n_325),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_438),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_441),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_400),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_442),
.A2(n_255),
.B1(n_242),
.B2(n_230),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_522),
.Y(n_596)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_504),
.B(n_397),
.Y(n_597)
);

INVx8_ASAP7_75t_L g598 ( 
.A(n_449),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_530),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_472),
.B(n_263),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_530),
.Y(n_601)
);

NAND3xp33_ASAP7_75t_L g602 ( 
.A(n_462),
.B(n_239),
.C(n_205),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_451),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_462),
.B(n_442),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_583),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_529),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_532),
.B(n_543),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_498),
.B(n_160),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_477),
.B(n_421),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_487),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_543),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_477),
.B(n_421),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_546),
.B(n_271),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_568),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_487),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_568),
.B(n_444),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_514),
.B(n_414),
.Y(n_617)
);

INVx1_ASAP7_75t_SL g618 ( 
.A(n_504),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_459),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_514),
.B(n_414),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_516),
.A2(n_381),
.B1(n_426),
.B2(n_285),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_534),
.B(n_414),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_546),
.B(n_283),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_534),
.B(n_511),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_511),
.B(n_415),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_539),
.B(n_415),
.Y(n_626)
);

INVxp33_ASAP7_75t_L g627 ( 
.A(n_468),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_453),
.B(n_169),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_516),
.A2(n_381),
.B1(n_426),
.B2(n_295),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_548),
.Y(n_630)
);

O2A1O1Ixp33_ASAP7_75t_L g631 ( 
.A1(n_567),
.A2(n_445),
.B(n_444),
.C(n_418),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_526),
.B(n_415),
.Y(n_632)
);

O2A1O1Ixp5_ASAP7_75t_L g633 ( 
.A1(n_447),
.A2(n_392),
.B(n_385),
.C(n_387),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_452),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_516),
.A2(n_381),
.B1(n_445),
.B2(n_418),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_548),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_489),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_463),
.B(n_454),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_541),
.B(n_381),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_489),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_550),
.B(n_381),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_550),
.B(n_413),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_475),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_552),
.B(n_413),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_552),
.B(n_413),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_447),
.B(n_413),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_513),
.B(n_169),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_569),
.B(n_363),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_560),
.B(n_575),
.Y(n_649)
);

OAI221xp5_ASAP7_75t_L g650 ( 
.A1(n_505),
.A2(n_567),
.B1(n_585),
.B2(n_528),
.C(n_535),
.Y(n_650)
);

INVx4_ASAP7_75t_L g651 ( 
.A(n_450),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_560),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_449),
.A2(n_267),
.B1(n_175),
.B2(n_176),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_575),
.B(n_413),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_582),
.Y(n_655)
);

INVxp33_ASAP7_75t_L g656 ( 
.A(n_468),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_457),
.B(n_413),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_497),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_566),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_516),
.A2(n_417),
.B1(n_419),
.B2(n_187),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_457),
.A2(n_264),
.B1(n_175),
.B2(n_176),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_582),
.B(n_413),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_587),
.Y(n_663)
);

BUFx6f_ASAP7_75t_SL g664 ( 
.A(n_517),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_587),
.B(n_416),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_557),
.A2(n_392),
.B(n_385),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_592),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_497),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_592),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_458),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_458),
.B(n_416),
.Y(n_671)
);

NAND3xp33_ASAP7_75t_L g672 ( 
.A(n_496),
.B(n_206),
.C(n_212),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_461),
.B(n_416),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_461),
.B(n_416),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_577),
.B(n_416),
.Y(n_675)
);

INVx4_ASAP7_75t_L g676 ( 
.A(n_450),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_566),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_581),
.A2(n_392),
.B(n_385),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_510),
.B(n_171),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_503),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_455),
.B(n_416),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_503),
.Y(n_682)
);

NAND2xp33_ASAP7_75t_L g683 ( 
.A(n_449),
.B(n_171),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_525),
.B(n_179),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_538),
.B(n_416),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_577),
.B(n_179),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_485),
.B(n_180),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_450),
.A2(n_185),
.B1(n_180),
.B2(n_181),
.Y(n_688)
);

INVx8_ASAP7_75t_L g689 ( 
.A(n_449),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_452),
.B(n_181),
.Y(n_690)
);

INVxp33_ASAP7_75t_L g691 ( 
.A(n_595),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_474),
.B(n_185),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_515),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_538),
.B(n_508),
.Y(n_694)
);

HB1xp67_ASAP7_75t_L g695 ( 
.A(n_538),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_508),
.B(n_402),
.Y(n_696)
);

O2A1O1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_494),
.A2(n_581),
.B(n_589),
.C(n_578),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_SL g698 ( 
.A(n_529),
.B(n_517),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_509),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_589),
.A2(n_419),
.B1(n_187),
.B2(n_276),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_509),
.B(n_430),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_519),
.B(n_430),
.Y(n_702)
);

NAND3xp33_ASAP7_75t_L g703 ( 
.A(n_553),
.B(n_259),
.C(n_221),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_519),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_L g705 ( 
.A(n_471),
.B(n_264),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_561),
.B(n_363),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_471),
.A2(n_184),
.B1(n_188),
.B2(n_287),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_495),
.B(n_562),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_517),
.B(n_368),
.Y(n_709)
);

NOR3xp33_ASAP7_75t_L g710 ( 
.A(n_466),
.B(n_352),
.C(n_347),
.Y(n_710)
);

INVx1_ASAP7_75t_SL g711 ( 
.A(n_506),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_467),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_475),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_474),
.B(n_266),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_520),
.B(n_430),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_555),
.A2(n_394),
.B(n_387),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_571),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_467),
.B(n_395),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_571),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_490),
.B(n_266),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_476),
.B(n_395),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_580),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_476),
.B(n_478),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_512),
.B(n_267),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_478),
.B(n_395),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_580),
.B(n_351),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_479),
.B(n_395),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_479),
.B(n_400),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_591),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_502),
.B(n_273),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_482),
.B(n_400),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_482),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_494),
.B(n_400),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_471),
.B(n_400),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_533),
.B(n_273),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_470),
.B(n_275),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_490),
.A2(n_492),
.B1(n_450),
.B2(n_570),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_591),
.Y(n_738)
);

INVx1_ASAP7_75t_SL g739 ( 
.A(n_500),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_499),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_492),
.B(n_278),
.Y(n_741)
);

A2O1A1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_586),
.A2(n_351),
.B(n_352),
.C(n_355),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_574),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_570),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_471),
.B(n_464),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_545),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_499),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_507),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_507),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_471),
.A2(n_188),
.B1(n_268),
.B2(n_281),
.Y(n_750)
);

BUFx5_ASAP7_75t_L g751 ( 
.A(n_563),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_471),
.B(n_400),
.Y(n_752)
);

O2A1O1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_588),
.A2(n_330),
.B(n_329),
.C(n_394),
.Y(n_753)
);

INVxp67_ASAP7_75t_SL g754 ( 
.A(n_518),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_471),
.B(n_400),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_518),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_521),
.Y(n_757)
);

NAND3xp33_ASAP7_75t_L g758 ( 
.A(n_480),
.B(n_235),
.C(n_241),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_464),
.B(n_394),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_521),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_523),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_464),
.B(n_387),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_603),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_619),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_606),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_708),
.B(n_491),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_615),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_615),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_708),
.B(n_545),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_638),
.A2(n_563),
.B1(n_554),
.B2(n_448),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_624),
.B(n_743),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_596),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_R g773 ( 
.A(n_643),
.B(n_500),
.Y(n_773)
);

BUFx2_ASAP7_75t_L g774 ( 
.A(n_713),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_614),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_SL g776 ( 
.A1(n_691),
.A2(n_281),
.B1(n_268),
.B2(n_276),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_638),
.B(n_278),
.Y(n_777)
);

NOR3xp33_ASAP7_75t_SL g778 ( 
.A(n_672),
.B(n_287),
.C(n_297),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_626),
.B(n_563),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_614),
.B(n_456),
.Y(n_780)
);

OAI21xp5_ASAP7_75t_L g781 ( 
.A1(n_639),
.A2(n_563),
.B(n_593),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_599),
.Y(n_782)
);

NOR2x2_ASAP7_75t_L g783 ( 
.A(n_738),
.B(n_515),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_659),
.B(n_456),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_618),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_616),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_625),
.B(n_563),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_627),
.B(n_280),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_634),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_604),
.B(n_709),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_632),
.B(n_601),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_724),
.A2(n_563),
.B1(n_448),
.B2(n_590),
.Y(n_792)
);

NOR3xp33_ASAP7_75t_SL g793 ( 
.A(n_602),
.B(n_302),
.C(n_301),
.Y(n_793)
);

NAND2x1p5_ASAP7_75t_L g794 ( 
.A(n_746),
.B(n_465),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_687),
.B(n_679),
.Y(n_795)
);

NAND2xp33_ASAP7_75t_L g796 ( 
.A(n_746),
.B(n_527),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_611),
.Y(n_797)
);

A2O1A1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_679),
.A2(n_542),
.B(n_593),
.C(n_590),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_670),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_680),
.Y(n_800)
);

INVx1_ASAP7_75t_SL g801 ( 
.A(n_711),
.Y(n_801)
);

AND2x4_ASAP7_75t_L g802 ( 
.A(n_677),
.B(n_456),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_649),
.B(n_523),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_723),
.B(n_524),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_682),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_744),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_687),
.A2(n_448),
.B1(n_584),
.B2(n_524),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_630),
.B(n_531),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_650),
.A2(n_551),
.B1(n_584),
.B2(n_531),
.Y(n_809)
);

INVx5_ASAP7_75t_L g810 ( 
.A(n_746),
.Y(n_810)
);

AOI21xp33_ASAP7_75t_L g811 ( 
.A1(n_647),
.A2(n_542),
.B(n_576),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_706),
.Y(n_812)
);

CKINVDCx16_ASAP7_75t_R g813 ( 
.A(n_664),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_648),
.B(n_329),
.Y(n_814)
);

INVx5_ASAP7_75t_L g815 ( 
.A(n_746),
.Y(n_815)
);

OR2x2_ASAP7_75t_SL g816 ( 
.A(n_597),
.B(n_330),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_699),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_636),
.B(n_652),
.Y(n_818)
);

A2O1A1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_647),
.A2(n_537),
.B(n_547),
.C(n_576),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_616),
.B(n_456),
.Y(n_820)
);

INVxp67_ASAP7_75t_SL g821 ( 
.A(n_634),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_695),
.B(n_282),
.Y(n_822)
);

NOR2x1_ASAP7_75t_R g823 ( 
.A(n_693),
.B(n_297),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_704),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_695),
.B(n_744),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_655),
.B(n_537),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_663),
.B(n_547),
.Y(n_827)
);

NAND2x1p5_ASAP7_75t_L g828 ( 
.A(n_651),
.B(n_465),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_656),
.B(n_282),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_605),
.Y(n_830)
);

BUFx2_ASAP7_75t_L g831 ( 
.A(n_739),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_694),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_610),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_637),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_667),
.B(n_549),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_SL g836 ( 
.A1(n_608),
.A2(n_594),
.B(n_465),
.C(n_486),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_669),
.B(n_549),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_726),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_712),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_684),
.B(n_481),
.Y(n_840)
);

NOR2x1_ASAP7_75t_L g841 ( 
.A(n_758),
.B(n_551),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_608),
.B(n_628),
.Y(n_842)
);

INVxp67_ASAP7_75t_L g843 ( 
.A(n_735),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_732),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_598),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_640),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_658),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_598),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_628),
.B(n_730),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_684),
.A2(n_559),
.B1(n_556),
.B2(n_558),
.Y(n_850)
);

BUFx2_ASAP7_75t_L g851 ( 
.A(n_717),
.Y(n_851)
);

INVx4_ASAP7_75t_L g852 ( 
.A(n_598),
.Y(n_852)
);

AOI21xp33_ASAP7_75t_L g853 ( 
.A1(n_700),
.A2(n_559),
.B(n_556),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_668),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_719),
.B(n_481),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_722),
.B(n_481),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_740),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_749),
.Y(n_858)
);

INVx5_ASAP7_75t_L g859 ( 
.A(n_689),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_730),
.B(n_288),
.Y(n_860)
);

AO22x1_ASAP7_75t_L g861 ( 
.A1(n_736),
.A2(n_245),
.B1(n_250),
.B2(n_254),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_685),
.A2(n_540),
.B(n_488),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_729),
.B(n_484),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_736),
.B(n_288),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_600),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_747),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_617),
.B(n_484),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_607),
.Y(n_868)
);

BUFx12f_ASAP7_75t_L g869 ( 
.A(n_664),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_607),
.B(n_558),
.Y(n_870)
);

INVx4_ASAP7_75t_L g871 ( 
.A(n_689),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_609),
.B(n_612),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_735),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_651),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_620),
.B(n_564),
.Y(n_875)
);

INVx4_ASAP7_75t_L g876 ( 
.A(n_689),
.Y(n_876)
);

INVxp67_ASAP7_75t_L g877 ( 
.A(n_698),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_676),
.B(n_292),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_622),
.B(n_564),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_600),
.B(n_565),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_700),
.B(n_565),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_676),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_710),
.B(n_293),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_737),
.A2(n_594),
.B1(n_486),
.B2(n_484),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_748),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_R g886 ( 
.A(n_683),
.B(n_293),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_641),
.B(n_594),
.Y(n_887)
);

AOI22xp5_ASAP7_75t_L g888 ( 
.A1(n_613),
.A2(n_501),
.B1(n_486),
.B2(n_572),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_728),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_686),
.B(n_460),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_703),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_756),
.Y(n_892)
);

OAI21xp33_ASAP7_75t_L g893 ( 
.A1(n_742),
.A2(n_572),
.B(n_536),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_707),
.A2(n_501),
.B1(n_536),
.B2(n_572),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_731),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_653),
.B(n_579),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_635),
.B(n_501),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_701),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_702),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_715),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_757),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_707),
.A2(n_536),
.B1(n_579),
.B2(n_527),
.Y(n_902)
);

INVx5_ASAP7_75t_L g903 ( 
.A(n_751),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_635),
.B(n_579),
.Y(n_904)
);

NAND2x1p5_ASAP7_75t_L g905 ( 
.A(n_675),
.B(n_460),
.Y(n_905)
);

OAI221xp5_ASAP7_75t_L g906 ( 
.A1(n_660),
.A2(n_750),
.B1(n_742),
.B2(n_631),
.C(n_690),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_760),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_761),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_718),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_686),
.B(n_460),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_633),
.Y(n_911)
);

AO21x1_ASAP7_75t_L g912 ( 
.A1(n_697),
.A2(n_473),
.B(n_488),
.Y(n_912)
);

AO22x2_ASAP7_75t_L g913 ( 
.A1(n_661),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_721),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_725),
.Y(n_915)
);

BUFx2_ASAP7_75t_L g916 ( 
.A(n_688),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_671),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_660),
.B(n_674),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_690),
.B(n_573),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_R g920 ( 
.A(n_705),
.B(n_51),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_642),
.B(n_579),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_727),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_613),
.A2(n_573),
.B1(n_544),
.B2(n_540),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_750),
.B(n_579),
.Y(n_924)
);

NOR2x1p5_ASAP7_75t_L g925 ( 
.A(n_745),
.B(n_527),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_644),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_645),
.Y(n_927)
);

INVx5_ASAP7_75t_L g928 ( 
.A(n_751),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_654),
.Y(n_929)
);

AOI22xp5_ASAP7_75t_L g930 ( 
.A1(n_623),
.A2(n_573),
.B1(n_544),
.B2(n_540),
.Y(n_930)
);

OAI221xp5_ASAP7_75t_L g931 ( 
.A1(n_692),
.A2(n_714),
.B1(n_720),
.B2(n_741),
.C(n_629),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_662),
.B(n_527),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_720),
.B(n_527),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_665),
.B(n_544),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_696),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_681),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_646),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_741),
.B(n_488),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_621),
.B(n_629),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_621),
.B(n_473),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_759),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_762),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_623),
.B(n_473),
.Y(n_943)
);

INVxp67_ASAP7_75t_L g944 ( 
.A(n_675),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_646),
.A2(n_469),
.B1(n_493),
.B2(n_483),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_657),
.B(n_0),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_785),
.Y(n_947)
);

BUFx12f_ASAP7_75t_L g948 ( 
.A(n_869),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_849),
.A2(n_673),
.B1(n_657),
.B2(n_755),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_767),
.Y(n_950)
);

INVx4_ASAP7_75t_L g951 ( 
.A(n_845),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_795),
.B(n_673),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_R g953 ( 
.A(n_765),
.B(n_733),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_772),
.Y(n_954)
);

NOR2xp67_ASAP7_75t_L g955 ( 
.A(n_843),
.B(n_734),
.Y(n_955)
);

OAI21xp33_ASAP7_75t_L g956 ( 
.A1(n_860),
.A2(n_753),
.B(n_754),
.Y(n_956)
);

BUFx12f_ASAP7_75t_L g957 ( 
.A(n_774),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_842),
.A2(n_716),
.B(n_666),
.C(n_678),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_873),
.B(n_752),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_939),
.A2(n_751),
.B1(n_493),
.B2(n_483),
.Y(n_960)
);

OAI21xp33_ASAP7_75t_L g961 ( 
.A1(n_790),
.A2(n_1),
.B(n_2),
.Y(n_961)
);

BUFx12f_ASAP7_75t_L g962 ( 
.A(n_764),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_872),
.A2(n_493),
.B(n_483),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_812),
.B(n_5),
.Y(n_964)
);

INVxp67_ASAP7_75t_L g965 ( 
.A(n_801),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_768),
.Y(n_966)
);

OAI22xp33_ASAP7_75t_L g967 ( 
.A1(n_838),
.A2(n_751),
.B1(n_493),
.B2(n_483),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_797),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_903),
.A2(n_751),
.B(n_493),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_903),
.A2(n_751),
.B(n_483),
.Y(n_970)
);

BUFx5_ASAP7_75t_L g971 ( 
.A(n_820),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_820),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_771),
.B(n_832),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_782),
.Y(n_974)
);

CKINVDCx16_ASAP7_75t_R g975 ( 
.A(n_773),
.Y(n_975)
);

OAI21x1_ASAP7_75t_L g976 ( 
.A1(n_862),
.A2(n_469),
.B(n_147),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_903),
.A2(n_469),
.B(n_134),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_770),
.A2(n_11),
.B(n_12),
.C(n_14),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_801),
.B(n_15),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_845),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_903),
.A2(n_469),
.B(n_133),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_816),
.B(n_16),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_928),
.A2(n_123),
.B(n_118),
.Y(n_983)
);

CKINVDCx20_ASAP7_75t_R g984 ( 
.A(n_813),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_799),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_771),
.B(n_115),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_SL g987 ( 
.A1(n_766),
.A2(n_113),
.B(n_103),
.C(n_75),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_800),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_814),
.B(n_16),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_877),
.B(n_19),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_898),
.B(n_73),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_R g992 ( 
.A(n_845),
.B(n_848),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_931),
.A2(n_19),
.B(n_21),
.C(n_22),
.Y(n_993)
);

CKINVDCx20_ASAP7_75t_R g994 ( 
.A(n_831),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_928),
.A2(n_71),
.B(n_70),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_928),
.A2(n_63),
.B(n_60),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_788),
.B(n_24),
.Y(n_997)
);

NAND2xp33_ASAP7_75t_SL g998 ( 
.A(n_806),
.B(n_25),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_865),
.A2(n_906),
.B(n_918),
.C(n_868),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_783),
.Y(n_1000)
);

AND2x4_ASAP7_75t_L g1001 ( 
.A(n_825),
.B(n_26),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_775),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_829),
.B(n_29),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_928),
.A2(n_31),
.B(n_32),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_874),
.A2(n_33),
.B(n_35),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_874),
.A2(n_46),
.B(n_37),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_939),
.A2(n_33),
.B1(n_40),
.B2(n_43),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_899),
.B(n_43),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_SL g1009 ( 
.A1(n_776),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_777),
.A2(n_864),
.B(n_918),
.C(n_769),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_900),
.B(n_791),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_791),
.A2(n_818),
.B(n_822),
.C(n_946),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_810),
.B(n_815),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_882),
.A2(n_872),
.B(n_796),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_805),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_818),
.B(n_935),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_904),
.A2(n_940),
.B1(n_792),
.B2(n_916),
.Y(n_1017)
);

INVx4_ASAP7_75t_L g1018 ( 
.A(n_848),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_824),
.B(n_817),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_926),
.B(n_927),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_808),
.Y(n_1021)
);

OAI22x1_ASAP7_75t_L g1022 ( 
.A1(n_851),
.A2(n_825),
.B1(n_883),
.B2(n_786),
.Y(n_1022)
);

NAND2xp33_ASAP7_75t_SL g1023 ( 
.A(n_806),
.B(n_778),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_909),
.B(n_914),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_878),
.A2(n_891),
.B(n_944),
.C(n_881),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_808),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_915),
.B(n_922),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_806),
.B(n_775),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_775),
.B(n_793),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_848),
.Y(n_1030)
);

O2A1O1Ixp5_ASAP7_75t_SL g1031 ( 
.A1(n_811),
.A2(n_933),
.B(n_853),
.C(n_896),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_810),
.B(n_815),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_889),
.B(n_895),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_763),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_917),
.B(n_941),
.Y(n_1035)
);

AOI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_890),
.A2(n_910),
.B1(n_919),
.B2(n_938),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_866),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_781),
.A2(n_870),
.B(n_887),
.Y(n_1038)
);

O2A1O1Ixp5_ASAP7_75t_L g1039 ( 
.A1(n_836),
.A2(n_924),
.B(n_912),
.C(n_840),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_830),
.Y(n_1040)
);

NOR2xp67_ASAP7_75t_L g1041 ( 
.A(n_839),
.B(n_844),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_882),
.A2(n_887),
.B(n_934),
.Y(n_1042)
);

OA22x2_ASAP7_75t_L g1043 ( 
.A1(n_913),
.A2(n_937),
.B1(n_904),
.B2(n_893),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_826),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_934),
.A2(n_810),
.B(n_815),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_852),
.B(n_871),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_833),
.Y(n_1047)
);

BUFx2_ASAP7_75t_L g1048 ( 
.A(n_823),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_885),
.Y(n_1049)
);

O2A1O1Ixp5_ASAP7_75t_L g1050 ( 
.A1(n_798),
.A2(n_819),
.B(n_811),
.C(n_853),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_917),
.B(n_942),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_841),
.A2(n_779),
.B1(n_787),
.B2(n_925),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_929),
.B(n_804),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_810),
.B(n_815),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_787),
.A2(n_943),
.B(n_921),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_780),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_921),
.A2(n_932),
.B(n_781),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_779),
.A2(n_881),
.B(n_807),
.C(n_880),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_936),
.A2(n_846),
.B1(n_847),
.B2(n_834),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_826),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_861),
.B(n_789),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_932),
.A2(n_803),
.B(n_804),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_803),
.B(n_875),
.Y(n_1063)
);

INVx4_ASAP7_75t_L g1064 ( 
.A(n_852),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_854),
.A2(n_892),
.B1(n_907),
.B2(n_901),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_827),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_940),
.A2(n_897),
.B1(n_902),
.B2(n_821),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_875),
.B(n_879),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_880),
.A2(n_870),
.B(n_863),
.C(n_855),
.Y(n_1069)
);

NAND2x1_ASAP7_75t_L g1070 ( 
.A(n_871),
.B(n_876),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_879),
.A2(n_867),
.B(n_897),
.Y(n_1071)
);

INVx1_ASAP7_75t_SL g1072 ( 
.A(n_780),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_886),
.B(n_908),
.Y(n_1073)
);

HB1xp67_ASAP7_75t_L g1074 ( 
.A(n_857),
.Y(n_1074)
);

BUFx12f_ASAP7_75t_L g1075 ( 
.A(n_876),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_827),
.Y(n_1076)
);

OR2x6_ASAP7_75t_L g1077 ( 
.A(n_784),
.B(n_802),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_859),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_789),
.B(n_784),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_894),
.A2(n_913),
.B1(n_809),
.B2(n_837),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_858),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_913),
.A2(n_837),
.B1(n_835),
.B2(n_856),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_923),
.A2(n_930),
.B(n_835),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_850),
.A2(n_884),
.B(n_888),
.C(n_911),
.Y(n_1084)
);

NOR2xp67_ASAP7_75t_SL g1085 ( 
.A(n_859),
.B(n_920),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_802),
.B(n_905),
.Y(n_1086)
);

BUFx8_ASAP7_75t_L g1087 ( 
.A(n_859),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_905),
.B(n_794),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_859),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_828),
.A2(n_794),
.B(n_945),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_828),
.A2(n_928),
.B(n_903),
.Y(n_1091)
);

NAND3xp33_ASAP7_75t_SL g1092 ( 
.A(n_873),
.B(n_849),
.C(n_795),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_801),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1011),
.B(n_973),
.Y(n_1094)
);

NOR2x1_ASAP7_75t_L g1095 ( 
.A(n_994),
.B(n_1064),
.Y(n_1095)
);

INVx1_ASAP7_75t_SL g1096 ( 
.A(n_947),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1016),
.B(n_952),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_962),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1021),
.B(n_1026),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1044),
.B(n_1060),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_989),
.B(n_1093),
.Y(n_1101)
);

INVxp67_ASAP7_75t_L g1102 ( 
.A(n_965),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_976),
.A2(n_1055),
.B(n_1042),
.Y(n_1103)
);

OAI21xp33_ASAP7_75t_L g1104 ( 
.A1(n_997),
.A2(n_1003),
.B(n_990),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1066),
.B(n_1076),
.Y(n_1105)
);

INVx2_ASAP7_75t_SL g1106 ( 
.A(n_1040),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_1036),
.A2(n_1027),
.B1(n_1024),
.B2(n_1080),
.Y(n_1107)
);

INVx4_ASAP7_75t_L g1108 ( 
.A(n_980),
.Y(n_1108)
);

INVxp67_ASAP7_75t_SL g1109 ( 
.A(n_1053),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_1092),
.B(n_959),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1020),
.B(n_1033),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_974),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_975),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_1057),
.A2(n_1038),
.B(n_1090),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1063),
.B(n_1068),
.Y(n_1115)
);

INVx2_ASAP7_75t_SL g1116 ( 
.A(n_1028),
.Y(n_1116)
);

AOI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1071),
.A2(n_1062),
.B(n_1083),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1063),
.B(n_1068),
.Y(n_1118)
);

INVx2_ASAP7_75t_SL g1119 ( 
.A(n_1002),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_1014),
.A2(n_1091),
.B(n_1050),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_SL g1121 ( 
.A(n_1085),
.B(n_1087),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1058),
.A2(n_956),
.B(n_999),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1045),
.A2(n_1039),
.B(n_970),
.Y(n_1123)
);

OA21x2_ASAP7_75t_L g1124 ( 
.A1(n_963),
.A2(n_1084),
.B(n_960),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_SL g1125 ( 
.A1(n_993),
.A2(n_978),
.B(n_986),
.C(n_991),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_969),
.A2(n_963),
.B(n_1031),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_953),
.B(n_1073),
.Y(n_1127)
);

NOR2xp67_ASAP7_75t_L g1128 ( 
.A(n_1074),
.B(n_1075),
.Y(n_1128)
);

OR2x6_ASAP7_75t_L g1129 ( 
.A(n_1077),
.B(n_1046),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1015),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_958),
.A2(n_1017),
.B(n_1069),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_960),
.A2(n_1086),
.B(n_991),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1086),
.A2(n_1052),
.B(n_977),
.Y(n_1133)
);

INVxp67_ASAP7_75t_SL g1134 ( 
.A(n_1035),
.Y(n_1134)
);

OR2x6_ASAP7_75t_L g1135 ( 
.A(n_1077),
.B(n_1046),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_980),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_981),
.A2(n_986),
.B(n_1025),
.Y(n_1137)
);

BUFx8_ASAP7_75t_L g1138 ( 
.A(n_1000),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1012),
.B(n_1017),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1019),
.B(n_1051),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_1010),
.A2(n_1061),
.B(n_1008),
.C(n_961),
.Y(n_1141)
);

BUFx3_ASAP7_75t_L g1142 ( 
.A(n_980),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_1001),
.B(n_1041),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_955),
.A2(n_1080),
.B(n_949),
.C(n_1088),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1072),
.B(n_988),
.Y(n_1145)
);

OA21x2_ASAP7_75t_L g1146 ( 
.A1(n_1082),
.A2(n_1067),
.B(n_1006),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_1047),
.B(n_1072),
.Y(n_1147)
);

OAI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1067),
.A2(n_1082),
.B(n_1043),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1043),
.A2(n_1005),
.B(n_1004),
.Y(n_1149)
);

NAND3xp33_ASAP7_75t_SL g1150 ( 
.A(n_982),
.B(n_979),
.C(n_998),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1029),
.B(n_964),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_950),
.B(n_966),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_1022),
.B(n_985),
.Y(n_1153)
);

AO31x2_ASAP7_75t_L g1154 ( 
.A1(n_1007),
.A2(n_996),
.A3(n_995),
.B(n_983),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_SL g1155 ( 
.A(n_1087),
.B(n_1009),
.Y(n_1155)
);

OA21x2_ASAP7_75t_L g1156 ( 
.A1(n_1065),
.A2(n_1059),
.B(n_1034),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_968),
.A2(n_1077),
.B1(n_1007),
.B2(n_1037),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1049),
.Y(n_1158)
);

AOI211x1_ASAP7_75t_L g1159 ( 
.A1(n_1079),
.A2(n_1032),
.B(n_1054),
.C(n_1013),
.Y(n_1159)
);

NAND3xp33_ASAP7_75t_L g1160 ( 
.A(n_1023),
.B(n_1081),
.C(n_987),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_972),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_967),
.A2(n_1070),
.B(n_972),
.Y(n_1162)
);

AO22x2_ASAP7_75t_L g1163 ( 
.A1(n_951),
.A2(n_1018),
.B1(n_1064),
.B2(n_1078),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1089),
.A2(n_971),
.B(n_992),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_1056),
.Y(n_1165)
);

NOR2xp67_ASAP7_75t_L g1166 ( 
.A(n_951),
.B(n_1018),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_971),
.B(n_1056),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1056),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1089),
.A2(n_1030),
.B(n_971),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_971),
.B(n_1030),
.Y(n_1170)
);

NOR2x1_ASAP7_75t_SL g1171 ( 
.A(n_1089),
.B(n_1030),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1048),
.B(n_984),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_971),
.A2(n_976),
.B(n_1055),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_994),
.Y(n_1174)
);

OAI22x1_ASAP7_75t_L g1175 ( 
.A1(n_997),
.A2(n_873),
.B1(n_849),
.B2(n_1003),
.Y(n_1175)
);

AO31x2_ASAP7_75t_L g1176 ( 
.A1(n_960),
.A2(n_1058),
.A3(n_1082),
.B(n_1083),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1062),
.A2(n_928),
.B(n_903),
.Y(n_1177)
);

INVx8_ASAP7_75t_L g1178 ( 
.A(n_1077),
.Y(n_1178)
);

BUFx12f_ASAP7_75t_L g1179 ( 
.A(n_948),
.Y(n_1179)
);

NAND3xp33_ASAP7_75t_L g1180 ( 
.A(n_997),
.B(n_849),
.C(n_860),
.Y(n_1180)
);

O2A1O1Ixp5_ASAP7_75t_L g1181 ( 
.A1(n_997),
.A2(n_849),
.B(n_795),
.C(n_842),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1011),
.B(n_973),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_976),
.A2(n_1055),
.B(n_1042),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_954),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_976),
.A2(n_1055),
.B(n_1042),
.Y(n_1185)
);

AO21x2_ASAP7_75t_L g1186 ( 
.A1(n_1036),
.A2(n_1083),
.B(n_963),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1062),
.A2(n_928),
.B(n_903),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1011),
.B(n_973),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_976),
.A2(n_1055),
.B(n_1042),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1011),
.B(n_973),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_976),
.A2(n_1055),
.B(n_1042),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_954),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1031),
.A2(n_795),
.B(n_849),
.Y(n_1193)
);

O2A1O1Ixp5_ASAP7_75t_SL g1194 ( 
.A1(n_1007),
.A2(n_842),
.B(n_766),
.C(n_1082),
.Y(n_1194)
);

O2A1O1Ixp5_ASAP7_75t_L g1195 ( 
.A1(n_997),
.A2(n_849),
.B(n_795),
.C(n_842),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1011),
.B(n_973),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_976),
.A2(n_1055),
.B(n_1042),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_954),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_975),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1062),
.A2(n_928),
.B(n_903),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_R g1201 ( 
.A(n_975),
.B(n_606),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_989),
.B(n_790),
.Y(n_1202)
);

NAND2xp33_ASAP7_75t_L g1203 ( 
.A(n_971),
.B(n_795),
.Y(n_1203)
);

O2A1O1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_997),
.A2(n_849),
.B(n_795),
.C(n_842),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1062),
.A2(n_928),
.B(n_903),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1093),
.B(n_698),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1093),
.B(n_698),
.Y(n_1207)
);

INVx4_ASAP7_75t_L g1208 ( 
.A(n_980),
.Y(n_1208)
);

AOI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_997),
.A2(n_849),
.B1(n_873),
.B2(n_860),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1093),
.B(n_698),
.Y(n_1210)
);

AOI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_997),
.A2(n_849),
.B1(n_873),
.B2(n_860),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_980),
.Y(n_1212)
);

OA21x2_ASAP7_75t_L g1213 ( 
.A1(n_1039),
.A2(n_1050),
.B(n_1083),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_980),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1062),
.A2(n_928),
.B(n_903),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1011),
.B(n_973),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_989),
.B(n_790),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1062),
.A2(n_928),
.B(n_903),
.Y(n_1218)
);

AOI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1042),
.A2(n_1071),
.B(n_1057),
.Y(n_1219)
);

OR2x6_ASAP7_75t_L g1220 ( 
.A(n_957),
.B(n_1093),
.Y(n_1220)
);

AOI211x1_ASAP7_75t_L g1221 ( 
.A1(n_973),
.A2(n_906),
.B(n_795),
.C(n_650),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1011),
.B(n_973),
.Y(n_1222)
);

AOI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1042),
.A2(n_1071),
.B(n_1057),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1031),
.A2(n_795),
.B(n_849),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1031),
.A2(n_795),
.B(n_849),
.Y(n_1225)
);

O2A1O1Ixp5_ASAP7_75t_SL g1226 ( 
.A1(n_1007),
.A2(n_842),
.B(n_766),
.C(n_1082),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_989),
.B(n_790),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_976),
.A2(n_1055),
.B(n_1042),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1062),
.A2(n_928),
.B(n_903),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_994),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_976),
.A2(n_1055),
.B(n_1042),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1011),
.B(n_973),
.Y(n_1232)
);

AO21x2_ASAP7_75t_L g1233 ( 
.A1(n_1036),
.A2(n_1083),
.B(n_963),
.Y(n_1233)
);

NAND2x1p5_ASAP7_75t_L g1234 ( 
.A(n_1095),
.B(n_1164),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1173),
.A2(n_1123),
.B(n_1103),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1183),
.A2(n_1189),
.B(n_1185),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1112),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1180),
.A2(n_1211),
.B(n_1209),
.Y(n_1238)
);

OAI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1104),
.A2(n_1195),
.B(n_1181),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1191),
.A2(n_1228),
.B(n_1197),
.Y(n_1240)
);

INVx2_ASAP7_75t_SL g1241 ( 
.A(n_1220),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1231),
.A2(n_1114),
.B(n_1120),
.Y(n_1242)
);

AOI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1122),
.A2(n_1139),
.B(n_1117),
.Y(n_1243)
);

AO31x2_ASAP7_75t_L g1244 ( 
.A1(n_1144),
.A2(n_1107),
.A3(n_1141),
.B(n_1157),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1094),
.B(n_1182),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1204),
.A2(n_1110),
.B(n_1225),
.Y(n_1246)
);

INVxp67_ASAP7_75t_SL g1247 ( 
.A(n_1115),
.Y(n_1247)
);

INVx2_ASAP7_75t_SL g1248 ( 
.A(n_1220),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1094),
.A2(n_1190),
.B1(n_1222),
.B2(n_1232),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1130),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1177),
.A2(n_1205),
.B(n_1200),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_1178),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1178),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_R g1254 ( 
.A(n_1113),
.B(n_1199),
.Y(n_1254)
);

AO21x2_ASAP7_75t_L g1255 ( 
.A1(n_1193),
.A2(n_1224),
.B(n_1225),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1129),
.B(n_1135),
.Y(n_1256)
);

AOI221xp5_ASAP7_75t_L g1257 ( 
.A1(n_1175),
.A2(n_1150),
.B1(n_1125),
.B2(n_1221),
.C(n_1224),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1219),
.A2(n_1223),
.B(n_1187),
.Y(n_1258)
);

AOI221xp5_ASAP7_75t_L g1259 ( 
.A1(n_1193),
.A2(n_1131),
.B1(n_1155),
.B2(n_1148),
.C(n_1217),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1182),
.B(n_1188),
.Y(n_1260)
);

NAND2xp33_ASAP7_75t_L g1261 ( 
.A(n_1115),
.B(n_1118),
.Y(n_1261)
);

INVx5_ASAP7_75t_L g1262 ( 
.A(n_1129),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1129),
.B(n_1135),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1202),
.B(n_1227),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1188),
.A2(n_1190),
.B1(n_1196),
.B2(n_1232),
.Y(n_1265)
);

AOI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1215),
.A2(n_1218),
.B(n_1229),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1126),
.A2(n_1132),
.B(n_1133),
.Y(n_1267)
);

OR2x2_ASAP7_75t_L g1268 ( 
.A(n_1196),
.B(n_1216),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1136),
.Y(n_1269)
);

BUFx12f_ASAP7_75t_L g1270 ( 
.A(n_1179),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1137),
.A2(n_1131),
.B(n_1162),
.Y(n_1271)
);

INVx6_ASAP7_75t_L g1272 ( 
.A(n_1108),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1155),
.A2(n_1097),
.B1(n_1109),
.B2(n_1148),
.Y(n_1273)
);

OA21x2_ASAP7_75t_L g1274 ( 
.A1(n_1149),
.A2(n_1118),
.B(n_1097),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1149),
.A2(n_1226),
.B(n_1194),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1216),
.B(n_1222),
.Y(n_1276)
);

AOI21xp33_ASAP7_75t_L g1277 ( 
.A1(n_1111),
.A2(n_1134),
.B(n_1140),
.Y(n_1277)
);

AO21x2_ASAP7_75t_L g1278 ( 
.A1(n_1186),
.A2(n_1233),
.B(n_1203),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1135),
.Y(n_1279)
);

INVx3_ASAP7_75t_L g1280 ( 
.A(n_1108),
.Y(n_1280)
);

AOI221xp5_ASAP7_75t_L g1281 ( 
.A1(n_1111),
.A2(n_1206),
.B1(n_1210),
.B2(n_1207),
.C(n_1102),
.Y(n_1281)
);

AO21x2_ASAP7_75t_L g1282 ( 
.A1(n_1186),
.A2(n_1233),
.B(n_1160),
.Y(n_1282)
);

A2O1A1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1099),
.A2(n_1105),
.B(n_1100),
.C(n_1198),
.Y(n_1283)
);

AOI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1127),
.A2(n_1151),
.B1(n_1143),
.B2(n_1153),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1213),
.A2(n_1124),
.B(n_1169),
.Y(n_1285)
);

INVx2_ASAP7_75t_SL g1286 ( 
.A(n_1220),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1184),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1213),
.A2(n_1099),
.B(n_1100),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1192),
.Y(n_1289)
);

NAND2x1p5_ASAP7_75t_L g1290 ( 
.A(n_1156),
.B(n_1166),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1124),
.A2(n_1146),
.B(n_1105),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1146),
.A2(n_1152),
.B(n_1156),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1158),
.Y(n_1293)
);

BUFx3_ASAP7_75t_L g1294 ( 
.A(n_1142),
.Y(n_1294)
);

INVx6_ASAP7_75t_L g1295 ( 
.A(n_1208),
.Y(n_1295)
);

NAND2x1p5_ASAP7_75t_L g1296 ( 
.A(n_1208),
.B(n_1096),
.Y(n_1296)
);

AO21x2_ASAP7_75t_L g1297 ( 
.A1(n_1170),
.A2(n_1167),
.B(n_1161),
.Y(n_1297)
);

NOR2xp67_ASAP7_75t_L g1298 ( 
.A(n_1106),
.B(n_1116),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_SL g1299 ( 
.A1(n_1201),
.A2(n_1121),
.B1(n_1147),
.B2(n_1101),
.Y(n_1299)
);

INVx1_ASAP7_75t_SL g1300 ( 
.A(n_1096),
.Y(n_1300)
);

AOI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1163),
.A2(n_1145),
.B(n_1168),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1119),
.B(n_1165),
.Y(n_1302)
);

AOI221xp5_ASAP7_75t_L g1303 ( 
.A1(n_1159),
.A2(n_1172),
.B1(n_1230),
.B2(n_1174),
.C(n_1098),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1154),
.A2(n_1176),
.B(n_1128),
.Y(n_1304)
);

NAND2x1p5_ASAP7_75t_L g1305 ( 
.A(n_1212),
.B(n_1214),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1163),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1171),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1154),
.A2(n_1176),
.B(n_1212),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_SL g1309 ( 
.A1(n_1212),
.A2(n_1214),
.B(n_1138),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1180),
.A2(n_849),
.B(n_795),
.Y(n_1310)
);

NAND3xp33_ASAP7_75t_L g1311 ( 
.A(n_1180),
.B(n_849),
.C(n_1209),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1173),
.A2(n_1123),
.B(n_1103),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_1157),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1178),
.Y(n_1314)
);

AOI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1209),
.A2(n_849),
.B1(n_1211),
.B2(n_1104),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1202),
.B(n_1217),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1209),
.A2(n_1211),
.B1(n_873),
.B2(n_1180),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1157),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1112),
.Y(n_1319)
);

OA21x2_ASAP7_75t_L g1320 ( 
.A1(n_1131),
.A2(n_1039),
.B(n_1126),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1094),
.B(n_1182),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1112),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1173),
.A2(n_1123),
.B(n_1103),
.Y(n_1323)
);

INVx3_ASAP7_75t_L g1324 ( 
.A(n_1178),
.Y(n_1324)
);

AND2x4_ASAP7_75t_L g1325 ( 
.A(n_1129),
.B(n_1135),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_1094),
.B(n_1182),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1157),
.Y(n_1327)
);

OAI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1209),
.A2(n_1211),
.B1(n_1180),
.B2(n_1155),
.Y(n_1328)
);

OA21x2_ASAP7_75t_L g1329 ( 
.A1(n_1131),
.A2(n_1039),
.B(n_1126),
.Y(n_1329)
);

INVx4_ASAP7_75t_SL g1330 ( 
.A(n_1129),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1112),
.Y(n_1331)
);

AO21x2_ASAP7_75t_L g1332 ( 
.A1(n_1193),
.A2(n_1225),
.B(n_1224),
.Y(n_1332)
);

A2O1A1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1180),
.A2(n_849),
.B(n_1204),
.C(n_795),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1180),
.A2(n_849),
.B1(n_1104),
.B2(n_1003),
.Y(n_1334)
);

NAND3xp33_ASAP7_75t_SL g1335 ( 
.A(n_1209),
.B(n_1211),
.C(n_1180),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1173),
.A2(n_1123),
.B(n_1103),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1112),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1202),
.B(n_1217),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_SL g1339 ( 
.A1(n_1149),
.A2(n_1012),
.B(n_1025),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1173),
.A2(n_1123),
.B(n_1103),
.Y(n_1340)
);

INVx1_ASAP7_75t_SL g1341 ( 
.A(n_1096),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1173),
.A2(n_1123),
.B(n_1103),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1202),
.B(n_1217),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1173),
.A2(n_1123),
.B(n_1103),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1129),
.B(n_1135),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1112),
.Y(n_1346)
);

OAI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1209),
.A2(n_1211),
.B1(n_1180),
.B2(n_1155),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1173),
.A2(n_1123),
.B(n_1103),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1173),
.A2(n_1123),
.B(n_1103),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1112),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1173),
.A2(n_1123),
.B(n_1103),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1180),
.B(n_1104),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1094),
.B(n_1182),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1094),
.B(n_1182),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1173),
.A2(n_1123),
.B(n_1103),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1173),
.A2(n_1123),
.B(n_1103),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1112),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_SL g1358 ( 
.A1(n_1155),
.A2(n_849),
.B1(n_1009),
.B2(n_1180),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1173),
.A2(n_1123),
.B(n_1103),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1173),
.A2(n_1123),
.B(n_1103),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1094),
.B(n_1182),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1308),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1264),
.B(n_1316),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1358),
.A2(n_1315),
.B1(n_1334),
.B2(n_1311),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1276),
.B(n_1245),
.Y(n_1365)
);

O2A1O1Ixp5_ASAP7_75t_L g1366 ( 
.A1(n_1246),
.A2(n_1310),
.B(n_1333),
.C(n_1238),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1338),
.B(n_1343),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1276),
.B(n_1260),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_1254),
.Y(n_1369)
);

O2A1O1Ixp5_ASAP7_75t_L g1370 ( 
.A1(n_1333),
.A2(n_1347),
.B(n_1328),
.C(n_1352),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1268),
.B(n_1321),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1358),
.A2(n_1334),
.B1(n_1284),
.B2(n_1273),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1352),
.B(n_1326),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1353),
.B(n_1247),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1330),
.B(n_1256),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_SL g1376 ( 
.A1(n_1249),
.A2(n_1265),
.B(n_1283),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1302),
.B(n_1281),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1354),
.B(n_1361),
.Y(n_1378)
);

O2A1O1Ixp5_ASAP7_75t_L g1379 ( 
.A1(n_1328),
.A2(n_1347),
.B(n_1239),
.C(n_1317),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1273),
.B(n_1299),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1299),
.B(n_1237),
.Y(n_1381)
);

BUFx3_ASAP7_75t_L g1382 ( 
.A(n_1269),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_1297),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_SL g1384 ( 
.A1(n_1283),
.A2(n_1247),
.B(n_1335),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1261),
.B(n_1277),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1259),
.A2(n_1303),
.B1(n_1341),
.B2(n_1300),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1298),
.A2(n_1257),
.B1(n_1296),
.B2(n_1286),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1319),
.B(n_1322),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1322),
.B(n_1331),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1331),
.B(n_1263),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1263),
.B(n_1325),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1261),
.B(n_1335),
.Y(n_1392)
);

BUFx12f_ASAP7_75t_L g1393 ( 
.A(n_1270),
.Y(n_1393)
);

O2A1O1Ixp33_ASAP7_75t_L g1394 ( 
.A1(n_1339),
.A2(n_1241),
.B(n_1248),
.C(n_1318),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1244),
.B(n_1313),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_SL g1396 ( 
.A1(n_1263),
.A2(n_1345),
.B(n_1274),
.Y(n_1396)
);

OA21x2_ASAP7_75t_L g1397 ( 
.A1(n_1275),
.A2(n_1271),
.B(n_1267),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1296),
.Y(n_1398)
);

A2O1A1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1313),
.A2(n_1318),
.B(n_1327),
.C(n_1288),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1337),
.B(n_1346),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1251),
.A2(n_1278),
.B(n_1274),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1244),
.B(n_1327),
.Y(n_1402)
);

O2A1O1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1309),
.A2(n_1234),
.B(n_1289),
.C(n_1287),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1330),
.B(n_1262),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1250),
.Y(n_1405)
);

OA21x2_ASAP7_75t_L g1406 ( 
.A1(n_1267),
.A2(n_1258),
.B(n_1291),
.Y(n_1406)
);

AND2x4_ASAP7_75t_L g1407 ( 
.A(n_1330),
.B(n_1262),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1262),
.A2(n_1279),
.B1(n_1307),
.B2(n_1306),
.Y(n_1408)
);

O2A1O1Ixp5_ASAP7_75t_L g1409 ( 
.A1(n_1243),
.A2(n_1301),
.B(n_1266),
.C(n_1314),
.Y(n_1409)
);

OA21x2_ASAP7_75t_L g1410 ( 
.A1(n_1258),
.A2(n_1285),
.B(n_1242),
.Y(n_1410)
);

INVx2_ASAP7_75t_SL g1411 ( 
.A(n_1269),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1350),
.B(n_1357),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1293),
.B(n_1274),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_SL g1414 ( 
.A1(n_1279),
.A2(n_1234),
.B(n_1290),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1244),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_SL g1416 ( 
.A1(n_1279),
.A2(n_1290),
.B(n_1294),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_1294),
.Y(n_1417)
);

NAND2x1p5_ASAP7_75t_L g1418 ( 
.A(n_1262),
.B(n_1279),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_1254),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1252),
.B(n_1314),
.Y(n_1420)
);

BUFx12f_ASAP7_75t_L g1421 ( 
.A(n_1270),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1304),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_1272),
.Y(n_1423)
);

A2O1A1Ixp33_ASAP7_75t_L g1424 ( 
.A1(n_1292),
.A2(n_1324),
.B(n_1253),
.C(n_1252),
.Y(n_1424)
);

OA21x2_ASAP7_75t_L g1425 ( 
.A1(n_1235),
.A2(n_1360),
.B(n_1356),
.Y(n_1425)
);

CKINVDCx20_ASAP7_75t_R g1426 ( 
.A(n_1272),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_SL g1427 ( 
.A1(n_1272),
.A2(n_1295),
.B1(n_1305),
.B2(n_1280),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1295),
.A2(n_1280),
.B1(n_1320),
.B2(n_1329),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1278),
.A2(n_1282),
.B(n_1236),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1282),
.Y(n_1430)
);

NOR2xp67_ASAP7_75t_L g1431 ( 
.A(n_1295),
.B(n_1329),
.Y(n_1431)
);

NAND2xp33_ASAP7_75t_SL g1432 ( 
.A(n_1255),
.B(n_1332),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1320),
.A2(n_1329),
.B1(n_1332),
.B2(n_1255),
.Y(n_1433)
);

AOI21x1_ASAP7_75t_SL g1434 ( 
.A1(n_1320),
.A2(n_1359),
.B(n_1349),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1236),
.A2(n_1240),
.B(n_1312),
.Y(n_1435)
);

NOR2x1_ASAP7_75t_SL g1436 ( 
.A(n_1323),
.B(n_1348),
.Y(n_1436)
);

A2O1A1Ixp33_ASAP7_75t_L g1437 ( 
.A1(n_1336),
.A2(n_1312),
.B(n_1340),
.C(n_1342),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1340),
.B(n_1342),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1344),
.B(n_1351),
.Y(n_1439)
);

AOI221x1_ASAP7_75t_SL g1440 ( 
.A1(n_1355),
.A2(n_1104),
.B1(n_1180),
.B2(n_1311),
.C(n_1352),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1355),
.B(n_1264),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1268),
.B(n_1321),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1358),
.A2(n_1209),
.B1(n_1211),
.B2(n_873),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_SL g1444 ( 
.A1(n_1333),
.A2(n_849),
.B(n_795),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1269),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1276),
.B(n_1245),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1358),
.A2(n_1209),
.B1(n_1211),
.B2(n_873),
.Y(n_1447)
);

CKINVDCx20_ASAP7_75t_R g1448 ( 
.A(n_1254),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1413),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1441),
.B(n_1415),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1429),
.A2(n_1401),
.B(n_1434),
.Y(n_1451)
);

OA21x2_ASAP7_75t_L g1452 ( 
.A1(n_1409),
.A2(n_1399),
.B(n_1437),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1375),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1383),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1383),
.Y(n_1455)
);

AOI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1435),
.A2(n_1433),
.B(n_1430),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1406),
.A2(n_1397),
.B(n_1422),
.Y(n_1457)
);

INVx3_ASAP7_75t_L g1458 ( 
.A(n_1438),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1397),
.B(n_1439),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1362),
.B(n_1395),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1425),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1362),
.B(n_1402),
.Y(n_1462)
);

OA21x2_ASAP7_75t_L g1463 ( 
.A1(n_1399),
.A2(n_1437),
.B(n_1424),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1431),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1425),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1428),
.Y(n_1466)
);

OA21x2_ASAP7_75t_L g1467 ( 
.A1(n_1424),
.A2(n_1366),
.B(n_1379),
.Y(n_1467)
);

OA21x2_ASAP7_75t_L g1468 ( 
.A1(n_1370),
.A2(n_1385),
.B(n_1392),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1374),
.Y(n_1469)
);

CKINVDCx20_ASAP7_75t_R g1470 ( 
.A(n_1419),
.Y(n_1470)
);

BUFx12f_ASAP7_75t_L g1471 ( 
.A(n_1393),
.Y(n_1471)
);

AO21x2_ASAP7_75t_L g1472 ( 
.A1(n_1376),
.A2(n_1436),
.B(n_1384),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1364),
.B(n_1443),
.Y(n_1473)
);

AO21x2_ASAP7_75t_L g1474 ( 
.A1(n_1444),
.A2(n_1396),
.B(n_1372),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1410),
.Y(n_1475)
);

AOI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1432),
.A2(n_1414),
.B(n_1416),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1378),
.B(n_1446),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1405),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1390),
.B(n_1373),
.Y(n_1479)
);

INVx2_ASAP7_75t_SL g1480 ( 
.A(n_1404),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1365),
.B(n_1368),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1408),
.Y(n_1482)
);

OR2x6_ASAP7_75t_L g1483 ( 
.A(n_1404),
.B(n_1407),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1388),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1440),
.B(n_1442),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1418),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1381),
.B(n_1389),
.Y(n_1487)
);

INVxp67_ASAP7_75t_L g1488 ( 
.A(n_1371),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1375),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1454),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1459),
.B(n_1391),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1459),
.B(n_1398),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1459),
.B(n_1363),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1458),
.B(n_1407),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1459),
.B(n_1367),
.Y(n_1495)
);

NOR2x1p5_ASAP7_75t_L g1496 ( 
.A(n_1485),
.B(n_1380),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1450),
.B(n_1412),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1450),
.B(n_1400),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1469),
.B(n_1386),
.Y(n_1499)
);

NOR2x1_ASAP7_75t_L g1500 ( 
.A(n_1472),
.B(n_1394),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1450),
.B(n_1375),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1450),
.B(n_1377),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1451),
.A2(n_1457),
.B(n_1456),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1473),
.B(n_1387),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1454),
.Y(n_1505)
);

INVxp67_ASAP7_75t_L g1506 ( 
.A(n_1478),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1483),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1473),
.B(n_1447),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1449),
.B(n_1403),
.Y(n_1509)
);

AND2x4_ASAP7_75t_L g1510 ( 
.A(n_1458),
.B(n_1420),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1469),
.B(n_1382),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1458),
.B(n_1382),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1508),
.A2(n_1474),
.B1(n_1468),
.B2(n_1467),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1491),
.B(n_1488),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1508),
.B(n_1485),
.Y(n_1515)
);

OAI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1504),
.A2(n_1485),
.B(n_1468),
.Y(n_1516)
);

NOR2x1_ASAP7_75t_L g1517 ( 
.A(n_1509),
.B(n_1472),
.Y(n_1517)
);

OAI221xp5_ASAP7_75t_L g1518 ( 
.A1(n_1504),
.A2(n_1488),
.B1(n_1468),
.B2(n_1467),
.C(n_1481),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1491),
.B(n_1453),
.Y(n_1519)
);

OAI31xp33_ASAP7_75t_L g1520 ( 
.A1(n_1496),
.A2(n_1482),
.A3(n_1466),
.B(n_1476),
.Y(n_1520)
);

OAI211xp5_ASAP7_75t_L g1521 ( 
.A1(n_1509),
.A2(n_1467),
.B(n_1468),
.C(n_1466),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1492),
.B(n_1449),
.Y(n_1522)
);

NAND3xp33_ASAP7_75t_L g1523 ( 
.A(n_1500),
.B(n_1468),
.C(n_1467),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1491),
.B(n_1489),
.Y(n_1524)
);

INVx3_ASAP7_75t_L g1525 ( 
.A(n_1510),
.Y(n_1525)
);

OR2x6_ASAP7_75t_L g1526 ( 
.A(n_1500),
.B(n_1476),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1496),
.A2(n_1474),
.B1(n_1468),
.B2(n_1467),
.Y(n_1527)
);

OAI21xp33_ASAP7_75t_L g1528 ( 
.A1(n_1499),
.A2(n_1477),
.B(n_1481),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1502),
.B(n_1468),
.Y(n_1529)
);

AOI221xp5_ASAP7_75t_L g1530 ( 
.A1(n_1499),
.A2(n_1481),
.B1(n_1477),
.B2(n_1474),
.C(n_1502),
.Y(n_1530)
);

AOI221xp5_ASAP7_75t_L g1531 ( 
.A1(n_1499),
.A2(n_1477),
.B1(n_1474),
.B2(n_1449),
.C(n_1482),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1490),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_L g1533 ( 
.A(n_1511),
.B(n_1479),
.Y(n_1533)
);

NOR2x1_ASAP7_75t_L g1534 ( 
.A(n_1511),
.B(n_1472),
.Y(n_1534)
);

AO21x2_ASAP7_75t_L g1535 ( 
.A1(n_1503),
.A2(n_1461),
.B(n_1465),
.Y(n_1535)
);

AOI221xp5_ASAP7_75t_L g1536 ( 
.A1(n_1502),
.A2(n_1474),
.B1(n_1482),
.B2(n_1479),
.C(n_1487),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1493),
.B(n_1495),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1493),
.B(n_1453),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1490),
.Y(n_1539)
);

OAI221xp5_ASAP7_75t_L g1540 ( 
.A1(n_1507),
.A2(n_1467),
.B1(n_1480),
.B2(n_1464),
.C(n_1411),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1493),
.B(n_1479),
.Y(n_1541)
);

OAI211xp5_ASAP7_75t_L g1542 ( 
.A1(n_1511),
.A2(n_1467),
.B(n_1463),
.C(n_1452),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_SL g1543 ( 
.A1(n_1496),
.A2(n_1474),
.B1(n_1472),
.B2(n_1463),
.Y(n_1543)
);

NAND4xp25_ASAP7_75t_L g1544 ( 
.A(n_1492),
.B(n_1462),
.C(n_1460),
.D(n_1455),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1501),
.A2(n_1470),
.B1(n_1426),
.B2(n_1423),
.Y(n_1545)
);

OAI31xp33_ASAP7_75t_L g1546 ( 
.A1(n_1507),
.A2(n_1486),
.A3(n_1427),
.B(n_1464),
.Y(n_1546)
);

OAI211xp5_ASAP7_75t_L g1547 ( 
.A1(n_1506),
.A2(n_1463),
.B(n_1452),
.C(n_1478),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1507),
.B(n_1483),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1495),
.B(n_1484),
.Y(n_1549)
);

BUFx6f_ASAP7_75t_L g1550 ( 
.A(n_1494),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_1512),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1495),
.A2(n_1472),
.B1(n_1471),
.B2(n_1470),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1532),
.Y(n_1553)
);

NOR2x1_ASAP7_75t_L g1554 ( 
.A(n_1523),
.B(n_1526),
.Y(n_1554)
);

INVx2_ASAP7_75t_SL g1555 ( 
.A(n_1550),
.Y(n_1555)
);

INVx4_ASAP7_75t_SL g1556 ( 
.A(n_1526),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1535),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1539),
.Y(n_1558)
);

NAND3xp33_ASAP7_75t_SL g1559 ( 
.A(n_1520),
.B(n_1419),
.C(n_1448),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1549),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1535),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1537),
.B(n_1507),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1522),
.Y(n_1563)
);

BUFx3_ASAP7_75t_L g1564 ( 
.A(n_1526),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1534),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1528),
.B(n_1497),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1550),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1541),
.Y(n_1568)
);

INVx4_ASAP7_75t_L g1569 ( 
.A(n_1550),
.Y(n_1569)
);

INVxp67_ASAP7_75t_SL g1570 ( 
.A(n_1517),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1514),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1529),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1533),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1533),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1544),
.Y(n_1575)
);

INVx4_ASAP7_75t_SL g1576 ( 
.A(n_1550),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1538),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1516),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1519),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1525),
.Y(n_1580)
);

OA21x2_ASAP7_75t_L g1581 ( 
.A1(n_1547),
.A2(n_1475),
.B(n_1461),
.Y(n_1581)
);

AND2x4_ASAP7_75t_SL g1582 ( 
.A(n_1548),
.B(n_1483),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1525),
.Y(n_1583)
);

BUFx3_ASAP7_75t_L g1584 ( 
.A(n_1540),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1576),
.B(n_1524),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1575),
.B(n_1518),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1553),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1575),
.B(n_1515),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1553),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1578),
.B(n_1515),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1576),
.B(n_1501),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1576),
.B(n_1543),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1576),
.B(n_1543),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1576),
.B(n_1527),
.Y(n_1594)
);

NAND2x1p5_ASAP7_75t_L g1595 ( 
.A(n_1554),
.B(n_1463),
.Y(n_1595)
);

NAND2x1_ASAP7_75t_L g1596 ( 
.A(n_1554),
.B(n_1527),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1578),
.A2(n_1530),
.B1(n_1531),
.B2(n_1536),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1573),
.B(n_1521),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1557),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1576),
.B(n_1552),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1559),
.A2(n_1513),
.B1(n_1552),
.B2(n_1546),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1558),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1582),
.B(n_1551),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1582),
.B(n_1510),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1582),
.B(n_1510),
.Y(n_1605)
);

NAND4xp25_ASAP7_75t_L g1606 ( 
.A(n_1584),
.B(n_1513),
.C(n_1542),
.D(n_1545),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1556),
.B(n_1582),
.Y(n_1607)
);

AND2x2_ASAP7_75t_SL g1608 ( 
.A(n_1581),
.B(n_1463),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1573),
.B(n_1497),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1562),
.B(n_1567),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1558),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1562),
.B(n_1510),
.Y(n_1612)
);

AOI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1559),
.A2(n_1452),
.B(n_1483),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1574),
.B(n_1497),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1574),
.B(n_1568),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1563),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1563),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1557),
.Y(n_1618)
);

NAND4xp25_ASAP7_75t_L g1619 ( 
.A(n_1584),
.B(n_1460),
.C(n_1462),
.D(n_1455),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1566),
.B(n_1498),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1568),
.B(n_1505),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1571),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1566),
.B(n_1498),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1556),
.B(n_1501),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1567),
.B(n_1510),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1602),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1591),
.B(n_1556),
.Y(n_1627)
);

INVx1_ASAP7_75t_SL g1628 ( 
.A(n_1585),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1610),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1602),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1587),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1591),
.B(n_1556),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1610),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1599),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1587),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1589),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1599),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1611),
.Y(n_1638)
);

AOI32xp33_ASAP7_75t_L g1639 ( 
.A1(n_1597),
.A2(n_1584),
.A3(n_1564),
.B1(n_1570),
.B2(n_1565),
.Y(n_1639)
);

OAI21xp33_ASAP7_75t_L g1640 ( 
.A1(n_1606),
.A2(n_1584),
.B(n_1564),
.Y(n_1640)
);

OAI21xp33_ASAP7_75t_L g1641 ( 
.A1(n_1590),
.A2(n_1586),
.B(n_1596),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1611),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1615),
.B(n_1572),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1588),
.B(n_1571),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1586),
.B(n_1577),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1589),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1598),
.B(n_1577),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1591),
.B(n_1556),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1598),
.B(n_1579),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1620),
.B(n_1471),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1622),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1615),
.B(n_1572),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_L g1653 ( 
.A(n_1623),
.B(n_1471),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1622),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1616),
.B(n_1560),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1616),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1600),
.B(n_1556),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1617),
.B(n_1560),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1618),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1617),
.B(n_1621),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1631),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1635),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1657),
.B(n_1632),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1640),
.B(n_1609),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1628),
.Y(n_1665)
);

NOR2xp67_ASAP7_75t_L g1666 ( 
.A(n_1632),
.B(n_1607),
.Y(n_1666)
);

CKINVDCx16_ASAP7_75t_R g1667 ( 
.A(n_1657),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1632),
.B(n_1600),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1629),
.Y(n_1669)
);

AO21x1_ASAP7_75t_L g1670 ( 
.A1(n_1646),
.A2(n_1596),
.B(n_1570),
.Y(n_1670)
);

INVx3_ASAP7_75t_L g1671 ( 
.A(n_1627),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1627),
.B(n_1607),
.Y(n_1672)
);

INVxp67_ASAP7_75t_SL g1673 ( 
.A(n_1636),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1641),
.B(n_1614),
.Y(n_1674)
);

AOI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1650),
.A2(n_1601),
.B1(n_1593),
.B2(n_1592),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1660),
.Y(n_1676)
);

INVx1_ASAP7_75t_SL g1677 ( 
.A(n_1648),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1639),
.B(n_1619),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1629),
.B(n_1621),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1644),
.B(n_1594),
.Y(n_1680)
);

INVx3_ASAP7_75t_L g1681 ( 
.A(n_1648),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1653),
.B(n_1393),
.Y(n_1682)
);

NAND2xp33_ASAP7_75t_R g1683 ( 
.A(n_1645),
.B(n_1369),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1633),
.B(n_1607),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1633),
.B(n_1647),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1663),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1678),
.A2(n_1595),
.B1(n_1608),
.B2(n_1564),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1670),
.B(n_1624),
.Y(n_1688)
);

AOI222xp33_ASAP7_75t_L g1689 ( 
.A1(n_1673),
.A2(n_1646),
.B1(n_1608),
.B2(n_1649),
.C1(n_1656),
.C2(n_1642),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1670),
.A2(n_1593),
.B1(n_1592),
.B2(n_1594),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1663),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1667),
.B(n_1651),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_SL g1693 ( 
.A1(n_1674),
.A2(n_1595),
.B1(n_1608),
.B2(n_1564),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1661),
.Y(n_1694)
);

OAI21xp33_ASAP7_75t_L g1695 ( 
.A1(n_1675),
.A2(n_1595),
.B(n_1654),
.Y(n_1695)
);

AOI21xp33_ASAP7_75t_L g1696 ( 
.A1(n_1683),
.A2(n_1660),
.B(n_1643),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1661),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1665),
.B(n_1656),
.Y(n_1698)
);

OA22x2_ASAP7_75t_L g1699 ( 
.A1(n_1677),
.A2(n_1624),
.B1(n_1565),
.B2(n_1638),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1662),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1682),
.B(n_1421),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1666),
.A2(n_1680),
.B1(n_1664),
.B2(n_1681),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1685),
.B(n_1643),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1662),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1703),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1698),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1694),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1697),
.Y(n_1708)
);

INVx3_ASAP7_75t_L g1709 ( 
.A(n_1686),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1700),
.B(n_1676),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1704),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1692),
.B(n_1685),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1691),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1701),
.B(n_1672),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1689),
.B(n_1676),
.Y(n_1715)
);

AOI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1715),
.A2(n_1688),
.B(n_1689),
.Y(n_1716)
);

AOI221xp5_ASAP7_75t_L g1717 ( 
.A1(n_1715),
.A2(n_1696),
.B1(n_1702),
.B2(n_1695),
.C(n_1687),
.Y(n_1717)
);

OAI32xp33_ASAP7_75t_L g1718 ( 
.A1(n_1706),
.A2(n_1687),
.A3(n_1671),
.B1(n_1681),
.B2(n_1668),
.Y(n_1718)
);

AOI221xp5_ASAP7_75t_L g1719 ( 
.A1(n_1705),
.A2(n_1690),
.B1(n_1693),
.B2(n_1681),
.C(n_1671),
.Y(n_1719)
);

NOR3xp33_ASAP7_75t_SL g1720 ( 
.A(n_1713),
.B(n_1369),
.C(n_1699),
.Y(n_1720)
);

OAI211xp5_ASAP7_75t_L g1721 ( 
.A1(n_1709),
.A2(n_1671),
.B(n_1668),
.C(n_1672),
.Y(n_1721)
);

AOI322xp5_ASAP7_75t_L g1722 ( 
.A1(n_1707),
.A2(n_1684),
.A3(n_1669),
.B1(n_1630),
.B2(n_1638),
.C1(n_1626),
.C2(n_1561),
.Y(n_1722)
);

OAI21xp33_ASAP7_75t_L g1723 ( 
.A1(n_1714),
.A2(n_1684),
.B(n_1669),
.Y(n_1723)
);

AOI322xp5_ASAP7_75t_L g1724 ( 
.A1(n_1708),
.A2(n_1630),
.A3(n_1626),
.B1(n_1557),
.B2(n_1561),
.C1(n_1624),
.C2(n_1659),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1709),
.Y(n_1725)
);

NOR4xp25_ASAP7_75t_L g1726 ( 
.A(n_1710),
.B(n_1679),
.C(n_1637),
.D(n_1634),
.Y(n_1726)
);

OAI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1716),
.A2(n_1712),
.B(n_1710),
.Y(n_1727)
);

O2A1O1Ixp33_ASAP7_75t_L g1728 ( 
.A1(n_1718),
.A2(n_1711),
.B(n_1679),
.C(n_1637),
.Y(n_1728)
);

AOI221xp5_ASAP7_75t_L g1729 ( 
.A1(n_1717),
.A2(n_1659),
.B1(n_1634),
.B2(n_1618),
.C(n_1613),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1725),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1721),
.B(n_1652),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1731),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1727),
.B(n_1723),
.Y(n_1733)
);

INVxp67_ASAP7_75t_L g1734 ( 
.A(n_1730),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1728),
.B(n_1720),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1729),
.B(n_1726),
.Y(n_1736)
);

OAI21xp33_ASAP7_75t_L g1737 ( 
.A1(n_1731),
.A2(n_1719),
.B(n_1722),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1732),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1733),
.Y(n_1739)
);

OAI21xp5_ASAP7_75t_SL g1740 ( 
.A1(n_1735),
.A2(n_1724),
.B(n_1652),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1737),
.A2(n_1658),
.B1(n_1655),
.B2(n_1581),
.Y(n_1741)
);

AOI221xp5_ASAP7_75t_L g1742 ( 
.A1(n_1736),
.A2(n_1658),
.B1(n_1655),
.B2(n_1561),
.C(n_1585),
.Y(n_1742)
);

NOR3xp33_ASAP7_75t_L g1743 ( 
.A(n_1738),
.B(n_1739),
.C(n_1740),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1742),
.B(n_1734),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1741),
.A2(n_1471),
.B1(n_1581),
.B2(n_1569),
.Y(n_1745)
);

INVx2_ASAP7_75t_SL g1746 ( 
.A(n_1744),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1746),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1747),
.A2(n_1743),
.B1(n_1745),
.B2(n_1421),
.Y(n_1748)
);

BUFx2_ASAP7_75t_L g1749 ( 
.A(n_1747),
.Y(n_1749)
);

OAI21xp5_ASAP7_75t_SL g1750 ( 
.A1(n_1748),
.A2(n_1448),
.B(n_1603),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1749),
.A2(n_1569),
.B1(n_1603),
.B2(n_1555),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1750),
.Y(n_1752)
);

NAND2x1_ASAP7_75t_SL g1753 ( 
.A(n_1751),
.B(n_1569),
.Y(n_1753)
);

OAI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1752),
.A2(n_1567),
.B1(n_1555),
.B2(n_1580),
.Y(n_1754)
);

NAND4xp75_ASAP7_75t_L g1755 ( 
.A(n_1754),
.B(n_1753),
.C(n_1417),
.D(n_1445),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1755),
.B(n_1625),
.Y(n_1756)
);

AOI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1756),
.A2(n_1567),
.B1(n_1555),
.B2(n_1569),
.Y(n_1757)
);

AOI221xp5_ASAP7_75t_L g1758 ( 
.A1(n_1757),
.A2(n_1569),
.B1(n_1625),
.B2(n_1583),
.C(n_1580),
.Y(n_1758)
);

AOI211xp5_ASAP7_75t_L g1759 ( 
.A1(n_1758),
.A2(n_1605),
.B(n_1604),
.C(n_1612),
.Y(n_1759)
);


endmodule