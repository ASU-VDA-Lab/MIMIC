module fake_jpeg_12997_n_180 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_180);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_31),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_21),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx24_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_7),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_6),
.B(n_1),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_1),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_9),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_11),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_51),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_58),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_66),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

CKINVDCx6p67_ASAP7_75t_R g92 ( 
.A(n_83),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_27),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_84),
.B(n_85),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_0),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_0),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_88),
.B(n_89),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_2),
.Y(n_89)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_90),
.Y(n_94)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_69),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_97),
.C(n_79),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_79),
.B(n_74),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_100),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_71),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_80),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_104),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_90),
.B(n_78),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_81),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_75),
.Y(n_121)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_10),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_59),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_12),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_109),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_62),
.B1(n_65),
.B2(n_72),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_111),
.B1(n_115),
.B2(n_116),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_94),
.A2(n_73),
.B1(n_66),
.B2(n_55),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_63),
.C(n_67),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_126),
.C(n_124),
.Y(n_138)
);

AND2x6_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_38),
.Y(n_113)
);

AND2x6_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_14),
.Y(n_133)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_61),
.B1(n_64),
.B2(n_56),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_56),
.B1(n_73),
.B2(n_55),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_92),
.Y(n_117)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_118),
.A2(n_120),
.B1(n_122),
.B2(n_26),
.Y(n_147)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_121),
.B(n_18),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_92),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_70),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

NAND2x1p5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_58),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_35),
.C(n_39),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_138),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_131),
.B(n_133),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_17),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_142),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_148),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_20),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_143),
.Y(n_149)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_22),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_147),
.Y(n_162)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_124),
.B(n_28),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_136),
.A2(n_29),
.B(n_33),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_150),
.A2(n_135),
.B(n_128),
.Y(n_168)
);

NOR2x1_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_34),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_145),
.Y(n_167)
);

A2O1A1O1Ixp25_ASAP7_75t_L g169 ( 
.A1(n_153),
.A2(n_134),
.B(n_137),
.C(n_140),
.D(n_150),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_132),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_157),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_43),
.B1(n_45),
.B2(n_48),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_129),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_161)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_161),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_158),
.B(n_155),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_167),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_139),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_168),
.Y(n_172)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_169),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_151),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_173),
.Y(n_175)
);

AOI321xp33_ASAP7_75t_L g174 ( 
.A1(n_171),
.A2(n_162),
.A3(n_166),
.B1(n_165),
.B2(n_159),
.C(n_164),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_175),
.B(n_174),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_176),
.A2(n_172),
.B1(n_170),
.B2(n_160),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_177),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_152),
.B(n_149),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_179),
.B(n_156),
.Y(n_180)
);


endmodule