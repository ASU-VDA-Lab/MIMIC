module fake_jpeg_3313_n_55 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_55);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx13_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_11),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_23),
.A2(n_19),
.B1(n_18),
.B2(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_21),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_22),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_25),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_28),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_29),
.A2(n_18),
.B1(n_23),
.B2(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_23),
.B1(n_24),
.B2(n_21),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_33),
.A2(n_34),
.B1(n_19),
.B2(n_20),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

AOI322xp5_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_20),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_26),
.C(n_16),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_38),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_39),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_19),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_33),
.B(n_34),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_12),
.B(n_13),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_44),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_43),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_46),
.Y(n_51)
);

MAJx2_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_14),
.C(n_15),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_42),
.B1(n_9),
.B2(n_10),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_47),
.Y(n_52)
);

OAI21x1_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_53),
.B(n_50),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_8),
.Y(n_53)
);

AOI21x1_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_9),
.B(n_10),
.Y(n_55)
);


endmodule