module fake_netlist_1_7298_n_923 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_923);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_923;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_911;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_171;
wire n_567;
wire n_809;
wire n_888;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_921;
wire n_543;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_482;
wire n_394;
wire n_243;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_900;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_622;
wire n_549;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_446;
wire n_420;
wire n_423;
wire n_165;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_716;
wire n_653;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_200;
wire n_208;
wire n_573;
wire n_898;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_733;
wire n_861;
wire n_899;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_721;
wire n_438;
wire n_134;
wire n_656;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_912;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_123;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_916;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_86), .Y(n_110) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_13), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_71), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_17), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_102), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_94), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_69), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_46), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_15), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_57), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_22), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_24), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_62), .Y(n_122) );
BUFx2_ASAP7_75t_L g123 ( .A(n_67), .Y(n_123) );
BUFx10_ASAP7_75t_L g124 ( .A(n_64), .Y(n_124) );
CKINVDCx16_ASAP7_75t_R g125 ( .A(n_22), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_70), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_39), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_52), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_84), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_43), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_17), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_27), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_61), .Y(n_133) );
CKINVDCx14_ASAP7_75t_R g134 ( .A(n_8), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_93), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_76), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_63), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_95), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_99), .Y(n_139) );
BUFx2_ASAP7_75t_L g140 ( .A(n_11), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g141 ( .A(n_82), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_50), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_45), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_91), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_3), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_21), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_38), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_27), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_72), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_4), .Y(n_150) );
BUFx3_ASAP7_75t_L g151 ( .A(n_58), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_83), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_79), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_25), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_114), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_131), .Y(n_156) );
INVx5_ASAP7_75t_L g157 ( .A(n_114), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_131), .Y(n_158) );
INVx4_ASAP7_75t_L g159 ( .A(n_111), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_123), .B(n_0), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_140), .B(n_0), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_114), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_151), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_123), .B(n_1), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_151), .Y(n_165) );
AND2x4_ASAP7_75t_L g166 ( .A(n_151), .B(n_1), .Y(n_166) );
INVx5_ASAP7_75t_L g167 ( .A(n_124), .Y(n_167) );
HB1xp67_ASAP7_75t_L g168 ( .A(n_134), .Y(n_168) );
BUFx12f_ASAP7_75t_L g169 ( .A(n_124), .Y(n_169) );
BUFx3_ASAP7_75t_L g170 ( .A(n_124), .Y(n_170) );
INVx5_ASAP7_75t_L g171 ( .A(n_124), .Y(n_171) );
BUFx8_ASAP7_75t_SL g172 ( .A(n_140), .Y(n_172) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_111), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_113), .B(n_2), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_111), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_111), .Y(n_176) );
AND2x6_ASAP7_75t_L g177 ( .A(n_131), .B(n_109), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_111), .Y(n_178) );
OAI22xp33_ASAP7_75t_SL g179 ( .A1(n_164), .A2(n_125), .B1(n_118), .B2(n_146), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_167), .B(n_135), .Y(n_180) );
INVx3_ASAP7_75t_L g181 ( .A(n_166), .Y(n_181) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_161), .A2(n_134), .B1(n_125), .B2(n_141), .Y(n_182) );
OAI22xp33_ASAP7_75t_SL g183 ( .A1(n_164), .A2(n_154), .B1(n_132), .B2(n_127), .Y(n_183) );
OAI22xp33_ASAP7_75t_SL g184 ( .A1(n_160), .A2(n_121), .B1(n_148), .B2(n_150), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_159), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_168), .B(n_113), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_167), .B(n_135), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_168), .B(n_120), .Y(n_188) );
OAI22xp33_ASAP7_75t_L g189 ( .A1(n_160), .A2(n_120), .B1(n_145), .B2(n_147), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_159), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_161), .A2(n_141), .B1(n_145), .B2(n_147), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_168), .B(n_110), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_161), .A2(n_112), .B1(n_115), .B2(n_111), .Y(n_193) );
AND2x4_ASAP7_75t_L g194 ( .A(n_170), .B(n_142), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_159), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_159), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_166), .Y(n_197) );
AO22x2_ASAP7_75t_L g198 ( .A1(n_166), .A2(n_142), .B1(n_149), .B2(n_116), .Y(n_198) );
INVx1_ASAP7_75t_SL g199 ( .A(n_170), .Y(n_199) );
AO22x2_ASAP7_75t_L g200 ( .A1(n_166), .A2(n_149), .B1(n_116), .B2(n_4), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_166), .Y(n_201) );
OAI22xp33_ASAP7_75t_L g202 ( .A1(n_160), .A2(n_153), .B1(n_152), .B2(n_144), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_166), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_161), .A2(n_143), .B1(n_139), .B2(n_138), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_159), .Y(n_205) );
OAI22xp5_ASAP7_75t_SL g206 ( .A1(n_174), .A2(n_137), .B1(n_136), .B2(n_133), .Y(n_206) );
OAI22xp33_ASAP7_75t_SL g207 ( .A1(n_174), .A2(n_130), .B1(n_129), .B2(n_128), .Y(n_207) );
XNOR2xp5_ASAP7_75t_SL g208 ( .A(n_172), .B(n_2), .Y(n_208) );
OAI22xp33_ASAP7_75t_SL g209 ( .A1(n_174), .A2(n_126), .B1(n_122), .B2(n_119), .Y(n_209) );
OAI22xp33_ASAP7_75t_L g210 ( .A1(n_169), .A2(n_117), .B1(n_5), .B2(n_6), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_159), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_170), .B(n_3), .Y(n_212) );
OAI22xp33_ASAP7_75t_SL g213 ( .A1(n_170), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_166), .Y(n_214) );
OAI22xp5_ASAP7_75t_SL g215 ( .A1(n_172), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_215) );
OAI22xp33_ASAP7_75t_SL g216 ( .A1(n_170), .A2(n_171), .B1(n_167), .B2(n_166), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_159), .Y(n_217) );
OA22x2_ASAP7_75t_L g218 ( .A1(n_156), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_218) );
OAI22xp33_ASAP7_75t_L g219 ( .A1(n_169), .A2(n_10), .B1(n_12), .B2(n_13), .Y(n_219) );
OR2x6_ASAP7_75t_L g220 ( .A(n_169), .B(n_12), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_155), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_169), .B(n_44), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g223 ( .A1(n_169), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_167), .B(n_14), .Y(n_224) );
INVx2_ASAP7_75t_SL g225 ( .A(n_167), .Y(n_225) );
OAI22xp5_ASAP7_75t_SL g226 ( .A1(n_156), .A2(n_16), .B1(n_18), .B2(n_19), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_220), .B(n_167), .Y(n_227) );
CKINVDCx11_ASAP7_75t_R g228 ( .A(n_220), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_225), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_181), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_181), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_181), .Y(n_232) );
BUFx6f_ASAP7_75t_SL g233 ( .A(n_220), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_197), .Y(n_234) );
XNOR2xp5_ASAP7_75t_L g235 ( .A(n_182), .B(n_18), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_221), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_220), .B(n_167), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_197), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_203), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_203), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_214), .Y(n_241) );
XNOR2x2_ASAP7_75t_L g242 ( .A(n_200), .B(n_156), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_225), .Y(n_243) );
BUFx3_ASAP7_75t_L g244 ( .A(n_214), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_201), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_198), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g247 ( .A(n_208), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_198), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_186), .B(n_167), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_186), .B(n_167), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_198), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_192), .B(n_167), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_198), .Y(n_253) );
OR2x6_ASAP7_75t_L g254 ( .A(n_200), .B(n_158), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_194), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_221), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_194), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_194), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_218), .Y(n_259) );
XNOR2xp5_ASAP7_75t_L g260 ( .A(n_193), .B(n_19), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_188), .B(n_167), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_188), .B(n_167), .Y(n_262) );
BUFx3_ASAP7_75t_L g263 ( .A(n_199), .Y(n_263) );
OAI21xp5_ASAP7_75t_L g264 ( .A1(n_185), .A2(n_162), .B(n_163), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_218), .Y(n_265) );
BUFx2_ASAP7_75t_L g266 ( .A(n_200), .Y(n_266) );
XNOR2x2_ASAP7_75t_L g267 ( .A(n_200), .B(n_158), .Y(n_267) );
INVxp67_ASAP7_75t_SL g268 ( .A(n_189), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_191), .B(n_171), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_202), .B(n_171), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_218), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_224), .B(n_171), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_224), .Y(n_273) );
INVxp33_ASAP7_75t_L g274 ( .A(n_206), .Y(n_274) );
NOR2xp33_ASAP7_75t_SL g275 ( .A(n_216), .B(n_171), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_212), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_185), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_204), .B(n_171), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_222), .B(n_171), .Y(n_279) );
XOR2xp5_ASAP7_75t_L g280 ( .A(n_208), .B(n_20), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_190), .Y(n_281) );
XOR2xp5_ASAP7_75t_L g282 ( .A(n_215), .B(n_20), .Y(n_282) );
AND2x6_ASAP7_75t_SL g283 ( .A(n_179), .B(n_158), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_190), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_180), .A2(n_162), .B(n_163), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_195), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_207), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_195), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_223), .B(n_171), .Y(n_289) );
XOR2xp5_ASAP7_75t_L g290 ( .A(n_184), .B(n_21), .Y(n_290) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_226), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_196), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_232), .Y(n_293) );
INVxp67_ASAP7_75t_L g294 ( .A(n_233), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_227), .B(n_171), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_227), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_232), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_268), .B(n_171), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_244), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_244), .Y(n_300) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_263), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_263), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_227), .B(n_171), .Y(n_303) );
BUFx3_ASAP7_75t_L g304 ( .A(n_263), .Y(n_304) );
INVx1_ASAP7_75t_SL g305 ( .A(n_228), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_227), .B(n_171), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_232), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_268), .B(n_183), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_234), .B(n_209), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_277), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_237), .B(n_180), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_277), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_237), .Y(n_313) );
INVx1_ASAP7_75t_SL g314 ( .A(n_237), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g315 ( .A1(n_254), .A2(n_177), .B1(n_219), .B2(n_213), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_244), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_230), .Y(n_317) );
AND2x2_ASAP7_75t_SL g318 ( .A(n_266), .B(n_162), .Y(n_318) );
INVx1_ASAP7_75t_SL g319 ( .A(n_237), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_230), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_231), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_229), .Y(n_322) );
BUFx3_ASAP7_75t_L g323 ( .A(n_229), .Y(n_323) );
OR2x2_ASAP7_75t_SL g324 ( .A(n_246), .B(n_162), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_233), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_234), .B(n_210), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_277), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_231), .Y(n_328) );
OAI21xp5_ASAP7_75t_L g329 ( .A1(n_285), .A2(n_217), .B(n_211), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_238), .B(n_187), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_238), .B(n_187), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_288), .Y(n_332) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_233), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_239), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_229), .Y(n_335) );
BUFx3_ASAP7_75t_L g336 ( .A(n_229), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_288), .Y(n_337) );
INVx3_ASAP7_75t_L g338 ( .A(n_229), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_239), .Y(n_339) );
AND2x2_ASAP7_75t_SL g340 ( .A(n_266), .B(n_162), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_240), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_288), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_240), .B(n_196), .Y(n_343) );
BUFx3_ASAP7_75t_L g344 ( .A(n_229), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_241), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_241), .B(n_205), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_249), .B(n_163), .Y(n_347) );
BUFx6f_ASAP7_75t_SL g348 ( .A(n_318), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_339), .B(n_245), .Y(n_349) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_301), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_313), .B(n_249), .Y(n_351) );
NOR2xp33_ASAP7_75t_SL g352 ( .A(n_318), .B(n_233), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_305), .Y(n_353) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_302), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_339), .B(n_245), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_310), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_310), .Y(n_357) );
INVx5_ASAP7_75t_L g358 ( .A(n_302), .Y(n_358) );
BUFx4f_ASAP7_75t_L g359 ( .A(n_313), .Y(n_359) );
INVx3_ASAP7_75t_L g360 ( .A(n_302), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_339), .B(n_250), .Y(n_361) );
BUFx12f_ASAP7_75t_L g362 ( .A(n_325), .Y(n_362) );
INVx1_ASAP7_75t_SL g363 ( .A(n_302), .Y(n_363) );
AND2x2_ASAP7_75t_SL g364 ( .A(n_318), .B(n_340), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_339), .B(n_250), .Y(n_365) );
NAND2x1p5_ASAP7_75t_L g366 ( .A(n_314), .B(n_259), .Y(n_366) );
AND2x4_ASAP7_75t_L g367 ( .A(n_313), .B(n_296), .Y(n_367) );
NAND2x1p5_ASAP7_75t_L g368 ( .A(n_314), .B(n_259), .Y(n_368) );
INVxp67_ASAP7_75t_SL g369 ( .A(n_302), .Y(n_369) );
BUFx12f_ASAP7_75t_L g370 ( .A(n_325), .Y(n_370) );
CKINVDCx11_ASAP7_75t_R g371 ( .A(n_305), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_326), .B(n_274), .Y(n_372) );
AO21x2_ASAP7_75t_L g373 ( .A1(n_315), .A2(n_248), .B(n_251), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_341), .B(n_265), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_341), .B(n_265), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_313), .B(n_261), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_341), .B(n_271), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_304), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_341), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_334), .Y(n_380) );
NOR2x1_ASAP7_75t_L g381 ( .A(n_309), .B(n_271), .Y(n_381) );
BUFx3_ASAP7_75t_L g382 ( .A(n_358), .Y(n_382) );
BUFx2_ASAP7_75t_SL g383 ( .A(n_358), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g384 ( .A(n_358), .B(n_304), .Y(n_384) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_354), .Y(n_385) );
BUFx8_ASAP7_75t_L g386 ( .A(n_348), .Y(n_386) );
BUFx2_ASAP7_75t_SL g387 ( .A(n_358), .Y(n_387) );
BUFx2_ASAP7_75t_L g388 ( .A(n_369), .Y(n_388) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_354), .Y(n_389) );
BUFx3_ASAP7_75t_L g390 ( .A(n_358), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_356), .Y(n_391) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_364), .A2(n_254), .B1(n_318), .B2(n_340), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_379), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_371), .Y(n_394) );
BUFx2_ASAP7_75t_L g395 ( .A(n_369), .Y(n_395) );
BUFx12f_ASAP7_75t_L g396 ( .A(n_371), .Y(n_396) );
CKINVDCx11_ASAP7_75t_R g397 ( .A(n_362), .Y(n_397) );
BUFx3_ASAP7_75t_L g398 ( .A(n_358), .Y(n_398) );
BUFx3_ASAP7_75t_L g399 ( .A(n_358), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_379), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_356), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_379), .Y(n_402) );
INVx1_ASAP7_75t_SL g403 ( .A(n_356), .Y(n_403) );
INVx8_ASAP7_75t_L g404 ( .A(n_348), .Y(n_404) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_354), .Y(n_405) );
INVx3_ASAP7_75t_L g406 ( .A(n_358), .Y(n_406) );
CKINVDCx16_ASAP7_75t_R g407 ( .A(n_352), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_380), .Y(n_408) );
AND2x4_ASAP7_75t_L g409 ( .A(n_356), .B(n_304), .Y(n_409) );
NAND2x1p5_ASAP7_75t_L g410 ( .A(n_358), .B(n_304), .Y(n_410) );
OR2x2_ASAP7_75t_SL g411 ( .A(n_348), .B(n_333), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_408), .Y(n_412) );
OAI21xp5_ASAP7_75t_SL g413 ( .A1(n_392), .A2(n_280), .B(n_305), .Y(n_413) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_385), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_392), .A2(n_348), .B1(n_364), .B2(n_372), .Y(n_415) );
AOI22xp33_ASAP7_75t_SL g416 ( .A1(n_407), .A2(n_352), .B1(n_348), .B2(n_364), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_407), .A2(n_372), .B1(n_348), .B2(n_364), .Y(n_417) );
NAND2x1p5_ASAP7_75t_L g418 ( .A(n_406), .B(n_358), .Y(n_418) );
AOI22xp33_ASAP7_75t_SL g419 ( .A1(n_383), .A2(n_364), .B1(n_242), .B2(n_267), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_408), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_391), .Y(n_421) );
OAI21xp33_ASAP7_75t_SL g422 ( .A1(n_403), .A2(n_254), .B(n_248), .Y(n_422) );
BUFx12f_ASAP7_75t_L g423 ( .A(n_397), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_386), .A2(n_254), .B1(n_260), .B2(n_315), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_391), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_391), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_401), .Y(n_427) );
INVx3_ASAP7_75t_L g428 ( .A(n_382), .Y(n_428) );
BUFx8_ASAP7_75t_L g429 ( .A(n_396), .Y(n_429) );
BUFx3_ASAP7_75t_L g430 ( .A(n_382), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_401), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_386), .A2(n_260), .B1(n_254), .B2(n_235), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_386), .A2(n_235), .B1(n_290), .B2(n_340), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_401), .B(n_357), .Y(n_434) );
BUFx8_ASAP7_75t_L g435 ( .A(n_396), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_393), .Y(n_436) );
AOI22xp33_ASAP7_75t_SL g437 ( .A1(n_383), .A2(n_267), .B1(n_242), .B2(n_340), .Y(n_437) );
BUFx3_ASAP7_75t_L g438 ( .A(n_382), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_386), .A2(n_290), .B1(n_340), .B2(n_318), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_396), .Y(n_440) );
INVx6_ASAP7_75t_L g441 ( .A(n_386), .Y(n_441) );
BUFx3_ASAP7_75t_L g442 ( .A(n_382), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_386), .A2(n_340), .B1(n_318), .B2(n_291), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_388), .A2(n_349), .B1(n_355), .B2(n_315), .Y(n_444) );
OAI21xp5_ASAP7_75t_L g445 ( .A1(n_403), .A2(n_308), .B(n_309), .Y(n_445) );
AOI22xp33_ASAP7_75t_SL g446 ( .A1(n_383), .A2(n_333), .B1(n_247), .B2(n_370), .Y(n_446) );
OAI21xp5_ASAP7_75t_SL g447 ( .A1(n_406), .A2(n_280), .B(n_282), .Y(n_447) );
CKINVDCx11_ASAP7_75t_R g448 ( .A(n_396), .Y(n_448) );
INVx3_ASAP7_75t_L g449 ( .A(n_390), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_393), .Y(n_450) );
INVx6_ASAP7_75t_L g451 ( .A(n_390), .Y(n_451) );
INVx2_ASAP7_75t_SL g452 ( .A(n_390), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_404), .A2(n_287), .B1(n_308), .B2(n_373), .Y(n_453) );
BUFx12f_ASAP7_75t_L g454 ( .A(n_397), .Y(n_454) );
INVx2_ASAP7_75t_SL g455 ( .A(n_390), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_404), .A2(n_308), .B1(n_373), .B2(n_376), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_424), .A2(n_404), .B1(n_373), .B2(n_387), .Y(n_457) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_424), .A2(n_411), .B1(n_388), .B2(n_395), .Y(n_458) );
INVx4_ASAP7_75t_L g459 ( .A(n_441), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_421), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_421), .Y(n_461) );
AOI22xp33_ASAP7_75t_SL g462 ( .A1(n_441), .A2(n_404), .B1(n_387), .B2(n_398), .Y(n_462) );
AOI22xp33_ASAP7_75t_SL g463 ( .A1(n_441), .A2(n_404), .B1(n_387), .B2(n_398), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_444), .A2(n_282), .B1(n_373), .B2(n_404), .Y(n_464) );
BUFx4f_ASAP7_75t_SL g465 ( .A(n_423), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_415), .A2(n_404), .B1(n_373), .B2(n_351), .Y(n_466) );
CKINVDCx11_ASAP7_75t_R g467 ( .A(n_423), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_432), .A2(n_411), .B1(n_388), .B2(n_395), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_439), .A2(n_373), .B1(n_351), .B2(n_376), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_433), .A2(n_376), .B1(n_351), .B2(n_365), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_421), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_443), .A2(n_376), .B1(n_351), .B2(n_365), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_412), .Y(n_473) );
OAI22xp33_ASAP7_75t_L g474 ( .A1(n_413), .A2(n_394), .B1(n_395), .B2(n_399), .Y(n_474) );
BUFx2_ASAP7_75t_L g475 ( .A(n_422), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_453), .A2(n_376), .B1(n_351), .B2(n_365), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_427), .Y(n_477) );
BUFx4f_ASAP7_75t_SL g478 ( .A(n_423), .Y(n_478) );
BUFx3_ASAP7_75t_L g479 ( .A(n_430), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_417), .A2(n_376), .B1(n_351), .B2(n_365), .Y(n_480) );
AOI22xp33_ASAP7_75t_SL g481 ( .A1(n_441), .A2(n_398), .B1(n_399), .B2(n_406), .Y(n_481) );
OAI22xp33_ASAP7_75t_SL g482 ( .A1(n_441), .A2(n_394), .B1(n_353), .B2(n_384), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_416), .A2(n_411), .B1(n_398), .B2(n_399), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_417), .A2(n_399), .B1(n_406), .B2(n_410), .Y(n_484) );
INVx4_ASAP7_75t_SL g485 ( .A(n_451), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_412), .Y(n_486) );
BUFx12f_ASAP7_75t_L g487 ( .A(n_429), .Y(n_487) );
OAI21xp5_ASAP7_75t_SL g488 ( .A1(n_447), .A2(n_294), .B(n_333), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_419), .A2(n_361), .B1(n_381), .B2(n_309), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_427), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_434), .B(n_400), .Y(n_491) );
AOI22xp33_ASAP7_75t_SL g492 ( .A1(n_429), .A2(n_406), .B1(n_370), .B2(n_362), .Y(n_492) );
OAI22xp5_ASAP7_75t_SL g493 ( .A1(n_454), .A2(n_353), .B1(n_362), .B2(n_370), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_437), .A2(n_410), .B1(n_380), .B2(n_349), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_446), .A2(n_410), .B1(n_380), .B2(n_355), .Y(n_495) );
OAI22xp5_ASAP7_75t_SL g496 ( .A1(n_454), .A2(n_370), .B1(n_362), .B2(n_294), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_454), .B(n_283), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_456), .A2(n_410), .B1(n_294), .B2(n_301), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_429), .A2(n_361), .B1(n_381), .B2(n_402), .Y(n_499) );
INVx5_ASAP7_75t_L g500 ( .A(n_451), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_429), .A2(n_361), .B1(n_381), .B2(n_402), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_427), .B(n_385), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_418), .A2(n_410), .B1(n_301), .B2(n_400), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_434), .B(n_361), .Y(n_504) );
BUFx4f_ASAP7_75t_SL g505 ( .A(n_435), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_431), .B(n_409), .Y(n_506) );
BUFx4f_ASAP7_75t_SL g507 ( .A(n_435), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_420), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_435), .A2(n_367), .B1(n_409), .B2(n_359), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_420), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_435), .A2(n_367), .B1(n_409), .B2(n_359), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_418), .A2(n_455), .B1(n_452), .B2(n_451), .Y(n_512) );
OAI21xp5_ASAP7_75t_SL g513 ( .A1(n_418), .A2(n_269), .B(n_326), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_431), .B(n_409), .Y(n_514) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_422), .A2(n_326), .B(n_289), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_452), .A2(n_269), .B1(n_289), .B2(n_278), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_431), .B(n_409), .Y(n_517) );
INVx3_ASAP7_75t_L g518 ( .A(n_428), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_430), .A2(n_367), .B1(n_409), .B2(n_359), .Y(n_519) );
BUFx2_ASAP7_75t_L g520 ( .A(n_430), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_436), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_455), .A2(n_253), .B1(n_251), .B2(n_246), .Y(n_522) );
CKINVDCx14_ASAP7_75t_R g523 ( .A(n_448), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_436), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_438), .A2(n_442), .B1(n_445), .B2(n_451), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_438), .A2(n_367), .B1(n_359), .B2(n_345), .Y(n_526) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_414), .Y(n_527) );
CKINVDCx5p33_ASAP7_75t_R g528 ( .A(n_440), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_450), .B(n_357), .Y(n_529) );
OR2x2_ASAP7_75t_SL g530 ( .A(n_451), .B(n_385), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_425), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_464), .A2(n_442), .B1(n_438), .B2(n_449), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_464), .A2(n_442), .B1(n_449), .B2(n_428), .Y(n_533) );
OAI22xp33_ASAP7_75t_L g534 ( .A1(n_495), .A2(n_449), .B1(n_428), .B2(n_426), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_474), .A2(n_449), .B1(n_428), .B2(n_450), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_473), .B(n_425), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_513), .A2(n_426), .B1(n_350), .B2(n_357), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_457), .A2(n_350), .B1(n_177), .B2(n_384), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_458), .A2(n_177), .B1(n_378), .B2(n_253), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_468), .A2(n_466), .B1(n_475), .B2(n_480), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_475), .A2(n_177), .B1(n_378), .B2(n_360), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_469), .A2(n_177), .B1(n_378), .B2(n_360), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_473), .Y(n_543) );
INVxp67_ASAP7_75t_L g544 ( .A(n_520), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_494), .A2(n_177), .B1(n_378), .B2(n_360), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_489), .A2(n_324), .B1(n_357), .B2(n_366), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_497), .A2(n_177), .B1(n_360), .B2(n_354), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_472), .A2(n_177), .B1(n_360), .B2(n_354), .Y(n_548) );
AOI22xp33_ASAP7_75t_SL g549 ( .A1(n_505), .A2(n_414), .B1(n_405), .B2(n_389), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_470), .A2(n_177), .B1(n_360), .B2(n_354), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_515), .A2(n_177), .B1(n_354), .B2(n_367), .Y(n_551) );
OAI222xp33_ASAP7_75t_L g552 ( .A1(n_459), .A2(n_366), .B1(n_368), .B2(n_363), .C1(n_163), .C2(n_314), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_462), .A2(n_324), .B1(n_366), .B2(n_368), .Y(n_553) );
OAI222xp33_ASAP7_75t_L g554 ( .A1(n_459), .A2(n_366), .B1(n_368), .B2(n_363), .C1(n_163), .C2(n_319), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_486), .B(n_283), .Y(n_555) );
OAI211xp5_ASAP7_75t_SL g556 ( .A1(n_467), .A2(n_178), .B(n_273), .C(n_276), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_487), .A2(n_345), .B1(n_334), .B2(n_375), .Y(n_557) );
AOI221xp5_ASAP7_75t_L g558 ( .A1(n_482), .A2(n_273), .B1(n_178), .B2(n_165), .C(n_155), .Y(n_558) );
OAI222xp33_ASAP7_75t_L g559 ( .A1(n_459), .A2(n_366), .B1(n_368), .B2(n_319), .C1(n_375), .C2(n_374), .Y(n_559) );
OAI22xp33_ASAP7_75t_L g560 ( .A1(n_507), .A2(n_359), .B1(n_368), .B2(n_389), .Y(n_560) );
AOI22xp33_ASAP7_75t_SL g561 ( .A1(n_487), .A2(n_414), .B1(n_405), .B2(n_389), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_492), .A2(n_324), .B1(n_359), .B2(n_389), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_486), .B(n_385), .Y(n_563) );
INVx2_ASAP7_75t_SL g564 ( .A(n_479), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_506), .B(n_414), .Y(n_565) );
AOI22xp33_ASAP7_75t_SL g566 ( .A1(n_483), .A2(n_414), .B1(n_405), .B2(n_389), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_508), .B(n_385), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_476), .A2(n_177), .B1(n_354), .B2(n_367), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_463), .A2(n_324), .B1(n_405), .B2(n_389), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_508), .B(n_510), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_499), .A2(n_177), .B1(n_354), .B2(n_389), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_510), .B(n_385), .Y(n_572) );
NOR3xp33_ASAP7_75t_L g573 ( .A(n_488), .B(n_178), .C(n_276), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_501), .A2(n_177), .B1(n_405), .B2(n_389), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_484), .A2(n_177), .B1(n_405), .B2(n_385), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_516), .A2(n_334), .B1(n_345), .B2(n_374), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_503), .A2(n_377), .B1(n_320), .B2(n_321), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_504), .A2(n_405), .B1(n_385), .B2(n_414), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_498), .A2(n_405), .B1(n_304), .B2(n_377), .Y(n_579) );
OAI221xp5_ASAP7_75t_SL g580 ( .A1(n_523), .A2(n_298), .B1(n_178), .B2(n_319), .C(n_347), .Y(n_580) );
AOI22xp33_ASAP7_75t_SL g581 ( .A1(n_465), .A2(n_275), .B1(n_296), .B2(n_313), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_521), .B(n_347), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_520), .A2(n_347), .B1(n_311), .B2(n_296), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_519), .A2(n_347), .B1(n_311), .B2(n_296), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_481), .B(n_155), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_521), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g587 ( .A1(n_509), .A2(n_312), .B1(n_327), .B2(n_332), .Y(n_587) );
AOI22xp33_ASAP7_75t_SL g588 ( .A1(n_478), .A2(n_275), .B1(n_296), .B2(n_295), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_511), .A2(n_311), .B1(n_296), .B2(n_317), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_524), .B(n_23), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_526), .A2(n_337), .B1(n_310), .B2(n_312), .Y(n_591) );
AOI22xp33_ASAP7_75t_SL g592 ( .A1(n_479), .A2(n_296), .B1(n_295), .B2(n_303), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_493), .A2(n_328), .B1(n_321), .B2(n_320), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_525), .A2(n_517), .B1(n_514), .B2(n_506), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_514), .A2(n_311), .B1(n_317), .B2(n_320), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_517), .A2(n_311), .B1(n_317), .B2(n_321), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_530), .A2(n_312), .B1(n_310), .B2(n_342), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_467), .A2(n_311), .B1(n_328), .B2(n_298), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_530), .A2(n_312), .B1(n_310), .B2(n_342), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_524), .B(n_460), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_496), .A2(n_311), .B1(n_328), .B2(n_298), .Y(n_601) );
NAND2xp5_ASAP7_75t_SL g602 ( .A(n_500), .B(n_155), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_500), .A2(n_512), .B1(n_461), .B2(n_491), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_518), .A2(n_311), .B1(n_155), .B2(n_165), .Y(n_604) );
OA21x2_ASAP7_75t_L g605 ( .A1(n_471), .A2(n_264), .B(n_178), .Y(n_605) );
OAI21xp33_ASAP7_75t_SL g606 ( .A1(n_531), .A2(n_306), .B(n_303), .Y(n_606) );
AOI22xp33_ASAP7_75t_SL g607 ( .A1(n_500), .A2(n_303), .B1(n_306), .B2(n_295), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_518), .A2(n_155), .B1(n_165), .B2(n_293), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_531), .B(n_23), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_518), .A2(n_155), .B1(n_165), .B2(n_293), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_471), .B(n_155), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_500), .A2(n_155), .B1(n_165), .B2(n_293), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_522), .A2(n_155), .B1(n_165), .B2(n_293), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_502), .A2(n_155), .B1(n_165), .B2(n_293), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_502), .A2(n_165), .B1(n_297), .B2(n_307), .Y(n_615) );
AOI21xp5_ASAP7_75t_SL g616 ( .A1(n_529), .A2(n_327), .B(n_342), .Y(n_616) );
AOI222xp33_ASAP7_75t_L g617 ( .A1(n_528), .A2(n_337), .B1(n_332), .B2(n_327), .C1(n_342), .C2(n_165), .Y(n_617) );
NAND3xp33_ASAP7_75t_SL g618 ( .A(n_528), .B(n_24), .C(n_25), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_502), .A2(n_165), .B1(n_297), .B2(n_307), .Y(n_619) );
AOI22xp33_ASAP7_75t_SL g620 ( .A1(n_477), .A2(n_295), .B1(n_306), .B2(n_303), .Y(n_620) );
NAND3xp33_ASAP7_75t_SL g621 ( .A(n_477), .B(n_26), .C(n_28), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_490), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_485), .A2(n_165), .B1(n_297), .B2(n_307), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_485), .A2(n_307), .B1(n_297), .B2(n_299), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_485), .A2(n_307), .B1(n_297), .B2(n_299), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_485), .A2(n_316), .B1(n_299), .B2(n_300), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_490), .A2(n_316), .B1(n_300), .B2(n_257), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_527), .A2(n_316), .B1(n_300), .B2(n_257), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_527), .A2(n_327), .B1(n_332), .B2(n_337), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_527), .A2(n_255), .B1(n_258), .B2(n_332), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_527), .A2(n_337), .B1(n_342), .B2(n_258), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_527), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_464), .A2(n_337), .B1(n_255), .B2(n_343), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_565), .B(n_173), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_565), .B(n_173), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_600), .B(n_173), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_600), .B(n_26), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_543), .B(n_28), .Y(n_638) );
NOR2xp33_ASAP7_75t_SL g639 ( .A(n_580), .B(n_322), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_543), .B(n_173), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_586), .B(n_173), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_586), .B(n_173), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_622), .B(n_173), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_622), .B(n_173), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_573), .A2(n_175), .B1(n_176), .B2(n_173), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_594), .B(n_173), .Y(n_646) );
NAND3xp33_ASAP7_75t_L g647 ( .A(n_558), .B(n_173), .C(n_175), .Y(n_647) );
NAND3xp33_ASAP7_75t_L g648 ( .A(n_617), .B(n_175), .C(n_176), .Y(n_648) );
NAND3xp33_ASAP7_75t_L g649 ( .A(n_617), .B(n_175), .C(n_176), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_570), .B(n_175), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_555), .B(n_29), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_537), .B(n_29), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_537), .B(n_30), .Y(n_653) );
AOI21xp5_ASAP7_75t_SL g654 ( .A1(n_562), .A2(n_306), .B(n_270), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_544), .B(n_175), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_533), .B(n_175), .Y(n_656) );
NAND3xp33_ASAP7_75t_L g657 ( .A(n_616), .B(n_175), .C(n_176), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_593), .A2(n_346), .B1(n_343), .B2(n_262), .Y(n_658) );
OAI221xp5_ASAP7_75t_L g659 ( .A1(n_593), .A2(n_175), .B1(n_176), .B2(n_329), .C(n_264), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_633), .A2(n_176), .B1(n_175), .B2(n_323), .Y(n_660) );
NAND2xp5_ASAP7_75t_SL g661 ( .A(n_561), .B(n_157), .Y(n_661) );
OAI21xp5_ASAP7_75t_L g662 ( .A1(n_618), .A2(n_157), .B(n_285), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_540), .B(n_30), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_536), .B(n_564), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_564), .B(n_31), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_633), .B(n_31), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_549), .B(n_157), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_632), .B(n_176), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_557), .A2(n_346), .B1(n_343), .B2(n_157), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_590), .B(n_32), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_532), .B(n_32), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_563), .B(n_176), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_577), .B(n_33), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_567), .B(n_176), .Y(n_674) );
AOI221xp5_ASAP7_75t_L g675 ( .A1(n_534), .A2(n_176), .B1(n_157), .B2(n_261), .C(n_329), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_603), .B(n_33), .Y(n_676) );
AND2x2_ASAP7_75t_SL g677 ( .A(n_535), .B(n_270), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_557), .B(n_34), .Y(n_678) );
NAND3xp33_ASAP7_75t_L g679 ( .A(n_616), .B(n_176), .C(n_157), .Y(n_679) );
OAI221xp5_ASAP7_75t_SL g680 ( .A1(n_606), .A2(n_330), .B1(n_331), .B2(n_36), .C(n_37), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_621), .A2(n_157), .B1(n_329), .B2(n_330), .C(n_331), .Y(n_681) );
AOI221xp5_ASAP7_75t_L g682 ( .A1(n_546), .A2(n_157), .B1(n_330), .B2(n_331), .C(n_37), .Y(n_682) );
NAND4xp25_ASAP7_75t_L g683 ( .A(n_547), .B(n_252), .C(n_35), .D(n_36), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_577), .B(n_34), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_609), .B(n_35), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g686 ( .A1(n_546), .A2(n_157), .B1(n_39), .B2(n_40), .C(n_41), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_588), .A2(n_346), .B1(n_157), .B2(n_336), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_572), .B(n_38), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_556), .B(n_40), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_576), .B(n_41), .Y(n_690) );
OAI21xp5_ASAP7_75t_SL g691 ( .A1(n_581), .A2(n_42), .B(n_279), .Y(n_691) );
NAND2xp33_ASAP7_75t_SL g692 ( .A(n_569), .B(n_42), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_576), .B(n_582), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_566), .B(n_157), .Y(n_694) );
NAND3xp33_ASAP7_75t_L g695 ( .A(n_541), .B(n_157), .C(n_279), .Y(n_695) );
OAI21xp5_ASAP7_75t_L g696 ( .A1(n_606), .A2(n_272), .B(n_338), .Y(n_696) );
NAND4xp25_ASAP7_75t_L g697 ( .A(n_601), .B(n_272), .C(n_284), .D(n_281), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_611), .B(n_47), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_607), .A2(n_344), .B1(n_336), .B2(n_323), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_611), .B(n_48), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_579), .B(n_49), .Y(n_701) );
OAI21xp33_ASAP7_75t_L g702 ( .A1(n_545), .A2(n_344), .B(n_336), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_553), .A2(n_344), .B1(n_336), .B2(n_323), .Y(n_703) );
NOR2xp33_ASAP7_75t_SL g704 ( .A(n_553), .B(n_344), .Y(n_704) );
NAND3xp33_ASAP7_75t_L g705 ( .A(n_574), .B(n_344), .C(n_336), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_598), .A2(n_338), .B1(n_335), .B2(n_323), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_597), .B(n_51), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_578), .B(n_53), .Y(n_708) );
AOI221xp5_ASAP7_75t_L g709 ( .A1(n_539), .A2(n_281), .B1(n_284), .B2(n_286), .C(n_292), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_599), .B(n_54), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_595), .B(n_55), .Y(n_711) );
OR2x6_ASAP7_75t_L g712 ( .A(n_585), .B(n_323), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_592), .A2(n_322), .B1(n_338), .B2(n_335), .Y(n_713) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_631), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_620), .A2(n_322), .B1(n_338), .B2(n_335), .Y(n_715) );
NOR2xp33_ASAP7_75t_R g716 ( .A(n_624), .B(n_56), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_596), .B(n_59), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_559), .B(n_60), .Y(n_718) );
OAI221xp5_ASAP7_75t_SL g719 ( .A1(n_551), .A2(n_322), .B1(n_335), .B2(n_338), .C(n_292), .Y(n_719) );
OAI221xp5_ASAP7_75t_SL g720 ( .A1(n_538), .A2(n_322), .B1(n_335), .B2(n_338), .C(n_286), .Y(n_720) );
AOI211xp5_ASAP7_75t_L g721 ( .A1(n_560), .A2(n_338), .B(n_335), .C(n_68), .Y(n_721) );
NAND2x1_ASAP7_75t_L g722 ( .A(n_605), .B(n_335), .Y(n_722) );
AOI21xp33_ASAP7_75t_L g723 ( .A1(n_568), .A2(n_65), .B(n_66), .Y(n_723) );
AOI221xp5_ASAP7_75t_L g724 ( .A1(n_542), .A2(n_256), .B1(n_236), .B2(n_217), .C(n_211), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_575), .B(n_73), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_631), .B(n_74), .Y(n_726) );
OAI221xp5_ASAP7_75t_SL g727 ( .A1(n_589), .A2(n_75), .B1(n_77), .B2(n_78), .C(n_80), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_583), .B(n_81), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_602), .B(n_85), .Y(n_729) );
OAI21xp33_ASAP7_75t_L g730 ( .A1(n_571), .A2(n_236), .B(n_256), .Y(n_730) );
OAI221xp5_ASAP7_75t_SL g731 ( .A1(n_550), .A2(n_87), .B1(n_88), .B2(n_89), .C(n_90), .Y(n_731) );
AND2x2_ASAP7_75t_L g732 ( .A(n_625), .B(n_92), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_629), .B(n_96), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_627), .B(n_97), .Y(n_734) );
NOR3xp33_ASAP7_75t_L g735 ( .A(n_552), .B(n_256), .C(n_236), .Y(n_735) );
AND2x4_ASAP7_75t_L g736 ( .A(n_636), .B(n_623), .Y(n_736) );
NAND3xp33_ASAP7_75t_L g737 ( .A(n_692), .B(n_604), .C(n_548), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_635), .B(n_614), .Y(n_738) );
NAND3xp33_ASAP7_75t_L g739 ( .A(n_692), .B(n_612), .C(n_610), .Y(n_739) );
NOR3xp33_ASAP7_75t_L g740 ( .A(n_663), .B(n_554), .C(n_591), .Y(n_740) );
OR2x2_ASAP7_75t_L g741 ( .A(n_635), .B(n_587), .Y(n_741) );
NAND3xp33_ASAP7_75t_L g742 ( .A(n_704), .B(n_608), .C(n_619), .Y(n_742) );
AOI221xp5_ASAP7_75t_L g743 ( .A1(n_651), .A2(n_584), .B1(n_626), .B2(n_613), .C(n_615), .Y(n_743) );
AO21x2_ASAP7_75t_L g744 ( .A1(n_655), .A2(n_628), .B(n_630), .Y(n_744) );
NAND4xp25_ASAP7_75t_L g745 ( .A(n_678), .B(n_98), .C(n_100), .D(n_101), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_650), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_655), .B(n_103), .Y(n_747) );
NAND3xp33_ASAP7_75t_L g748 ( .A(n_686), .B(n_243), .C(n_105), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_672), .B(n_104), .Y(n_749) );
NOR3xp33_ASAP7_75t_L g750 ( .A(n_683), .B(n_106), .C(n_107), .Y(n_750) );
OAI211xp5_ASAP7_75t_SL g751 ( .A1(n_691), .A2(n_108), .B(n_205), .C(n_243), .Y(n_751) );
INVx3_ASAP7_75t_L g752 ( .A(n_722), .Y(n_752) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_677), .A2(n_243), .B1(n_639), .B2(n_676), .Y(n_753) );
NOR3xp33_ASAP7_75t_SL g754 ( .A(n_680), .B(n_243), .C(n_662), .Y(n_754) );
NAND3xp33_ASAP7_75t_L g755 ( .A(n_718), .B(n_243), .C(n_665), .Y(n_755) );
NAND3xp33_ASAP7_75t_L g756 ( .A(n_657), .B(n_243), .C(n_721), .Y(n_756) );
NOR2x1_ASAP7_75t_L g757 ( .A(n_661), .B(n_667), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_640), .Y(n_758) );
NAND3xp33_ASAP7_75t_L g759 ( .A(n_646), .B(n_637), .C(n_714), .Y(n_759) );
INVx1_ASAP7_75t_SL g760 ( .A(n_700), .Y(n_760) );
OAI211xp5_ASAP7_75t_L g761 ( .A1(n_716), .A2(n_654), .B(n_697), .C(n_661), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g762 ( .A1(n_677), .A2(n_693), .B1(n_689), .B2(n_653), .Y(n_762) );
AO21x2_ASAP7_75t_L g763 ( .A1(n_638), .A2(n_668), .B(n_641), .Y(n_763) );
AND2x2_ASAP7_75t_L g764 ( .A(n_672), .B(n_674), .Y(n_764) );
NAND2xp5_ASAP7_75t_SL g765 ( .A(n_716), .B(n_667), .Y(n_765) );
NAND2xp5_ASAP7_75t_SL g766 ( .A(n_694), .B(n_679), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_652), .B(n_671), .Y(n_767) );
NAND3xp33_ASAP7_75t_L g768 ( .A(n_646), .B(n_670), .C(n_703), .Y(n_768) );
OR2x2_ASAP7_75t_L g769 ( .A(n_674), .B(n_688), .Y(n_769) );
NOR3xp33_ASAP7_75t_SL g770 ( .A(n_648), .B(n_649), .C(n_673), .Y(n_770) );
NAND3xp33_ASAP7_75t_L g771 ( .A(n_685), .B(n_681), .C(n_682), .Y(n_771) );
NAND3xp33_ASAP7_75t_L g772 ( .A(n_675), .B(n_656), .C(n_694), .Y(n_772) );
NOR3xp33_ASAP7_75t_SL g773 ( .A(n_684), .B(n_727), .C(n_666), .Y(n_773) );
NOR3xp33_ASAP7_75t_L g774 ( .A(n_690), .B(n_658), .C(n_731), .Y(n_774) );
OR2x2_ASAP7_75t_L g775 ( .A(n_642), .B(n_643), .Y(n_775) );
OR2x2_ASAP7_75t_L g776 ( .A(n_644), .B(n_712), .Y(n_776) );
NOR2xp33_ASAP7_75t_L g777 ( .A(n_669), .B(n_656), .Y(n_777) );
OR2x2_ASAP7_75t_L g778 ( .A(n_712), .B(n_700), .Y(n_778) );
NAND3xp33_ASAP7_75t_L g779 ( .A(n_645), .B(n_647), .C(n_695), .Y(n_779) );
NAND3xp33_ASAP7_75t_L g780 ( .A(n_705), .B(n_659), .C(n_660), .Y(n_780) );
AND2x4_ASAP7_75t_SL g781 ( .A(n_712), .B(n_699), .Y(n_781) );
XNOR2xp5_ASAP7_75t_L g782 ( .A(n_706), .B(n_715), .Y(n_782) );
AOI221x1_ASAP7_75t_SL g783 ( .A1(n_687), .A2(n_702), .B1(n_713), .B2(n_728), .C(n_726), .Y(n_783) );
NOR3xp33_ASAP7_75t_L g784 ( .A(n_711), .B(n_717), .C(n_701), .Y(n_784) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_712), .Y(n_785) );
AND2x4_ASAP7_75t_L g786 ( .A(n_708), .B(n_729), .Y(n_786) );
AND2x4_ASAP7_75t_L g787 ( .A(n_698), .B(n_725), .Y(n_787) );
NAND4xp75_ASAP7_75t_L g788 ( .A(n_725), .B(n_732), .C(n_707), .D(n_710), .Y(n_788) );
OAI211xp5_ASAP7_75t_L g789 ( .A1(n_720), .A2(n_719), .B(n_723), .C(n_696), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g790 ( .A(n_734), .B(n_733), .Y(n_790) );
AND2x2_ASAP7_75t_L g791 ( .A(n_735), .B(n_730), .Y(n_791) );
NAND3xp33_ASAP7_75t_L g792 ( .A(n_709), .B(n_692), .C(n_663), .Y(n_792) );
AND2x2_ASAP7_75t_L g793 ( .A(n_724), .B(n_634), .Y(n_793) );
BUFx3_ASAP7_75t_L g794 ( .A(n_636), .Y(n_794) );
NAND3xp33_ASAP7_75t_L g795 ( .A(n_692), .B(n_663), .C(n_704), .Y(n_795) );
BUFx2_ASAP7_75t_L g796 ( .A(n_636), .Y(n_796) );
NOR2xp33_ASAP7_75t_L g797 ( .A(n_663), .B(n_651), .Y(n_797) );
AND2x4_ASAP7_75t_L g798 ( .A(n_664), .B(n_564), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_677), .A2(n_573), .B1(n_692), .B2(n_540), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_664), .Y(n_800) );
AO21x2_ASAP7_75t_L g801 ( .A1(n_636), .A2(n_635), .B(n_634), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_664), .Y(n_802) );
NAND3xp33_ASAP7_75t_L g803 ( .A(n_692), .B(n_663), .C(n_704), .Y(n_803) );
OA211x2_ASAP7_75t_L g804 ( .A1(n_704), .A2(n_661), .B(n_667), .C(n_694), .Y(n_804) );
BUFx2_ASAP7_75t_L g805 ( .A(n_636), .Y(n_805) );
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_761), .A2(n_799), .B1(n_801), .B2(n_774), .Y(n_806) );
AND2x2_ASAP7_75t_L g807 ( .A(n_800), .B(n_802), .Y(n_807) );
NAND4xp75_ASAP7_75t_SL g808 ( .A(n_791), .B(n_777), .C(n_767), .D(n_790), .Y(n_808) );
INVx2_ASAP7_75t_SL g809 ( .A(n_798), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_801), .Y(n_810) );
AND2x2_ASAP7_75t_L g811 ( .A(n_798), .B(n_796), .Y(n_811) );
BUFx3_ASAP7_75t_L g812 ( .A(n_794), .Y(n_812) );
INVx2_ASAP7_75t_L g813 ( .A(n_805), .Y(n_813) );
XOR2xp5_ASAP7_75t_L g814 ( .A(n_782), .B(n_769), .Y(n_814) );
INVx1_ASAP7_75t_SL g815 ( .A(n_760), .Y(n_815) );
INVx4_ASAP7_75t_L g816 ( .A(n_752), .Y(n_816) );
HB1xp67_ASAP7_75t_L g817 ( .A(n_785), .Y(n_817) );
NAND4xp75_ASAP7_75t_SL g818 ( .A(n_777), .B(n_767), .C(n_790), .D(n_797), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_763), .B(n_746), .Y(n_819) );
NAND4xp75_ASAP7_75t_L g820 ( .A(n_804), .B(n_757), .C(n_765), .D(n_773), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_759), .B(n_758), .Y(n_821) );
INVx1_ASAP7_75t_SL g822 ( .A(n_778), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_764), .B(n_785), .Y(n_823) );
XOR2xp5_ASAP7_75t_L g824 ( .A(n_762), .B(n_788), .Y(n_824) );
INVx1_ASAP7_75t_SL g825 ( .A(n_781), .Y(n_825) );
NAND4xp75_ASAP7_75t_SL g826 ( .A(n_797), .B(n_783), .C(n_761), .D(n_793), .Y(n_826) );
HB1xp67_ASAP7_75t_L g827 ( .A(n_775), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g828 ( .A1(n_799), .A2(n_774), .B1(n_750), .B2(n_792), .Y(n_828) );
HB1xp67_ASAP7_75t_L g829 ( .A(n_752), .Y(n_829) );
INVx5_ASAP7_75t_L g830 ( .A(n_747), .Y(n_830) );
XNOR2xp5_ASAP7_75t_L g831 ( .A(n_753), .B(n_768), .Y(n_831) );
INVx2_ASAP7_75t_SL g832 ( .A(n_776), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g833 ( .A1(n_795), .A2(n_803), .B1(n_755), .B2(n_786), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_741), .Y(n_834) );
NAND2xp33_ASAP7_75t_R g835 ( .A(n_754), .B(n_773), .Y(n_835) );
INVx2_ASAP7_75t_L g836 ( .A(n_736), .Y(n_836) );
AND2x2_ASAP7_75t_SL g837 ( .A(n_750), .B(n_786), .Y(n_837) );
NAND4xp75_ASAP7_75t_L g838 ( .A(n_766), .B(n_770), .C(n_754), .D(n_743), .Y(n_838) );
AND2x2_ASAP7_75t_L g839 ( .A(n_736), .B(n_738), .Y(n_839) );
NAND4xp25_ASAP7_75t_L g840 ( .A(n_771), .B(n_740), .C(n_737), .D(n_772), .Y(n_840) );
AND2x2_ASAP7_75t_L g841 ( .A(n_787), .B(n_744), .Y(n_841) );
AND2x2_ASAP7_75t_L g842 ( .A(n_787), .B(n_744), .Y(n_842) );
NAND4xp75_ASAP7_75t_L g843 ( .A(n_770), .B(n_743), .C(n_749), .D(n_751), .Y(n_843) );
NAND4xp75_ASAP7_75t_SL g844 ( .A(n_751), .B(n_789), .C(n_745), .D(n_740), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_756), .Y(n_845) );
NOR4xp25_ASAP7_75t_L g846 ( .A(n_789), .B(n_739), .C(n_780), .D(n_779), .Y(n_846) );
XOR2x2_ASAP7_75t_L g847 ( .A(n_784), .B(n_748), .Y(n_847) );
CKINVDCx16_ASAP7_75t_R g848 ( .A(n_835), .Y(n_848) );
AOI22xp5_ASAP7_75t_L g849 ( .A1(n_806), .A2(n_742), .B1(n_784), .B2(n_828), .Y(n_849) );
XOR2x2_ASAP7_75t_L g850 ( .A(n_826), .B(n_818), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_836), .Y(n_851) );
INVx1_ASAP7_75t_SL g852 ( .A(n_812), .Y(n_852) );
INVx2_ASAP7_75t_L g853 ( .A(n_836), .Y(n_853) );
XNOR2xp5_ASAP7_75t_L g854 ( .A(n_814), .B(n_824), .Y(n_854) );
AND2x2_ASAP7_75t_L g855 ( .A(n_841), .B(n_842), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_810), .Y(n_856) );
INVx2_ASAP7_75t_L g857 ( .A(n_813), .Y(n_857) );
XNOR2xp5_ASAP7_75t_L g858 ( .A(n_814), .B(n_824), .Y(n_858) );
AND2x2_ASAP7_75t_L g859 ( .A(n_841), .B(n_842), .Y(n_859) );
INVx2_ASAP7_75t_SL g860 ( .A(n_812), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_807), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_810), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_807), .Y(n_863) );
XOR2x2_ASAP7_75t_L g864 ( .A(n_808), .B(n_820), .Y(n_864) );
INVx2_ASAP7_75t_L g865 ( .A(n_813), .Y(n_865) );
INVx2_ASAP7_75t_L g866 ( .A(n_811), .Y(n_866) );
INVxp67_ASAP7_75t_L g867 ( .A(n_820), .Y(n_867) );
XOR2x2_ASAP7_75t_L g868 ( .A(n_838), .B(n_828), .Y(n_868) );
INVx1_ASAP7_75t_SL g869 ( .A(n_825), .Y(n_869) );
AOI22xp5_ASAP7_75t_L g870 ( .A1(n_806), .A2(n_838), .B1(n_840), .B2(n_833), .Y(n_870) );
INVxp67_ASAP7_75t_L g871 ( .A(n_840), .Y(n_871) );
INVx1_ASAP7_75t_SL g872 ( .A(n_811), .Y(n_872) );
XNOR2xp5_ASAP7_75t_L g873 ( .A(n_846), .B(n_847), .Y(n_873) );
AOI22x1_ASAP7_75t_L g874 ( .A1(n_848), .A2(n_816), .B1(n_831), .B2(n_829), .Y(n_874) );
OA22x2_ASAP7_75t_L g875 ( .A1(n_870), .A2(n_831), .B1(n_816), .B2(n_809), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_863), .Y(n_876) );
AO22x2_ASAP7_75t_L g877 ( .A1(n_871), .A2(n_843), .B1(n_844), .B2(n_816), .Y(n_877) );
BUFx3_ASAP7_75t_L g878 ( .A(n_860), .Y(n_878) );
XOR2x2_ASAP7_75t_L g879 ( .A(n_854), .B(n_843), .Y(n_879) );
OA22x2_ASAP7_75t_L g880 ( .A1(n_873), .A2(n_809), .B1(n_817), .B2(n_845), .Y(n_880) );
OAI22x1_ASAP7_75t_L g881 ( .A1(n_873), .A2(n_815), .B1(n_845), .B2(n_830), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_863), .Y(n_882) );
INVx2_ASAP7_75t_L g883 ( .A(n_860), .Y(n_883) );
INVx1_ASAP7_75t_SL g884 ( .A(n_852), .Y(n_884) );
OAI22xp5_ASAP7_75t_SL g885 ( .A1(n_854), .A2(n_837), .B1(n_830), .B2(n_847), .Y(n_885) );
XNOR2x1_ASAP7_75t_L g886 ( .A(n_868), .B(n_839), .Y(n_886) );
OA22x2_ASAP7_75t_L g887 ( .A1(n_849), .A2(n_839), .B1(n_832), .B2(n_834), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_861), .Y(n_888) );
OA22x2_ASAP7_75t_L g889 ( .A1(n_858), .A2(n_832), .B1(n_834), .B2(n_822), .Y(n_889) );
AOI22xp5_ASAP7_75t_L g890 ( .A1(n_885), .A2(n_868), .B1(n_858), .B2(n_867), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_884), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_884), .Y(n_892) );
INVx2_ASAP7_75t_L g893 ( .A(n_878), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_883), .Y(n_894) );
INVx3_ASAP7_75t_L g895 ( .A(n_877), .Y(n_895) );
OA22x2_ASAP7_75t_L g896 ( .A1(n_885), .A2(n_869), .B1(n_859), .B2(n_855), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_888), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_876), .Y(n_898) );
AOI22xp5_ASAP7_75t_L g899 ( .A1(n_890), .A2(n_877), .B1(n_875), .B2(n_879), .Y(n_899) );
AOI221xp5_ASAP7_75t_L g900 ( .A1(n_895), .A2(n_881), .B1(n_859), .B2(n_855), .C(n_875), .Y(n_900) );
OAI322xp33_ASAP7_75t_L g901 ( .A1(n_896), .A2(n_880), .A3(n_889), .B1(n_887), .B2(n_886), .C1(n_874), .C2(n_872), .Y(n_901) );
AOI311xp33_ASAP7_75t_L g902 ( .A1(n_891), .A2(n_880), .A3(n_889), .B(n_850), .C(n_887), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_892), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_903), .Y(n_904) );
OAI22xp33_ASAP7_75t_L g905 ( .A1(n_899), .A2(n_896), .B1(n_893), .B2(n_895), .Y(n_905) );
OAI22xp5_ASAP7_75t_L g906 ( .A1(n_900), .A2(n_893), .B1(n_895), .B2(n_894), .Y(n_906) );
OAI22xp5_ASAP7_75t_L g907 ( .A1(n_905), .A2(n_897), .B1(n_898), .B2(n_902), .Y(n_907) );
AOI31xp33_ASAP7_75t_L g908 ( .A1(n_906), .A2(n_901), .A3(n_850), .B(n_864), .Y(n_908) );
AOI31xp33_ASAP7_75t_L g909 ( .A1(n_904), .A2(n_864), .A3(n_862), .B(n_856), .Y(n_909) );
INVxp67_ASAP7_75t_SL g910 ( .A(n_907), .Y(n_910) );
AO22x2_ASAP7_75t_L g911 ( .A1(n_908), .A2(n_882), .B1(n_856), .B2(n_862), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_911), .Y(n_912) );
HB1xp67_ASAP7_75t_L g913 ( .A(n_910), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_913), .Y(n_914) );
INVx2_ASAP7_75t_L g915 ( .A(n_912), .Y(n_915) );
AO22x2_ASAP7_75t_L g916 ( .A1(n_915), .A2(n_912), .B1(n_914), .B2(n_909), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_916), .Y(n_917) );
AOI31xp33_ASAP7_75t_L g918 ( .A1(n_917), .A2(n_915), .A3(n_821), .B(n_819), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_918), .Y(n_919) );
AO22x2_ASAP7_75t_L g920 ( .A1(n_919), .A2(n_866), .B1(n_865), .B2(n_857), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_920), .Y(n_921) );
AOI221xp5_ASAP7_75t_L g922 ( .A1(n_921), .A2(n_866), .B1(n_865), .B2(n_857), .C(n_851), .Y(n_922) );
AOI211xp5_ASAP7_75t_L g923 ( .A1(n_922), .A2(n_827), .B(n_823), .C(n_853), .Y(n_923) );
endmodule