module fake_jpeg_20878_n_313 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_25),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_8),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_30),
.B(n_8),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_44),
.B(n_15),
.Y(n_79)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_0),
.Y(n_46)
);

AOI21xp33_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_25),
.B(n_24),
.Y(n_69)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_20),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx4f_ASAP7_75t_SL g115 ( 
.A(n_50),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_46),
.A2(n_28),
.B1(n_35),
.B2(n_22),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_48),
.A2(n_28),
.B1(n_35),
.B2(n_36),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_55),
.A2(n_48),
.B1(n_45),
.B2(n_47),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_35),
.B1(n_28),
.B2(n_19),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_56),
.A2(n_71),
.B1(n_73),
.B2(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_32),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_57),
.B(n_13),
.Y(n_119)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_82),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_68),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_41),
.A2(n_28),
.B1(n_36),
.B2(n_19),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_65),
.B(n_69),
.Y(n_118)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_21),
.Y(n_68)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_42),
.A2(n_19),
.B1(n_23),
.B2(n_24),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_22),
.B1(n_32),
.B2(n_38),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_38),
.B1(n_23),
.B2(n_24),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_46),
.A2(n_23),
.B1(n_27),
.B2(n_34),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_77),
.A2(n_80),
.B1(n_20),
.B2(n_31),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_43),
.A2(n_27),
.B(n_34),
.C(n_21),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_78),
.B(n_79),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_47),
.A2(n_37),
.B1(n_31),
.B2(n_29),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_48),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_SL g84 ( 
.A(n_62),
.B(n_51),
.C(n_78),
.Y(n_84)
);

AND2x4_ASAP7_75t_L g138 ( 
.A(n_84),
.B(n_33),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_86),
.A2(n_61),
.B1(n_82),
.B2(n_53),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_44),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_96),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_43),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_50),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_99),
.B(n_101),
.Y(n_151)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_20),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_46),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_114),
.Y(n_120)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_61),
.A2(n_20),
.B1(n_21),
.B2(n_31),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_20),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_106),
.B(n_112),
.Y(n_129)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_111),
.A2(n_1),
.B1(n_2),
.B2(n_37),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_20),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_113),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_65),
.B(n_21),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_65),
.B(n_33),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_116),
.B(n_119),
.Y(n_136)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_118),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_127),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_80),
.B(n_70),
.C(n_66),
.Y(n_126)
);

O2A1O1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_126),
.A2(n_151),
.B(n_150),
.C(n_130),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_52),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_53),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_130),
.B(n_141),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_92),
.A2(n_67),
.B1(n_58),
.B2(n_63),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_131),
.A2(n_126),
.B1(n_151),
.B2(n_138),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_133),
.A2(n_139),
.B(n_149),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_134),
.A2(n_137),
.B1(n_107),
.B2(n_108),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_37),
.B1(n_31),
.B2(n_29),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_138),
.B(n_2),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_98),
.A2(n_33),
.B(n_29),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_98),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_84),
.A2(n_37),
.B1(n_29),
.B2(n_26),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_144),
.A2(n_153),
.B1(n_117),
.B2(n_103),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_92),
.B(n_26),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_146),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_83),
.B(n_26),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_26),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_97),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_150),
.B(n_152),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_83),
.B(n_90),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_100),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_155),
.A2(n_158),
.B1(n_170),
.B2(n_171),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_157),
.A2(n_159),
.B1(n_164),
.B2(n_185),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_85),
.B1(n_108),
.B2(n_87),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_145),
.A2(n_87),
.B1(n_93),
.B2(n_91),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_91),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_123),
.Y(n_162)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_109),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_163),
.Y(n_202)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_121),
.B(n_109),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_168),
.B(n_169),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_88),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_85),
.B1(n_89),
.B2(n_110),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_149),
.A2(n_89),
.B1(n_88),
.B2(n_113),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_124),
.Y(n_172)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_124),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_173),
.B(n_174),
.Y(n_214)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

MAJx2_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_11),
.C(n_16),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_175),
.A2(n_146),
.B(n_138),
.Y(n_189)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_176),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_147),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_177),
.B(n_178),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_135),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_120),
.B(n_99),
.C(n_115),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_144),
.Y(n_200)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_181),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_182),
.A2(n_134),
.B1(n_122),
.B2(n_143),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_126),
.A2(n_10),
.B1(n_17),
.B2(n_3),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_184),
.A2(n_155),
.B1(n_122),
.B2(n_183),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_120),
.A2(n_115),
.B1(n_105),
.B2(n_1),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_186),
.A2(n_139),
.B(n_137),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_SL g236 ( 
.A(n_189),
.B(n_197),
.C(n_199),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_165),
.A2(n_138),
.B1(n_132),
.B2(n_133),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_190),
.A2(n_195),
.B(n_175),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

BUFx24_ASAP7_75t_SL g194 ( 
.A(n_166),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_205),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_136),
.B(n_152),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_L g197 ( 
.A1(n_180),
.A2(n_136),
.B(n_127),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_167),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_142),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_135),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_172),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_173),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_208),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_207),
.A2(n_157),
.B1(n_159),
.B2(n_185),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_174),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_212),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_179),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_140),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_213),
.A2(n_176),
.B(n_180),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_168),
.C(n_156),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_235),
.C(n_189),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_165),
.B1(n_158),
.B2(n_170),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_217),
.A2(n_223),
.B1(n_237),
.B2(n_188),
.Y(n_244)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_218),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_220),
.A2(n_233),
.B1(n_198),
.B2(n_191),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_156),
.Y(n_221)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_192),
.A2(n_184),
.B1(n_183),
.B2(n_169),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_209),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_225),
.B(n_227),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_234),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_186),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_228),
.B(n_229),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_195),
.B(n_186),
.Y(n_229)
);

NAND5xp2_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_142),
.C(n_153),
.D(n_154),
.E(n_140),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_230),
.A2(n_213),
.B(n_208),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_231),
.B(n_232),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_154),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_143),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_201),
.B(n_125),
.C(n_148),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_188),
.A2(n_148),
.B1(n_5),
.B2(n_6),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_239),
.A2(n_244),
.B1(n_246),
.B2(n_249),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_230),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_234),
.C(n_229),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_217),
.A2(n_213),
.B1(n_187),
.B2(n_206),
.Y(n_246)
);

A2O1A1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_216),
.A2(n_202),
.B(n_203),
.C(n_190),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_253),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_223),
.A2(n_205),
.B1(n_204),
.B2(n_196),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_210),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_236),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_204),
.C(n_196),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_221),
.C(n_219),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_226),
.A2(n_210),
.B(n_193),
.Y(n_253)
);

OAI21xp33_ASAP7_75t_L g254 ( 
.A1(n_225),
.A2(n_193),
.B(n_198),
.Y(n_254)
);

NAND3xp33_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_228),
.C(n_227),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_255),
.A2(n_237),
.B1(n_224),
.B2(n_233),
.Y(n_257)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_256),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_257),
.A2(n_244),
.B1(n_247),
.B2(n_252),
.Y(n_275)
);

OAI21xp33_ASAP7_75t_R g259 ( 
.A1(n_240),
.A2(n_236),
.B(n_218),
.Y(n_259)
);

AO22x1_ASAP7_75t_L g273 ( 
.A1(n_259),
.A2(n_262),
.B1(n_248),
.B2(n_253),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_260),
.B(n_265),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_235),
.C(n_216),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_266),
.C(n_272),
.Y(n_276)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_238),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_271),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_243),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_269),
.A2(n_238),
.B1(n_191),
.B2(n_6),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_222),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_270),
.B(n_263),
.Y(n_281)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_247),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_281),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_269),
.B1(n_259),
.B2(n_258),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_274),
.A2(n_283),
.B1(n_17),
.B2(n_8),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_275),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_284),
.Y(n_288)
);

NOR2x1_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_268),
.Y(n_280)
);

MAJx2_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_4),
.C(n_5),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_261),
.A2(n_219),
.B(n_251),
.Y(n_283)
);

OAI221xp5_ASAP7_75t_L g285 ( 
.A1(n_284),
.A2(n_260),
.B1(n_272),
.B2(n_258),
.C(n_10),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_287),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_278),
.A2(n_276),
.B1(n_283),
.B2(n_280),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_291),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_4),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_293),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_4),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_274),
.C(n_279),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_298),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_282),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_282),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_300),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_277),
.Y(n_300)
);

AO21x1_ASAP7_75t_L g301 ( 
.A1(n_296),
.A2(n_294),
.B(n_287),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_301),
.A2(n_304),
.B(n_305),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_297),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_288),
.C(n_275),
.Y(n_305)
);

OA21x2_ASAP7_75t_SL g306 ( 
.A1(n_303),
.A2(n_273),
.B(n_11),
.Y(n_306)
);

NOR2xp67_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_15),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_302),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_307),
.B(n_308),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_309),
.B(n_310),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_15),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_17),
.Y(n_313)
);


endmodule