module fake_jpeg_9332_n_50 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

AOI21xp33_ASAP7_75t_L g7 ( 
.A1(n_0),
.A2(n_1),
.B(n_5),
.Y(n_7)
);

INVx5_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_8),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_15),
.B(n_19),
.Y(n_22)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_20),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_17),
.Y(n_25)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_4),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_10),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_27),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_18),
.B1(n_16),
.B2(n_10),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_25),
.C(n_12),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_15),
.B1(n_20),
.B2(n_17),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_31),
.B(n_13),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_23),
.B(n_19),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_32),
.B(n_26),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_36),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_14),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_35),
.Y(n_38)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_R g39 ( 
.A(n_37),
.B(n_7),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_11),
.B1(n_30),
.B2(n_24),
.Y(n_42)
);

A2O1A1O1Ixp25_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_28),
.B(n_25),
.C(n_24),
.D(n_17),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_41),
.B(n_9),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_11),
.C(n_13),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_43),
.B(n_44),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_38),
.B1(n_40),
.B2(n_30),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_44),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_45),
.C(n_13),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_6),
.Y(n_50)
);


endmodule