module real_aes_8077_n_286 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_286);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_286;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_905;
wire n_503;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_792;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_919;
wire n_461;
wire n_908;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_289;
wire n_462;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_356;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_892;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_468;
wire n_755;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_298;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_671;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_642;
wire n_869;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_756;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_915;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_926;
wire n_922;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_314;
wire n_753;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_0), .A2(n_161), .B1(n_544), .B2(n_790), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_1), .A2(n_75), .B1(n_368), .B2(n_567), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_2), .A2(n_51), .B1(n_330), .B2(n_335), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g577 ( .A(n_3), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_4), .Y(n_749) );
AOI22xp33_ASAP7_75t_SL g762 ( .A1(n_5), .A2(n_279), .B1(n_669), .B2(n_670), .Y(n_762) );
AOI22xp33_ASAP7_75t_SL g607 ( .A1(n_6), .A2(n_106), .B1(n_458), .B2(n_512), .Y(n_607) );
AOI22xp33_ASAP7_75t_SL g509 ( .A1(n_7), .A2(n_32), .B1(n_510), .B2(n_512), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g839 ( .A1(n_8), .A2(n_128), .B1(n_330), .B2(n_642), .Y(n_839) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_9), .Y(n_797) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_10), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_11), .A2(n_43), .B1(n_564), .B2(n_566), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g387 ( .A1(n_12), .A2(n_388), .B1(n_437), .B2(n_438), .Y(n_387) );
INVx1_ASAP7_75t_L g437 ( .A(n_12), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_13), .A2(n_222), .B1(n_544), .B2(n_546), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_14), .Y(n_736) );
INVx1_ASAP7_75t_L g742 ( .A(n_15), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g613 ( .A(n_16), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_17), .A2(n_236), .B1(n_368), .B2(n_371), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_18), .A2(n_100), .B1(n_425), .B2(n_727), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_19), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_20), .A2(n_34), .B1(n_335), .B2(n_700), .Y(n_882) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_21), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_22), .A2(n_147), .B1(n_471), .B2(n_474), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_23), .A2(n_133), .B1(n_380), .B2(n_494), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_24), .A2(n_130), .B1(n_570), .B2(n_640), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_25), .A2(n_276), .B1(n_352), .B2(n_357), .Y(n_351) );
AO22x2_ASAP7_75t_L g322 ( .A1(n_26), .A2(n_93), .B1(n_313), .B2(n_318), .Y(n_322) );
INVx1_ASAP7_75t_L g862 ( .A(n_26), .Y(n_862) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_27), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_28), .A2(n_251), .B1(n_330), .B2(n_335), .Y(n_329) );
AOI211xp5_ASAP7_75t_L g286 ( .A1(n_29), .A2(n_287), .B(n_295), .C(n_864), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_30), .A2(n_66), .B1(n_561), .B2(n_562), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_31), .A2(n_181), .B1(n_422), .B2(n_564), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g838 ( .A1(n_33), .A2(n_269), .B1(n_512), .B2(n_551), .Y(n_838) );
AOI22xp33_ASAP7_75t_SL g610 ( .A1(n_35), .A2(n_47), .B1(n_309), .B2(n_453), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_36), .A2(n_136), .B1(n_564), .B2(n_672), .Y(n_671) );
AOI22xp33_ASAP7_75t_SL g504 ( .A1(n_37), .A2(n_203), .B1(n_323), .B2(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g341 ( .A(n_38), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_39), .B(n_738), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g909 ( .A(n_40), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_41), .A2(n_164), .B1(n_331), .B2(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g731 ( .A(n_42), .Y(n_731) );
AO22x2_ASAP7_75t_L g320 ( .A1(n_44), .A2(n_95), .B1(n_313), .B2(n_314), .Y(n_320) );
INVx1_ASAP7_75t_L g863 ( .A(n_44), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_45), .A2(n_211), .B1(n_432), .B2(n_435), .Y(n_431) );
AOI22xp33_ASAP7_75t_SL g506 ( .A1(n_46), .A2(n_104), .B1(n_330), .B2(n_507), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_48), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_49), .Y(n_469) );
INVx1_ASAP7_75t_L g575 ( .A(n_50), .Y(n_575) );
AOI22xp33_ASAP7_75t_SL g636 ( .A1(n_52), .A2(n_205), .B1(n_365), .B2(n_368), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g842 ( .A(n_53), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_54), .B(n_346), .Y(n_345) );
CKINVDCx20_ASAP7_75t_R g891 ( .A(n_55), .Y(n_891) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_56), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g836 ( .A1(n_57), .A2(n_218), .B1(n_672), .B2(n_728), .Y(n_836) );
AOI22xp5_ASAP7_75t_L g759 ( .A1(n_58), .A2(n_92), .B1(n_364), .B2(n_365), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g869 ( .A(n_59), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_60), .A2(n_112), .B1(n_423), .B2(n_436), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_61), .A2(n_240), .B1(n_383), .B2(n_407), .Y(n_655) );
AOI22xp33_ASAP7_75t_SL g668 ( .A1(n_62), .A2(n_243), .B1(n_669), .B2(n_670), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_63), .A2(n_173), .B1(n_561), .B2(n_725), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_64), .A2(n_175), .B1(n_357), .B2(n_473), .Y(n_604) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_65), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_67), .A2(n_80), .B1(n_786), .B2(n_788), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_68), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_69), .A2(n_90), .B1(n_407), .B2(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_70), .B(n_738), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g875 ( .A(n_71), .Y(n_875) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_72), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g846 ( .A1(n_73), .A2(n_137), .B1(n_380), .B2(n_404), .Y(n_846) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_74), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g916 ( .A(n_76), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_77), .A2(n_234), .B1(n_570), .B2(n_571), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_78), .A2(n_129), .B1(n_364), .B2(n_422), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_79), .A2(n_193), .B1(n_790), .B2(n_881), .Y(n_914) );
CKINVDCx20_ASAP7_75t_R g845 ( .A(n_81), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_82), .A2(n_197), .B1(n_371), .B2(n_510), .Y(n_722) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_83), .A2(n_105), .B1(n_425), .B2(n_452), .Y(n_572) );
AOI222xp33_ASAP7_75t_L g374 ( .A1(n_84), .A2(n_160), .B1(n_170), .B2(n_375), .C1(n_379), .C2(n_383), .Y(n_374) );
CKINVDCx20_ASAP7_75t_R g886 ( .A(n_85), .Y(n_886) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_86), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g903 ( .A(n_87), .Y(n_903) );
AOI211xp5_ASAP7_75t_L g901 ( .A1(n_88), .A2(n_624), .B(n_902), .C(n_906), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_89), .A2(n_199), .B1(n_368), .B2(n_642), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_91), .A2(n_151), .B1(n_358), .B2(n_482), .Y(n_843) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_94), .Y(n_536) );
AOI22xp33_ASAP7_75t_SL g501 ( .A1(n_96), .A2(n_265), .B1(n_473), .B2(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_97), .B(n_774), .Y(n_773) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_98), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_99), .A2(n_172), .B1(n_699), .B2(n_700), .Y(n_698) );
INVx1_ASAP7_75t_L g294 ( .A(n_101), .Y(n_294) );
INVx1_ASAP7_75t_L g414 ( .A(n_102), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_103), .A2(n_202), .B1(n_452), .B2(n_454), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_107), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_108), .A2(n_208), .B1(n_642), .B2(n_913), .Y(n_912) );
INVx1_ASAP7_75t_L g290 ( .A(n_109), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_110), .A2(n_174), .B1(n_362), .B2(n_365), .Y(n_361) );
INVx1_ASAP7_75t_L g409 ( .A(n_111), .Y(n_409) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_113), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_114), .A2(n_198), .B1(n_449), .B2(n_450), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_115), .A2(n_253), .B1(n_484), .B2(n_485), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_116), .A2(n_278), .B1(n_381), .B2(n_494), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_117), .Y(n_813) );
AOI22xp5_ASAP7_75t_L g834 ( .A1(n_118), .A2(n_246), .B1(n_640), .B2(n_835), .Y(n_834) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_119), .Y(n_817) );
AOI22xp33_ASAP7_75t_SL g633 ( .A1(n_120), .A2(n_124), .B1(n_357), .B2(n_494), .Y(n_633) );
OA22x2_ASAP7_75t_L g618 ( .A1(n_121), .A2(n_619), .B1(n_620), .B2(n_643), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_121), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_122), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_123), .A2(n_239), .B1(n_702), .B2(n_705), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_125), .B(n_659), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_126), .A2(n_231), .B1(n_371), .B2(n_570), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_127), .B(n_500), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_131), .A2(n_132), .B1(n_307), .B2(n_323), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_134), .A2(n_214), .B1(n_480), .B2(n_776), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_135), .A2(n_138), .B1(n_428), .B2(n_429), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_139), .B(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_140), .B(n_602), .Y(n_601) );
CKINVDCx20_ASAP7_75t_R g841 ( .A(n_141), .Y(n_841) );
XNOR2x2_ASAP7_75t_L g444 ( .A(n_142), .B(n_445), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_143), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_144), .B(n_484), .Y(n_904) );
AND2x2_ASAP7_75t_L g293 ( .A(n_145), .B(n_294), .Y(n_293) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_146), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_148), .B(n_474), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_149), .A2(n_718), .B1(n_743), .B2(n_744), .Y(n_717) );
INVx1_ASAP7_75t_L g743 ( .A(n_149), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_150), .B(n_630), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_152), .A2(n_219), .B1(n_452), .B2(n_696), .Y(n_695) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_153), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g920 ( .A(n_154), .Y(n_920) );
CKINVDCx20_ASAP7_75t_R g907 ( .A(n_155), .Y(n_907) );
CKINVDCx20_ASAP7_75t_R g582 ( .A(n_156), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_157), .Y(n_778) );
AND2x6_ASAP7_75t_L g289 ( .A(n_158), .B(n_290), .Y(n_289) );
HB1xp67_ASAP7_75t_L g856 ( .A(n_158), .Y(n_856) );
AO22x2_ASAP7_75t_L g312 ( .A1(n_159), .A2(n_235), .B1(n_313), .B2(n_314), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_162), .A2(n_194), .B1(n_432), .B2(n_549), .Y(n_548) );
CKINVDCx16_ASAP7_75t_R g899 ( .A(n_163), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_165), .A2(n_188), .B1(n_561), .B2(n_725), .Y(n_724) );
AOI22xp33_ASAP7_75t_SL g477 ( .A1(n_166), .A2(n_247), .B1(n_478), .B2(n_480), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_167), .B(n_485), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g580 ( .A(n_168), .Y(n_580) );
CKINVDCx20_ASAP7_75t_R g652 ( .A(n_169), .Y(n_652) );
INVx1_ASAP7_75t_L g552 ( .A(n_171), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_176), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_177), .Y(n_456) );
AOI22xp33_ASAP7_75t_SL g641 ( .A1(n_178), .A2(n_266), .B1(n_331), .B2(n_642), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_179), .A2(n_190), .B1(n_358), .B2(n_627), .Y(n_660) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_180), .Y(n_808) );
AOI22xp33_ASAP7_75t_SL g639 ( .A1(n_182), .A2(n_259), .B1(n_428), .B2(n_640), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g880 ( .A1(n_183), .A2(n_215), .B1(n_309), .B2(n_881), .Y(n_880) );
CKINVDCx20_ASAP7_75t_R g587 ( .A(n_184), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_185), .A2(n_285), .B1(n_664), .B2(n_665), .Y(n_663) );
INVx1_ASAP7_75t_L g680 ( .A(n_186), .Y(n_680) );
AO22x2_ASAP7_75t_L g317 ( .A1(n_187), .A2(n_255), .B1(n_313), .B2(n_318), .Y(n_317) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_189), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_191), .A2(n_224), .B1(n_480), .B2(n_776), .Y(n_775) );
AOI22xp5_ASAP7_75t_L g865 ( .A1(n_192), .A2(n_866), .B1(n_892), .B2(n_893), .Y(n_865) );
CKINVDCx20_ASAP7_75t_R g892 ( .A(n_192), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_195), .A2(n_281), .B1(n_432), .B2(n_825), .Y(n_824) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_196), .A2(n_557), .B1(n_591), .B2(n_592), .Y(n_556) );
INVx1_ASAP7_75t_L g591 ( .A(n_196), .Y(n_591) );
AOI22xp5_ASAP7_75t_SL g674 ( .A1(n_200), .A2(n_675), .B1(n_707), .B2(n_708), .Y(n_674) );
INVx1_ASAP7_75t_L g708 ( .A(n_200), .Y(n_708) );
INVx1_ASAP7_75t_L g922 ( .A(n_201), .Y(n_922) );
AOI22xp5_ASAP7_75t_L g804 ( .A1(n_204), .A2(n_805), .B1(n_827), .B2(n_828), .Y(n_804) );
INVx1_ASAP7_75t_L g827 ( .A(n_204), .Y(n_827) );
AOI22xp33_ASAP7_75t_SL g637 ( .A1(n_206), .A2(n_237), .B1(n_453), .B2(n_612), .Y(n_637) );
CKINVDCx20_ASAP7_75t_R g872 ( .A(n_207), .Y(n_872) );
AOI22xp33_ASAP7_75t_SL g513 ( .A1(n_209), .A2(n_248), .B1(n_450), .B2(n_514), .Y(n_513) );
AOI22xp33_ASAP7_75t_SL g626 ( .A1(n_210), .A2(n_258), .B1(n_380), .B2(n_627), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_212), .A2(n_233), .B1(n_380), .B2(n_494), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g395 ( .A(n_213), .Y(n_395) );
INVx1_ASAP7_75t_L g687 ( .A(n_216), .Y(n_687) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_217), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_220), .Y(n_771) );
CKINVDCx20_ASAP7_75t_R g870 ( .A(n_221), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_223), .A2(n_245), .B1(n_323), .B2(n_696), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_225), .A2(n_262), .B1(n_514), .B2(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_226), .B(n_346), .Y(n_657) );
AOI22xp33_ASAP7_75t_SL g493 ( .A1(n_227), .A2(n_263), .B1(n_407), .B2(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_228), .B(n_499), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g890 ( .A(n_229), .Y(n_890) );
INVx1_ASAP7_75t_L g678 ( .A(n_230), .Y(n_678) );
CKINVDCx20_ASAP7_75t_R g918 ( .A(n_232), .Y(n_918) );
NOR2xp33_ASAP7_75t_L g860 ( .A(n_235), .B(n_861), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_238), .B(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_241), .A2(n_273), .B1(n_323), .B2(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g831 ( .A(n_242), .Y(n_831) );
INVx1_ASAP7_75t_L g764 ( .A(n_244), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_249), .Y(n_673) );
INVx1_ASAP7_75t_L g684 ( .A(n_250), .Y(n_684) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_252), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_254), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g859 ( .A(n_255), .Y(n_859) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_256), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_257), .A2(n_270), .B1(n_365), .B2(n_551), .Y(n_550) );
AOI211xp5_ASAP7_75t_L g769 ( .A1(n_260), .A2(n_624), .B(n_770), .C(n_777), .Y(n_769) );
INVx1_ASAP7_75t_L g690 ( .A(n_261), .Y(n_690) );
CKINVDCx20_ASAP7_75t_R g884 ( .A(n_264), .Y(n_884) );
INVx1_ASAP7_75t_L g313 ( .A(n_267), .Y(n_313) );
INVx1_ASAP7_75t_L g315 ( .A(n_267), .Y(n_315) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_268), .Y(n_391) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_271), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g598 ( .A(n_272), .Y(n_598) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_274), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_275), .Y(n_530) );
INVx1_ASAP7_75t_L g691 ( .A(n_277), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_280), .Y(n_779) );
CKINVDCx20_ASAP7_75t_R g876 ( .A(n_282), .Y(n_876) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_283), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_284), .Y(n_401) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
HB1xp67_ASAP7_75t_L g855 ( .A(n_290), .Y(n_855) );
OAI21xp5_ASAP7_75t_L g925 ( .A1(n_291), .A2(n_854), .B(n_926), .Y(n_925) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_292), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_517), .B1(n_849), .B2(n_850), .C(n_851), .Y(n_295) );
INVx1_ASAP7_75t_L g850 ( .A(n_296), .Y(n_850) );
OAI22xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_298), .B1(n_440), .B2(n_516), .Y(n_296) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
BUFx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OAI22xp5_ASAP7_75t_SL g299 ( .A1(n_300), .A2(n_301), .B1(n_387), .B2(n_439), .Y(n_299) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
XOR2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_386), .Y(n_303) );
NAND4xp75_ASAP7_75t_L g304 ( .A(n_305), .B(n_340), .C(n_360), .D(n_374), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_329), .Y(n_305) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx3_ASAP7_75t_L g428 ( .A(n_308), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_308), .A2(n_461), .B1(n_462), .B2(n_463), .Y(n_460) );
INVx2_ASAP7_75t_L g505 ( .A(n_308), .Y(n_505) );
INVx2_ASAP7_75t_L g669 ( .A(n_308), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g915 ( .A1(n_308), .A2(n_916), .B1(n_917), .B2(n_918), .Y(n_915) );
INVx6_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
BUFx3_ASAP7_75t_L g551 ( .A(n_309), .Y(n_551) );
BUFx3_ASAP7_75t_L g561 ( .A(n_309), .Y(n_561) );
BUFx3_ASAP7_75t_L g704 ( .A(n_309), .Y(n_704) );
AND2x4_ASAP7_75t_L g309 ( .A(n_310), .B(n_319), .Y(n_309) );
AND2x6_ASAP7_75t_L g364 ( .A(n_310), .B(n_349), .Y(n_364) );
AND2x2_ASAP7_75t_L g370 ( .A(n_310), .B(n_332), .Y(n_370) );
AND2x6_ASAP7_75t_L g377 ( .A(n_310), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_316), .Y(n_310) );
AND2x2_ASAP7_75t_L g334 ( .A(n_311), .B(n_317), .Y(n_334) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g327 ( .A(n_312), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_312), .B(n_317), .Y(n_339) );
AND2x2_ASAP7_75t_L g356 ( .A(n_312), .B(n_322), .Y(n_356) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g318 ( .A(n_315), .Y(n_318) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g328 ( .A(n_317), .Y(n_328) );
INVx1_ASAP7_75t_L g355 ( .A(n_317), .Y(n_355) );
AND2x2_ASAP7_75t_L g326 ( .A(n_319), .B(n_327), .Y(n_326) );
NAND2x1p5_ASAP7_75t_L g344 ( .A(n_319), .B(n_334), .Y(n_344) );
AND2x6_ASAP7_75t_L g486 ( .A(n_319), .B(n_334), .Y(n_486) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx2_ASAP7_75t_L g333 ( .A(n_320), .Y(n_333) );
INVx1_ASAP7_75t_L g338 ( .A(n_320), .Y(n_338) );
OR2x2_ASAP7_75t_L g350 ( .A(n_320), .B(n_321), .Y(n_350) );
AND2x2_ASAP7_75t_L g378 ( .A(n_320), .B(n_322), .Y(n_378) );
AND2x2_ASAP7_75t_L g332 ( .A(n_321), .B(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx3_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
BUFx3_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx4_ASAP7_75t_L g453 ( .A(n_325), .Y(n_453) );
INVx3_ASAP7_75t_L g670 ( .A(n_325), .Y(n_670) );
INVx5_ASAP7_75t_L g728 ( .A(n_325), .Y(n_728) );
INVx1_ASAP7_75t_L g881 ( .A(n_325), .Y(n_881) );
INVx8_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g366 ( .A(n_327), .B(n_332), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_327), .B(n_332), .Y(n_465) );
INVx1_ASAP7_75t_L g385 ( .A(n_328), .Y(n_385) );
BUFx3_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_331), .Y(n_434) );
INVx2_ASAP7_75t_L g565 ( .A(n_331), .Y(n_565) );
BUFx3_ASAP7_75t_L g700 ( .A(n_331), .Y(n_700) );
AND2x4_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
AND2x4_ASAP7_75t_L g372 ( .A(n_332), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g354 ( .A(n_333), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g413 ( .A(n_333), .Y(n_413) );
AND2x4_ASAP7_75t_L g348 ( .A(n_334), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g394 ( .A(n_334), .Y(n_394) );
BUFx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx4f_ASAP7_75t_SL g425 ( .A(n_336), .Y(n_425) );
BUFx2_ASAP7_75t_L g454 ( .A(n_336), .Y(n_454) );
BUFx2_ASAP7_75t_L g507 ( .A(n_336), .Y(n_507) );
BUFx2_ASAP7_75t_L g696 ( .A(n_336), .Y(n_696) );
INVx6_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g546 ( .A(n_337), .Y(n_546) );
INVx1_ASAP7_75t_SL g612 ( .A(n_337), .Y(n_612) );
INVx1_ASAP7_75t_SL g790 ( .A(n_337), .Y(n_790) );
OR2x6_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_L g359 ( .A(n_338), .Y(n_359) );
INVx1_ASAP7_75t_L g373 ( .A(n_339), .Y(n_373) );
OA211x2_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_342), .B(n_345), .C(n_351), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_342), .A2(n_575), .B1(n_576), .B2(n_577), .Y(n_574) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g681 ( .A(n_343), .Y(n_681) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx3_ASAP7_75t_L g398 ( .A(n_344), .Y(n_398) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g484 ( .A(n_347), .Y(n_484) );
INVx5_ASAP7_75t_L g500 ( .A(n_347), .Y(n_500) );
INVx2_ASAP7_75t_L g602 ( .A(n_347), .Y(n_602) );
INVx4_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g393 ( .A(n_350), .B(n_394), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_352), .Y(n_812) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_353), .Y(n_404) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_353), .Y(n_473) );
BUFx4f_ASAP7_75t_SL g627 ( .A(n_353), .Y(n_627) );
BUFx2_ASAP7_75t_L g686 ( .A(n_353), .Y(n_686) );
AND2x4_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g382 ( .A(n_355), .Y(n_382) );
AND2x4_ASAP7_75t_L g358 ( .A(n_356), .B(n_359), .Y(n_358) );
AND2x4_ASAP7_75t_L g381 ( .A(n_356), .B(n_382), .Y(n_381) );
NAND2x1p5_ASAP7_75t_L g412 ( .A(n_356), .B(n_413), .Y(n_412) );
BUFx3_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g479 ( .A(n_358), .Y(n_479) );
BUFx2_ASAP7_75t_L g502 ( .A(n_358), .Y(n_502) );
BUFx2_ASAP7_75t_L g776 ( .A(n_358), .Y(n_776) );
AND2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_367), .Y(n_360) );
INVx2_ASAP7_75t_L g889 ( .A(n_362), .Y(n_889) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx5_ASAP7_75t_SL g458 ( .A(n_363), .Y(n_458) );
INVx4_ASAP7_75t_L g664 ( .A(n_363), .Y(n_664) );
INVx2_ASAP7_75t_L g699 ( .A(n_363), .Y(n_699) );
INVx11_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx11_ASAP7_75t_L g511 ( .A(n_364), .Y(n_511) );
INVx1_ASAP7_75t_L g430 ( .A(n_365), .Y(n_430) );
BUFx2_ASAP7_75t_L g562 ( .A(n_365), .Y(n_562) );
BUFx3_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx3_ASAP7_75t_L g512 ( .A(n_366), .Y(n_512) );
BUFx3_ASAP7_75t_L g665 ( .A(n_366), .Y(n_665) );
INVx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx3_ASAP7_75t_L g835 ( .A(n_369), .Y(n_835) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_370), .Y(n_423) );
BUFx2_ASAP7_75t_SL g514 ( .A(n_370), .Y(n_514) );
BUFx3_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx3_ASAP7_75t_L g436 ( .A(n_372), .Y(n_436) );
BUFx2_ASAP7_75t_SL g450 ( .A(n_372), .Y(n_450) );
BUFx2_ASAP7_75t_SL g542 ( .A(n_372), .Y(n_542) );
BUFx3_ASAP7_75t_L g567 ( .A(n_372), .Y(n_567) );
BUFx2_ASAP7_75t_L g642 ( .A(n_372), .Y(n_642) );
AND2x2_ASAP7_75t_L g672 ( .A(n_373), .B(n_413), .Y(n_672) );
INVx2_ASAP7_75t_L g683 ( .A(n_375), .Y(n_683) );
INVx4_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx2_ASAP7_75t_L g531 ( .A(n_376), .Y(n_531) );
OAI21xp5_ASAP7_75t_SL g751 ( .A1(n_376), .A2(n_752), .B(n_753), .Y(n_751) );
INVx4_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g400 ( .A(n_377), .Y(n_400) );
INVx2_ASAP7_75t_L g468 ( .A(n_377), .Y(n_468) );
INVx2_ASAP7_75t_SL g579 ( .A(n_377), .Y(n_579) );
BUFx3_ASAP7_75t_L g624 ( .A(n_377), .Y(n_624) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_377), .Y(n_654) );
AND2x4_ASAP7_75t_L g384 ( .A(n_378), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g417 ( .A(n_378), .Y(n_417) );
BUFx4f_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g782 ( .A(n_380), .Y(n_782) );
BUFx12f_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_381), .Y(n_407) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_381), .Y(n_475) );
BUFx2_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_384), .Y(n_482) );
BUFx2_ASAP7_75t_SL g494 ( .A(n_384), .Y(n_494) );
INVx1_ASAP7_75t_L g418 ( .A(n_385), .Y(n_418) );
INVx1_ASAP7_75t_L g439 ( .A(n_387), .Y(n_439) );
INVx2_ASAP7_75t_L g438 ( .A(n_388), .Y(n_438) );
AND2x2_ASAP7_75t_SL g388 ( .A(n_389), .B(n_419), .Y(n_388) );
NOR3xp33_ASAP7_75t_L g389 ( .A(n_390), .B(n_399), .C(n_408), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_392), .B1(n_395), .B2(n_396), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_392), .A2(n_681), .B1(n_749), .B2(n_750), .Y(n_748) );
BUFx3_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g527 ( .A(n_393), .Y(n_527) );
BUFx6f_ASAP7_75t_L g732 ( .A(n_393), .Y(n_732) );
OAI221xp5_ASAP7_75t_L g840 ( .A1(n_393), .A2(n_398), .B1(n_841), .B2(n_842), .C(n_843), .Y(n_840) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_396), .A2(n_525), .B1(n_526), .B2(n_528), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g807 ( .A1(n_396), .A2(n_679), .B1(n_808), .B2(n_809), .Y(n_807) );
OAI22xp5_ASAP7_75t_SL g868 ( .A1(n_396), .A2(n_679), .B1(n_869), .B2(n_870), .Y(n_868) );
OAI211xp5_ASAP7_75t_L g902 ( .A1(n_396), .A2(n_903), .B(n_904), .C(n_905), .Y(n_902) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_398), .A2(n_731), .B1(n_732), .B2(n_733), .Y(n_730) );
BUFx3_ASAP7_75t_L g772 ( .A(n_398), .Y(n_772) );
OAI221xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B1(n_402), .B2(n_405), .C(n_406), .Y(n_399) );
OAI21xp5_ASAP7_75t_SL g491 ( .A1(n_400), .A2(n_492), .B(n_493), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_402), .A2(n_412), .B1(n_755), .B2(n_756), .Y(n_754) );
INVx2_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_SL g581 ( .A(n_403), .Y(n_581) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g908 ( .A(n_404), .Y(n_908) );
INVx2_ASAP7_75t_L g585 ( .A(n_407), .Y(n_585) );
BUFx3_ASAP7_75t_L g738 ( .A(n_407), .Y(n_738) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B1(n_414), .B2(n_415), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_410), .A2(n_535), .B1(n_536), .B2(n_537), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_410), .A2(n_590), .B1(n_816), .B2(n_817), .Y(n_815) );
INVx3_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g588 ( .A(n_411), .Y(n_588) );
INVx4_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_412), .A2(n_537), .B1(n_690), .B2(n_691), .Y(n_689) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_412), .Y(n_741) );
BUFx3_ASAP7_75t_L g877 ( .A(n_412), .Y(n_877) );
BUFx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
CKINVDCx16_ASAP7_75t_R g538 ( .A(n_416), .Y(n_538) );
OR2x6_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_420), .B(n_426), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_424), .Y(n_420) );
BUFx3_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_423), .Y(n_449) );
BUFx3_ASAP7_75t_L g570 ( .A(n_423), .Y(n_570) );
INVx3_ASAP7_75t_L g787 ( .A(n_423), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_431), .Y(n_426) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx4_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_433), .A2(n_456), .B1(n_457), .B2(n_459), .Y(n_455) );
INVx3_ASAP7_75t_L g913 ( .A(n_433), .Y(n_913) );
INVx4_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g826 ( .A(n_436), .Y(n_826) );
INVx1_ASAP7_75t_L g516 ( .A(n_440), .Y(n_516) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B1(n_487), .B2(n_488), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_446), .B(n_466), .Y(n_445) );
NOR3xp33_ASAP7_75t_L g446 ( .A(n_447), .B(n_455), .C(n_460), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_451), .Y(n_447) );
INVx1_ASAP7_75t_SL g921 ( .A(n_449), .Y(n_921) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g545 ( .A(n_453), .Y(n_545) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_458), .Y(n_788) );
OAI22xp5_ASAP7_75t_L g888 ( .A1(n_463), .A2(n_889), .B1(n_890), .B2(n_891), .Y(n_888) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g795 ( .A(n_464), .Y(n_795) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_476), .Y(n_466) );
OAI21xp5_ASAP7_75t_SL g467 ( .A1(n_468), .A2(n_469), .B(n_470), .Y(n_467) );
OAI21xp5_ASAP7_75t_SL g597 ( .A1(n_468), .A2(n_598), .B(n_599), .Y(n_597) );
INVx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx4_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx2_ASAP7_75t_L g533 ( .A(n_473), .Y(n_533) );
BUFx4f_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_483), .Y(n_476) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
BUFx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx2_ASAP7_75t_L g497 ( .A(n_486), .Y(n_497) );
INVx1_ASAP7_75t_SL g631 ( .A(n_486), .Y(n_631) );
BUFx4f_ASAP7_75t_L g659 ( .A(n_486), .Y(n_659) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
XOR2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_515), .Y(n_488) );
NAND3x1_ASAP7_75t_L g489 ( .A(n_490), .B(n_503), .C(n_508), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_491), .B(n_495), .Y(n_490) );
NAND3xp33_ASAP7_75t_L g495 ( .A(n_496), .B(n_498), .C(n_501), .Y(n_495) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_506), .Y(n_503) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_513), .Y(n_508) );
INVx4_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_SL g549 ( .A(n_511), .Y(n_549) );
INVx3_ASAP7_75t_L g571 ( .A(n_511), .Y(n_571) );
INVx4_ASAP7_75t_L g640 ( .A(n_511), .Y(n_640) );
BUFx3_ASAP7_75t_L g725 ( .A(n_512), .Y(n_725) );
INVx1_ASAP7_75t_L g885 ( .A(n_514), .Y(n_885) );
INVxp67_ASAP7_75t_L g849 ( .A(n_517), .Y(n_849) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B1(n_712), .B2(n_713), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_616), .B1(n_710), .B2(n_711), .Y(n_519) );
INVx1_ASAP7_75t_L g710 ( .A(n_520), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_553), .B1(n_554), .B2(n_615), .Y(n_520) );
INVx1_ASAP7_75t_L g615 ( .A(n_521), .Y(n_615) );
XOR2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_552), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_539), .Y(n_522) );
NOR3xp33_ASAP7_75t_L g523 ( .A(n_524), .B(n_529), .C(n_534), .Y(n_523) );
INVx1_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g576 ( .A(n_527), .Y(n_576) );
INVx2_ASAP7_75t_L g679 ( .A(n_527), .Y(n_679) );
OAI21xp33_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B(n_532), .Y(n_529) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g590 ( .A(n_538), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_540), .B(n_547), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
INVx1_ASAP7_75t_SL g887 ( .A(n_542), .Y(n_887) );
INVx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
OAI22xp5_ASAP7_75t_SL g554 ( .A1(n_555), .A2(n_593), .B1(n_594), .B2(n_614), .Y(n_554) );
INVx2_ASAP7_75t_L g614 ( .A(n_555), .Y(n_614) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g592 ( .A(n_557), .Y(n_592) );
AND2x2_ASAP7_75t_SL g557 ( .A(n_558), .B(n_573), .Y(n_557) );
NOR2xp33_ASAP7_75t_SL g558 ( .A(n_559), .B(n_568), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .Y(n_559) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_565), .A2(n_797), .B1(n_798), .B2(n_799), .Y(n_796) );
INVx1_ASAP7_75t_L g799 ( .A(n_566), .Y(n_799) );
BUFx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_572), .Y(n_568) );
INVx1_ASAP7_75t_L g917 ( .A(n_571), .Y(n_917) );
NOR3xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_578), .C(n_586), .Y(n_573) );
OAI221xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_580), .B1(n_581), .B2(n_582), .C(n_583), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_581), .A2(n_778), .B1(n_779), .B2(n_780), .Y(n_777) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_588), .B1(n_589), .B2(n_590), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_590), .A2(n_740), .B1(n_741), .B2(n_742), .Y(n_739) );
INVx3_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
XOR2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_613), .Y(n_594) );
NAND2x1_ASAP7_75t_SL g595 ( .A(n_596), .B(n_605), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_600), .Y(n_596) );
NAND3xp33_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .C(n_604), .Y(n_600) );
BUFx2_ASAP7_75t_L g774 ( .A(n_602), .Y(n_774) );
NOR2x1_ASAP7_75t_L g605 ( .A(n_606), .B(n_609), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_L g711 ( .A(n_616), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_644), .B1(n_645), .B2(n_709), .Y(n_616) );
INVx1_ASAP7_75t_L g709 ( .A(n_617), .Y(n_709) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g643 ( .A(n_620), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_621), .B(n_634), .Y(n_620) );
NOR2xp67_ASAP7_75t_L g621 ( .A(n_622), .B(n_628), .Y(n_621) );
OAI21xp5_ASAP7_75t_SL g622 ( .A1(n_623), .A2(n_625), .B(n_626), .Y(n_622) );
OAI21xp5_ASAP7_75t_SL g844 ( .A1(n_623), .A2(n_845), .B(n_846), .Y(n_844) );
OAI21xp33_ASAP7_75t_L g871 ( .A1(n_623), .A2(n_872), .B(n_873), .Y(n_871) );
INVx3_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND3xp33_ASAP7_75t_L g628 ( .A(n_629), .B(n_632), .C(n_633), .Y(n_628) );
INVx1_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
NOR2x1_ASAP7_75t_L g634 ( .A(n_635), .B(n_638), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_641), .Y(n_638) );
INVx4_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
XOR2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_674), .Y(n_645) );
INVx2_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
INVx3_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
XOR2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_673), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_650), .B(n_661), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_656), .Y(n_650) );
OAI21xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B(n_655), .Y(n_651) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND3xp33_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .C(n_660), .Y(n_656) );
NOR2x1_ASAP7_75t_L g661 ( .A(n_662), .B(n_667), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_666), .Y(n_662) );
INVx1_ASAP7_75t_L g706 ( .A(n_665), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_671), .Y(n_667) );
INVxp67_ASAP7_75t_L g793 ( .A(n_669), .Y(n_793) );
INVx1_ASAP7_75t_SL g707 ( .A(n_675), .Y(n_707) );
AND2x2_ASAP7_75t_SL g675 ( .A(n_676), .B(n_692), .Y(n_675) );
NOR3xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_682), .C(n_689), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B1(n_680), .B2(n_681), .Y(n_677) );
OAI221xp5_ASAP7_75t_SL g682 ( .A1(n_683), .A2(n_684), .B1(n_685), .B2(n_687), .C(n_688), .Y(n_682) );
OAI221xp5_ASAP7_75t_SL g734 ( .A1(n_683), .A2(n_685), .B1(n_735), .B2(n_736), .C(n_737), .Y(n_734) );
OAI221xp5_ASAP7_75t_SL g810 ( .A1(n_683), .A2(n_811), .B1(n_812), .B2(n_813), .C(n_814), .Y(n_810) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_697), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_698), .B(n_701), .Y(n_697) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx3_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
OAI22xp5_ASAP7_75t_SL g713 ( .A1(n_714), .A2(n_802), .B1(n_847), .B2(n_848), .Y(n_713) );
INVx1_ASAP7_75t_L g847 ( .A(n_714), .Y(n_847) );
OAI22xp5_ASAP7_75t_SL g714 ( .A1(n_715), .A2(n_766), .B1(n_800), .B2(n_801), .Y(n_714) );
INVx1_ASAP7_75t_L g800 ( .A(n_715), .Y(n_800) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_717), .B1(n_745), .B2(n_765), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g744 ( .A(n_718), .Y(n_744) );
AND2x2_ASAP7_75t_SL g718 ( .A(n_719), .B(n_729), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_723), .Y(n_719) );
NAND2xp33_ASAP7_75t_SL g720 ( .A(n_721), .B(n_722), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_724), .B(n_726), .Y(n_723) );
BUFx6f_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NOR3xp33_ASAP7_75t_L g729 ( .A(n_730), .B(n_734), .C(n_739), .Y(n_729) );
INVx1_ASAP7_75t_L g765 ( .A(n_745), .Y(n_765) );
XOR2x2_ASAP7_75t_L g745 ( .A(n_746), .B(n_764), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_757), .Y(n_746) );
NOR3xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_751), .C(n_754), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_758), .B(n_761), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .Y(n_761) );
INVx2_ASAP7_75t_L g801 ( .A(n_766), .Y(n_801) );
XNOR2x1_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
AND2x2_ASAP7_75t_L g768 ( .A(n_769), .B(n_783), .Y(n_768) );
OAI211xp5_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_772), .B(n_773), .C(n_775), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g906 ( .A1(n_780), .A2(n_907), .B1(n_908), .B2(n_909), .Y(n_906) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx3_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
NOR3xp33_ASAP7_75t_L g783 ( .A(n_784), .B(n_791), .C(n_796), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_785), .B(n_789), .Y(n_784) );
INVx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_793), .B1(n_794), .B2(n_795), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_795), .A2(n_920), .B1(n_921), .B2(n_922), .Y(n_919) );
INVx2_ASAP7_75t_L g848 ( .A(n_802), .Y(n_848) );
OAI22xp5_ASAP7_75t_SL g802 ( .A1(n_803), .A2(n_804), .B1(n_829), .B2(n_830), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx2_ASAP7_75t_L g828 ( .A(n_805), .Y(n_828) );
AND2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_818), .Y(n_805) );
NOR3xp33_ASAP7_75t_L g806 ( .A(n_807), .B(n_810), .C(n_815), .Y(n_806) );
OAI22xp33_ASAP7_75t_L g874 ( .A1(n_812), .A2(n_875), .B1(n_876), .B2(n_877), .Y(n_874) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_819), .B(n_822), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .Y(n_822) );
INVx2_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx2_ASAP7_75t_SL g829 ( .A(n_830), .Y(n_829) );
XNOR2x2_ASAP7_75t_L g830 ( .A(n_831), .B(n_832), .Y(n_830) );
NOR4xp75_ASAP7_75t_L g832 ( .A(n_833), .B(n_837), .C(n_840), .D(n_844), .Y(n_832) );
NAND2xp5_ASAP7_75t_SL g833 ( .A(n_834), .B(n_836), .Y(n_833) );
NAND2xp5_ASAP7_75t_SL g837 ( .A(n_838), .B(n_839), .Y(n_837) );
INVx1_ASAP7_75t_SL g851 ( .A(n_852), .Y(n_851) );
NOR2x1_ASAP7_75t_L g852 ( .A(n_853), .B(n_857), .Y(n_852) );
OR2x2_ASAP7_75t_SL g923 ( .A(n_853), .B(n_858), .Y(n_923) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_854), .B(n_856), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_854), .B(n_895), .Y(n_894) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_855), .B(n_895), .Y(n_926) );
CKINVDCx16_ASAP7_75t_R g895 ( .A(n_856), .Y(n_895) );
CKINVDCx20_ASAP7_75t_R g857 ( .A(n_858), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_859), .B(n_860), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_862), .B(n_863), .Y(n_861) );
OAI222xp33_ASAP7_75t_L g864 ( .A1(n_865), .A2(n_894), .B1(n_896), .B2(n_899), .C1(n_923), .C2(n_924), .Y(n_864) );
INVx2_ASAP7_75t_SL g893 ( .A(n_866), .Y(n_893) );
AND2x2_ASAP7_75t_L g866 ( .A(n_867), .B(n_878), .Y(n_866) );
NOR3xp33_ASAP7_75t_L g867 ( .A(n_868), .B(n_871), .C(n_874), .Y(n_867) );
NOR3xp33_ASAP7_75t_L g878 ( .A(n_879), .B(n_883), .C(n_888), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_880), .B(n_882), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g883 ( .A1(n_884), .A2(n_885), .B1(n_886), .B2(n_887), .Y(n_883) );
INVx1_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
INVx2_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
XNOR2xp5_ASAP7_75t_L g898 ( .A(n_899), .B(n_900), .Y(n_898) );
AND2x2_ASAP7_75t_L g900 ( .A(n_901), .B(n_910), .Y(n_900) );
NOR3xp33_ASAP7_75t_L g910 ( .A(n_911), .B(n_915), .C(n_919), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_912), .B(n_914), .Y(n_911) );
CKINVDCx16_ASAP7_75t_R g924 ( .A(n_925), .Y(n_924) );
endmodule