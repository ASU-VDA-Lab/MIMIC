module fake_jpeg_3511_n_74 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_74);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_74;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_73;
wire n_59;
wire n_71;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_24;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_21),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_28),
.B(n_0),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_36),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_10),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_26),
.Y(n_42)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_25),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_29),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_30),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_51),
.Y(n_57)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_48),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_32),
.B1(n_34),
.B2(n_29),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_49),
.A2(n_36),
.B1(n_28),
.B2(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_9),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_33),
.C(n_30),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_24),
.C(n_23),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_59),
.C(n_1),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_24),
.B(n_40),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_52),
.B(n_53),
.C(n_3),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_17),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_11),
.C(n_20),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_52),
.B(n_7),
.Y(n_60)
);

MAJx2_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_61),
.C(n_65),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_SL g61 ( 
.A(n_57),
.B(n_0),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_SL g68 ( 
.A1(n_63),
.A2(n_64),
.B(n_66),
.C(n_5),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_5),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_60),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_67),
.B1(n_69),
.B2(n_6),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_6),
.Y(n_72)
);

FAx1_ASAP7_75t_SL g73 ( 
.A(n_72),
.B(n_13),
.CI(n_16),
.CON(n_73),
.SN(n_73)
);

O2A1O1Ixp33_ASAP7_75t_SL g74 ( 
.A1(n_73),
.A2(n_22),
.B(n_18),
.C(n_19),
.Y(n_74)
);


endmodule