module fake_netlist_1_7563_n_1185 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_182, n_166, n_162, n_186, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_92, n_11, n_25, n_30, n_59, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_96, n_39, n_1185, n_1186);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_96;
input n_39;
output n_1185;
output n_1186;
wire n_1173;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_1092;
wire n_963;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_1158;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_1022;
wire n_918;
wire n_252;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_1122;
wire n_528;
wire n_383;
wire n_288;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_1175;
wire n_853;
wire n_1161;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_1177;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_1185;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_1163;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_857;
wire n_786;
wire n_345;
wire n_360;
wire n_1090;
wire n_236;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_1179;
wire n_222;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1174;
wire n_246;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1024;
wire n_1016;
wire n_1078;
wire n_572;
wire n_1017;
wire n_324;
wire n_1097;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_1169;
wire n_652;
wire n_975;
wire n_279;
wire n_303;
wire n_1060;
wire n_968;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_1011;
wire n_1025;
wire n_1132;
wire n_880;
wire n_1101;
wire n_1159;
wire n_630;
wire n_1155;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_1180;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_844;
wire n_818;
wire n_1160;
wire n_1184;
wire n_230;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_828;
wire n_767;
wire n_1063;
wire n_293;
wire n_1138;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_1171;
wire n_665;
wire n_571;
wire n_1154;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_950;
wire n_460;
wire n_1046;
wire n_478;
wire n_243;
wire n_415;
wire n_235;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_1076;
wire n_268;
wire n_882;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_1145;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_1167;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_1157;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_1147;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_1178;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_224;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_996;
wire n_1176;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_446;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_666;
wire n_799;
wire n_1089;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_1181;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_716;
wire n_653;
wire n_899;
wire n_260;
wire n_806;
wire n_881;
wire n_539;
wire n_1055;
wire n_1066;
wire n_974;
wire n_1153;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_1144;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_1152;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_1149;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_1170;
wire n_419;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_1125;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_955;
wire n_1133;
wire n_429;
wire n_488;
wire n_233;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_553;
wire n_440;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1131;
wire n_1102;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_1069;
wire n_1021;
wire n_1123;
wire n_811;
wire n_972;
wire n_1039;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_1156;
wire n_221;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_912;
wire n_947;
wire n_1043;
wire n_1141;
wire n_378;
wire n_582;
wire n_924;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_272;
wire n_1172;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1142;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1117;
wire n_1040;
wire n_1165;
wire n_994;
wire n_930;
wire n_1182;
wire n_424;
wire n_714;
wire n_1143;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_1168;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_581;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1164;
wire n_1038;
wire n_341;
wire n_1162;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_1150;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_1104;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_287;
wire n_1146;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_1137;
wire n_781;
wire n_916;
wire n_421;
wire n_1148;
wire n_709;
wire n_739;
wire n_1166;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_257;
wire n_992;
wire n_1127;
wire n_269;
INVx1_ASAP7_75t_L g221 ( .A(n_83), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_113), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_122), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_168), .Y(n_224) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_110), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_165), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_146), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_187), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_92), .Y(n_229) );
INVxp67_ASAP7_75t_L g230 ( .A(n_216), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_116), .Y(n_231) );
INVx1_ASAP7_75t_SL g232 ( .A(n_26), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_74), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_125), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_177), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_42), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_21), .Y(n_237) );
INVxp67_ASAP7_75t_SL g238 ( .A(n_211), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_139), .Y(n_239) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_203), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_189), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_148), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_42), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_1), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_32), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_173), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_214), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g248 ( .A(n_19), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_204), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_121), .Y(n_250) );
INVx1_ASAP7_75t_SL g251 ( .A(n_155), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_17), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_28), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_154), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_69), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_152), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_119), .Y(n_257) );
CKINVDCx14_ASAP7_75t_R g258 ( .A(n_219), .Y(n_258) );
INVx1_ASAP7_75t_SL g259 ( .A(n_1), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_186), .Y(n_260) );
CKINVDCx16_ASAP7_75t_R g261 ( .A(n_201), .Y(n_261) );
INVx1_ASAP7_75t_SL g262 ( .A(n_162), .Y(n_262) );
INVx2_ASAP7_75t_SL g263 ( .A(n_29), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_120), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_0), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_196), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_183), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_127), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_19), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_157), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_105), .Y(n_271) );
BUFx5_ASAP7_75t_L g272 ( .A(n_141), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_124), .Y(n_273) );
BUFx8_ASAP7_75t_SL g274 ( .A(n_218), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_171), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_202), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_104), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_10), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_108), .Y(n_279) );
CKINVDCx20_ASAP7_75t_R g280 ( .A(n_129), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_8), .Y(n_281) );
CKINVDCx20_ASAP7_75t_R g282 ( .A(n_18), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_107), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_21), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_220), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_175), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_118), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_161), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_106), .Y(n_289) );
CKINVDCx16_ASAP7_75t_R g290 ( .A(n_140), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_82), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_197), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_169), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_159), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_115), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_55), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_103), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_138), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_185), .Y(n_299) );
BUFx3_ASAP7_75t_L g300 ( .A(n_207), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_41), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_163), .Y(n_302) );
CKINVDCx16_ASAP7_75t_R g303 ( .A(n_178), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_209), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_208), .Y(n_305) );
CKINVDCx20_ASAP7_75t_R g306 ( .A(n_199), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_164), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_172), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_56), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_184), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_206), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_131), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_52), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_126), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_114), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_117), .Y(n_316) );
NOR2xp67_ASAP7_75t_L g317 ( .A(n_6), .B(n_195), .Y(n_317) );
CKINVDCx20_ASAP7_75t_R g318 ( .A(n_200), .Y(n_318) );
NOR2xp67_ASAP7_75t_L g319 ( .A(n_2), .B(n_50), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_10), .Y(n_320) );
INVx1_ASAP7_75t_SL g321 ( .A(n_74), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_132), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_5), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_9), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_213), .Y(n_325) );
INVxp33_ASAP7_75t_L g326 ( .A(n_123), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_133), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_156), .Y(n_328) );
CKINVDCx16_ASAP7_75t_R g329 ( .A(n_198), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_31), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_11), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_77), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_160), .Y(n_333) );
CKINVDCx20_ASAP7_75t_R g334 ( .A(n_176), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_93), .Y(n_335) );
CKINVDCx20_ASAP7_75t_R g336 ( .A(n_212), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_48), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_153), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_73), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_48), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_7), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_47), .Y(n_342) );
BUFx3_ASAP7_75t_L g343 ( .A(n_205), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_174), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_158), .Y(n_345) );
CKINVDCx20_ASAP7_75t_R g346 ( .A(n_65), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_58), .Y(n_347) );
BUFx3_ASAP7_75t_L g348 ( .A(n_5), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_22), .Y(n_349) );
CKINVDCx16_ASAP7_75t_R g350 ( .A(n_130), .Y(n_350) );
INVxp67_ASAP7_75t_SL g351 ( .A(n_217), .Y(n_351) );
BUFx10_ASAP7_75t_L g352 ( .A(n_136), .Y(n_352) );
BUFx10_ASAP7_75t_L g353 ( .A(n_33), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_190), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_188), .Y(n_355) );
BUFx10_ASAP7_75t_L g356 ( .A(n_54), .Y(n_356) );
CKINVDCx20_ASAP7_75t_R g357 ( .A(n_151), .Y(n_357) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_182), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_100), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_166), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_91), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_87), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_210), .Y(n_363) );
INVx6_ASAP7_75t_L g364 ( .A(n_352), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_284), .Y(n_365) );
INVx6_ASAP7_75t_L g366 ( .A(n_352), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_284), .Y(n_367) );
BUFx6f_ASAP7_75t_L g368 ( .A(n_240), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_309), .Y(n_369) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_240), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_272), .Y(n_371) );
INVx3_ASAP7_75t_L g372 ( .A(n_352), .Y(n_372) );
OAI21x1_ASAP7_75t_L g373 ( .A1(n_256), .A2(n_97), .B(n_96), .Y(n_373) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_240), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_263), .B(n_0), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_272), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_272), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_272), .Y(n_378) );
INVxp33_ASAP7_75t_SL g379 ( .A(n_279), .Y(n_379) );
CKINVDCx20_ASAP7_75t_R g380 ( .A(n_236), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_348), .B(n_2), .Y(n_381) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_240), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_348), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_309), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_274), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_320), .Y(n_386) );
OA21x2_ASAP7_75t_L g387 ( .A1(n_256), .A2(n_99), .B(n_98), .Y(n_387) );
INVx6_ASAP7_75t_L g388 ( .A(n_272), .Y(n_388) );
BUFx2_ASAP7_75t_L g389 ( .A(n_274), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_272), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_320), .Y(n_391) );
AND2x6_ASAP7_75t_L g392 ( .A(n_300), .B(n_101), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_327), .B(n_3), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_272), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_257), .B(n_3), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_302), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_222), .Y(n_397) );
CKINVDCx6p67_ASAP7_75t_R g398 ( .A(n_261), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_221), .B(n_4), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_326), .B(n_6), .Y(n_400) );
INVx3_ASAP7_75t_L g401 ( .A(n_296), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_302), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_223), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_302), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_302), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_371), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_371), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_395), .A2(n_229), .B1(n_243), .B2(n_237), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_398), .A2(n_267), .B1(n_280), .B2(n_226), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_389), .B(n_232), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_395), .A2(n_244), .B1(n_252), .B2(n_245), .Y(n_411) );
INVx3_ASAP7_75t_L g412 ( .A(n_395), .Y(n_412) );
INVx3_ASAP7_75t_L g413 ( .A(n_395), .Y(n_413) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_368), .Y(n_414) );
BUFx2_ASAP7_75t_L g415 ( .A(n_389), .Y(n_415) );
INVx2_ASAP7_75t_SL g416 ( .A(n_364), .Y(n_416) );
INVx3_ASAP7_75t_L g417 ( .A(n_395), .Y(n_417) );
INVx2_ASAP7_75t_SL g418 ( .A(n_364), .Y(n_418) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_372), .B(n_290), .Y(n_419) );
INVx3_ASAP7_75t_L g420 ( .A(n_381), .Y(n_420) );
BUFx2_ASAP7_75t_L g421 ( .A(n_398), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_376), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g423 ( .A(n_372), .B(n_303), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g424 ( .A(n_372), .B(n_329), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_376), .Y(n_425) );
INVx2_ASAP7_75t_SL g426 ( .A(n_364), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_372), .B(n_326), .Y(n_427) );
AND2x6_ASAP7_75t_L g428 ( .A(n_381), .B(n_300), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_377), .Y(n_429) );
OR2x6_ASAP7_75t_L g430 ( .A(n_400), .B(n_319), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_377), .Y(n_431) );
INVx8_ASAP7_75t_L g432 ( .A(n_392), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_364), .B(n_350), .Y(n_433) );
OR2x6_ASAP7_75t_L g434 ( .A(n_400), .B(n_253), .Y(n_434) );
NAND3xp33_ASAP7_75t_L g435 ( .A(n_397), .B(n_234), .C(n_231), .Y(n_435) );
INVx2_ASAP7_75t_SL g436 ( .A(n_364), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_378), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_378), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_366), .B(n_230), .Y(n_439) );
NOR3xp33_ASAP7_75t_L g440 ( .A(n_393), .B(n_321), .C(n_259), .Y(n_440) );
NOR2xp33_ASAP7_75t_SL g441 ( .A(n_392), .B(n_226), .Y(n_441) );
INVx3_ASAP7_75t_L g442 ( .A(n_381), .Y(n_442) );
OR2x6_ASAP7_75t_L g443 ( .A(n_400), .B(n_269), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_381), .A2(n_379), .B1(n_398), .B2(n_280), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_397), .B(n_289), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_366), .B(n_403), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_390), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_366), .B(n_289), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_390), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_366), .B(n_258), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_366), .B(n_277), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_380), .Y(n_452) );
INVx4_ASAP7_75t_L g453 ( .A(n_388), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_427), .B(n_383), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_420), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_419), .B(n_403), .Y(n_456) );
INVxp67_ASAP7_75t_SL g457 ( .A(n_412), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_432), .A2(n_373), .B(n_387), .Y(n_458) );
NOR2xp33_ASAP7_75t_SL g459 ( .A(n_441), .B(n_267), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_420), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_446), .B(n_393), .Y(n_461) );
BUFx3_ASAP7_75t_L g462 ( .A(n_421), .Y(n_462) );
NOR2x1p5_ASAP7_75t_L g463 ( .A(n_410), .B(n_385), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_423), .B(n_375), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_433), .B(n_399), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_432), .A2(n_373), .B(n_387), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_442), .A2(n_394), .B(n_373), .C(n_399), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_413), .A2(n_392), .B1(n_388), .B2(n_394), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_441), .B(n_224), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_434), .B(n_388), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_434), .B(n_388), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_424), .B(n_365), .Y(n_472) );
OR2x2_ASAP7_75t_SL g473 ( .A(n_410), .B(n_236), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_434), .B(n_258), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_413), .Y(n_475) );
AND2x4_ASAP7_75t_L g476 ( .A(n_443), .B(n_306), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_415), .B(n_353), .Y(n_477) );
AOI22xp33_ASAP7_75t_SL g478 ( .A1(n_409), .A2(n_248), .B1(n_346), .B2(n_282), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_408), .B(n_225), .Y(n_479) );
OR2x6_ASAP7_75t_L g480 ( .A(n_443), .B(n_291), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_443), .B(n_365), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_439), .B(n_367), .Y(n_482) );
NAND3xp33_ASAP7_75t_SL g483 ( .A(n_444), .B(n_318), .C(n_306), .Y(n_483) );
OAI22xp33_ASAP7_75t_L g484 ( .A1(n_444), .A2(n_334), .B1(n_336), .B2(n_318), .Y(n_484) );
OR2x6_ASAP7_75t_L g485 ( .A(n_430), .B(n_301), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_428), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_451), .B(n_367), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_411), .B(n_227), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_417), .A2(n_392), .B1(n_394), .B2(n_384), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_417), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_430), .A2(n_357), .B1(n_233), .B2(n_265), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_448), .B(n_369), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_417), .A2(n_384), .B(n_386), .C(n_369), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_445), .B(n_386), .Y(n_494) );
BUFx3_ASAP7_75t_L g495 ( .A(n_416), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_430), .A2(n_278), .B1(n_281), .B2(n_255), .Y(n_496) );
AND2x4_ASAP7_75t_L g497 ( .A(n_430), .B(n_391), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_450), .B(n_228), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_442), .A2(n_324), .B1(n_331), .B2(n_313), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_418), .B(n_235), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_418), .B(n_239), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_428), .A2(n_392), .B1(n_323), .B2(n_330), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_426), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_406), .B(n_241), .Y(n_504) );
AOI22xp5_ASAP7_75t_SL g505 ( .A1(n_452), .A2(n_248), .B1(n_346), .B2(n_282), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_435), .A2(n_392), .B1(n_332), .B2(n_337), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_436), .B(n_356), .Y(n_507) );
OAI22xp33_ASAP7_75t_L g508 ( .A1(n_435), .A2(n_335), .B1(n_342), .B2(n_341), .Y(n_508) );
INVx2_ASAP7_75t_SL g509 ( .A(n_432), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_447), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_447), .B(n_453), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_453), .B(n_242), .Y(n_512) );
NAND2xp33_ASAP7_75t_L g513 ( .A(n_407), .B(n_283), .Y(n_513) );
OR2x6_ASAP7_75t_L g514 ( .A(n_407), .B(n_349), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_422), .B(n_293), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_425), .A2(n_362), .B1(n_387), .B2(n_296), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_429), .A2(n_387), .B1(n_296), .B2(n_246), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_429), .A2(n_296), .B1(n_247), .B2(n_250), .Y(n_518) );
BUFx12f_ASAP7_75t_L g519 ( .A(n_414), .Y(n_519) );
NOR2x1p5_ASAP7_75t_L g520 ( .A(n_431), .B(n_339), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_437), .B(n_249), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_437), .A2(n_340), .B1(n_361), .B2(n_347), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_438), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_449), .B(n_254), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_458), .A2(n_351), .B(n_238), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_480), .A2(n_260), .B1(n_266), .B2(n_264), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_466), .A2(n_271), .B(n_268), .Y(n_527) );
O2A1O1Ixp33_ASAP7_75t_L g528 ( .A1(n_454), .A2(n_275), .B(n_285), .C(n_273), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_461), .B(n_298), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_480), .A2(n_287), .B1(n_292), .B2(n_286), .Y(n_530) );
INVx4_ASAP7_75t_L g531 ( .A(n_480), .Y(n_531) );
O2A1O1Ixp33_ASAP7_75t_L g532 ( .A1(n_508), .A2(n_295), .B(n_297), .C(n_294), .Y(n_532) );
BUFx2_ASAP7_75t_L g533 ( .A(n_476), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_SL g534 ( .A1(n_501), .A2(n_401), .B(n_402), .C(n_396), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_476), .A2(n_305), .B1(n_308), .B2(n_299), .Y(n_535) );
BUFx8_ASAP7_75t_L g536 ( .A(n_462), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_464), .B(n_304), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_467), .A2(n_325), .B(n_322), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_459), .B(n_307), .Y(n_539) );
NOR3xp33_ASAP7_75t_L g540 ( .A(n_483), .B(n_262), .C(n_251), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_490), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_481), .B(n_310), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_470), .B(n_312), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_471), .A2(n_344), .B(n_338), .Y(n_544) );
OAI21xp33_ASAP7_75t_L g545 ( .A1(n_456), .A2(n_315), .B(n_314), .Y(n_545) );
BUFx3_ASAP7_75t_L g546 ( .A(n_497), .Y(n_546) );
OAI22x1_ASAP7_75t_L g547 ( .A1(n_491), .A2(n_328), .B1(n_333), .B2(n_316), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_511), .A2(n_359), .B(n_345), .Y(n_548) );
AND2x4_ASAP7_75t_L g549 ( .A(n_497), .B(n_317), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_457), .A2(n_276), .B(n_270), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_456), .B(n_354), .Y(n_551) );
BUFx2_ASAP7_75t_L g552 ( .A(n_514), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_457), .A2(n_288), .B(n_276), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_472), .A2(n_311), .B1(n_355), .B2(n_288), .Y(n_554) );
A2O1A1Ixp33_ASAP7_75t_L g555 ( .A1(n_493), .A2(n_355), .B(n_360), .C(n_311), .Y(n_555) );
O2A1O1Ixp33_ASAP7_75t_L g556 ( .A1(n_508), .A2(n_360), .B(n_401), .C(n_363), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_486), .B(n_343), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_477), .B(n_9), .Y(n_558) );
A2O1A1Ixp33_ASAP7_75t_L g559 ( .A1(n_494), .A2(n_401), .B(n_402), .C(n_396), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_460), .A2(n_404), .B(n_402), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_494), .B(n_11), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_486), .B(n_358), .Y(n_562) );
NOR2xp33_ASAP7_75t_R g563 ( .A(n_502), .B(n_12), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_507), .B(n_12), .Y(n_564) );
OAI21xp33_ASAP7_75t_L g565 ( .A1(n_474), .A2(n_405), .B(n_404), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_492), .A2(n_405), .B(n_404), .Y(n_566) );
BUFx6f_ASAP7_75t_L g567 ( .A(n_519), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_510), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_517), .A2(n_414), .B(n_370), .Y(n_569) );
AO32x1_ASAP7_75t_L g570 ( .A1(n_503), .A2(n_382), .A3(n_374), .B1(n_370), .B2(n_368), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_520), .B(n_13), .Y(n_571) );
NAND2x1p5_ASAP7_75t_L g572 ( .A(n_463), .B(n_13), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_496), .B(n_14), .Y(n_573) );
O2A1O1Ixp33_ASAP7_75t_L g574 ( .A1(n_479), .A2(n_16), .B(n_14), .C(n_15), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_485), .B(n_15), .Y(n_575) );
NOR3xp33_ASAP7_75t_L g576 ( .A(n_484), .B(n_16), .C(n_17), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_516), .A2(n_382), .B(n_374), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_516), .A2(n_382), .B(n_374), .Y(n_578) );
BUFx2_ASAP7_75t_L g579 ( .A(n_485), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_499), .A2(n_382), .B1(n_374), .B2(n_23), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_515), .A2(n_382), .B(n_102), .Y(n_581) );
NOR3xp33_ASAP7_75t_L g582 ( .A(n_484), .B(n_20), .C(n_22), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_482), .A2(n_25), .B1(n_23), .B2(n_24), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_488), .B(n_487), .Y(n_584) );
OR2x6_ASAP7_75t_L g585 ( .A(n_509), .B(n_24), .Y(n_585) );
NOR2xp33_ASAP7_75t_SL g586 ( .A(n_522), .B(n_27), .Y(n_586) );
INVxp67_ASAP7_75t_L g587 ( .A(n_505), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_473), .B(n_29), .Y(n_588) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_504), .Y(n_589) );
O2A1O1Ixp5_ASAP7_75t_SL g590 ( .A1(n_521), .A2(n_111), .B(n_112), .C(n_109), .Y(n_590) );
INVx3_ASAP7_75t_SL g591 ( .A(n_500), .Y(n_591) );
NOR2xp67_ASAP7_75t_L g592 ( .A(n_501), .B(n_30), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_498), .B(n_31), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_523), .B(n_32), .Y(n_594) );
NAND3xp33_ASAP7_75t_L g595 ( .A(n_506), .B(n_33), .C(n_34), .Y(n_595) );
AND2x2_ASAP7_75t_SL g596 ( .A(n_478), .B(n_34), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_512), .A2(n_35), .B1(n_36), .B2(n_37), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_512), .B(n_35), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_504), .B(n_36), .Y(n_599) );
O2A1O1Ixp33_ASAP7_75t_L g600 ( .A1(n_524), .A2(n_37), .B(n_38), .C(n_39), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_495), .B(n_38), .Y(n_601) );
A2O1A1Ixp33_ASAP7_75t_L g602 ( .A1(n_489), .A2(n_40), .B(n_41), .C(n_43), .Y(n_602) );
NAND3xp33_ASAP7_75t_L g603 ( .A(n_506), .B(n_40), .C(n_44), .Y(n_603) );
AO21x1_ASAP7_75t_L g604 ( .A1(n_469), .A2(n_44), .B(n_45), .Y(n_604) );
BUFx2_ASAP7_75t_L g605 ( .A(n_513), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_521), .A2(n_46), .B1(n_47), .B2(n_49), .Y(n_606) );
INVx3_ASAP7_75t_L g607 ( .A(n_518), .Y(n_607) );
BUFx8_ASAP7_75t_L g608 ( .A(n_518), .Y(n_608) );
INVxp67_ASAP7_75t_L g609 ( .A(n_489), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_468), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_476), .B(n_46), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_465), .B(n_49), .Y(n_612) );
AND2x4_ASAP7_75t_L g613 ( .A(n_480), .B(n_51), .Y(n_613) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_480), .Y(n_614) );
O2A1O1Ixp33_ASAP7_75t_L g615 ( .A1(n_454), .A2(n_52), .B(n_53), .C(n_54), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_475), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_459), .A2(n_53), .B1(n_55), .B2(n_56), .Y(n_617) );
OR2x2_ASAP7_75t_SL g618 ( .A(n_483), .B(n_57), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_480), .A2(n_57), .B1(n_58), .B2(n_59), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_459), .A2(n_59), .B1(n_60), .B2(n_61), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_459), .A2(n_60), .B1(n_61), .B2(n_62), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_459), .A2(n_62), .B1(n_63), .B2(n_64), .Y(n_622) );
AND2x4_ASAP7_75t_L g623 ( .A(n_480), .B(n_63), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_459), .B(n_64), .Y(n_624) );
BUFx6f_ASAP7_75t_L g625 ( .A(n_519), .Y(n_625) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_480), .Y(n_626) );
O2A1O1Ixp33_ASAP7_75t_L g627 ( .A1(n_454), .A2(n_65), .B(n_66), .C(n_67), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_455), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_465), .B(n_67), .Y(n_629) );
NAND2x1_ASAP7_75t_L g630 ( .A(n_480), .B(n_128), .Y(n_630) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_459), .B(n_68), .Y(n_631) );
BUFx3_ASAP7_75t_L g632 ( .A(n_462), .Y(n_632) );
AND2x4_ASAP7_75t_L g633 ( .A(n_480), .B(n_69), .Y(n_633) );
A2O1A1Ixp33_ASAP7_75t_L g634 ( .A1(n_456), .A2(n_70), .B(n_71), .C(n_72), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_613), .A2(n_70), .B1(n_71), .B2(n_72), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_612), .Y(n_636) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_567), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_533), .B(n_73), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_568), .Y(n_639) );
AO31x2_ASAP7_75t_L g640 ( .A1(n_538), .A2(n_75), .A3(n_76), .B(n_78), .Y(n_640) );
OAI22x1_ASAP7_75t_L g641 ( .A1(n_613), .A2(n_75), .B1(n_76), .B2(n_78), .Y(n_641) );
INVx4_ASAP7_75t_L g642 ( .A(n_567), .Y(n_642) );
BUFx2_ASAP7_75t_L g643 ( .A(n_536), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_535), .B(n_79), .Y(n_644) );
OAI21x1_ASAP7_75t_L g645 ( .A1(n_578), .A2(n_167), .B(n_215), .Y(n_645) );
AND2x6_ASAP7_75t_L g646 ( .A(n_623), .B(n_80), .Y(n_646) );
BUFx6f_ASAP7_75t_L g647 ( .A(n_567), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_596), .B(n_81), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_623), .B(n_82), .Y(n_649) );
INVx1_ASAP7_75t_SL g650 ( .A(n_625), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_579), .B(n_83), .Y(n_651) );
BUFx10_ASAP7_75t_L g652 ( .A(n_625), .Y(n_652) );
BUFx2_ASAP7_75t_L g653 ( .A(n_536), .Y(n_653) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_625), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_552), .B(n_84), .Y(n_655) );
INVxp67_ASAP7_75t_SL g656 ( .A(n_633), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_558), .B(n_85), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_629), .Y(n_658) );
NOR2xp67_ASAP7_75t_L g659 ( .A(n_531), .B(n_614), .Y(n_659) );
A2O1A1Ixp33_ASAP7_75t_L g660 ( .A1(n_556), .A2(n_548), .B(n_544), .C(n_532), .Y(n_660) );
NOR2xp67_ASAP7_75t_L g661 ( .A(n_531), .B(n_150), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_626), .B(n_86), .Y(n_662) );
INVx3_ASAP7_75t_SL g663 ( .A(n_632), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_546), .B(n_88), .Y(n_664) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_588), .A2(n_88), .B1(n_89), .B2(n_90), .C(n_91), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_611), .B(n_89), .Y(n_666) );
BUFx2_ASAP7_75t_L g667 ( .A(n_585), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_587), .B(n_90), .Y(n_668) );
AO31x2_ASAP7_75t_L g669 ( .A1(n_604), .A2(n_92), .A3(n_93), .B(n_94), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_628), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_576), .A2(n_94), .B1(n_95), .B2(n_134), .Y(n_671) );
A2O1A1Ixp33_ASAP7_75t_L g672 ( .A1(n_592), .A2(n_95), .B(n_135), .C(n_137), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_541), .Y(n_673) );
BUFx3_ASAP7_75t_L g674 ( .A(n_572), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_616), .Y(n_675) );
AO31x2_ASAP7_75t_L g676 ( .A1(n_555), .A2(n_142), .A3(n_143), .B(n_144), .Y(n_676) );
OAI21x1_ASAP7_75t_L g677 ( .A1(n_590), .A2(n_145), .B(n_147), .Y(n_677) );
OAI21x1_ASAP7_75t_L g678 ( .A1(n_581), .A2(n_149), .B(n_170), .Y(n_678) );
INVx1_ASAP7_75t_SL g679 ( .A(n_585), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_585), .A2(n_179), .B1(n_180), .B2(n_181), .Y(n_680) );
BUFx3_ASAP7_75t_L g681 ( .A(n_591), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_601), .Y(n_682) );
NOR2x1_ASAP7_75t_SL g683 ( .A(n_526), .B(n_191), .Y(n_683) );
INVx2_ASAP7_75t_SL g684 ( .A(n_571), .Y(n_684) );
BUFx10_ASAP7_75t_L g685 ( .A(n_571), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_573), .B(n_192), .Y(n_686) );
NOR3xp33_ASAP7_75t_L g687 ( .A(n_582), .B(n_193), .C(n_194), .Y(n_687) );
AOI221xp5_ASAP7_75t_SL g688 ( .A1(n_609), .A2(n_610), .B1(n_550), .B2(n_553), .C(n_615), .Y(n_688) );
A2O1A1Ixp33_ASAP7_75t_L g689 ( .A1(n_561), .A2(n_627), .B(n_598), .C(n_574), .Y(n_689) );
INVxp67_ASAP7_75t_L g690 ( .A(n_586), .Y(n_690) );
NAND3xp33_ASAP7_75t_L g691 ( .A(n_540), .B(n_580), .C(n_600), .Y(n_691) );
INVxp67_ASAP7_75t_SL g692 ( .A(n_608), .Y(n_692) );
CKINVDCx9p33_ASAP7_75t_R g693 ( .A(n_618), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_549), .B(n_564), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_594), .Y(n_695) );
INVxp67_ASAP7_75t_L g696 ( .A(n_575), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g697 ( .A1(n_584), .A2(n_529), .B(n_557), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_549), .B(n_537), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_607), .A2(n_530), .B1(n_605), .B2(n_620), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_608), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_547), .B(n_563), .Y(n_701) );
AOI21xp5_ASAP7_75t_L g702 ( .A1(n_551), .A2(n_542), .B(n_565), .Y(n_702) );
INVx4_ASAP7_75t_L g703 ( .A(n_589), .Y(n_703) );
OAI21x1_ASAP7_75t_L g704 ( .A1(n_566), .A2(n_562), .B(n_560), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_599), .Y(n_705) );
AO31x2_ASAP7_75t_L g706 ( .A1(n_559), .A2(n_602), .A3(n_583), .B(n_597), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_554), .B(n_593), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_543), .A2(n_570), .B(n_545), .Y(n_708) );
AOI21xp5_ASAP7_75t_SL g709 ( .A1(n_617), .A2(n_622), .B(n_621), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_617), .A2(n_620), .B1(n_622), .B2(n_621), .Y(n_710) );
O2A1O1Ixp33_ASAP7_75t_L g711 ( .A1(n_624), .A2(n_631), .B(n_539), .C(n_595), .Y(n_711) );
A2O1A1Ixp33_ASAP7_75t_L g712 ( .A1(n_606), .A2(n_528), .B(n_525), .C(n_556), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_603), .B(n_570), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_570), .A2(n_466), .B(n_458), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_596), .B(n_476), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_533), .B(n_476), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_596), .B(n_476), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_612), .Y(n_718) );
O2A1O1Ixp33_ASAP7_75t_SL g719 ( .A1(n_630), .A2(n_534), .B(n_555), .C(n_467), .Y(n_719) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_567), .Y(n_720) );
INVx4_ASAP7_75t_L g721 ( .A(n_567), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_596), .B(n_476), .Y(n_722) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_527), .A2(n_466), .B(n_458), .Y(n_723) );
AOI221xp5_ASAP7_75t_L g724 ( .A1(n_588), .A2(n_484), .B1(n_535), .B2(n_440), .C(n_483), .Y(n_724) );
OAI21xp33_ASAP7_75t_L g725 ( .A1(n_612), .A2(n_465), .B(n_459), .Y(n_725) );
INVx3_ASAP7_75t_L g726 ( .A(n_567), .Y(n_726) );
AOI221xp5_ASAP7_75t_L g727 ( .A1(n_588), .A2(n_484), .B1(n_535), .B2(n_440), .C(n_483), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_612), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_612), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_527), .A2(n_466), .B(n_458), .Y(n_730) );
AO31x2_ASAP7_75t_L g731 ( .A1(n_538), .A2(n_467), .A3(n_527), .B(n_569), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_552), .B(n_454), .Y(n_732) );
AO31x2_ASAP7_75t_L g733 ( .A1(n_538), .A2(n_467), .A3(n_527), .B(n_569), .Y(n_733) );
BUFx12f_ASAP7_75t_L g734 ( .A(n_536), .Y(n_734) );
O2A1O1Ixp33_ASAP7_75t_L g735 ( .A1(n_555), .A2(n_528), .B(n_634), .C(n_532), .Y(n_735) );
AO31x2_ASAP7_75t_L g736 ( .A1(n_538), .A2(n_467), .A3(n_527), .B(n_569), .Y(n_736) );
AO31x2_ASAP7_75t_L g737 ( .A1(n_538), .A2(n_467), .A3(n_527), .B(n_569), .Y(n_737) );
AO31x2_ASAP7_75t_L g738 ( .A1(n_538), .A2(n_467), .A3(n_527), .B(n_569), .Y(n_738) );
NOR2xp67_ASAP7_75t_L g739 ( .A(n_531), .B(n_613), .Y(n_739) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_567), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_536), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_552), .B(n_454), .Y(n_742) );
AOI221x1_ASAP7_75t_L g743 ( .A1(n_538), .A2(n_527), .B1(n_569), .B2(n_578), .C(n_577), .Y(n_743) );
OR2x2_ASAP7_75t_L g744 ( .A(n_533), .B(n_409), .Y(n_744) );
OAI21xp5_ASAP7_75t_L g745 ( .A1(n_527), .A2(n_525), .B(n_467), .Y(n_745) );
OAI21xp5_ASAP7_75t_L g746 ( .A1(n_527), .A2(n_525), .B(n_467), .Y(n_746) );
AO32x2_ASAP7_75t_L g747 ( .A1(n_597), .A2(n_583), .A3(n_619), .B1(n_535), .B2(n_526), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_533), .B(n_476), .Y(n_748) );
BUFx2_ASAP7_75t_L g749 ( .A(n_536), .Y(n_749) );
OR2x2_ASAP7_75t_L g750 ( .A(n_533), .B(n_409), .Y(n_750) );
O2A1O1Ixp33_ASAP7_75t_L g751 ( .A1(n_555), .A2(n_528), .B(n_634), .C(n_532), .Y(n_751) );
AOI21xp5_ASAP7_75t_L g752 ( .A1(n_527), .A2(n_466), .B(n_458), .Y(n_752) );
AOI21xp5_ASAP7_75t_L g753 ( .A1(n_527), .A2(n_466), .B(n_458), .Y(n_753) );
O2A1O1Ixp33_ASAP7_75t_SL g754 ( .A1(n_630), .A2(n_534), .B(n_555), .C(n_467), .Y(n_754) );
AO31x2_ASAP7_75t_L g755 ( .A1(n_538), .A2(n_467), .A3(n_527), .B(n_569), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g756 ( .A1(n_527), .A2(n_466), .B(n_458), .Y(n_756) );
AOI221xp5_ASAP7_75t_SL g757 ( .A1(n_538), .A2(n_555), .B1(n_556), .B2(n_532), .C(n_528), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_568), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_533), .B(n_476), .Y(n_759) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_567), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_552), .B(n_454), .Y(n_761) );
O2A1O1Ixp33_ASAP7_75t_SL g762 ( .A1(n_630), .A2(n_534), .B(n_555), .C(n_467), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_639), .Y(n_763) );
NOR2x1_ASAP7_75t_L g764 ( .A(n_741), .B(n_642), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_758), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g766 ( .A1(n_714), .A2(n_730), .B(n_723), .Y(n_766) );
AOI21xp5_ASAP7_75t_L g767 ( .A1(n_752), .A2(n_756), .B(n_753), .Y(n_767) );
NOR2xp33_ASAP7_75t_SL g768 ( .A(n_646), .B(n_739), .Y(n_768) );
AOI21xp5_ASAP7_75t_L g769 ( .A1(n_713), .A2(n_754), .B(n_719), .Y(n_769) );
INVx3_ASAP7_75t_L g770 ( .A(n_647), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_673), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_675), .Y(n_772) );
AO31x2_ASAP7_75t_L g773 ( .A1(n_743), .A2(n_689), .A3(n_708), .B(n_702), .Y(n_773) );
AND2x2_ASAP7_75t_L g774 ( .A(n_715), .B(n_717), .Y(n_774) );
AO31x2_ASAP7_75t_L g775 ( .A1(n_712), .A2(n_699), .A3(n_672), .B(n_660), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_710), .A2(n_656), .B1(n_635), .B2(n_739), .Y(n_776) );
AOI21xp5_ASAP7_75t_L g777 ( .A1(n_762), .A2(n_746), .B(n_745), .Y(n_777) );
INVx3_ASAP7_75t_L g778 ( .A(n_652), .Y(n_778) );
OAI21xp5_ASAP7_75t_L g779 ( .A1(n_688), .A2(n_691), .B(n_697), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_635), .Y(n_780) );
OAI21x1_ASAP7_75t_SL g781 ( .A1(n_683), .A2(n_680), .B(n_710), .Y(n_781) );
AND2x4_ASAP7_75t_L g782 ( .A(n_642), .B(n_721), .Y(n_782) );
A2O1A1Ixp33_ASAP7_75t_L g783 ( .A1(n_735), .A2(n_751), .B(n_725), .C(n_658), .Y(n_783) );
AND2x4_ASAP7_75t_L g784 ( .A(n_721), .B(n_659), .Y(n_784) );
AO21x2_ASAP7_75t_L g785 ( .A1(n_725), .A2(n_677), .B(n_709), .Y(n_785) );
OAI21x1_ASAP7_75t_L g786 ( .A1(n_645), .A2(n_704), .B(n_678), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_722), .B(n_732), .Y(n_787) );
BUFx6f_ASAP7_75t_L g788 ( .A(n_652), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_641), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_705), .B(n_636), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g791 ( .A(n_696), .B(n_744), .Y(n_791) );
INVx3_ASAP7_75t_L g792 ( .A(n_726), .Y(n_792) );
AND2x2_ASAP7_75t_L g793 ( .A(n_742), .B(n_761), .Y(n_793) );
BUFx3_ASAP7_75t_L g794 ( .A(n_663), .Y(n_794) );
BUFx8_ASAP7_75t_L g795 ( .A(n_734), .Y(n_795) );
BUFx6f_ASAP7_75t_L g796 ( .A(n_726), .Y(n_796) );
A2O1A1Ixp33_ASAP7_75t_L g797 ( .A1(n_718), .A2(n_728), .B(n_729), .C(n_711), .Y(n_797) );
BUFx2_ASAP7_75t_L g798 ( .A(n_637), .Y(n_798) );
INVx2_ASAP7_75t_SL g799 ( .A(n_650), .Y(n_799) );
HB1xp67_ASAP7_75t_L g800 ( .A(n_650), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_670), .Y(n_801) );
AND2x2_ASAP7_75t_L g802 ( .A(n_692), .B(n_716), .Y(n_802) );
OAI21xp5_ASAP7_75t_L g803 ( .A1(n_688), .A2(n_691), .B(n_707), .Y(n_803) );
BUFx2_ASAP7_75t_SL g804 ( .A(n_700), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_695), .B(n_724), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_748), .B(n_759), .Y(n_806) );
OR2x2_ASAP7_75t_L g807 ( .A(n_750), .B(n_654), .Y(n_807) );
AOI22xp5_ASAP7_75t_L g808 ( .A1(n_727), .A2(n_644), .B1(n_698), .B2(n_648), .Y(n_808) );
NAND2x1p5_ASAP7_75t_L g809 ( .A(n_659), .B(n_679), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g810 ( .A(n_684), .B(n_694), .Y(n_810) );
NAND2x1p5_ASAP7_75t_L g811 ( .A(n_679), .B(n_667), .Y(n_811) );
AND2x2_ASAP7_75t_L g812 ( .A(n_649), .B(n_720), .Y(n_812) );
NAND2x1p5_ASAP7_75t_L g813 ( .A(n_674), .B(n_681), .Y(n_813) );
BUFx12f_ASAP7_75t_L g814 ( .A(n_643), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_757), .B(n_682), .Y(n_815) );
OAI21x1_ASAP7_75t_SL g816 ( .A1(n_703), .A2(n_657), .B(n_671), .Y(n_816) );
INVx2_ASAP7_75t_L g817 ( .A(n_640), .Y(n_817) );
HB1xp67_ASAP7_75t_L g818 ( .A(n_760), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_662), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_655), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_693), .Y(n_821) );
OAI21x1_ASAP7_75t_SL g822 ( .A1(n_671), .A2(n_686), .B(n_666), .Y(n_822) );
AO31x2_ASAP7_75t_L g823 ( .A1(n_731), .A2(n_737), .A3(n_733), .B(n_755), .Y(n_823) );
AND2x2_ASAP7_75t_L g824 ( .A(n_740), .B(n_685), .Y(n_824) );
OAI21xp5_ASAP7_75t_L g825 ( .A1(n_687), .A2(n_690), .B(n_661), .Y(n_825) );
BUFx2_ASAP7_75t_SL g826 ( .A(n_653), .Y(n_826) );
BUFx2_ASAP7_75t_L g827 ( .A(n_749), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_706), .B(n_701), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_706), .B(n_736), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_706), .B(n_731), .Y(n_830) );
AOI21xp5_ASAP7_75t_L g831 ( .A1(n_665), .A2(n_638), .B(n_664), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_731), .B(n_736), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_669), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_669), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_669), .Y(n_835) );
AOI21xp5_ASAP7_75t_L g836 ( .A1(n_737), .A2(n_738), .B(n_755), .Y(n_836) );
AOI21xp5_ASAP7_75t_SL g837 ( .A1(n_651), .A2(n_668), .B(n_747), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_685), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_676), .Y(n_839) );
AND2x2_ASAP7_75t_L g840 ( .A(n_715), .B(n_476), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_639), .Y(n_841) );
NAND2x1p5_ASAP7_75t_L g842 ( .A(n_739), .B(n_531), .Y(n_842) );
NOR2x1_ASAP7_75t_L g843 ( .A(n_741), .B(n_642), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_639), .Y(n_844) );
INVxp67_ASAP7_75t_L g845 ( .A(n_637), .Y(n_845) );
CKINVDCx16_ASAP7_75t_R g846 ( .A(n_734), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_639), .Y(n_847) );
OR2x2_ASAP7_75t_L g848 ( .A(n_650), .B(n_476), .Y(n_848) );
AND2x4_ASAP7_75t_L g849 ( .A(n_739), .B(n_531), .Y(n_849) );
INVx6_ASAP7_75t_L g850 ( .A(n_652), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_639), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_639), .Y(n_852) );
OAI22xp5_ASAP7_75t_L g853 ( .A1(n_710), .A2(n_656), .B1(n_635), .B2(n_613), .Y(n_853) );
INVx2_ASAP7_75t_SL g854 ( .A(n_652), .Y(n_854) );
AOI221xp5_ASAP7_75t_L g855 ( .A1(n_724), .A2(n_484), .B1(n_727), .B2(n_588), .C(n_576), .Y(n_855) );
NOR2xp33_ASAP7_75t_L g856 ( .A(n_696), .B(n_484), .Y(n_856) );
OR2x6_ASAP7_75t_L g857 ( .A(n_739), .B(n_531), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_639), .Y(n_858) );
INVx3_ASAP7_75t_L g859 ( .A(n_647), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_639), .Y(n_860) );
NOR2xp33_ASAP7_75t_SL g861 ( .A(n_646), .B(n_613), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_639), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_639), .Y(n_863) );
AOI21xp5_ASAP7_75t_L g864 ( .A1(n_714), .A2(n_730), .B(n_723), .Y(n_864) );
AOI21xp5_ASAP7_75t_L g865 ( .A1(n_714), .A2(n_730), .B(n_723), .Y(n_865) );
AND2x4_ASAP7_75t_L g866 ( .A(n_739), .B(n_531), .Y(n_866) );
CKINVDCx20_ASAP7_75t_R g867 ( .A(n_741), .Y(n_867) );
BUFx12f_ASAP7_75t_L g868 ( .A(n_734), .Y(n_868) );
OAI21xp5_ASAP7_75t_L g869 ( .A1(n_723), .A2(n_752), .B(n_730), .Y(n_869) );
INVx4_ASAP7_75t_L g870 ( .A(n_857), .Y(n_870) );
INVx3_ASAP7_75t_L g871 ( .A(n_842), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_771), .Y(n_872) );
OR2x6_ASAP7_75t_L g873 ( .A(n_853), .B(n_776), .Y(n_873) );
OR2x2_ASAP7_75t_L g874 ( .A(n_780), .B(n_828), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_815), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_793), .B(n_805), .Y(n_876) );
BUFx4f_ASAP7_75t_SL g877 ( .A(n_795), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_805), .B(n_855), .Y(n_878) );
BUFx2_ASAP7_75t_SL g879 ( .A(n_849), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_772), .Y(n_880) );
AO21x2_ASAP7_75t_L g881 ( .A1(n_779), .A2(n_864), .B(n_766), .Y(n_881) );
INVx2_ASAP7_75t_SL g882 ( .A(n_788), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_817), .Y(n_883) );
AO21x2_ASAP7_75t_L g884 ( .A1(n_779), .A2(n_865), .B(n_777), .Y(n_884) );
AND2x2_ASAP7_75t_L g885 ( .A(n_787), .B(n_861), .Y(n_885) );
BUFx2_ASAP7_75t_L g886 ( .A(n_809), .Y(n_886) );
BUFx3_ASAP7_75t_L g887 ( .A(n_794), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_855), .B(n_808), .Y(n_888) );
BUFx3_ASAP7_75t_L g889 ( .A(n_788), .Y(n_889) );
INVx1_ASAP7_75t_SL g890 ( .A(n_850), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_833), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_834), .Y(n_892) );
HB1xp67_ASAP7_75t_L g893 ( .A(n_800), .Y(n_893) );
OA21x2_ASAP7_75t_L g894 ( .A1(n_767), .A2(n_869), .B(n_777), .Y(n_894) );
AO21x2_ASAP7_75t_L g895 ( .A1(n_769), .A2(n_767), .B(n_869), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_808), .B(n_856), .Y(n_896) );
AND2x2_ASAP7_75t_L g897 ( .A(n_763), .B(n_765), .Y(n_897) );
INVx2_ASAP7_75t_SL g898 ( .A(n_850), .Y(n_898) );
AND2x2_ASAP7_75t_L g899 ( .A(n_841), .B(n_844), .Y(n_899) );
BUFx3_ASAP7_75t_L g900 ( .A(n_782), .Y(n_900) );
BUFx2_ASAP7_75t_L g901 ( .A(n_809), .Y(n_901) );
HB1xp67_ASAP7_75t_SL g902 ( .A(n_795), .Y(n_902) );
HB1xp67_ASAP7_75t_L g903 ( .A(n_818), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_835), .Y(n_904) );
HB1xp67_ASAP7_75t_L g905 ( .A(n_798), .Y(n_905) );
AND2x2_ASAP7_75t_L g906 ( .A(n_847), .B(n_851), .Y(n_906) );
AO21x2_ASAP7_75t_L g907 ( .A1(n_803), .A2(n_836), .B(n_839), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_852), .Y(n_908) );
HB1xp67_ASAP7_75t_L g909 ( .A(n_848), .Y(n_909) );
OR2x6_ASAP7_75t_L g910 ( .A(n_781), .B(n_816), .Y(n_910) );
OR2x2_ASAP7_75t_L g911 ( .A(n_829), .B(n_830), .Y(n_911) );
OR2x6_ASAP7_75t_L g912 ( .A(n_842), .B(n_837), .Y(n_912) );
HB1xp67_ASAP7_75t_L g913 ( .A(n_812), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_829), .Y(n_914) );
AND2x2_ASAP7_75t_L g915 ( .A(n_858), .B(n_860), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_862), .Y(n_916) );
INVx2_ASAP7_75t_L g917 ( .A(n_773), .Y(n_917) );
INVx2_ASAP7_75t_SL g918 ( .A(n_764), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_863), .Y(n_919) );
INVx2_ASAP7_75t_SL g920 ( .A(n_843), .Y(n_920) );
INVx2_ASAP7_75t_L g921 ( .A(n_773), .Y(n_921) );
INVx4_ASAP7_75t_L g922 ( .A(n_784), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_789), .A2(n_831), .B1(n_822), .B2(n_791), .Y(n_923) );
INVx2_ASAP7_75t_SL g924 ( .A(n_778), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_830), .Y(n_925) );
OR2x2_ASAP7_75t_L g926 ( .A(n_807), .B(n_823), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_806), .B(n_790), .Y(n_927) );
INVx2_ASAP7_75t_SL g928 ( .A(n_778), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_832), .Y(n_929) );
BUFx3_ASAP7_75t_L g930 ( .A(n_813), .Y(n_930) );
INVx2_ASAP7_75t_L g931 ( .A(n_823), .Y(n_931) );
OAI22xp5_ASAP7_75t_L g932 ( .A1(n_797), .A2(n_831), .B1(n_821), .B2(n_820), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_823), .Y(n_933) );
HB1xp67_ASAP7_75t_L g934 ( .A(n_845), .Y(n_934) );
AND2x2_ASAP7_75t_L g935 ( .A(n_774), .B(n_801), .Y(n_935) );
AND2x2_ASAP7_75t_L g936 ( .A(n_873), .B(n_775), .Y(n_936) );
AND2x2_ASAP7_75t_L g937 ( .A(n_873), .B(n_775), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_891), .Y(n_938) );
OR2x2_ASAP7_75t_L g939 ( .A(n_926), .B(n_874), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_891), .Y(n_940) );
HB1xp67_ASAP7_75t_L g941 ( .A(n_903), .Y(n_941) );
AND2x4_ASAP7_75t_L g942 ( .A(n_910), .B(n_785), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_892), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_892), .Y(n_944) );
INVx1_ASAP7_75t_L g945 ( .A(n_904), .Y(n_945) );
AND2x2_ASAP7_75t_L g946 ( .A(n_873), .B(n_783), .Y(n_946) );
INVx1_ASAP7_75t_L g947 ( .A(n_904), .Y(n_947) );
HB1xp67_ASAP7_75t_L g948 ( .A(n_905), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_873), .A2(n_840), .B1(n_802), .B2(n_819), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_933), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_933), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_896), .B(n_799), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_929), .Y(n_953) );
INVx1_ASAP7_75t_SL g954 ( .A(n_887), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_914), .Y(n_955) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_876), .B(n_888), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_935), .B(n_770), .Y(n_957) );
INVx1_ASAP7_75t_L g958 ( .A(n_914), .Y(n_958) );
INVx4_ASAP7_75t_R g959 ( .A(n_902), .Y(n_959) );
BUFx2_ASAP7_75t_L g960 ( .A(n_886), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_925), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_925), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_927), .B(n_811), .Y(n_963) );
BUFx3_ASAP7_75t_L g964 ( .A(n_900), .Y(n_964) );
AND2x2_ASAP7_75t_L g965 ( .A(n_935), .B(n_859), .Y(n_965) );
INVx4_ASAP7_75t_L g966 ( .A(n_870), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_883), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g968 ( .A(n_878), .B(n_810), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_885), .A2(n_827), .B1(n_768), .B2(n_826), .Y(n_969) );
INVxp67_ASAP7_75t_SL g970 ( .A(n_893), .Y(n_970) );
AND2x2_ASAP7_75t_L g971 ( .A(n_875), .B(n_825), .Y(n_971) );
INVx2_ASAP7_75t_SL g972 ( .A(n_922), .Y(n_972) );
AND2x4_ASAP7_75t_L g973 ( .A(n_912), .B(n_786), .Y(n_973) );
INVx1_ASAP7_75t_SL g974 ( .A(n_887), .Y(n_974) );
BUFx3_ASAP7_75t_L g975 ( .A(n_922), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_897), .B(n_796), .Y(n_976) );
OAI22xp5_ASAP7_75t_L g977 ( .A1(n_879), .A2(n_866), .B1(n_867), .B2(n_813), .Y(n_977) );
BUFx2_ASAP7_75t_L g978 ( .A(n_901), .Y(n_978) );
NOR2x1p5_ASAP7_75t_L g979 ( .A(n_870), .B(n_868), .Y(n_979) );
NOR2x1_ASAP7_75t_L g980 ( .A(n_870), .B(n_792), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_899), .B(n_824), .Y(n_981) );
AND2x2_ASAP7_75t_L g982 ( .A(n_936), .B(n_931), .Y(n_982) );
BUFx2_ASAP7_75t_L g983 ( .A(n_960), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_936), .B(n_931), .Y(n_984) );
AND2x2_ASAP7_75t_L g985 ( .A(n_937), .B(n_917), .Y(n_985) );
AND2x2_ASAP7_75t_L g986 ( .A(n_937), .B(n_917), .Y(n_986) );
OR2x2_ASAP7_75t_L g987 ( .A(n_939), .B(n_911), .Y(n_987) );
NOR2x1_ASAP7_75t_L g988 ( .A(n_975), .B(n_912), .Y(n_988) );
HB1xp67_ASAP7_75t_L g989 ( .A(n_941), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_956), .B(n_872), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_950), .Y(n_991) );
AND2x2_ASAP7_75t_L g992 ( .A(n_946), .B(n_921), .Y(n_992) );
HB1xp67_ASAP7_75t_L g993 ( .A(n_948), .Y(n_993) );
NOR2xp33_ASAP7_75t_L g994 ( .A(n_954), .B(n_877), .Y(n_994) );
NAND2xp5_ASAP7_75t_L g995 ( .A(n_957), .B(n_913), .Y(n_995) );
OR2x2_ASAP7_75t_L g996 ( .A(n_939), .B(n_911), .Y(n_996) );
NOR2xp33_ASAP7_75t_L g997 ( .A(n_974), .B(n_814), .Y(n_997) );
AND2x4_ASAP7_75t_L g998 ( .A(n_973), .B(n_881), .Y(n_998) );
AND2x2_ASAP7_75t_L g999 ( .A(n_971), .B(n_907), .Y(n_999) );
INVx4_ASAP7_75t_L g1000 ( .A(n_966), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_971), .B(n_907), .Y(n_1001) );
HB1xp67_ASAP7_75t_L g1002 ( .A(n_970), .Y(n_1002) );
NAND2xp5_ASAP7_75t_L g1003 ( .A(n_957), .B(n_909), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_965), .B(n_906), .Y(n_1004) );
AND2x4_ASAP7_75t_L g1005 ( .A(n_973), .B(n_884), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_951), .Y(n_1006) );
NOR2xp33_ASAP7_75t_L g1007 ( .A(n_981), .B(n_846), .Y(n_1007) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_965), .B(n_906), .Y(n_1008) );
AND2x4_ASAP7_75t_L g1009 ( .A(n_973), .B(n_884), .Y(n_1009) );
HB1xp67_ASAP7_75t_L g1010 ( .A(n_960), .Y(n_1010) );
INVxp67_ASAP7_75t_SL g1011 ( .A(n_964), .Y(n_1011) );
AOI33xp33_ASAP7_75t_L g1012 ( .A1(n_949), .A2(n_923), .A3(n_919), .B1(n_916), .B2(n_908), .B3(n_880), .Y(n_1012) );
AND2x4_ASAP7_75t_L g1013 ( .A(n_973), .B(n_884), .Y(n_1013) );
AND2x2_ASAP7_75t_L g1014 ( .A(n_938), .B(n_907), .Y(n_1014) );
AND2x2_ASAP7_75t_L g1015 ( .A(n_938), .B(n_894), .Y(n_1015) );
INVx3_ASAP7_75t_L g1016 ( .A(n_966), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_940), .B(n_894), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_951), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_940), .B(n_943), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_943), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_944), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_952), .B(n_915), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_944), .Y(n_1023) );
AND2x2_ASAP7_75t_L g1024 ( .A(n_945), .B(n_894), .Y(n_1024) );
INVxp67_ASAP7_75t_SL g1025 ( .A(n_964), .Y(n_1025) );
NOR2x1_ASAP7_75t_L g1026 ( .A(n_975), .B(n_912), .Y(n_1026) );
INVx3_ASAP7_75t_L g1027 ( .A(n_966), .Y(n_1027) );
HB1xp67_ASAP7_75t_L g1028 ( .A(n_978), .Y(n_1028) );
AND2x4_ASAP7_75t_L g1029 ( .A(n_1005), .B(n_1009), .Y(n_1029) );
AND2x4_ASAP7_75t_L g1030 ( .A(n_1005), .B(n_942), .Y(n_1030) );
OR2x2_ASAP7_75t_L g1031 ( .A(n_987), .B(n_953), .Y(n_1031) );
NAND2xp33_ASAP7_75t_L g1032 ( .A(n_988), .B(n_979), .Y(n_1032) );
INVxp67_ASAP7_75t_SL g1033 ( .A(n_1002), .Y(n_1033) );
INVx2_ASAP7_75t_L g1034 ( .A(n_991), .Y(n_1034) );
INVx1_ASAP7_75t_L g1035 ( .A(n_1020), .Y(n_1035) );
NAND2xp5_ASAP7_75t_L g1036 ( .A(n_989), .B(n_955), .Y(n_1036) );
NAND2x1p5_ASAP7_75t_L g1037 ( .A(n_1000), .B(n_966), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_992), .B(n_999), .Y(n_1038) );
NAND2xp5_ASAP7_75t_L g1039 ( .A(n_993), .B(n_955), .Y(n_1039) );
INVx2_ASAP7_75t_SL g1040 ( .A(n_1000), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1020), .Y(n_1041) );
HB1xp67_ASAP7_75t_L g1042 ( .A(n_983), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_1022), .B(n_958), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_999), .B(n_947), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_1001), .B(n_958), .Y(n_1045) );
BUFx2_ASAP7_75t_L g1046 ( .A(n_1000), .Y(n_1046) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_1019), .B(n_961), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1021), .Y(n_1048) );
OR2x2_ASAP7_75t_L g1049 ( .A(n_987), .B(n_961), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_1001), .B(n_962), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1023), .Y(n_1051) );
AND2x4_ASAP7_75t_L g1052 ( .A(n_1005), .B(n_942), .Y(n_1052) );
AOI22xp5_ASAP7_75t_L g1053 ( .A1(n_1000), .A2(n_977), .B1(n_932), .B2(n_885), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_1019), .B(n_962), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_982), .B(n_895), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1023), .Y(n_1056) );
BUFx2_ASAP7_75t_L g1057 ( .A(n_1011), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_982), .B(n_895), .Y(n_1058) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_1004), .B(n_976), .Y(n_1059) );
INVxp33_ASAP7_75t_L g1060 ( .A(n_994), .Y(n_1060) );
OR2x2_ASAP7_75t_L g1061 ( .A(n_996), .B(n_967), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_984), .B(n_895), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_1008), .B(n_976), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1006), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1018), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1018), .Y(n_1066) );
NAND2xp5_ASAP7_75t_L g1067 ( .A(n_1044), .B(n_1015), .Y(n_1067) );
NAND2xp5_ASAP7_75t_L g1068 ( .A(n_1044), .B(n_1015), .Y(n_1068) );
INVx1_ASAP7_75t_L g1069 ( .A(n_1036), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_1045), .B(n_1017), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1039), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1033), .Y(n_1072) );
OR2x2_ASAP7_75t_L g1073 ( .A(n_1038), .B(n_996), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1061), .Y(n_1074) );
NOR2xp33_ASAP7_75t_L g1075 ( .A(n_1060), .B(n_1007), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1038), .B(n_985), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_1055), .B(n_985), .Y(n_1077) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_1055), .B(n_986), .Y(n_1078) );
NAND2xp5_ASAP7_75t_L g1079 ( .A(n_1045), .B(n_1017), .Y(n_1079) );
INVx2_ASAP7_75t_L g1080 ( .A(n_1034), .Y(n_1080) );
INVx2_ASAP7_75t_L g1081 ( .A(n_1034), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1061), .Y(n_1082) );
NAND2xp5_ASAP7_75t_L g1083 ( .A(n_1050), .B(n_1024), .Y(n_1083) );
NAND2xp5_ASAP7_75t_L g1084 ( .A(n_1050), .B(n_1024), .Y(n_1084) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1035), .Y(n_1085) );
NOR2xp33_ASAP7_75t_L g1086 ( .A(n_1043), .B(n_1031), .Y(n_1086) );
NOR2xp33_ASAP7_75t_L g1087 ( .A(n_1031), .B(n_990), .Y(n_1087) );
AOI22xp5_ASAP7_75t_L g1088 ( .A1(n_1053), .A2(n_968), .B1(n_986), .B2(n_979), .Y(n_1088) );
INVxp33_ASAP7_75t_L g1089 ( .A(n_1037), .Y(n_1089) );
NOR2x1_ASAP7_75t_L g1090 ( .A(n_1032), .B(n_988), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_1047), .B(n_1014), .Y(n_1091) );
NAND3xp33_ASAP7_75t_L g1092 ( .A(n_1042), .B(n_1028), .C(n_1010), .Y(n_1092) );
AND2x4_ASAP7_75t_L g1093 ( .A(n_1029), .B(n_998), .Y(n_1093) );
INVx1_ASAP7_75t_SL g1094 ( .A(n_1046), .Y(n_1094) );
NAND2xp5_ASAP7_75t_L g1095 ( .A(n_1054), .B(n_1014), .Y(n_1095) );
INVx1_ASAP7_75t_SL g1096 ( .A(n_1046), .Y(n_1096) );
AND2x4_ASAP7_75t_L g1097 ( .A(n_1029), .B(n_998), .Y(n_1097) );
AND2x4_ASAP7_75t_L g1098 ( .A(n_1029), .B(n_998), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_1058), .B(n_1005), .Y(n_1099) );
INVx1_ASAP7_75t_L g1100 ( .A(n_1035), .Y(n_1100) );
AOI21xp33_ASAP7_75t_SL g1101 ( .A1(n_1037), .A2(n_997), .B(n_959), .Y(n_1101) );
OAI22xp33_ASAP7_75t_L g1102 ( .A1(n_1089), .A2(n_1040), .B1(n_1037), .B2(n_1053), .Y(n_1102) );
INVx2_ASAP7_75t_L g1103 ( .A(n_1080), .Y(n_1103) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1081), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1081), .Y(n_1105) );
AOI211xp5_ASAP7_75t_L g1106 ( .A1(n_1101), .A2(n_1040), .B(n_1057), .C(n_975), .Y(n_1106) );
AOI221x1_ASAP7_75t_L g1107 ( .A1(n_1092), .A2(n_1027), .B1(n_1016), .B2(n_1064), .C(n_1056), .Y(n_1107) );
NOR3xp33_ASAP7_75t_SL g1108 ( .A(n_1075), .B(n_959), .C(n_1003), .Y(n_1108) );
INVx1_ASAP7_75t_SL g1109 ( .A(n_1094), .Y(n_1109) );
INVx1_ASAP7_75t_SL g1110 ( .A(n_1096), .Y(n_1110) );
OAI21xp5_ASAP7_75t_L g1111 ( .A1(n_1090), .A2(n_1026), .B(n_1057), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_1099), .B(n_1058), .Y(n_1112) );
NOR2xp33_ASAP7_75t_L g1113 ( .A(n_1069), .B(n_1071), .Y(n_1113) );
INVx2_ASAP7_75t_SL g1114 ( .A(n_1093), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_1099), .B(n_1062), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1085), .Y(n_1116) );
OAI21xp5_ASAP7_75t_L g1117 ( .A1(n_1089), .A2(n_1026), .B(n_1016), .Y(n_1117) );
NAND2xp5_ASAP7_75t_SL g1118 ( .A(n_1088), .B(n_1016), .Y(n_1118) );
INVx2_ASAP7_75t_L g1119 ( .A(n_1100), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1074), .Y(n_1120) );
AOI331xp33_ASAP7_75t_L g1121 ( .A1(n_1075), .A2(n_969), .A3(n_1065), .B1(n_1064), .B2(n_1066), .B3(n_1051), .C1(n_1048), .Y(n_1121) );
NAND2xp5_ASAP7_75t_L g1122 ( .A(n_1086), .B(n_1062), .Y(n_1122) );
OAI21xp33_ASAP7_75t_L g1123 ( .A1(n_1072), .A2(n_1012), .B(n_1049), .Y(n_1123) );
INVx2_ASAP7_75t_L g1124 ( .A(n_1093), .Y(n_1124) );
OR2x2_ASAP7_75t_L g1125 ( .A(n_1122), .B(n_1073), .Y(n_1125) );
OAI221xp5_ASAP7_75t_L g1126 ( .A1(n_1123), .A2(n_1106), .B1(n_1111), .B2(n_1117), .C(n_1108), .Y(n_1126) );
OAI21xp33_ASAP7_75t_L g1127 ( .A1(n_1123), .A2(n_1087), .B(n_1086), .Y(n_1127) );
INVx2_ASAP7_75t_L g1128 ( .A(n_1103), .Y(n_1128) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1116), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_1112), .B(n_1077), .Y(n_1130) );
AOI222xp33_ASAP7_75t_L g1131 ( .A1(n_1113), .A2(n_1087), .B1(n_1082), .B2(n_1077), .C1(n_1078), .C2(n_995), .Y(n_1131) );
AOI21xp5_ASAP7_75t_L g1132 ( .A1(n_1106), .A2(n_1097), .B(n_1093), .Y(n_1132) );
NOR2x1_ASAP7_75t_L g1133 ( .A(n_1102), .B(n_1027), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1116), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g1135 ( .A1(n_1118), .A2(n_1013), .B1(n_1009), .B2(n_998), .Y(n_1135) );
A2O1A1Ixp33_ASAP7_75t_SL g1136 ( .A1(n_1120), .A2(n_838), .B(n_792), .C(n_871), .Y(n_1136) );
O2A1O1Ixp33_ASAP7_75t_L g1137 ( .A1(n_1109), .A2(n_918), .B(n_920), .C(n_934), .Y(n_1137) );
OAI31xp33_ASAP7_75t_L g1138 ( .A1(n_1110), .A2(n_1098), .A3(n_1097), .B(n_1029), .Y(n_1138) );
INVx2_ASAP7_75t_L g1139 ( .A(n_1103), .Y(n_1139) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1120), .Y(n_1140) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1119), .Y(n_1141) );
AOI211xp5_ASAP7_75t_L g1142 ( .A1(n_1114), .A2(n_1098), .B(n_1097), .C(n_1052), .Y(n_1142) );
OAI221xp5_ASAP7_75t_L g1143 ( .A1(n_1114), .A2(n_1095), .B1(n_1091), .B2(n_1049), .C(n_1084), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_1121), .B(n_1112), .Y(n_1144) );
OAI21xp5_ASAP7_75t_SL g1145 ( .A1(n_1107), .A2(n_1027), .B(n_1098), .Y(n_1145) );
AOI221xp5_ASAP7_75t_L g1146 ( .A1(n_1115), .A2(n_1078), .B1(n_1083), .B2(n_1079), .C(n_1067), .Y(n_1146) );
OAI21xp33_ASAP7_75t_L g1147 ( .A1(n_1124), .A2(n_1070), .B(n_1068), .Y(n_1147) );
NAND2xp5_ASAP7_75t_L g1148 ( .A(n_1115), .B(n_1076), .Y(n_1148) );
NAND4xp25_ASAP7_75t_L g1149 ( .A(n_1107), .B(n_963), .C(n_983), .D(n_1052), .Y(n_1149) );
AOI211xp5_ASAP7_75t_L g1150 ( .A1(n_1124), .A2(n_1030), .B(n_1052), .C(n_1009), .Y(n_1150) );
OAI211xp5_ASAP7_75t_L g1151 ( .A1(n_1124), .A2(n_922), .B(n_1025), .C(n_972), .Y(n_1151) );
AOI221xp5_ASAP7_75t_L g1152 ( .A1(n_1119), .A2(n_1063), .B1(n_1059), .B2(n_1052), .C(n_1030), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1153 ( .A(n_1119), .B(n_1041), .Y(n_1153) );
NAND4xp25_ASAP7_75t_L g1154 ( .A(n_1138), .B(n_1126), .C(n_1144), .D(n_1142), .Y(n_1154) );
NAND5xp2_ASAP7_75t_L g1155 ( .A(n_1145), .B(n_1150), .C(n_1137), .D(n_1132), .E(n_1135), .Y(n_1155) );
NAND3xp33_ASAP7_75t_L g1156 ( .A(n_1133), .B(n_1149), .C(n_1135), .Y(n_1156) );
NAND2xp5_ASAP7_75t_SL g1157 ( .A(n_1151), .B(n_1127), .Y(n_1157) );
NOR3xp33_ASAP7_75t_L g1158 ( .A(n_1136), .B(n_890), .C(n_898), .Y(n_1158) );
AOI21xp5_ASAP7_75t_L g1159 ( .A1(n_1136), .A2(n_1131), .B(n_1143), .Y(n_1159) );
AOI221xp5_ASAP7_75t_L g1160 ( .A1(n_1152), .A2(n_1146), .B1(n_1147), .B2(n_1140), .C(n_1129), .Y(n_1160) );
NAND2xp5_ASAP7_75t_L g1161 ( .A(n_1130), .B(n_1134), .Y(n_1161) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1161), .Y(n_1162) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1157), .Y(n_1163) );
AND2x4_ASAP7_75t_L g1164 ( .A(n_1158), .B(n_1130), .Y(n_1164) );
OA22x2_ASAP7_75t_L g1165 ( .A1(n_1154), .A2(n_804), .B1(n_1139), .B2(n_1128), .Y(n_1165) );
NAND2xp5_ASAP7_75t_SL g1166 ( .A(n_1156), .B(n_1128), .Y(n_1166) );
NAND2xp5_ASAP7_75t_L g1167 ( .A(n_1159), .B(n_1125), .Y(n_1167) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1163), .Y(n_1168) );
NAND2xp5_ASAP7_75t_L g1169 ( .A(n_1167), .B(n_1160), .Y(n_1169) );
AND2x4_ASAP7_75t_L g1170 ( .A(n_1162), .B(n_1148), .Y(n_1170) );
NAND3x1_ASAP7_75t_L g1171 ( .A(n_1165), .B(n_1155), .C(n_871), .Y(n_1171) );
NOR3xp33_ASAP7_75t_L g1172 ( .A(n_1166), .B(n_898), .C(n_854), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1168), .Y(n_1173) );
INVx1_ASAP7_75t_SL g1174 ( .A(n_1170), .Y(n_1174) );
INVx2_ASAP7_75t_SL g1175 ( .A(n_1169), .Y(n_1175) );
XNOR2xp5_ASAP7_75t_L g1176 ( .A(n_1171), .B(n_1164), .Y(n_1176) );
INVx2_ASAP7_75t_L g1177 ( .A(n_1174), .Y(n_1177) );
AO22x1_ASAP7_75t_L g1178 ( .A1(n_1175), .A2(n_1172), .B1(n_1164), .B2(n_930), .Y(n_1178) );
OAI22xp5_ASAP7_75t_L g1179 ( .A1(n_1177), .A2(n_1176), .B1(n_1173), .B2(n_1139), .Y(n_1179) );
HB1xp67_ASAP7_75t_L g1180 ( .A(n_1178), .Y(n_1180) );
NAND3xp33_ASAP7_75t_L g1181 ( .A(n_1179), .B(n_1141), .C(n_889), .Y(n_1181) );
AOI22xp33_ASAP7_75t_L g1182 ( .A1(n_1180), .A2(n_1153), .B1(n_1105), .B2(n_1104), .Y(n_1182) );
OA21x2_ASAP7_75t_L g1183 ( .A1(n_1181), .A2(n_928), .B(n_924), .Y(n_1183) );
OAI21x1_ASAP7_75t_L g1184 ( .A1(n_1182), .A2(n_871), .B(n_980), .Y(n_1184) );
UNKNOWN g1185 ( );
AOI21xp5_ASAP7_75t_L g1186 ( .A1(n_1185), .A2(n_1184), .B(n_882), .Y(n_1186) );
endmodule