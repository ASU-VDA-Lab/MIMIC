module fake_jpeg_15551_n_349 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_349);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_349;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_6),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_36),
.B(n_40),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_L g45 ( 
.A1(n_18),
.A2(n_0),
.B(n_1),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_18),
.B(n_27),
.C(n_32),
.Y(n_53)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_16),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_47),
.B(n_48),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_23),
.B1(n_20),
.B2(n_31),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_56),
.B1(n_64),
.B2(n_67),
.Y(n_83)
);

OR2x2_ASAP7_75t_SL g77 ( 
.A(n_53),
.B(n_45),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_23),
.B1(n_20),
.B2(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_26),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_48),
.Y(n_97)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_23),
.B1(n_20),
.B2(n_31),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_38),
.B1(n_40),
.B2(n_49),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_65),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_78)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_29),
.B1(n_27),
.B2(n_30),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_38),
.A2(n_29),
.B1(n_27),
.B2(n_30),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_68),
.A2(n_33),
.B1(n_26),
.B2(n_25),
.Y(n_93)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_39),
.Y(n_84)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVxp33_ASAP7_75t_SL g75 ( 
.A(n_58),
.Y(n_75)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_74),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_76),
.B(n_92),
.Y(n_128)
);

NOR2xp67_ASAP7_75t_R g126 ( 
.A(n_77),
.B(n_100),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_78),
.A2(n_93),
.B1(n_102),
.B2(n_32),
.Y(n_120)
);

AOI22x1_ASAP7_75t_L g80 ( 
.A1(n_53),
.A2(n_49),
.B1(n_43),
.B2(n_40),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_80),
.A2(n_72),
.B1(n_63),
.B2(n_73),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_53),
.A2(n_29),
.B1(n_25),
.B2(n_26),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

AO22x1_ASAP7_75t_SL g88 ( 
.A1(n_65),
.A2(n_49),
.B1(n_43),
.B2(n_42),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_88),
.A2(n_95),
.B1(n_104),
.B2(n_110),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_74),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_94),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_52),
.A2(n_43),
.B1(n_25),
.B2(n_33),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

BUFx24_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

AOI21xp33_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_108),
.B(n_21),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_48),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_107),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_61),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_99),
.B(n_101),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_70),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_55),
.B(n_47),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_62),
.A2(n_47),
.B1(n_36),
.B2(n_32),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

FAx1_ASAP7_75t_SL g112 ( 
.A(n_103),
.B(n_50),
.CI(n_39),
.CON(n_112),
.SN(n_112)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_54),
.A2(n_33),
.B1(n_17),
.B2(n_34),
.Y(n_104)
);

BUFx24_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_54),
.B(n_21),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_42),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_62),
.A2(n_30),
.B1(n_21),
.B2(n_24),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_19),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_131),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_95),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_0),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_114),
.A2(n_118),
.B(n_119),
.Y(n_161)
);

NAND3xp33_ASAP7_75t_SL g167 ( 
.A(n_115),
.B(n_63),
.C(n_72),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_0),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_0),
.Y(n_119)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_17),
.C(n_19),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_121),
.B(n_104),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_122),
.A2(n_125),
.B1(n_132),
.B2(n_100),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_72),
.B1(n_63),
.B2(n_73),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_50),
.C(n_42),
.Y(n_131)
);

AO22x2_ASAP7_75t_L g132 ( 
.A1(n_83),
.A2(n_42),
.B1(n_57),
.B2(n_59),
.Y(n_132)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_94),
.B(n_59),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_136),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_59),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_139),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_141),
.B(n_153),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_144),
.A2(n_150),
.B1(n_166),
.B2(n_160),
.Y(n_176)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_151),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_147),
.A2(n_148),
.B(n_156),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_126),
.A2(n_105),
.B(n_87),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_149),
.B(n_121),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_88),
.B1(n_106),
.B2(n_86),
.Y(n_150)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_152),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_140),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_109),
.Y(n_155)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_134),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_89),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_163),
.Y(n_201)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_160),
.A2(n_168),
.B1(n_169),
.B2(n_173),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_85),
.Y(n_162)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_82),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_126),
.A2(n_113),
.B(n_118),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_165),
.A2(n_170),
.B(n_19),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_113),
.A2(n_88),
.B1(n_106),
.B2(n_96),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_167),
.B(n_41),
.Y(n_208)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_127),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_119),
.A2(n_24),
.B(n_78),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_171),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_130),
.A2(n_100),
.B1(n_79),
.B2(n_82),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_172),
.A2(n_79),
.B1(n_112),
.B2(n_24),
.Y(n_188)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_124),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_176),
.A2(n_190),
.B1(n_198),
.B2(n_199),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_131),
.C(n_111),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_177),
.B(n_178),
.C(n_187),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_117),
.C(n_123),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_152),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_183),
.B(n_141),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_184),
.B(n_193),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_143),
.A2(n_114),
.B1(n_118),
.B2(n_116),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_186),
.A2(n_159),
.B1(n_170),
.B2(n_169),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_149),
.B(n_125),
.C(n_112),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_114),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_194),
.C(n_161),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_143),
.A2(n_119),
.B1(n_116),
.B2(n_137),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_144),
.B(n_1),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_192),
.A2(n_197),
.B(n_203),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_154),
.B(n_138),
.C(n_107),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_146),
.B(n_138),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_195),
.B(n_41),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_148),
.A2(n_35),
.B(n_17),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_151),
.A2(n_138),
.B1(n_13),
.B2(n_14),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_145),
.A2(n_35),
.B1(n_91),
.B2(n_90),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_147),
.A2(n_35),
.B(n_3),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_145),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_204),
.A2(n_173),
.B1(n_171),
.B2(n_164),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_146),
.B(n_35),
.Y(n_205)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_157),
.B(n_2),
.Y(n_206)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_206),
.Y(n_215)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_163),
.Y(n_207)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_208),
.A2(n_155),
.B(n_162),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_156),
.Y(n_209)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_209),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_154),
.Y(n_212)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_212),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_153),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_213),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_191),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_216),
.B(n_218),
.Y(n_261)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_217),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_221),
.A2(n_192),
.B1(n_193),
.B2(n_189),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_180),
.A2(n_161),
.B(n_166),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_222),
.A2(n_197),
.B(n_192),
.Y(n_239)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_223),
.Y(n_241)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_224),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_237),
.C(n_2),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_150),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_226),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_185),
.B(n_158),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_227),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_179),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_229),
.A2(n_230),
.B1(n_234),
.B2(n_235),
.Y(n_238)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_231),
.A2(n_200),
.B1(n_182),
.B2(n_175),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_233),
.B(n_236),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_206),
.B(n_152),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

AOI322xp5_ASAP7_75t_L g236 ( 
.A1(n_196),
.A2(n_55),
.A3(n_107),
.B1(n_173),
.B2(n_15),
.C1(n_14),
.C2(n_12),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_184),
.B(n_15),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_239),
.B(n_222),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_247),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_220),
.A2(n_176),
.B1(n_174),
.B2(n_175),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_244),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_216),
.A2(n_198),
.B1(n_204),
.B2(n_190),
.Y(n_245)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_177),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_211),
.A2(n_187),
.B1(n_178),
.B2(n_196),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_251),
.A2(n_215),
.B1(n_230),
.B2(n_228),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_226),
.A2(n_203),
.B1(n_186),
.B2(n_194),
.Y(n_252)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_220),
.A2(n_195),
.B1(n_200),
.B2(n_5),
.Y(n_253)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_253),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_210),
.A2(n_10),
.B(n_3),
.Y(n_254)
);

OAI31xp33_ASAP7_75t_SL g283 ( 
.A1(n_254),
.A2(n_258),
.A3(n_5),
.B(n_8),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_257),
.C(n_259),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_219),
.B(n_2),
.C(n_3),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_210),
.A2(n_10),
.B(n_7),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_219),
.B(n_5),
.C(n_7),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_238),
.Y(n_263)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_263),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_279),
.Y(n_289)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_255),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_267),
.Y(n_291)
);

OAI21x1_ASAP7_75t_L g269 ( 
.A1(n_261),
.A2(n_221),
.B(n_218),
.Y(n_269)
);

XOR2x2_ASAP7_75t_L g300 ( 
.A(n_269),
.B(n_258),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_255),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_276),
.Y(n_288)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_240),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_275),
.Y(n_292)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_240),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_248),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_228),
.Y(n_298)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_248),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_214),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_232),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_225),
.C(n_233),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_281),
.C(n_256),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_212),
.C(n_209),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_283),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_250),
.Y(n_284)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_284),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_249),
.B(n_239),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_286),
.A2(n_254),
.B(n_283),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_290),
.C(n_294),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_259),
.C(n_246),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_262),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_298),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_266),
.B(n_252),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_273),
.A2(n_249),
.B1(n_243),
.B2(n_242),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_296),
.A2(n_300),
.B1(n_271),
.B2(n_264),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_246),
.C(n_241),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_215),
.C(n_214),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_278),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_292),
.Y(n_302)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_302),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_300),
.A2(n_268),
.B(n_271),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_303),
.A2(n_299),
.B(n_296),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_308),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_244),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_310),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_306),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_274),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_309),
.C(n_289),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_295),
.A2(n_274),
.B1(n_265),
.B2(n_241),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_223),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_311),
.B(n_260),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_288),
.B(n_235),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_314),
.B(n_224),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_297),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_290),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_313),
.A2(n_285),
.B1(n_294),
.B2(n_286),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_317),
.B(n_323),
.C(n_301),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_321),
.B(n_324),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_322),
.B(n_325),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_315),
.A2(n_287),
.B1(n_270),
.B2(n_260),
.Y(n_323)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_312),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_326),
.B(n_270),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_327),
.A2(n_307),
.B(n_279),
.Y(n_331)
);

NOR2x1_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_309),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_328),
.B(n_330),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_306),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_331),
.B(n_333),
.C(n_335),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_320),
.B(n_308),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_332),
.A2(n_336),
.B1(n_327),
.B2(n_237),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_318),
.B(n_301),
.Y(n_335)
);

A2O1A1O1Ixp25_ASAP7_75t_L g338 ( 
.A1(n_334),
.A2(n_332),
.B(n_318),
.C(n_329),
.D(n_324),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_338),
.B(n_339),
.Y(n_342)
);

AO21x1_ASAP7_75t_L g340 ( 
.A1(n_329),
.A2(n_5),
.B(n_8),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_340),
.B(n_9),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_337),
.A2(n_8),
.B(n_9),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_343),
.B(n_344),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_342),
.C(n_341),
.Y(n_346)
);

BUFx24_ASAP7_75t_SL g347 ( 
.A(n_346),
.Y(n_347)
);

AOI221xp5_ASAP7_75t_L g348 ( 
.A1(n_347),
.A2(n_9),
.B1(n_10),
.B2(n_340),
.C(n_342),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_9),
.Y(n_349)
);


endmodule