module real_jpeg_24807_n_29 (n_17, n_8, n_0, n_21, n_168, n_2, n_10, n_9, n_12, n_24, n_165, n_166, n_170, n_6, n_28, n_161, n_162, n_169, n_167, n_23, n_11, n_14, n_160, n_25, n_163, n_7, n_22, n_18, n_3, n_5, n_4, n_1, n_26, n_27, n_20, n_19, n_164, n_16, n_15, n_13, n_29);

input n_17;
input n_8;
input n_0;
input n_21;
input n_168;
input n_2;
input n_10;
input n_9;
input n_12;
input n_24;
input n_165;
input n_166;
input n_170;
input n_6;
input n_28;
input n_161;
input n_162;
input n_169;
input n_167;
input n_23;
input n_11;
input n_14;
input n_160;
input n_25;
input n_163;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_164;
input n_16;
input n_15;
input n_13;

output n_29;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_64;
wire n_47;
wire n_131;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_113;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g94 ( 
.A(n_0),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_2),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_3),
.A2(n_32),
.B(n_36),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_3),
.B(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_3),
.B(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_3),
.B(n_39),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_4),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_4),
.B(n_68),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_5),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_6),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_7),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_8),
.A2(n_30),
.B(n_158),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_8),
.B(n_33),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_9),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_10),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_11),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_12),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_15),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_15),
.B(n_127),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_16),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_18),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_18),
.B(n_99),
.Y(n_101)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_19),
.Y(n_33)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_20),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_21),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_21),
.B(n_77),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_22),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_22),
.B(n_61),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_23),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_24),
.B(n_66),
.C(n_143),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_25),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_25),
.B(n_147),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_26),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_26),
.B(n_132),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_27),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_28),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_28),
.B(n_117),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_37),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_34),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_34),
.B(n_153),
.Y(n_152)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_35),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_35),
.B(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_35),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_35),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_35),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_41),
.B(n_157),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_57),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_48),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_45),
.B(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_69),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_53),
.B(n_148),
.Y(n_147)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_54),
.Y(n_145)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B(n_156),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_150),
.B(n_155),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_146),
.B(n_149),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_70),
.B(n_142),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_136),
.B(n_141),
.Y(n_70)
);

OAI321xp33_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_126),
.A3(n_131),
.B1(n_134),
.B2(n_135),
.C(n_160),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_121),
.B(n_125),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_116),
.B(n_120),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_110),
.B(n_115),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_82),
.B(n_109),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_102),
.B(n_108),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_98),
.B(n_101),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_90),
.B(n_97),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_86),
.B(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_96),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_103),
.B(n_104),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_111),
.B(n_112),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_122),
.B(n_123),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_128),
.B(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_140),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_137),
.B(n_140),
.Y(n_141)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_154),
.Y(n_155)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_161),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_162),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_163),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_164),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_165),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_166),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_167),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_168),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_169),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_170),
.Y(n_133)
);


endmodule