module fake_jpeg_24826_n_322 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_14),
.Y(n_24)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_24),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_39),
.B(n_45),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_46),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_0),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_19),
.Y(n_82)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_36),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_50),
.B(n_60),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_45),
.A2(n_37),
.B1(n_26),
.B2(n_35),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_51),
.A2(n_59),
.B(n_65),
.Y(n_116)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_55),
.Y(n_89)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_37),
.B1(n_20),
.B2(n_27),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_56),
.A2(n_63),
.B1(n_67),
.B2(n_68),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_21),
.B1(n_37),
.B2(n_29),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_72),
.B(n_33),
.C(n_21),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_58),
.B(n_69),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_37),
.B1(n_30),
.B2(n_26),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_36),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_25),
.C(n_29),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_62),
.B(n_64),
.C(n_73),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_27),
.B1(n_31),
.B2(n_23),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_49),
.A2(n_36),
.B1(n_27),
.B2(n_23),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_35),
.B1(n_26),
.B2(n_30),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_31),
.B1(n_23),
.B2(n_22),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_35),
.B1(n_30),
.B2(n_22),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_79),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_40),
.A2(n_20),
.B1(n_22),
.B2(n_31),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_71),
.B(n_83),
.Y(n_104)
);

NAND2x1_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_33),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_40),
.B(n_33),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_40),
.A2(n_20),
.B1(n_25),
.B2(n_34),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_39),
.A2(n_25),
.B1(n_34),
.B2(n_38),
.Y(n_75)
);

OA22x2_ASAP7_75t_SL g117 ( 
.A1(n_75),
.A2(n_80),
.B1(n_18),
.B2(n_28),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_40),
.B(n_21),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_84),
.Y(n_94)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_42),
.A2(n_38),
.B1(n_34),
.B2(n_18),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_87),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_42),
.A2(n_32),
.B1(n_34),
.B2(n_38),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_19),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_42),
.B(n_19),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_85),
.B(n_1),
.Y(n_107)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_93),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_90),
.A2(n_86),
.B(n_54),
.Y(n_147)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_91),
.B(n_103),
.Y(n_144)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_11),
.C(n_17),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_96),
.Y(n_140)
);

INVx6_ASAP7_75t_SL g96 ( 
.A(n_55),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_97),
.B(n_100),
.Y(n_142)
);

OR2x2_ASAP7_75t_SL g98 ( 
.A(n_62),
.B(n_19),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_98),
.A2(n_99),
.B(n_101),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_60),
.A2(n_32),
.B(n_38),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

NOR2xp67_ASAP7_75t_L g101 ( 
.A(n_57),
.B(n_9),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_77),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_107),
.Y(n_146)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_108),
.B(n_109),
.Y(n_155)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_32),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_121),
.Y(n_131)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_117),
.A2(n_119),
.B1(n_52),
.B2(n_66),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_78),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_118),
.B(n_123),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_77),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_18),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_78),
.B(n_28),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_97),
.A2(n_76),
.B1(n_52),
.B2(n_66),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_125),
.A2(n_135),
.B1(n_152),
.B2(n_154),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_118),
.B(n_85),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_127),
.B(n_151),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_128),
.A2(n_129),
.B1(n_141),
.B2(n_147),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_117),
.A2(n_52),
.B1(n_87),
.B2(n_70),
.Y(n_129)
);

AO22x1_ASAP7_75t_L g132 ( 
.A1(n_117),
.A2(n_73),
.B1(n_84),
.B2(n_87),
.Y(n_132)
);

OAI32xp33_ASAP7_75t_L g164 ( 
.A1(n_132),
.A2(n_88),
.A3(n_123),
.B1(n_93),
.B2(n_98),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_73),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_153),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_92),
.B1(n_90),
.B2(n_102),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_91),
.A2(n_69),
.B1(n_86),
.B2(n_61),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_136),
.A2(n_148),
.B1(n_119),
.B2(n_93),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_53),
.C(n_54),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_156),
.Y(n_169)
);

OA21x2_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_18),
.B(n_79),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_103),
.B(n_10),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_143),
.B(n_150),
.Y(n_185)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_145),
.B(n_109),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_88),
.A2(n_79),
.B1(n_28),
.B2(n_3),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_114),
.Y(n_166)
);

NOR2x1_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_28),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_28),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_104),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_1),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_2),
.C(n_3),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_4),
.C(n_5),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_4),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_144),
.B(n_115),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_182),
.Y(n_200)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_161),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_138),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_162),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_SL g203 ( 
.A1(n_164),
.A2(n_173),
.B(n_131),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_147),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_172),
.Y(n_196)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_96),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_167),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_168),
.A2(n_132),
.B1(n_141),
.B2(n_139),
.Y(n_193)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_170),
.B(n_171),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_144),
.B(n_113),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_146),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_175),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_145),
.B(n_113),
.Y(n_175)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_125),
.B(n_89),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_178),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_124),
.B(n_94),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_179),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_135),
.A2(n_104),
.B1(n_94),
.B2(n_99),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_180),
.A2(n_181),
.B1(n_157),
.B2(n_140),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_132),
.A2(n_111),
.B1(n_89),
.B2(n_122),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_131),
.B(n_107),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_130),
.B(n_110),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_105),
.Y(n_215)
);

INVx3_ASAP7_75t_SL g184 ( 
.A(n_134),
.Y(n_184)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_143),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_186),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_134),
.Y(n_187)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_152),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_189),
.A2(n_137),
.B1(n_108),
.B2(n_100),
.Y(n_220)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_141),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_191),
.A2(n_190),
.B1(n_150),
.B2(n_170),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_185),
.B(n_153),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_192),
.B(n_213),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_193),
.A2(n_204),
.B(n_209),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_126),
.B(n_133),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_194),
.A2(n_163),
.B(n_169),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_198),
.A2(n_189),
.B1(n_160),
.B2(n_186),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_203),
.A2(n_205),
.B1(n_211),
.B2(n_185),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_191),
.A2(n_126),
.B1(n_156),
.B2(n_124),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_151),
.Y(n_207)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_164),
.A2(n_127),
.B(n_111),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_106),
.C(n_137),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_158),
.C(n_159),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_176),
.Y(n_222)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_168),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_220),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_159),
.Y(n_221)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_222),
.B(n_226),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_223),
.B(n_236),
.Y(n_260)
);

BUFx8_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_229),
.Y(n_251)
);

AOI21x1_ASAP7_75t_SL g226 ( 
.A1(n_198),
.A2(n_183),
.B(n_188),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_235),
.C(n_242),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_201),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_169),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_231),
.Y(n_247)
);

INVx13_ASAP7_75t_L g233 ( 
.A(n_202),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_234),
.Y(n_256)
);

AND2x6_ASAP7_75t_L g234 ( 
.A(n_194),
.B(n_169),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_180),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_177),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_237),
.Y(n_257)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_208),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_197),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_162),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_243),
.B(n_199),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_193),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_244),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_244),
.A2(n_216),
.B1(n_213),
.B2(n_205),
.Y(n_245)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_245),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_224),
.A2(n_163),
.B1(n_204),
.B2(n_218),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_248),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_224),
.A2(n_231),
.B1(n_234),
.B2(n_240),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_225),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_250),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_252),
.B(n_239),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_227),
.A2(n_218),
.B1(n_219),
.B2(n_217),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_SL g270 ( 
.A1(n_255),
.A2(n_253),
.B(n_247),
.C(n_259),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_226),
.A2(n_211),
.B1(n_201),
.B2(n_214),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_259),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_229),
.A2(n_219),
.B1(n_217),
.B2(n_212),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_223),
.A2(n_212),
.B1(n_199),
.B2(n_195),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_261),
.A2(n_233),
.B1(n_195),
.B2(n_210),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_228),
.C(n_242),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_272),
.C(n_275),
.Y(n_288)
);

NAND3xp33_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_238),
.C(n_172),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_269),
.Y(n_281)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_267),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_252),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_268),
.B(n_271),
.Y(n_287)
);

BUFx12_ASAP7_75t_L g269 ( 
.A(n_254),
.Y(n_269)
);

O2A1O1Ixp33_ASAP7_75t_L g291 ( 
.A1(n_270),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_251),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_235),
.C(n_230),
.Y(n_272)
);

OAI322xp33_ASAP7_75t_L g273 ( 
.A1(n_260),
.A2(n_232),
.A3(n_207),
.B1(n_221),
.B2(n_222),
.C1(n_215),
.C2(n_230),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_262),
.Y(n_289)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_274),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_210),
.C(n_192),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_173),
.C(n_225),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_276),
.B(n_6),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_4),
.Y(n_279)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_279),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_256),
.B1(n_246),
.B2(n_255),
.Y(n_282)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_282),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_277),
.A2(n_245),
.B1(n_258),
.B2(n_261),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_286),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_277),
.A2(n_257),
.B1(n_262),
.B2(n_184),
.Y(n_286)
);

OAI211xp5_ASAP7_75t_SL g298 ( 
.A1(n_289),
.A2(n_291),
.B(n_270),
.C(n_269),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_278),
.A2(n_250),
.B1(n_184),
.B2(n_108),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_276),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_292),
.B(n_279),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_294),
.B(n_300),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_264),
.C(n_275),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_299),
.C(n_284),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_298),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_272),
.C(n_280),
.Y(n_299)
);

NOR2xp67_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_270),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_282),
.A2(n_280),
.B(n_270),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_301),
.A2(n_283),
.B(n_293),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_303),
.A2(n_306),
.B(n_307),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_299),
.B(n_286),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_309),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_302),
.A2(n_287),
.B(n_290),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_296),
.A2(n_283),
.B1(n_285),
.B2(n_269),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_308),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_310),
.B(n_313),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_285),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_291),
.Y(n_314)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_297),
.A3(n_304),
.B1(n_307),
.B2(n_295),
.C1(n_289),
.C2(n_7),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_317),
.C(n_9),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_7),
.C(n_9),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_316),
.A2(n_312),
.B(n_13),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_318),
.A2(n_319),
.B(n_15),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_16),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_16),
.Y(n_322)
);


endmodule