module fake_jpeg_13272_n_164 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_20),
.B(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_30),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_36),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_48),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_28),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_16),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_38),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_6),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_0),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_69),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_71),
.B(n_0),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_75),
.B(n_54),
.Y(n_89)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_76),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_81),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_71),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_67),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_59),
.B1(n_70),
.B2(n_50),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_91),
.B1(n_80),
.B2(n_69),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_79),
.A2(n_70),
.B1(n_72),
.B2(n_55),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_65),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_25),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_65),
.B1(n_50),
.B2(n_72),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_93),
.A2(n_94),
.B1(n_52),
.B2(n_53),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_51),
.B1(n_55),
.B2(n_58),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_104),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_78),
.B1(n_81),
.B2(n_74),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_96),
.A2(n_98),
.B1(n_99),
.B2(n_112),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_SL g97 ( 
.A(n_82),
.B(n_64),
.C(n_51),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_113),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_60),
.B1(n_63),
.B2(n_62),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_105),
.Y(n_131)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_109),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_108),
.Y(n_125)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_110),
.Y(n_127)
);

NAND2x1_ASAP7_75t_SL g130 ( 
.A(n_111),
.B(n_10),
.Y(n_130)
);

AOI32xp33_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_56),
.A3(n_61),
.B1(n_57),
.B2(n_21),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_18),
.B1(n_49),
.B2(n_47),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_114),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_88),
.C(n_76),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_124),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_128),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_76),
.B1(n_7),
.B2(n_8),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_123),
.B1(n_126),
.B2(n_129),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_L g123 ( 
.A1(n_108),
.A2(n_76),
.B1(n_19),
.B2(n_24),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_17),
.C(n_44),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_96),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_33),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_109),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_42),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_134),
.A2(n_15),
.B1(n_16),
.B2(n_31),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_37),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_124),
.C(n_140),
.Y(n_151)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_139),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_131),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_141),
.B(n_144),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_35),
.B(n_39),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_SL g154 ( 
.A1(n_143),
.A2(n_145),
.B(n_146),
.C(n_147),
.Y(n_154)
);

OA22x2_ASAP7_75t_L g145 ( 
.A1(n_133),
.A2(n_43),
.B1(n_126),
.B2(n_123),
.Y(n_145)
);

AO22x1_ASAP7_75t_L g146 ( 
.A1(n_133),
.A2(n_121),
.B1(n_127),
.B2(n_132),
.Y(n_146)
);

OA21x2_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_129),
.B(n_135),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_115),
.A2(n_117),
.B1(n_125),
.B2(n_128),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_148),
.B(n_130),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_148),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_151),
.B(n_152),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_146),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_154),
.A2(n_147),
.B1(n_145),
.B2(n_136),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_157),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_155),
.A2(n_150),
.B(n_153),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_158),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_157),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_159),
.B(n_149),
.C(n_154),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_162),
.A2(n_142),
.B(n_145),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_141),
.Y(n_164)
);


endmodule