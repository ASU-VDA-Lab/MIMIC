module fake_jpeg_2450_n_182 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_182);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_182;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_22),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_27),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_0),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_1),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_56),
.C(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_2),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_67),
.B(n_63),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_65),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_69),
.B1(n_68),
.B2(n_64),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_76),
.B(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_59),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_47),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_81),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_70),
.B(n_47),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_74),
.A2(n_48),
.B1(n_50),
.B2(n_68),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_93),
.B1(n_82),
.B2(n_57),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_88),
.Y(n_107)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_93),
.B1(n_84),
.B2(n_65),
.Y(n_101)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_92),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_74),
.B(n_52),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_98),
.Y(n_102)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_59),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_48),
.B1(n_69),
.B2(n_55),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_73),
.A2(n_69),
.B1(n_60),
.B2(n_55),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_99),
.B(n_5),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_52),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_82),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_60),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_51),
.B(n_58),
.C(n_61),
.Y(n_99)
);

BUFx24_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_100),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_101),
.A2(n_105),
.B1(n_32),
.B2(n_23),
.Y(n_137)
);

OAI32xp33_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_64),
.A3(n_57),
.B1(n_53),
.B2(n_82),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_6),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_96),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_106),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_2),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_111),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_83),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_57),
.B(n_4),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_18),
.B(n_20),
.Y(n_136)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_116),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_95),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_118),
.B1(n_9),
.B2(n_10),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_3),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_115),
.B(n_15),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_87),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_118),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_120),
.A2(n_122),
.B1(n_126),
.B2(n_131),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_110),
.A2(n_11),
.B(n_12),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_124),
.A2(n_137),
.B(n_138),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_133),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_101),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_126)
);

OAI32xp33_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_13),
.A3(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_130),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_31),
.B1(n_43),
.B2(n_19),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_30),
.C(n_42),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_16),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_29),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

OA21x2_ASAP7_75t_L g138 ( 
.A1(n_100),
.A2(n_34),
.B(n_24),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_129),
.A2(n_117),
.B(n_100),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_121),
.B(n_108),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_143),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_120),
.A2(n_114),
.B1(n_113),
.B2(n_18),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_142),
.A2(n_44),
.B1(n_150),
.B2(n_151),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_123),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_127),
.A2(n_25),
.B(n_26),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_151),
.B(n_153),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_149),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_126),
.A2(n_35),
.B(n_38),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_134),
.B(n_39),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_145),
.B1(n_148),
.B2(n_146),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_40),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_138),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_144),
.C(n_142),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_140),
.A2(n_138),
.B1(n_131),
.B2(n_136),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_140),
.A2(n_122),
.B1(n_132),
.B2(n_41),
.Y(n_157)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_168),
.Y(n_173)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_161),
.Y(n_165)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_165),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_147),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_155),
.Y(n_171)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_169),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_144),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_171),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_164),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_174),
.A2(n_171),
.B(n_170),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_176),
.A2(n_175),
.B1(n_163),
.B2(n_156),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_166),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_172),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_179),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_180),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_158),
.Y(n_182)
);


endmodule