module real_jpeg_19981_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_0),
.A2(n_33),
.B1(n_35),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_0),
.A2(n_23),
.B1(n_24),
.B2(n_39),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_39),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_1),
.B(n_23),
.Y(n_22)
);

A2O1A1O1Ixp25_ASAP7_75t_L g54 ( 
.A1(n_1),
.A2(n_22),
.B(n_23),
.C(n_55),
.D(n_58),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_1),
.B(n_70),
.Y(n_69)
);

A2O1A1O1Ixp25_ASAP7_75t_L g90 ( 
.A1(n_1),
.A2(n_26),
.B(n_46),
.C(n_81),
.D(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_1),
.B(n_26),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_1),
.B(n_56),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_1),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_1),
.A2(n_106),
.B(n_107),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_44),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_2),
.A2(n_33),
.B1(n_35),
.B2(n_44),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_4),
.B(n_35),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_4),
.A2(n_32),
.B1(n_40),
.B2(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_4),
.B(n_38),
.Y(n_107)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_4),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_5),
.A2(n_33),
.B1(n_35),
.B2(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_5),
.Y(n_75)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_7),
.A2(n_33),
.B1(n_35),
.B2(n_52),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_72),
.Y(n_71)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_86),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_85),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_61),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_17),
.B(n_61),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_41),
.C(n_54),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_18),
.A2(n_19),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_30),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_20),
.B(n_30),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B1(n_27),
.B2(n_29),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_28),
.Y(n_29)
);

O2A1O1Ixp33_ASAP7_75t_SL g55 ( 
.A1(n_24),
.A2(n_28),
.B(n_29),
.C(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_57),
.Y(n_56)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_27),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_27),
.B(n_47),
.Y(n_48)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_36),
.B(n_37),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_33),
.A2(n_35),
.B1(n_47),
.B2(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_33),
.A2(n_48),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_35),
.B(n_47),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_35),
.B(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_36),
.A2(n_37),
.B(n_112),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_36),
.B(n_121),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_40),
.A2(n_111),
.B1(n_113),
.B2(n_114),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_41),
.A2(n_42),
.B1(n_54),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_45),
.B1(n_51),
.B2(n_53),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_43),
.A2(n_53),
.B(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_45),
.A2(n_51),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_46),
.B(n_103),
.Y(n_102)
);

CKINVDCx9p33_ASAP7_75t_R g50 ( 
.A(n_47),
.Y(n_50)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_53),
.B(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_54),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_60),
.A2(n_65),
.B(n_66),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_77),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_68),
.B2(n_76),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_68),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_84),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_78),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_130),
.B(n_136),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_108),
.B(n_129),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_96),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_89),
.B(n_96),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_90),
.A2(n_92),
.B1(n_93),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_91),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_104),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_101),
.C(n_104),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_106),
.B(n_107),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_105),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_118),
.B(n_128),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_116),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_110),
.B(n_116),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_123),
.B(n_127),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_120),
.B(n_122),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_131),
.B(n_132),
.Y(n_136)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);


endmodule