module fake_jpeg_1159_n_226 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_226);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_28),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_27),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_6),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_2),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_45),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_9),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

BUFx16f_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

BUFx10_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

BUFx24_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_59),
.B(n_0),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_88),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_56),
.B(n_0),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_84),
.B1(n_87),
.B2(n_86),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_91),
.B1(n_99),
.B2(n_65),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_71),
.B1(n_65),
.B2(n_63),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_81),
.A2(n_79),
.B1(n_73),
.B2(n_55),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_96),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_67),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_64),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_73),
.B1(n_79),
.B2(n_61),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_55),
.B1(n_75),
.B2(n_69),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_101),
.A2(n_83),
.B1(n_61),
.B2(n_69),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_102),
.A2(n_62),
.B1(n_58),
.B2(n_80),
.Y(n_133)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_114),
.Y(n_126)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_117),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_78),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_111),
.B(n_112),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_66),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_68),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_113),
.B(n_119),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_71),
.B1(n_66),
.B2(n_54),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_116),
.A2(n_89),
.B1(n_115),
.B2(n_108),
.Y(n_123)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_118),
.A2(n_100),
.B1(n_70),
.B2(n_74),
.Y(n_129)
);

AOI21xp33_ASAP7_75t_L g119 ( 
.A1(n_98),
.A2(n_83),
.B(n_80),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_123),
.A2(n_129),
.B1(n_131),
.B2(n_135),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_94),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_141),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_54),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_125),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_120),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_128),
.B(n_130),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_111),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_116),
.A2(n_63),
.B1(n_100),
.B2(n_80),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_110),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_136),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_76),
.B1(n_60),
.B2(n_62),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_58),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_76),
.C(n_60),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_24),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_150),
.Y(n_169)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_137),
.A2(n_72),
.B1(n_3),
.B2(n_4),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_147),
.A2(n_158),
.B1(n_139),
.B2(n_13),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_127),
.A2(n_72),
.B(n_5),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_148),
.A2(n_165),
.B(n_136),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_143),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_149),
.B(n_151),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_1),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_33),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_143),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_155),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_29),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_157),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_34),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_129),
.A2(n_72),
.B1(n_53),
.B2(n_52),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_133),
.A2(n_1),
.B1(n_7),
.B2(n_8),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_159),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_8),
.Y(n_160)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_121),
.B(n_10),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_162),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_10),
.B(n_11),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_164),
.A2(n_142),
.B(n_140),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_11),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_140),
.B(n_12),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_166),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_170),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

OA21x2_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_142),
.B(n_139),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_178),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_173),
.A2(n_177),
.B1(n_181),
.B2(n_183),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_167),
.A2(n_12),
.B(n_13),
.Y(n_175)
);

OA21x2_ASAP7_75t_L g198 ( 
.A1(n_175),
.A2(n_152),
.B(n_43),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_156),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_156),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_163),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_183)
);

AOI322xp5_ASAP7_75t_L g184 ( 
.A1(n_161),
.A2(n_40),
.A3(n_48),
.B1(n_46),
.B2(n_36),
.C1(n_37),
.C2(n_38),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_158),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_161),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_186),
.A2(n_187),
.B1(n_164),
.B2(n_157),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_161),
.A2(n_23),
.B1(n_39),
.B2(n_41),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_151),
.C(n_145),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_194),
.C(n_195),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_146),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_193),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_182),
.B(n_148),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_154),
.C(n_155),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_159),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_197),
.A2(n_198),
.B1(n_186),
.B2(n_177),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_201),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_196),
.A2(n_179),
.B1(n_152),
.B2(n_181),
.Y(n_201)
);

AO21x2_ASAP7_75t_L g202 ( 
.A1(n_199),
.A2(n_171),
.B(n_178),
.Y(n_202)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_202),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_196),
.A2(n_175),
.B1(n_172),
.B2(n_168),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_204),
.B(n_198),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_174),
.C(n_172),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_199),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_212),
.C(n_203),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_203),
.B(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_213),
.B(n_214),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_207),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_210),
.B(n_169),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_215),
.A2(n_217),
.B(n_187),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_218),
.B(n_219),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_216),
.A2(n_205),
.B1(n_206),
.B2(n_198),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_214),
.C(n_209),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_221),
.A2(n_208),
.B(n_189),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_222),
.A2(n_202),
.B1(n_208),
.B2(n_51),
.Y(n_223)
);

BUFx24_ASAP7_75t_SL g224 ( 
.A(n_223),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_202),
.C(n_42),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_202),
.Y(n_226)
);


endmodule