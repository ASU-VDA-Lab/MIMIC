module fake_jpeg_28791_n_411 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_411);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_411;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_46),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_47),
.B(n_51),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_20),
.B(n_0),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_27),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_54),
.B(n_56),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_20),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_17),
.B(n_1),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_57),
.B(n_59),
.Y(n_137)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_22),
.Y(n_58)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_17),
.B(n_2),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_25),
.B(n_3),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_60),
.B(n_61),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_16),
.B(n_3),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_27),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_63),
.B(n_66),
.Y(n_117)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_27),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_25),
.B(n_3),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

AND2x6_ASAP7_75t_L g72 ( 
.A(n_34),
.B(n_4),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_72),
.A2(n_83),
.B(n_5),
.C(n_6),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_27),
.Y(n_73)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

BUFx4f_ASAP7_75t_SL g82 ( 
.A(n_34),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_29),
.B(n_5),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_27),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_84),
.A2(n_30),
.B1(n_16),
.B2(n_33),
.Y(n_127)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_85),
.A2(n_86),
.B1(n_31),
.B2(n_37),
.Y(n_94)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_94),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_18),
.B1(n_43),
.B2(n_41),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_95),
.A2(n_128),
.B1(n_61),
.B2(n_84),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_58),
.A2(n_18),
.B1(n_43),
.B2(n_36),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_97),
.A2(n_103),
.B1(n_104),
.B2(n_112),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_50),
.A2(n_18),
.B1(n_29),
.B2(n_42),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_98),
.A2(n_101),
.B1(n_123),
.B2(n_124),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_53),
.A2(n_67),
.B1(n_62),
.B2(n_86),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_71),
.A2(n_43),
.B1(n_36),
.B2(n_31),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_75),
.A2(n_36),
.B1(n_37),
.B2(n_19),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_76),
.A2(n_36),
.B1(n_37),
.B2(n_19),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_64),
.A2(n_36),
.B1(n_37),
.B2(n_19),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_115),
.A2(n_119),
.B1(n_132),
.B2(n_136),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_54),
.A2(n_37),
.B1(n_41),
.B2(n_40),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_65),
.A2(n_42),
.B1(n_16),
.B2(n_30),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_45),
.A2(n_40),
.B1(n_38),
.B2(n_35),
.Y(n_124)
);

OA22x2_ASAP7_75t_L g180 ( 
.A1(n_127),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_57),
.A2(n_38),
.B1(n_35),
.B2(n_30),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_69),
.A2(n_28),
.B1(n_6),
.B2(n_7),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_129),
.A2(n_87),
.B1(n_102),
.B2(n_28),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_131),
.B(n_61),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_63),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_73),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_138),
.Y(n_227)
);

INVx4_ASAP7_75t_SL g139 ( 
.A(n_106),
.Y(n_139)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_139),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_92),
.Y(n_140)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_140),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_117),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_141),
.B(n_145),
.Y(n_200)
);

AOI21xp33_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_59),
.B(n_44),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_142),
.B(n_147),
.Y(n_196)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_143),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_L g144 ( 
.A1(n_92),
.A2(n_85),
.B1(n_74),
.B2(n_55),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_144),
.A2(n_148),
.B1(n_180),
.B2(n_113),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_127),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_91),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_146),
.B(n_158),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_46),
.Y(n_147)
);

AO22x1_ASAP7_75t_SL g148 ( 
.A1(n_95),
.A2(n_96),
.B1(n_122),
.B2(n_107),
.Y(n_148)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_149),
.Y(n_190)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_150),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_151),
.B(n_169),
.Y(n_205)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_109),
.Y(n_152)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_152),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_153),
.A2(n_168),
.B1(n_170),
.B2(n_179),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_82),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_163),
.Y(n_189)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_156),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_111),
.B(n_82),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_157),
.B(n_159),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_88),
.B(n_70),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_91),
.Y(n_159)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_89),
.Y(n_160)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_160),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_122),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_88),
.B(n_81),
.Y(n_165)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

AND2x2_ASAP7_75t_SL g166 ( 
.A(n_105),
.B(n_80),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_166),
.B(n_176),
.C(n_183),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_167),
.A2(n_139),
.B1(n_164),
.B2(n_140),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_87),
.B(n_79),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_131),
.A2(n_49),
.B1(n_78),
.B2(n_52),
.Y(n_170)
);

NAND3xp33_ASAP7_75t_SL g171 ( 
.A(n_133),
.B(n_77),
.C(n_10),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_171),
.B(n_172),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_102),
.B(n_9),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_110),
.Y(n_173)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_173),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_96),
.B(n_110),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_177),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_118),
.B(n_10),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_93),
.B(n_134),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_121),
.A2(n_93),
.B(n_108),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_178),
.A2(n_100),
.B(n_120),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_90),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_118),
.B(n_12),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_184),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_130),
.B(n_106),
.Y(n_182)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

AND2x2_ASAP7_75t_SL g183 ( 
.A(n_125),
.B(n_13),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_130),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_125),
.B(n_13),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_187),
.Y(n_217)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_134),
.Y(n_187)
);

AND2x6_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_114),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_188),
.B(n_216),
.Y(n_234)
);

OAI32xp33_ASAP7_75t_L g191 ( 
.A1(n_163),
.A2(n_145),
.A3(n_151),
.B1(n_154),
.B2(n_170),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_191),
.B(n_199),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_114),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_194),
.B(n_226),
.C(n_207),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_199),
.B(n_213),
.Y(n_258)
);

A2O1A1Ixp33_ASAP7_75t_L g206 ( 
.A1(n_148),
.A2(n_89),
.B(n_100),
.C(n_14),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_206),
.B(n_162),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_155),
.A2(n_120),
.B1(n_126),
.B2(n_108),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_210),
.A2(n_215),
.B1(n_222),
.B2(n_229),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_212),
.A2(n_230),
.B(n_215),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_155),
.A2(n_14),
.B1(n_126),
.B2(n_185),
.Y(n_215)
);

AND2x6_ASAP7_75t_L g216 ( 
.A(n_158),
.B(n_14),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_186),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_230),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_156),
.A2(n_144),
.B1(n_185),
.B2(n_180),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_220),
.A2(n_138),
.B1(n_167),
.B2(n_212),
.Y(n_246)
);

O2A1O1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_178),
.A2(n_180),
.B(n_175),
.C(n_177),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_221),
.A2(n_159),
.B(n_167),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_161),
.A2(n_174),
.B1(n_180),
.B2(n_141),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_183),
.B(n_187),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_183),
.A2(n_173),
.B1(n_143),
.B2(n_166),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_166),
.B(n_146),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_231),
.A2(n_190),
.B(n_198),
.Y(n_285)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_202),
.Y(n_232)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_232),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_200),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_233),
.B(n_237),
.Y(n_281)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_197),
.Y(n_236)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_236),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_223),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_197),
.Y(n_238)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_238),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_239),
.A2(n_253),
.B(n_225),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_205),
.A2(n_149),
.B1(n_162),
.B2(n_140),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_240),
.A2(n_243),
.B1(n_246),
.B2(n_256),
.Y(n_271)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_202),
.Y(n_241)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_241),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_227),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_242),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_205),
.A2(n_160),
.B1(n_184),
.B2(n_139),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_150),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_244),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_189),
.B(n_152),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_248),
.Y(n_275)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_247),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_189),
.B(n_167),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_227),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_249),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_250),
.B(n_251),
.Y(n_292)
);

MAJx2_ASAP7_75t_L g251 ( 
.A(n_207),
.B(n_205),
.C(n_219),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_252),
.B(n_254),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_193),
.B(n_217),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_193),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_255),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_221),
.A2(n_191),
.B1(n_222),
.B2(n_188),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_257),
.B(n_259),
.Y(n_296)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_208),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_225),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_260),
.Y(n_280)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_208),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_261),
.B(n_263),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_194),
.B(n_226),
.C(n_196),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_195),
.C(n_211),
.Y(n_282)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_192),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_195),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_265),
.B(n_266),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_217),
.B(n_204),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_204),
.A2(n_228),
.B1(n_210),
.B2(n_206),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_267),
.A2(n_225),
.B1(n_224),
.B2(n_201),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_264),
.A2(n_224),
.B1(n_229),
.B2(n_216),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_270),
.A2(n_284),
.B1(n_289),
.B2(n_241),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_273),
.A2(n_274),
.B1(n_271),
.B2(n_290),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_257),
.A2(n_258),
.B1(n_267),
.B2(n_253),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_276),
.B(n_279),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_233),
.B(n_237),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_288),
.C(n_251),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_264),
.A2(n_190),
.B1(n_211),
.B2(n_198),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_285),
.A2(n_295),
.B(n_243),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_248),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_290),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_250),
.B(n_203),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_258),
.A2(n_190),
.B1(n_203),
.B2(n_214),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_245),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_239),
.A2(n_214),
.B(n_256),
.Y(n_295)
);

NOR3xp33_ASAP7_75t_SL g299 ( 
.A(n_234),
.B(n_258),
.C(n_235),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_299),
.B(n_273),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_300),
.A2(n_303),
.B(n_306),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_272),
.B(n_255),
.Y(n_302)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_302),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_296),
.A2(n_231),
.B(n_240),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_297),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_305),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_296),
.A2(n_246),
.B(n_262),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_279),
.B(n_232),
.Y(n_307)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_307),
.Y(n_333)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_297),
.Y(n_308)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_308),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_271),
.A2(n_260),
.B1(n_254),
.B2(n_235),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_309),
.A2(n_321),
.B1(n_324),
.B2(n_295),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_310),
.B(n_312),
.C(n_314),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_311),
.B(n_315),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_251),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_277),
.Y(n_313)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_313),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_266),
.C(n_265),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_270),
.A2(n_261),
.B1(n_259),
.B2(n_242),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_247),
.C(n_252),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_316),
.B(n_275),
.C(n_287),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_272),
.B(n_249),
.Y(n_317)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_317),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_281),
.B(n_263),
.Y(n_318)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_318),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_277),
.Y(n_319)
);

INVx11_ASAP7_75t_L g337 ( 
.A(n_319),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_284),
.A2(n_236),
.B1(n_238),
.B2(n_289),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_320),
.A2(n_268),
.B1(n_269),
.B2(n_280),
.Y(n_326)
);

AOI221xp5_ASAP7_75t_L g341 ( 
.A1(n_322),
.A2(n_299),
.B1(n_276),
.B2(n_294),
.C(n_275),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_280),
.B(n_281),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_323),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_274),
.A2(n_286),
.B1(n_285),
.B2(n_298),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_287),
.B(n_298),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_325),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_326),
.A2(n_329),
.B1(n_341),
.B2(n_311),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_288),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_328),
.B(n_336),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_317),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_331),
.B(n_323),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_310),
.B(n_288),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_314),
.B(n_282),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_345),
.C(n_346),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_316),
.B(n_282),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_332),
.A2(n_321),
.B1(n_324),
.B2(n_309),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_348),
.A2(n_354),
.B1(n_358),
.B2(n_363),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_333),
.B(n_307),
.Y(n_349)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_349),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_350),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_327),
.B(n_318),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_352),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_326),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_335),
.B(n_302),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_353),
.B(n_355),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_332),
.A2(n_305),
.B1(n_308),
.B2(n_301),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_347),
.B(n_304),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_342),
.A2(n_300),
.B(n_301),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_356),
.B(n_357),
.Y(n_367)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_335),
.Y(n_357)
);

NOR3xp33_ASAP7_75t_SL g358 ( 
.A(n_343),
.B(n_299),
.C(n_304),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_360),
.A2(n_343),
.B1(n_329),
.B2(n_330),
.Y(n_378)
);

MAJx2_ASAP7_75t_L g361 ( 
.A(n_334),
.B(n_306),
.C(n_325),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_361),
.B(n_336),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_347),
.B(n_268),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_362),
.B(n_344),
.Y(n_370)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_342),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_334),
.B(n_315),
.C(n_303),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_364),
.B(n_338),
.C(n_346),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_365),
.B(n_328),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_366),
.B(n_369),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_370),
.B(n_362),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_360),
.A2(n_339),
.B1(n_340),
.B2(n_319),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_372),
.A2(n_378),
.B1(n_352),
.B2(n_320),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_365),
.B(n_345),
.Y(n_375)
);

XNOR2x1_ASAP7_75t_L g390 ( 
.A(n_375),
.B(n_359),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_377),
.B(n_379),
.C(n_359),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_364),
.B(n_330),
.Y(n_379)
);

AO21x1_ASAP7_75t_L g380 ( 
.A1(n_367),
.A2(n_353),
.B(n_355),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_380),
.B(n_382),
.Y(n_395)
);

OAI221xp5_ASAP7_75t_L g383 ( 
.A1(n_368),
.A2(n_371),
.B1(n_373),
.B2(n_356),
.C(n_354),
.Y(n_383)
);

AOI21x1_ASAP7_75t_SL g398 ( 
.A1(n_383),
.A2(n_337),
.B(n_283),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_384),
.B(n_386),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_376),
.A2(n_363),
.B1(n_357),
.B2(n_358),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_385),
.A2(n_269),
.B1(n_337),
.B2(n_313),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_374),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_387),
.B(n_389),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_370),
.A2(n_351),
.B(n_349),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_388),
.A2(n_379),
.B(n_361),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_378),
.B(n_348),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_390),
.B(n_369),
.C(n_377),
.Y(n_391)
);

MAJx2_ASAP7_75t_L g401 ( 
.A(n_391),
.B(n_387),
.C(n_388),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_392),
.B(n_398),
.Y(n_403)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_393),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_390),
.B(n_375),
.C(n_366),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_394),
.B(n_381),
.C(n_389),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_398),
.A2(n_380),
.B(n_293),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_399),
.B(n_403),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_401),
.B(n_402),
.Y(n_406)
);

AOI322xp5_ASAP7_75t_L g404 ( 
.A1(n_400),
.A2(n_397),
.A3(n_395),
.B1(n_393),
.B2(n_396),
.C1(n_293),
.C2(n_283),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_404),
.B(n_403),
.Y(n_407)
);

AOI321xp33_ASAP7_75t_SL g409 ( 
.A1(n_407),
.A2(n_408),
.A3(n_406),
.B1(n_394),
.B2(n_291),
.C(n_278),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_405),
.B(n_396),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_409),
.A2(n_278),
.B(n_291),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_410),
.B(n_408),
.Y(n_411)
);


endmodule