module fake_jpeg_13270_n_329 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_38),
.B(n_41),
.Y(n_72)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_16),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_31),
.Y(n_49)
);

CKINVDCx9p33_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_49),
.B(n_19),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_29),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_62),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_46),
.A2(n_28),
.B1(n_19),
.B2(n_25),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_45),
.B1(n_44),
.B2(n_36),
.Y(n_76)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_54),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_16),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_61),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_22),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_34),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_22),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_67),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_33),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_35),
.B1(n_24),
.B2(n_21),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_68),
.A2(n_25),
.B1(n_23),
.B2(n_30),
.Y(n_98)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_17),
.Y(n_78)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_34),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_75),
.B(n_32),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_76),
.A2(n_85),
.B1(n_73),
.B2(n_71),
.Y(n_135)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_47),
.B1(n_39),
.B2(n_44),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_79),
.A2(n_82),
.B1(n_113),
.B2(n_64),
.Y(n_116)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_47),
.B1(n_39),
.B2(n_44),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_70),
.A2(n_18),
.B1(n_26),
.B2(n_33),
.Y(n_85)
);

AO22x1_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_44),
.B1(n_36),
.B2(n_37),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_86),
.B(n_96),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_26),
.C(n_37),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_110),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_89),
.B(n_102),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_36),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_93),
.Y(n_139)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_70),
.Y(n_94)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_27),
.B1(n_36),
.B2(n_37),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_95),
.A2(n_98),
.B1(n_111),
.B2(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_67),
.B(n_32),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_100),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_73),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_56),
.B(n_74),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_109),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_52),
.B(n_19),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_28),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_104),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_55),
.B(n_28),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_55),
.B(n_27),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_107),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_56),
.B(n_11),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_66),
.B(n_0),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_48),
.B(n_12),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_48),
.B(n_12),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_57),
.B(n_1),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_57),
.A2(n_35),
.B1(n_30),
.B2(n_24),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_73),
.B(n_69),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_115),
.A2(n_100),
.B(n_93),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_140),
.Y(n_148)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

INVx3_ASAP7_75t_SL g123 ( 
.A(n_90),
.Y(n_123)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_123),
.Y(n_164)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

NAND2x1_ASAP7_75t_SL g126 ( 
.A(n_80),
.B(n_73),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_126),
.A2(n_143),
.B(n_115),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_99),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_129),
.B(n_136),
.Y(n_177)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_135),
.Y(n_175)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_138),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_84),
.A2(n_60),
.B1(n_21),
.B2(n_35),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_141),
.A2(n_113),
.B1(n_94),
.B2(n_60),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_101),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_133),
.A2(n_84),
.B1(n_98),
.B2(n_88),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_144),
.A2(n_155),
.B1(n_163),
.B2(n_171),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_146),
.B(n_168),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_126),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_147),
.B(n_165),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_143),
.B(n_142),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_149),
.B(n_151),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_89),
.C(n_91),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_157),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_122),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_92),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_153),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_124),
.A2(n_91),
.B1(n_87),
.B2(n_94),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_154),
.A2(n_1),
.B(n_2),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_133),
.A2(n_112),
.B1(n_109),
.B2(n_111),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_79),
.C(n_82),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_139),
.A2(n_87),
.B(n_96),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_154),
.B(n_149),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_110),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_166),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_161),
.A2(n_176),
.B1(n_119),
.B2(n_123),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_134),
.B(n_92),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_162),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_116),
.A2(n_86),
.B1(n_21),
.B2(n_30),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_126),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_131),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_124),
.B(n_86),
.C(n_83),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_128),
.A2(n_86),
.B1(n_24),
.B2(n_23),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_114),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_172),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_114),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_173),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_83),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_174),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_127),
.A2(n_25),
.B1(n_108),
.B2(n_106),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_167),
.Y(n_179)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_180),
.B(n_174),
.Y(n_218)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_151),
.A2(n_121),
.B1(n_125),
.B2(n_141),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_183),
.A2(n_191),
.B1(n_198),
.B2(n_201),
.Y(n_214)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_185),
.B(n_164),
.Y(n_225)
);

OA21x2_ASAP7_75t_L g189 ( 
.A1(n_171),
.A2(n_121),
.B(n_130),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_189),
.A2(n_200),
.B(n_147),
.Y(n_211)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_190),
.B(n_194),
.Y(n_236)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_195),
.Y(n_215)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_145),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_196),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_157),
.A2(n_123),
.B1(n_140),
.B2(n_132),
.Y(n_198)
);

OAI22x1_ASAP7_75t_L g200 ( 
.A1(n_175),
.A2(n_108),
.B1(n_119),
.B2(n_71),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_170),
.A2(n_138),
.B1(n_137),
.B2(n_118),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_166),
.A2(n_138),
.B1(n_136),
.B2(n_120),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_209),
.B1(n_164),
.B2(n_172),
.Y(n_224)
);

AOI21xp33_ASAP7_75t_SL g203 ( 
.A1(n_159),
.A2(n_14),
.B(n_13),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_203),
.B(n_205),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_1),
.Y(n_235)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_148),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_146),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_177),
.A2(n_15),
.B1(n_10),
.B2(n_9),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_182),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_226),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_213),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_187),
.C(n_184),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_229),
.C(n_231),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_199),
.A2(n_165),
.B(n_177),
.Y(n_213)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_186),
.A2(n_150),
.B1(n_161),
.B2(n_160),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_217),
.A2(n_224),
.B1(n_198),
.B2(n_183),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_184),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_189),
.A2(n_148),
.B1(n_144),
.B2(n_176),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_220),
.A2(n_186),
.B1(n_207),
.B2(n_189),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_162),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_222),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_173),
.Y(n_223)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_155),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_145),
.Y(n_228)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_178),
.B(n_148),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_206),
.B(n_152),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_230),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_180),
.B(n_163),
.Y(n_231)
);

OAI21xp33_ASAP7_75t_SL g238 ( 
.A1(n_232),
.A2(n_235),
.B(n_208),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_10),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_234),
.C(n_195),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_187),
.B(n_8),
.C(n_2),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_257),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_242),
.A2(n_256),
.B1(n_227),
.B2(n_221),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_243),
.B(n_233),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_216),
.A2(n_197),
.B(n_199),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_253),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_217),
.A2(n_231),
.B1(n_223),
.B2(n_201),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_251),
.A2(n_214),
.B1(n_234),
.B2(n_219),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_235),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_220),
.A2(n_199),
.B1(n_190),
.B2(n_179),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_215),
.Y(n_254)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_254),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_212),
.B(n_194),
.C(n_192),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_239),
.C(n_259),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_214),
.A2(n_200),
.B1(n_8),
.B2(n_3),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_236),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_236),
.Y(n_258)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_258),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_218),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_213),
.Y(n_262)
);

XNOR2x1_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_276),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_272),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_266),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_255),
.C(n_243),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_247),
.A2(n_221),
.B1(n_219),
.B2(n_227),
.Y(n_268)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_211),
.Y(n_270)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_270),
.Y(n_292)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_274),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_235),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_245),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_277),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_1),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_2),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_273),
.A2(n_251),
.B1(n_242),
.B2(n_240),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_285),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_284),
.B(n_287),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_244),
.C(n_241),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_269),
.A2(n_241),
.B(n_237),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_7),
.Y(n_303)
);

AOI322xp5_ASAP7_75t_L g287 ( 
.A1(n_263),
.A2(n_249),
.A3(n_246),
.B1(n_253),
.B2(n_237),
.C1(n_256),
.C2(n_252),
.Y(n_287)
);

INVx13_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_288),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_3),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_261),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_273),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_290),
.A2(n_269),
.B1(n_270),
.B2(n_267),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_285),
.B(n_262),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_297),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_283),
.Y(n_296)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_296),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_282),
.B(n_260),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_298),
.A2(n_280),
.B1(n_290),
.B2(n_278),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_300),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_276),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_276),
.C(n_6),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_289),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_304),
.Y(n_313)
);

XNOR2x1_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_279),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_306),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_296),
.A2(n_281),
.B1(n_278),
.B2(n_286),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_307),
.A2(n_308),
.B1(n_310),
.B2(n_311),
.Y(n_317)
);

OAI21xp33_ASAP7_75t_L g311 ( 
.A1(n_301),
.A2(n_279),
.B(n_288),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_311),
.A2(n_303),
.B1(n_304),
.B2(n_7),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_291),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_293),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_295),
.C(n_297),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_316),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_317),
.B(n_319),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_318),
.B(n_313),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_313),
.B(n_4),
.Y(n_319)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_322),
.Y(n_323)
);

OAI211xp5_ASAP7_75t_L g324 ( 
.A1(n_320),
.A2(n_315),
.B(n_318),
.C(n_314),
.Y(n_324)
);

AOI31xp33_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_321),
.A3(n_6),
.B(n_7),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_323),
.C(n_4),
.Y(n_326)
);

BUFx24_ASAP7_75t_SL g327 ( 
.A(n_326),
.Y(n_327)
);

OAI21xp33_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_4),
.B(n_6),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_6),
.Y(n_329)
);


endmodule