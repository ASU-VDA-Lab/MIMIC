module fake_jpeg_21860_n_139 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx8_ASAP7_75t_SL g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_0),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_22),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_30),
.B(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_16),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_24),
.B1(n_29),
.B2(n_18),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_49),
.B1(n_27),
.B2(n_26),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_45),
.B(n_14),
.Y(n_66)
);

AO22x1_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_15),
.B1(n_27),
.B2(n_20),
.Y(n_47)
);

OA21x2_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_35),
.B(n_36),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_33),
.A2(n_24),
.B1(n_27),
.B2(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_24),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_22),
.Y(n_54)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_67),
.B(n_16),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_68),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_22),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_34),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_70),
.C(n_41),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_69),
.B1(n_43),
.B2(n_23),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_37),
.B1(n_38),
.B2(n_20),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_46),
.B1(n_40),
.B2(n_37),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_66),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_39),
.A2(n_17),
.B1(n_26),
.B2(n_25),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_22),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_43),
.A2(n_19),
.B1(n_23),
.B2(n_21),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_34),
.C(n_25),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_71),
.A2(n_46),
.B1(n_39),
.B2(n_48),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_72),
.A2(n_76),
.B(n_53),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_81),
.B(n_84),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_82),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_34),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_70),
.C(n_61),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_56),
.Y(n_91)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_98),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_92),
.C(n_97),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_56),
.Y(n_92)
);

AOI221xp5_ASAP7_75t_L g104 ( 
.A1(n_93),
.A2(n_80),
.B1(n_76),
.B2(n_85),
.C(n_84),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_62),
.B1(n_58),
.B2(n_60),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_96),
.B1(n_77),
.B2(n_82),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_60),
.B1(n_55),
.B2(n_57),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_55),
.Y(n_97)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_100),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_73),
.B(n_66),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_79),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_106),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_103),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_88),
.A2(n_78),
.B1(n_86),
.B2(n_77),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_95),
.B1(n_72),
.B2(n_74),
.Y(n_117)
);

AO221x1_ASAP7_75t_L g106 ( 
.A1(n_99),
.A2(n_77),
.B1(n_71),
.B2(n_65),
.C(n_87),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_107),
.A2(n_109),
.B1(n_89),
.B2(n_90),
.Y(n_113)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_1),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_74),
.B1(n_73),
.B2(n_87),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_113),
.B(n_105),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_118),
.C(n_119),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_119),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_91),
.C(n_92),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_93),
.B(n_97),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_125),
.C(n_115),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_108),
.C(n_107),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_126),
.A2(n_116),
.B1(n_117),
.B2(n_109),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_129),
.C(n_127),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_130),
.A2(n_122),
.B(n_3),
.Y(n_132)
);

AOI222xp33_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_19),
.B1(n_111),
.B2(n_5),
.C1(n_6),
.C2(n_8),
.Y(n_131)
);

AO21x1_ASAP7_75t_SL g135 ( 
.A1(n_131),
.A2(n_6),
.B(n_8),
.Y(n_135)
);

AO21x1_ASAP7_75t_L g136 ( 
.A1(n_132),
.A2(n_134),
.B(n_135),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_9),
.Y(n_137)
);

OAI21x1_ASAP7_75t_SL g134 ( 
.A1(n_130),
.A2(n_1),
.B(n_5),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_12),
.Y(n_138)
);

AOI221xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_136),
.B1(n_10),
.B2(n_12),
.C(n_1),
.Y(n_139)
);


endmodule