module fake_jpeg_25271_n_256 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_256);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_14;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_16),
.B(n_6),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_27),
.Y(n_38)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_6),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_12),
.B1(n_11),
.B2(n_21),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_11),
.C(n_15),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_33),
.C(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

MAJx2_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_61),
.C(n_30),
.Y(n_69)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_47),
.B(n_48),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_25),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_52),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_25),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g81 ( 
.A(n_50),
.B(n_57),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_17),
.B1(n_18),
.B2(n_16),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_59),
.B1(n_26),
.B2(n_31),
.Y(n_68)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_25),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

AOI22x1_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_30),
.B1(n_26),
.B2(n_31),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_36),
.A2(n_27),
.B(n_19),
.Y(n_61)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_28),
.B1(n_33),
.B2(n_32),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_47),
.B1(n_53),
.B2(n_59),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_41),
.B1(n_31),
.B2(n_36),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_36),
.B1(n_35),
.B2(n_49),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_41),
.B1(n_26),
.B2(n_31),
.Y(n_75)
);

OA21x2_ASAP7_75t_L g96 ( 
.A1(n_75),
.A2(n_60),
.B(n_37),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_77),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_27),
.B(n_18),
.Y(n_77)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_54),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_74),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_83),
.B(n_87),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_56),
.B1(n_72),
.B2(n_71),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_66),
.Y(n_87)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_68),
.A2(n_57),
.B1(n_45),
.B2(n_33),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_90),
.A2(n_92),
.B1(n_94),
.B2(n_97),
.Y(n_104)
);

INVxp33_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_99),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_28),
.B1(n_32),
.B2(n_41),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_93),
.B(n_98),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_66),
.A2(n_39),
.B1(n_41),
.B2(n_48),
.Y(n_94)
);

BUFx4f_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVxp67_ASAP7_75t_SL g121 ( 
.A(n_95),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_78),
.B(n_72),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_69),
.A2(n_39),
.B1(n_56),
.B2(n_46),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

AO21x1_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_50),
.B(n_62),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_100),
.B(n_119),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_82),
.A2(n_70),
.B1(n_64),
.B2(n_62),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_102),
.A2(n_55),
.B1(n_95),
.B2(n_26),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_75),
.B(n_69),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_114),
.B(n_96),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_81),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_107),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_81),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_110),
.B(n_96),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_75),
.B(n_78),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_112),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_75),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_115),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_75),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_80),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_116),
.A2(n_98),
.B1(n_93),
.B2(n_82),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_71),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_39),
.Y(n_126)
);

OA22x2_ASAP7_75t_L g157 ( 
.A1(n_122),
.A2(n_121),
.B1(n_18),
.B2(n_17),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_123),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_142),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_114),
.A2(n_96),
.B1(n_82),
.B2(n_89),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_128),
.B1(n_131),
.B2(n_101),
.Y(n_156)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_70),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_141),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_95),
.B1(n_55),
.B2(n_60),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_133),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_95),
.B(n_2),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_24),
.C(n_29),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_137),
.C(n_143),
.Y(n_167)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_144),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_24),
.C(n_29),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_138)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_30),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_115),
.A2(n_20),
.B(n_19),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_24),
.C(n_29),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_112),
.A2(n_111),
.B(n_103),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_109),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_145),
.Y(n_159)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_103),
.B(n_30),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_30),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_24),
.C(n_29),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_149),
.C(n_132),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_37),
.C(n_40),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_155),
.B(n_166),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_156),
.A2(n_158),
.B1(n_164),
.B2(n_148),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_157),
.B(n_163),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_139),
.A2(n_21),
.B1(n_22),
.B2(n_20),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_136),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_125),
.A2(n_21),
.B1(n_22),
.B2(n_40),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_140),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_165),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_130),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_168),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_169),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_142),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_171),
.B(n_122),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_147),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_127),
.C(n_135),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_177),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_178),
.A2(n_188),
.B1(n_190),
.B2(n_161),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_172),
.A2(n_124),
.B1(n_137),
.B2(n_143),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_179),
.A2(n_183),
.B1(n_153),
.B2(n_157),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_151),
.Y(n_199)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_184),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_154),
.A2(n_128),
.B1(n_141),
.B2(n_135),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_40),
.C(n_11),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_11),
.C(n_15),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_186),
.B(n_189),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_160),
.A2(n_17),
.B1(n_12),
.B2(n_15),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_151),
.B(n_150),
.C(n_173),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_159),
.A2(n_15),
.B1(n_23),
.B2(n_11),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_193),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_187),
.A2(n_154),
.B1(n_170),
.B2(n_163),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_196),
.A2(n_197),
.B1(n_206),
.B2(n_23),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_187),
.A2(n_156),
.B1(n_162),
.B2(n_164),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_150),
.B(n_158),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_8),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_200),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_175),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_153),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_30),
.C(n_23),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_202),
.A2(n_203),
.B1(n_8),
.B2(n_2),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_176),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_183),
.B(n_157),
.Y(n_204)
);

FAx1_ASAP7_75t_SL g218 ( 
.A(n_204),
.B(n_30),
.CI(n_14),
.CON(n_218),
.SN(n_218)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_191),
.A2(n_23),
.B1(n_2),
.B2(n_3),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_205),
.B(n_8),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_177),
.A2(n_185),
.B1(n_179),
.B2(n_181),
.Y(n_206)
);

FAx1_ASAP7_75t_L g207 ( 
.A(n_204),
.B(n_186),
.CI(n_184),
.CON(n_207),
.SN(n_207)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_209),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_218),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_206),
.A2(n_14),
.B1(n_2),
.B2(n_3),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_213),
.A2(n_215),
.B1(n_196),
.B2(n_1),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_214),
.B(n_217),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_192),
.A2(n_14),
.B1(n_13),
.B2(n_1),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_14),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_200),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_225),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_203),
.Y(n_222)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_222),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_223),
.B(n_228),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_201),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_211),
.A2(n_194),
.B(n_199),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_219),
.A2(n_207),
.B1(n_209),
.B2(n_218),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_230),
.B(n_232),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_219),
.A2(n_207),
.B(n_216),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_222),
.A2(n_4),
.B(n_5),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_235),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_227),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_226),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_7),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_226),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_7),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_233),
.A2(n_4),
.B1(n_7),
.B2(n_9),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_239),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_231),
.B(n_4),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_234),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_243),
.A2(n_244),
.B(n_9),
.Y(n_245)
);

NOR2x1_ASAP7_75t_SL g244 ( 
.A(n_231),
.B(n_9),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_247),
.B(n_242),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_246),
.A2(n_248),
.B(n_229),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_241),
.Y(n_248)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_249),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_242),
.C(n_9),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_251),
.A2(n_10),
.B(n_1),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_10),
.Y(n_254)
);

NAND3xp33_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_10),
.C(n_1),
.Y(n_255)
);

FAx1_ASAP7_75t_SL g256 ( 
.A(n_255),
.B(n_252),
.CI(n_1),
.CON(n_256),
.SN(n_256)
);


endmodule