module fake_jpeg_5772_n_325 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_325);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_39),
.Y(n_100)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_40),
.B(n_46),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_15),
.B(n_13),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_41),
.B(n_43),
.Y(n_101)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_15),
.B(n_13),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_52),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_18),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_50),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_22),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_16),
.B(n_0),
.Y(n_51)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_51),
.B(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_35),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_53),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_57),
.Y(n_83)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_59),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_16),
.B(n_12),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_60),
.B(n_61),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_21),
.B(n_11),
.Y(n_62)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_63),
.B(n_71),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_26),
.B1(n_30),
.B2(n_20),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_64),
.A2(n_99),
.B1(n_103),
.B2(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_65),
.B(n_11),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_20),
.B1(n_17),
.B2(n_30),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_66),
.A2(n_69),
.B1(n_80),
.B2(n_84),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_60),
.A2(n_20),
.B1(n_17),
.B2(n_30),
.Y(n_69)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_73),
.Y(n_119)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_74),
.B(n_79),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_26),
.B1(n_17),
.B2(n_36),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_75),
.A2(n_27),
.B1(n_31),
.B2(n_25),
.Y(n_113)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_47),
.A2(n_26),
.B1(n_22),
.B2(n_37),
.Y(n_80)
);

BUFx10_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_40),
.A2(n_37),
.B1(n_23),
.B2(n_36),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_85),
.B(n_87),
.Y(n_139)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_90),
.B(n_97),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_50),
.A2(n_29),
.B1(n_28),
.B2(n_24),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_91),
.A2(n_110),
.B1(n_0),
.B2(n_1),
.Y(n_138)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_51),
.A2(n_28),
.B1(n_24),
.B2(n_23),
.Y(n_99)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_102),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_59),
.A2(n_29),
.B1(n_34),
.B2(n_21),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_104),
.B(n_105),
.Y(n_112)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_107),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_41),
.B(n_38),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_19),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_43),
.A2(n_32),
.B1(n_31),
.B2(n_27),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_49),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_44),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_111),
.B(n_0),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_125),
.B1(n_128),
.B2(n_131),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_65),
.A2(n_27),
.B1(n_31),
.B2(n_38),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_115),
.A2(n_136),
.B1(n_143),
.B2(n_116),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_38),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_141),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_84),
.A2(n_38),
.B(n_19),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_122),
.B(n_127),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_120),
.B(n_3),
.Y(n_163)
);

NAND2x1_ASAP7_75t_SL g122 ( 
.A(n_108),
.B(n_54),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_66),
.A2(n_32),
.B1(n_31),
.B2(n_27),
.Y(n_125)
);

AND2x4_ASAP7_75t_L g127 ( 
.A(n_69),
.B(n_32),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_80),
.A2(n_32),
.B1(n_19),
.B2(n_54),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_101),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_98),
.A2(n_68),
.B1(n_82),
.B2(n_87),
.Y(n_131)
);

NOR4xp25_ASAP7_75t_SL g132 ( 
.A(n_93),
.B(n_77),
.C(n_8),
.D(n_10),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_5),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_68),
.A2(n_7),
.B1(n_1),
.B2(n_2),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_138),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_67),
.B(n_0),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_3),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_85),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_143)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_144),
.B(n_151),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_145),
.B(n_162),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_106),
.B1(n_83),
.B2(n_89),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_147),
.A2(n_154),
.B1(n_168),
.B2(n_177),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_150),
.A2(n_159),
.B1(n_170),
.B2(n_173),
.Y(n_202)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_156),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_110),
.Y(n_153)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

AO21x2_ASAP7_75t_SL g154 ( 
.A1(n_127),
.A2(n_111),
.B(n_76),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_127),
.A2(n_89),
.B1(n_100),
.B2(n_70),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_94),
.C(n_88),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_112),
.C(n_142),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_76),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_158),
.A2(n_163),
.B(n_169),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_134),
.A2(n_70),
.B1(n_86),
.B2(n_100),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_114),
.B(n_74),
.Y(n_160)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_165),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_73),
.Y(n_164)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

NAND3xp33_ASAP7_75t_SL g165 ( 
.A(n_122),
.B(n_127),
.C(n_120),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_166),
.B(n_176),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_117),
.B(n_81),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_170),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_118),
.A2(n_72),
.B1(n_102),
.B2(n_107),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_5),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_6),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_172),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_121),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_6),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_136),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_135),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_175),
.Y(n_182)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_125),
.A2(n_86),
.B1(n_81),
.B2(n_7),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_178),
.B(n_179),
.Y(n_213)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_129),
.Y(n_179)
);

A2O1A1O1Ixp25_ASAP7_75t_L g180 ( 
.A1(n_148),
.A2(n_132),
.B(n_134),
.C(n_130),
.D(n_124),
.Y(n_180)
);

AOI221xp5_ASAP7_75t_L g238 ( 
.A1(n_180),
.A2(n_192),
.B1(n_156),
.B2(n_176),
.C(n_179),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_172),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_195),
.Y(n_219)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_186),
.B(n_198),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_199),
.C(n_205),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_149),
.B(n_112),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_196),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_146),
.A2(n_113),
.B1(n_124),
.B2(n_135),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_194),
.A2(n_144),
.B1(n_156),
.B2(n_176),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_175),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_149),
.B(n_141),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_154),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_148),
.B(n_119),
.C(n_123),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_202),
.A2(n_209),
.B1(n_163),
.B2(n_178),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_123),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_206),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_157),
.B(n_119),
.C(n_126),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_173),
.B(n_152),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_159),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_207),
.B(n_214),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_150),
.A2(n_133),
.B1(n_137),
.B2(n_6),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_154),
.B(n_168),
.C(n_147),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_211),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_154),
.A2(n_133),
.B1(n_7),
.B2(n_6),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_198),
.A2(n_154),
.B(n_174),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_215),
.A2(n_220),
.B(n_224),
.Y(n_245)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_216),
.B(n_226),
.Y(n_254)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_186),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_217),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_200),
.A2(n_158),
.B(n_169),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_210),
.A2(n_146),
.B1(n_177),
.B2(n_174),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_221),
.A2(n_225),
.B1(n_235),
.B2(n_194),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_158),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_182),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_229),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_151),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_166),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_236),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_193),
.B(n_169),
.Y(n_232)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

INVxp67_ASAP7_75t_SL g233 ( 
.A(n_213),
.Y(n_233)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_233),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_207),
.A2(n_161),
.B1(n_162),
.B2(n_137),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_184),
.A2(n_7),
.B(n_144),
.Y(n_236)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_237),
.Y(n_243)
);

OA21x2_ASAP7_75t_SL g251 ( 
.A1(n_238),
.A2(n_197),
.B(n_211),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_212),
.A2(n_179),
.B(n_206),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_231),
.C(n_227),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_240),
.A2(n_236),
.B1(n_215),
.B2(n_237),
.Y(n_265)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_248),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_221),
.A2(n_184),
.B1(n_185),
.B2(n_192),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_246),
.A2(n_252),
.B1(n_222),
.B2(n_232),
.Y(n_275)
);

NAND5xp2_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_181),
.C(n_202),
.D(n_180),
.E(n_214),
.Y(n_247)
);

BUFx24_ASAP7_75t_SL g270 ( 
.A(n_247),
.Y(n_270)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_217),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_249),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_260),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_234),
.A2(n_185),
.B1(n_181),
.B2(n_209),
.Y(n_252)
);

NAND3xp33_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_183),
.C(n_195),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_257),
.Y(n_272)
);

BUFx12f_ASAP7_75t_SL g257 ( 
.A(n_239),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_250),
.Y(n_266)
);

BUFx12_ASAP7_75t_L g259 ( 
.A(n_226),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_187),
.Y(n_263)
);

A2O1A1O1Ixp25_ASAP7_75t_L g260 ( 
.A1(n_231),
.A2(n_197),
.B(n_191),
.C(n_205),
.D(n_190),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_218),
.Y(n_261)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_256),
.B(n_187),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_264),
.B(n_267),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_265),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_274),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_242),
.B(n_189),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_218),
.Y(n_269)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_269),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_243),
.A2(n_222),
.B1(n_224),
.B2(n_216),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_241),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_230),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_276),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_223),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_277),
.B(n_287),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_254),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_279),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_275),
.A2(n_257),
.B(n_245),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_285),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_254),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_282),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_245),
.B(n_241),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_273),
.A2(n_246),
.B1(n_240),
.B2(n_252),
.Y(n_287)
);

NOR2xp67_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_247),
.Y(n_290)
);

AOI31xp33_ASAP7_75t_L g295 ( 
.A1(n_290),
.A2(n_260),
.A3(n_229),
.B(n_220),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_266),
.C(n_274),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_296),
.C(n_299),
.Y(n_303)
);

MAJx2_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_273),
.C(n_276),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_292),
.A2(n_287),
.B(n_284),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_224),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_282),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_285),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_223),
.C(n_262),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_225),
.C(n_268),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_288),
.A2(n_235),
.B1(n_201),
.B2(n_189),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_284),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_188),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_279),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_305),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_306),
.A2(n_308),
.B(n_310),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_286),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_293),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_300),
.C(n_294),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_280),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_303),
.A2(n_299),
.B(n_297),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_311),
.A2(n_291),
.B(n_292),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_313),
.A2(n_316),
.B(n_315),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_314),
.A2(n_278),
.B1(n_286),
.B2(n_201),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_307),
.A2(n_296),
.B(n_302),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_317),
.B(n_278),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_318),
.A2(n_319),
.B(n_312),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_320),
.A2(n_321),
.B(n_301),
.Y(n_322)
);

AO21x1_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_249),
.B(n_259),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_208),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_259),
.Y(n_325)
);


endmodule