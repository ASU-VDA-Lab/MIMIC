module fake_netlist_6_3642_n_4584 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_442, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_468, n_111, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_466, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_397, n_155, n_109, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_298, n_18, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_363, n_395, n_323, n_393, n_411, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_102, n_204, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_464, n_33, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_328, n_429, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_64, n_288, n_427, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_4584);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_468;
input n_111;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_466;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_397;
input n_155;
input n_109;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_102;
input n_204;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_464;
input n_33;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_328;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_64;
input n_288;
input n_427;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_4584;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_801;
wire n_4452;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_1234;
wire n_2576;
wire n_3254;
wire n_3684;
wire n_1199;
wire n_1674;
wire n_3392;
wire n_741;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_625;
wire n_1189;
wire n_3152;
wire n_4154;
wire n_3579;
wire n_1212;
wire n_4251;
wire n_726;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3773;
wire n_700;
wire n_3783;
wire n_4177;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_4127;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_4504;
wire n_3844;
wire n_4388;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_4395;
wire n_4099;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_3741;
wire n_4517;
wire n_4168;
wire n_783;
wire n_2451;
wire n_1738;
wire n_4490;
wire n_2243;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_798;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_509;
wire n_1342;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_2977;
wire n_3952;
wire n_1739;
wire n_2051;
wire n_4370;
wire n_2317;
wire n_1380;
wire n_3911;
wire n_2359;
wire n_480;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_4285;
wire n_3465;
wire n_1975;
wire n_1009;
wire n_1930;
wire n_1743;
wire n_2405;
wire n_3706;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_4092;
wire n_1724;
wire n_1032;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_4078;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_4249;
wire n_1264;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_3619;
wire n_4359;
wire n_4087;
wire n_1700;
wire n_4578;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_4302;
wire n_2291;
wire n_830;
wire n_2299;
wire n_3340;
wire n_4179;
wire n_873;
wire n_1371;
wire n_1285;
wire n_2974;
wire n_2886;
wire n_3946;
wire n_1985;
wire n_4213;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_4474;
wire n_852;
wire n_2509;
wire n_4065;
wire n_4026;
wire n_4531;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_3904;
wire n_4178;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_4273;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_4446;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_4029;
wire n_836;
wire n_3345;
wire n_2074;
wire n_4417;
wire n_2447;
wire n_522;
wire n_2919;
wire n_4501;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_3879;
wire n_4010;
wire n_2286;
wire n_1649;
wire n_4555;
wire n_2094;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1772;
wire n_1232;
wire n_1572;
wire n_3979;
wire n_616;
wire n_658;
wire n_4308;
wire n_1874;
wire n_4347;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2739;
wire n_3023;
wire n_822;
wire n_3232;
wire n_693;
wire n_1313;
wire n_2791;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_1056;
wire n_3877;
wire n_3316;
wire n_4325;
wire n_2212;
wire n_3929;
wire n_758;
wire n_516;
wire n_3494;
wire n_3063;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3048;
wire n_4311;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_4060;
wire n_1550;
wire n_2703;
wire n_491;
wire n_3998;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_772;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_666;
wire n_4187;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2603;
wire n_2058;
wire n_2660;
wire n_538;
wire n_3028;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_4164;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_1094;
wire n_953;
wire n_3624;
wire n_3077;
wire n_3737;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3655;
wire n_494;
wire n_539;
wire n_4556;
wire n_493;
wire n_3107;
wire n_4563;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_4117;
wire n_3948;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_4327;
wire n_1961;
wire n_3047;
wire n_4414;
wire n_1280;
wire n_3765;
wire n_713;
wire n_2655;
wire n_4125;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_4221;
wire n_1467;
wire n_3297;
wire n_4250;
wire n_976;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_3906;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_4262;
wire n_4392;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3963;
wire n_3368;
wire n_917;
wire n_574;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_907;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_2591;
wire n_3507;
wire n_4334;
wire n_659;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_4253;
wire n_913;
wire n_4110;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_4071;
wire n_4255;
wire n_4403;
wire n_3506;
wire n_4268;
wire n_3568;
wire n_3269;
wire n_4047;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_473;
wire n_1193;
wire n_1967;
wire n_3999;
wire n_1054;
wire n_3928;
wire n_559;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_4139;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_4549;
wire n_4575;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_3943;
wire n_4320;
wire n_4305;
wire n_564;
wire n_2397;
wire n_3931;
wire n_3884;
wire n_4349;
wire n_824;
wire n_686;
wire n_4102;
wire n_4297;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_3871;
wire n_2907;
wire n_577;
wire n_3438;
wire n_2735;
wire n_4141;
wire n_1843;
wire n_619;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_2778;
wire n_4227;
wire n_2850;
wire n_572;
wire n_4314;
wire n_813;
wire n_2080;
wire n_1909;
wire n_1481;
wire n_3822;
wire n_4163;
wire n_606;
wire n_1441;
wire n_818;
wire n_3373;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_1699;
wire n_3910;
wire n_916;
wire n_3934;
wire n_2093;
wire n_4033;
wire n_4415;
wire n_4296;
wire n_4009;
wire n_2633;
wire n_483;
wire n_3883;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_4507;
wire n_630;
wire n_2059;
wire n_4080;
wire n_2198;
wire n_3319;
wire n_541;
wire n_512;
wire n_2669;
wire n_2925;
wire n_3728;
wire n_4094;
wire n_4499;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_2522;
wire n_792;
wire n_476;
wire n_3949;
wire n_4364;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_4354;
wire n_2616;
wire n_3912;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_3923;
wire n_2529;
wire n_3900;
wire n_4393;
wire n_1162;
wire n_860;
wire n_1530;
wire n_3798;
wire n_788;
wire n_939;
wire n_3488;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_3732;
wire n_982;
wire n_4372;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_2832;
wire n_4581;
wire n_4226;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_932;
wire n_2831;
wire n_2998;
wire n_4318;
wire n_4366;
wire n_3446;
wire n_4158;
wire n_4377;
wire n_3317;
wire n_3857;
wire n_3978;
wire n_1876;
wire n_4107;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_4074;
wire n_3716;
wire n_1873;
wire n_4294;
wire n_905;
wire n_3630;
wire n_3518;
wire n_4445;
wire n_3824;
wire n_3859;
wire n_1866;
wire n_4013;
wire n_1680;
wire n_2692;
wire n_993;
wire n_3842;
wire n_689;
wire n_3248;
wire n_2031;
wire n_4544;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_4456;
wire n_3914;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_547;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_558;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_4032;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_634;
wire n_2355;
wire n_3927;
wire n_4147;
wire n_4477;
wire n_966;
wire n_3888;
wire n_4511;
wire n_2908;
wire n_3168;
wire n_764;
wire n_4468;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_4337;
wire n_4130;
wire n_4161;
wire n_2895;
wire n_2009;
wire n_4172;
wire n_692;
wire n_3403;
wire n_733;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_3882;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_487;
wire n_3055;
wire n_3092;
wire n_3492;
wire n_3966;
wire n_4369;
wire n_3895;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_4454;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_1014;
wire n_3734;
wire n_4331;
wire n_3686;
wire n_4520;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_4118;
wire n_4502;
wire n_882;
wire n_4503;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_586;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_2459;
wire n_3746;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_4375;
wire n_715;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_3935;
wire n_1265;
wire n_4277;
wire n_4526;
wire n_2711;
wire n_3490;
wire n_4291;
wire n_4199;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_4319;
wire n_3369;
wire n_3419;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_2878;
wire n_618;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_3875;
wire n_4478;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_3794;
wire n_674;
wire n_3247;
wire n_871;
wire n_3069;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_2641;
wire n_1664;
wire n_1722;
wire n_612;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_3933;
wire n_702;
wire n_2749;
wire n_2008;
wire n_3298;
wire n_2192;
wire n_3346;
wire n_2254;
wire n_2345;
wire n_3281;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_4467;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_3691;
wire n_4427;
wire n_780;
wire n_3861;
wire n_675;
wire n_2624;
wire n_4066;
wire n_903;
wire n_4386;
wire n_4485;
wire n_4146;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_4340;
wire n_3891;
wire n_2193;
wire n_3961;
wire n_2676;
wire n_1655;
wire n_3940;
wire n_4072;
wire n_4220;
wire n_4523;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_1654;
wire n_816;
wire n_4371;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3428;
wire n_3153;
wire n_3410;
wire n_4552;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_604;
wire n_4004;
wire n_2810;
wire n_2967;
wire n_2519;
wire n_2319;
wire n_4043;
wire n_825;
wire n_728;
wire n_4353;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_4292;
wire n_1588;
wire n_3785;
wire n_3942;
wire n_3997;
wire n_2963;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_4381;
wire n_1124;
wire n_1624;
wire n_3873;
wire n_3983;
wire n_515;
wire n_2096;
wire n_2980;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_598;
wire n_3434;
wire n_4510;
wire n_696;
wire n_1515;
wire n_4473;
wire n_961;
wire n_4356;
wire n_3510;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_593;
wire n_4169;
wire n_514;
wire n_4055;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_3271;
wire n_950;
wire n_4362;
wire n_4248;
wire n_2812;
wire n_4518;
wire n_484;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_4361;
wire n_2393;
wire n_1796;
wire n_1757;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_3889;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_3707;
wire n_2075;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_4367;
wire n_2763;
wire n_2762;
wire n_4070;
wire n_1987;
wire n_3545;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_3578;
wire n_3885;
wire n_881;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_760;
wire n_3993;
wire n_1546;
wire n_2583;
wire n_4560;
wire n_590;
wire n_4394;
wire n_4116;
wire n_2606;
wire n_4031;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_2431;
wire n_3073;
wire n_4018;
wire n_2987;
wire n_694;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_3696;
wire n_3780;
wire n_4082;
wire n_2078;
wire n_1634;
wire n_3252;
wire n_2932;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_524;
wire n_3253;
wire n_3337;
wire n_3431;
wire n_3209;
wire n_3450;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_4002;
wire n_2658;
wire n_4329;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_2750;
wire n_2558;
wire n_2893;
wire n_1523;
wire n_2775;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_3477;
wire n_4289;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_4288;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_495;
wire n_815;
wire n_3953;
wire n_1100;
wire n_585;
wire n_1487;
wire n_4435;
wire n_2691;
wire n_3421;
wire n_840;
wire n_2913;
wire n_3614;
wire n_874;
wire n_4471;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_4019;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_898;
wire n_4385;
wire n_1952;
wire n_865;
wire n_3616;
wire n_4228;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_4044;
wire n_3436;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_4191;
wire n_1364;
wire n_4322;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_3937;
wire n_615;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_4287;
wire n_1293;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_3941;
wire n_963;
wire n_639;
wire n_2767;
wire n_794;
wire n_3793;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_4576;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_3385;
wire n_4350;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_872;
wire n_1139;
wire n_1714;
wire n_3922;
wire n_3179;
wire n_718;
wire n_1018;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_4330;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_2897;
wire n_2537;
wire n_3970;
wire n_4389;
wire n_4483;
wire n_4345;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_1513;
wire n_2747;
wire n_3924;
wire n_3171;
wire n_1913;
wire n_791;
wire n_4216;
wire n_3608;
wire n_510;
wire n_837;
wire n_4540;
wire n_4315;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_4156;
wire n_3491;
wire n_4240;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_704;
wire n_2148;
wire n_4284;
wire n_4162;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_536;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2590;
wire n_2643;
wire n_3353;
wire n_3150;
wire n_3018;
wire n_3782;
wire n_3975;
wire n_1469;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_4011;
wire n_1835;
wire n_3470;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_4098;
wire n_4021;
wire n_4476;
wire n_765;
wire n_1492;
wire n_987;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_4058;
wire n_4103;
wire n_3104;
wire n_631;
wire n_720;
wire n_3435;
wire n_842;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_4022;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_4310;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_4481;
wire n_1246;
wire n_4528;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_4475;
wire n_899;
wire n_738;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_499;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_705;
wire n_3580;
wire n_3775;
wire n_3537;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_2335;
wire n_1529;
wire n_2473;
wire n_4443;
wire n_3887;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_684;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_4096;
wire n_1431;
wire n_4123;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_3835;
wire n_4286;
wire n_1809;
wire n_3119;
wire n_4280;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_4379;
wire n_3731;
wire n_1822;
wire n_486;
wire n_947;
wire n_2936;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_648;
wire n_657;
wire n_1049;
wire n_3223;
wire n_3996;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_4525;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_4097;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_4218;
wire n_4440;
wire n_4402;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_3880;
wire n_1849;
wire n_2848;
wire n_919;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_478;
wire n_4541;
wire n_4100;
wire n_2231;
wire n_3609;
wire n_929;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_4551;
wire n_4264;
wire n_4484;
wire n_2857;
wire n_3693;
wire n_4497;
wire n_3788;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_777;
wire n_4459;
wire n_1299;
wire n_4545;
wire n_2896;
wire n_526;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_4079;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_2368;
wire n_4464;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_4175;
wire n_998;
wire n_717;
wire n_3200;
wire n_1665;
wire n_3893;
wire n_4306;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_4224;
wire n_3390;
wire n_3656;
wire n_4339;
wire n_1178;
wire n_2127;
wire n_2338;
wire n_1424;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_4455;
wire n_3867;
wire n_4453;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_3559;
wire n_4514;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_4005;
wire n_1507;
wire n_2482;
wire n_552;
wire n_3810;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_4564;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_912;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_3201;
wire n_3633;
wire n_3447;
wire n_4487;
wire n_3971;
wire n_1142;
wire n_2849;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_2354;
wire n_2682;
wire n_1774;
wire n_3032;
wire n_3103;
wire n_3638;
wire n_4573;
wire n_2589;
wire n_4535;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_3393;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_2442;
wire n_3627;
wire n_1791;
wire n_1368;
wire n_3480;
wire n_3451;
wire n_1418;
wire n_1250;
wire n_958;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_4222;
wire n_2545;
wire n_3540;
wire n_3577;
wire n_4401;
wire n_889;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_4368;
wire n_1478;
wire n_589;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_819;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_3641;
wire n_767;
wire n_3591;
wire n_1314;
wire n_600;
wire n_964;
wire n_1837;
wire n_2218;
wire n_2788;
wire n_831;
wire n_4533;
wire n_477;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_954;
wire n_4419;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_4120;
wire n_1382;
wire n_1534;
wire n_3892;
wire n_1736;
wire n_1564;
wire n_4069;
wire n_2748;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_505;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_537;
wire n_2511;
wire n_3964;
wire n_1993;
wire n_2281;
wire n_4167;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_596;
wire n_3944;
wire n_3909;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_4223;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_4431;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_4387;
wire n_2618;
wire n_2357;
wire n_2025;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_970;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_3481;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_4299;
wire n_3033;
wire n_3724;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_3913;
wire n_4276;
wire n_511;
wire n_2990;
wire n_3847;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_4430;
wire n_2410;
wire n_2552;
wire n_3302;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_4348;
wire n_520;
wire n_1093;
wire n_4428;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3226;
wire n_3323;
wire n_3364;
wire n_4020;
wire n_4176;
wire n_4489;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_775;
wire n_4404;
wire n_651;
wire n_1153;
wire n_1618;
wire n_3407;
wire n_518;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_2384;
wire n_3894;
wire n_4261;
wire n_4204;
wire n_1745;
wire n_914;
wire n_759;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_4496;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_4063;
wire n_1625;
wire n_3986;
wire n_4237;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_4513;
wire n_1453;
wire n_2146;
wire n_4006;
wire n_2226;
wire n_2131;
wire n_488;
wire n_2502;
wire n_2801;
wire n_3646;
wire n_497;
wire n_2920;
wire n_4015;
wire n_773;
wire n_3547;
wire n_1901;
wire n_3869;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_4570;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1892;
wire n_1459;
wire n_1614;
wire n_3188;
wire n_3742;
wire n_4410;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_4034;
wire n_1617;
wire n_4056;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_3960;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_3175;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_848;
wire n_2732;
wire n_2928;
wire n_4206;
wire n_4448;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_3862;
wire n_4267;
wire n_1580;
wire n_2227;
wire n_4247;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_4180;
wire n_3205;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_3284;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2720;
wire n_1520;
wire n_496;
wire n_3126;
wire n_2204;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_2863;
wire n_3299;
wire n_3663;
wire n_4132;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_3360;
wire n_4438;
wire n_2135;
wire n_3956;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_4001;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_4149;
wire n_1331;
wire n_736;
wire n_613;
wire n_2627;
wire n_4355;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_3234;
wire n_4422;
wire n_3917;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_2993;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3016;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_4126;
wire n_1129;
wire n_4003;
wire n_3870;
wire n_554;
wire n_602;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_3751;
wire n_664;
wire n_1869;
wire n_2911;
wire n_3625;
wire n_3804;
wire n_1764;
wire n_4207;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_4113;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_793;
wire n_4470;
wire n_587;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_4546;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_3901;
wire n_1937;
wire n_4583;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_4014;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_4067;
wire n_4252;
wire n_4357;
wire n_607;
wire n_1551;
wire n_4028;
wire n_4509;
wire n_4054;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_3907;
wire n_2555;
wire n_4048;
wire n_4444;
wire n_3338;
wire n_4217;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_820;
wire n_2327;
wire n_951;
wire n_4374;
wire n_2201;
wire n_725;
wire n_952;
wire n_3919;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_2984;
wire n_575;
wire n_994;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_4024;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_3194;
wire n_3113;
wire n_3276;
wire n_1934;
wire n_3250;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_4214;
wire n_4582;
wire n_1728;
wire n_3973;
wire n_557;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_4338;
wire n_617;
wire n_3886;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_485;
wire n_1549;
wire n_4420;
wire n_1510;
wire n_892;
wire n_768;
wire n_3637;
wire n_4574;
wire n_3120;
wire n_1468;
wire n_3991;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3797;
wire n_3926;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_2598;
wire n_1916;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_4405;
wire n_610;
wire n_4304;
wire n_4234;
wire n_4413;
wire n_1669;
wire n_1403;
wire n_4558;
wire n_1852;
wire n_4488;
wire n_4101;
wire n_3548;
wire n_3767;
wire n_1024;
wire n_3864;
wire n_4036;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_3974;
wire n_2052;
wire n_1847;
wire n_3634;
wire n_2302;
wire n_517;
wire n_4211;
wire n_4182;
wire n_1667;
wire n_667;
wire n_1206;
wire n_3230;
wire n_4016;
wire n_621;
wire n_1037;
wire n_1397;
wire n_3268;
wire n_3236;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_3592;
wire n_2755;
wire n_3141;
wire n_923;
wire n_504;
wire n_1409;
wire n_4230;
wire n_1841;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_3967;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_4328;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_4274;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_4189;
wire n_4270;
wire n_4151;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_710;
wire n_1108;
wire n_1818;
wire n_3730;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_4124;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_4397;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_785;
wire n_4155;
wire n_2740;
wire n_746;
wire n_4238;
wire n_609;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2401;
wire n_2337;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_4472;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_4152;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_4406;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_4380;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_4398;
wire n_2498;
wire n_4219;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_3238;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3529;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_4192;
wire n_4109;
wire n_1443;
wire n_2392;
wire n_1272;
wire n_2894;
wire n_3424;
wire n_4038;
wire n_3957;
wire n_2790;
wire n_4131;
wire n_4565;
wire n_2808;
wire n_2037;
wire n_3710;
wire n_4195;
wire n_4159;
wire n_4567;
wire n_3784;
wire n_2298;
wire n_2326;
wire n_782;
wire n_1539;
wire n_490;
wire n_4554;
wire n_3594;
wire n_809;
wire n_1043;
wire n_3819;
wire n_4090;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_4165;
wire n_986;
wire n_2305;
wire n_2373;
wire n_1472;
wire n_2050;
wire n_2120;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_4174;
wire n_1870;
wire n_2964;
wire n_4144;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3501;
wire n_662;
wire n_3475;
wire n_4442;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3905;
wire n_4434;
wire n_3262;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_4008;
wire n_2244;
wire n_4290;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_3692;
wire n_4515;
wire n_3845;
wire n_1682;
wire n_2017;
wire n_4516;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_4258;
wire n_4547;
wire n_650;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_4548;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_3826;
wire n_1406;
wire n_3790;
wire n_3878;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_4323;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_4300;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_4553;
wire n_2882;
wire n_3675;
wire n_3666;
wire n_4017;
wire n_4260;
wire n_3320;
wire n_2541;
wire n_654;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_1823;
wire n_2479;
wire n_776;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_1974;
wire n_3988;
wire n_4122;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_482;
wire n_934;
wire n_1637;
wire n_2635;
wire n_3307;
wire n_3439;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_3588;
wire n_4209;
wire n_2871;
wire n_4279;
wire n_4135;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_3858;
wire n_1845;
wire n_4183;
wire n_4321;
wire n_1489;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_4128;
wire n_543;
wire n_2229;
wire n_1964;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_4145;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_4271;
wire n_1946;
wire n_1355;
wire n_4181;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_4040;
wire n_4561;
wire n_804;
wire n_4461;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_4111;
wire n_533;
wire n_2390;
wire n_4007;
wire n_806;
wire n_3712;
wire n_959;
wire n_879;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_4239;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_4184;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_4037;
wire n_1319;
wire n_523;
wire n_707;
wire n_2986;
wire n_1900;
wire n_3930;
wire n_3246;
wire n_799;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_3915;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_787;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_4571;
wire n_4343;
wire n_2835;
wire n_4530;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_4215;
wire n_1282;
wire n_2561;
wire n_550;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_3377;
wire n_2939;
wire n_560;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_4185;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_4378;
wire n_4407;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_4045;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_3762;
wire n_3469;
wire n_3932;
wire n_2266;
wire n_2960;
wire n_3958;
wire n_3005;
wire n_3985;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1029;
wire n_4196;
wire n_3779;
wire n_1447;
wire n_4519;
wire n_2388;
wire n_3984;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_4358;
wire n_1706;
wire n_4242;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_4524;
wire n_2653;
wire n_2417;
wire n_4232;
wire n_4190;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_4052;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_4084;
wire n_4469;
wire n_3558;
wire n_3899;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_4326;
wire n_3156;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_4572;
wire n_3207;
wire n_502;
wire n_2668;
wire n_672;
wire n_4424;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_3939;
wire n_1375;
wire n_1941;
wire n_3483;
wire n_3613;
wire n_3972;
wire n_4153;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_2398;
wire n_1725;
wire n_1928;
wire n_1559;
wire n_3743;
wire n_3855;
wire n_1872;
wire n_3091;
wire n_4317;
wire n_834;
wire n_4493;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_4269;
wire n_743;
wire n_766;
wire n_3124;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_4088;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_545;
wire n_3524;
wire n_2671;
wire n_489;
wire n_2888;
wire n_2761;
wire n_2793;
wire n_2715;
wire n_2923;
wire n_1804;
wire n_2885;
wire n_3711;
wire n_3776;
wire n_4235;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_4301;
wire n_3511;
wire n_2054;
wire n_4143;
wire n_4170;
wire n_729;
wire n_876;
wire n_774;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_660;
wire n_2062;
wire n_4539;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_4421;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_4498;
wire n_2070;
wire n_2588;
wire n_479;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_869;
wire n_1154;
wire n_4492;
wire n_3308;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_4423;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_897;
wire n_846;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_841;
wire n_1476;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_4376;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_3515;
wire n_1150;
wire n_4203;
wire n_3808;
wire n_1742;
wire n_3190;
wire n_4505;
wire n_1562;
wire n_1690;
wire n_4365;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1118;
wire n_1076;
wire n_4512;
wire n_2949;
wire n_3726;
wire n_1807;
wire n_1007;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_3758;
wire n_1879;
wire n_853;
wire n_695;
wire n_3806;
wire n_4081;
wire n_1542;
wire n_2587;
wire n_4542;
wire n_3199;
wire n_2931;
wire n_875;
wire n_680;
wire n_4462;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_3866;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_671;
wire n_3565;
wire n_1953;
wire n_4450;
wire n_4536;
wire n_4543;
wire n_933;
wire n_740;
wire n_703;
wire n_3343;
wire n_3303;
wire n_978;
wire n_4157;
wire n_2752;
wire n_4173;
wire n_3135;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_4229;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_3990;
wire n_751;
wire n_749;
wire n_3865;
wire n_1824;
wire n_3954;
wire n_1628;
wire n_4073;
wire n_1324;
wire n_3890;
wire n_1399;
wire n_2122;
wire n_4550;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_988;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_3658;
wire n_1516;
wire n_4534;
wire n_1536;
wire n_3846;
wire n_2186;
wire n_2163;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3951;
wire n_3034;
wire n_823;
wire n_4408;
wire n_4577;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_4439;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_3874;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2969;
wire n_2395;
wire n_935;
wire n_3027;
wire n_781;
wire n_789;
wire n_1554;
wire n_3231;
wire n_4083;
wire n_4494;
wire n_1130;
wire n_3083;
wire n_4212;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_4295;
wire n_1120;
wire n_832;
wire n_1583;
wire n_4480;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_2746;
wire n_2946;
wire n_4579;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_4225;
wire n_4171;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_747;
wire n_3541;
wire n_2565;
wire n_4023;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_721;
wire n_1461;
wire n_742;
wire n_3432;
wire n_535;
wire n_691;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_3860;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_4282;
wire n_1598;
wire n_3493;
wire n_4344;
wire n_2935;
wire n_4046;
wire n_3807;
wire n_863;
wire n_3015;
wire n_2175;
wire n_601;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_3701;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_3473;
wire n_4557;
wire n_895;
wire n_866;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_3739;
wire n_2284;
wire n_4432;
wire n_3898;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_4352;
wire n_744;
wire n_971;
wire n_4391;
wire n_4416;
wire n_2702;
wire n_3241;
wire n_946;
wire n_2906;
wire n_761;
wire n_1303;
wire n_2769;
wire n_4342;
wire n_4465;
wire n_3622;
wire n_4568;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_4095;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_4495;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_4436;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3897;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_4569;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1016;
wire n_4559;
wire n_1347;
wire n_4106;
wire n_795;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_4027;
wire n_4373;
wire n_1245;
wire n_838;
wire n_3215;
wire n_3969;
wire n_3336;
wire n_647;
wire n_4160;
wire n_4231;
wire n_844;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_3853;
wire n_2117;
wire n_2234;
wire n_4256;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_3553;
wire n_1561;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_3811;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_653;
wire n_2430;
wire n_1414;
wire n_3486;
wire n_4086;
wire n_752;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_4335;
wire n_3556;
wire n_2034;
wire n_576;
wire n_1028;
wire n_3836;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_563;
wire n_4068;
wire n_2032;
wire n_4409;
wire n_2744;
wire n_4309;
wire n_4363;
wire n_1011;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_4521;
wire n_2437;
wire n_2444;
wire n_839;
wire n_1215;
wire n_2743;
wire n_3962;
wire n_708;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_668;
wire n_4166;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_3699;
wire n_4243;
wire n_3204;
wire n_1104;
wire n_1058;
wire n_854;
wire n_3378;
wire n_4025;
wire n_2312;
wire n_498;
wire n_3404;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_3362;
wire n_3745;
wire n_4059;
wire n_1509;
wire n_4188;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_4121;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3256;
wire n_1276;
wire n_3802;
wire n_3868;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_2118;
wire n_4313;
wire n_2111;
wire n_2466;
wire n_3982;
wire n_4266;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2505;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_3796;
wire n_2999;
wire n_4115;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3697;
wire n_3643;
wire n_1584;
wire n_771;
wire n_2425;
wire n_475;
wire n_924;
wire n_3461;
wire n_3408;
wire n_1582;
wire n_492;
wire n_3680;
wire n_4265;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_2408;
wire n_4246;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_4532;
wire n_719;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_4383;
wire n_4491;
wire n_3098;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_2666;
wire n_4105;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_4244;
wire n_4486;
wire n_1816;
wire n_4064;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_4049;
wire n_829;
wire n_1156;
wire n_1362;
wire n_4259;
wire n_3123;
wire n_2600;
wire n_984;
wire n_3380;
wire n_1829;
wire n_503;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_868;
wire n_3038;
wire n_570;
wire n_859;
wire n_2033;
wire n_3086;
wire n_735;
wire n_4104;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_3285;
wire n_519;
wire n_4208;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_500;
wire n_3769;
wire n_1482;
wire n_4529;
wire n_3361;
wire n_981;
wire n_3596;
wire n_714;
wire n_3478;
wire n_4537;
wire n_3936;
wire n_1349;
wire n_4346;
wire n_4351;
wire n_4089;
wire n_1144;
wire n_2071;
wire n_3669;
wire n_3863;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_985;
wire n_4316;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_481;
wire n_3521;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_4437;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_4390;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_4061;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_4075;
wire n_3344;
wire n_2334;
wire n_4062;
wire n_3902;
wire n_3881;
wire n_3295;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_4396;
wire n_4508;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_3989;
wire n_2478;
wire n_2303;
wire n_1619;
wire n_756;
wire n_1981;
wire n_2285;
wire n_4233;
wire n_4451;
wire n_1606;
wire n_4332;
wire n_810;
wire n_4460;
wire n_1133;
wire n_4108;
wire n_635;
wire n_1194;
wire n_3374;
wire n_4429;
wire n_4506;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_4538;
wire n_2640;
wire n_3695;
wire n_4051;
wire n_1051;
wire n_3976;
wire n_4254;
wire n_1552;
wire n_2918;
wire n_583;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_4307;
wire n_2367;
wire n_3992;
wire n_3876;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_4303;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_4293;
wire n_941;
wire n_3552;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2578;
wire n_2363;
wire n_4562;
wire n_553;
wire n_849;
wire n_2662;
wire n_3147;
wire n_3116;
wire n_3383;
wire n_3709;
wire n_753;
wire n_3925;
wire n_4091;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_4186;
wire n_3187;
wire n_2540;
wire n_4412;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_4580;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_2879;
wire n_861;
wire n_3717;
wire n_857;
wire n_967;
wire n_4522;
wire n_4148;
wire n_571;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_4341;
wire n_1884;
wire n_2040;
wire n_679;
wire n_4057;
wire n_2968;
wire n_4336;
wire n_4201;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_4263;
wire n_1819;
wire n_2055;
wire n_1260;
wire n_3555;
wire n_1010;
wire n_3444;
wire n_4210;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_4447;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_3955;
wire n_1805;
wire n_2477;
wire n_1557;
wire n_2280;
wire n_1888;
wire n_1833;
wire n_3903;
wire n_730;
wire n_1311;
wire n_3945;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_4205;
wire n_2308;
wire n_3854;
wire n_2162;
wire n_3908;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_4278;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3950;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_4463;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_3833;
wire n_4281;
wire n_3815;
wire n_2774;
wire n_3896;
wire n_3039;
wire n_681;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3333;
wire n_3274;
wire n_3186;
wire n_640;
wire n_1322;
wire n_4129;
wire n_4457;
wire n_965;
wire n_1899;
wire n_1428;
wire n_4093;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_3965;
wire n_2632;
wire n_2579;
wire n_722;
wire n_4500;
wire n_862;
wire n_2105;
wire n_3079;
wire n_4360;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_540;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_3584;
wire n_4039;
wire n_3387;
wire n_2027;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_4566;
wire n_4197;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_629;
wire n_1621;
wire n_4275;
wire n_4482;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_4283;
wire n_900;
wire n_3504;
wire n_4194;
wire n_1449;
wire n_4426;
wire n_531;
wire n_827;
wire n_2912;
wire n_4272;
wire n_2659;
wire n_2930;
wire n_4425;
wire n_1025;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_4449;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_649;
wire n_4030;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_73),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_51),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_91),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_252),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_459),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_425),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_145),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_406),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_150),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_295),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_13),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_119),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_423),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_118),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_221),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_261),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_457),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_199),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_414),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_38),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_224),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_236),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_308),
.Y(n_495)
);

BUFx10_ASAP7_75t_L g496 ( 
.A(n_301),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_127),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_168),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_284),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_419),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_449),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_40),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_75),
.Y(n_503)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_194),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_428),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_283),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_291),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_332),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_61),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_342),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_248),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_41),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_118),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_285),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_7),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_188),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_297),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_249),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_470),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_81),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_396),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_392),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_298),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_409),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_288),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_312),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_205),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_90),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_209),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_69),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_268),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_228),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_365),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_399),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_410),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_304),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_226),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_97),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_217),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_325),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_382),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_15),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_448),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_417),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_30),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_360),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_277),
.Y(n_547)
);

CKINVDCx16_ASAP7_75t_R g548 ( 
.A(n_407),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_158),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_395),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_6),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_468),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_92),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_337),
.Y(n_554)
);

BUFx5_ASAP7_75t_L g555 ( 
.A(n_456),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_254),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_463),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_19),
.Y(n_558)
);

INVx1_ASAP7_75t_SL g559 ( 
.A(n_455),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_137),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_187),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_49),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_206),
.Y(n_563)
);

BUFx10_ASAP7_75t_L g564 ( 
.A(n_71),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_426),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_161),
.Y(n_566)
);

CKINVDCx16_ASAP7_75t_R g567 ( 
.A(n_293),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_257),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_186),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_452),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_413),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_464),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_28),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_349),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_444),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_227),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_194),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_412),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_115),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_96),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_462),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_438),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_352),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_401),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_52),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_443),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_40),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_111),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_385),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_451),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_64),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_222),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_55),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_203),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_97),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_415),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_230),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_299),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_179),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_404),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_77),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_20),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_113),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_273),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_126),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_139),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_132),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_45),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_108),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_231),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_104),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_275),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_177),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_101),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_233),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_228),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_328),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_104),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_453),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_439),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_245),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_343),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_287),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_77),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_289),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_232),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_430),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_388),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_250),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_313),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_54),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_286),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_127),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_146),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_48),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_454),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_368),
.Y(n_637)
);

CKINVDCx6p67_ASAP7_75t_R g638 ( 
.A(n_86),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_229),
.Y(n_639)
);

CKINVDCx16_ASAP7_75t_R g640 ( 
.A(n_54),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_317),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_122),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_8),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_150),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_355),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_402),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_115),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_52),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_113),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_375),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_222),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_379),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_331),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_32),
.Y(n_654)
);

BUFx10_ASAP7_75t_L g655 ( 
.A(n_387),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_373),
.Y(n_656)
);

BUFx5_ASAP7_75t_L g657 ( 
.A(n_148),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_408),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_266),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_157),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_152),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_227),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_69),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_460),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_323),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_176),
.Y(n_666)
);

BUFx10_ASAP7_75t_L g667 ( 
.A(n_201),
.Y(n_667)
);

BUFx10_ASAP7_75t_L g668 ( 
.A(n_278),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_225),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_339),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_122),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_201),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_424),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_422),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_99),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_281),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_400),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_442),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_256),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_91),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_10),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_215),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_15),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_134),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_467),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_315),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_447),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_220),
.Y(n_688)
);

CKINVDCx20_ASAP7_75t_R g689 ( 
.A(n_377),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_221),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_270),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_321),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_182),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_471),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_319),
.Y(n_695)
);

BUFx10_ASAP7_75t_L g696 ( 
.A(n_165),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_74),
.Y(n_697)
);

BUFx2_ASAP7_75t_SL g698 ( 
.A(n_296),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_133),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_465),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_441),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_153),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_160),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_212),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_73),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_357),
.Y(n_706)
);

INVx1_ASAP7_75t_SL g707 ( 
.A(n_204),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_28),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_34),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_10),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_8),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_243),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_420),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_187),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_96),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_71),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_461),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_440),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_182),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_466),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_158),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_458),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_23),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_30),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_12),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_36),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_384),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_144),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_348),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_207),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_184),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_326),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_167),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_380),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_445),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_271),
.Y(n_736)
);

CKINVDCx14_ASAP7_75t_R g737 ( 
.A(n_213),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_184),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_186),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_105),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_383),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_306),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_121),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_235),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_251),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_136),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_429),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_200),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_397),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_370),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_292),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_7),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_151),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_195),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_133),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_49),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_469),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_237),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_78),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_160),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_450),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_137),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_55),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_42),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_446),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_335),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_129),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_179),
.Y(n_768)
);

CKINVDCx14_ASAP7_75t_R g769 ( 
.A(n_51),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_3),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_50),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_106),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_437),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_389),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_143),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_76),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_371),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_262),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_282),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_196),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_161),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_116),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_369),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_92),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_311),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_83),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_81),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_390),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_63),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_93),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_191),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_224),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_238),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_433),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_25),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_391),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_334),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_11),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_381),
.Y(n_799)
);

INVx1_ASAP7_75t_SL g800 ( 
.A(n_431),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_196),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_86),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_411),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_93),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_657),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_657),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_657),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_657),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_577),
.Y(n_809)
);

INVxp67_ASAP7_75t_SL g810 ( 
.A(n_628),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_572),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_657),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_572),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_657),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_694),
.B(n_0),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_564),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_475),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_657),
.Y(n_818)
);

BUFx5_ASAP7_75t_L g819 ( 
.A(n_478),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_657),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_484),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_605),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_737),
.B(n_0),
.Y(n_823)
);

BUFx3_ASAP7_75t_L g824 ( 
.A(n_501),
.Y(n_824)
);

CKINVDCx16_ASAP7_75t_R g825 ( 
.A(n_640),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_531),
.Y(n_826)
);

NOR2xp67_ASAP7_75t_L g827 ( 
.A(n_558),
.B(n_1),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_534),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_605),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_605),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_572),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_769),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_605),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_605),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_483),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_564),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_486),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_490),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_638),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_555),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_497),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_572),
.Y(n_842)
);

INVx1_ASAP7_75t_SL g843 ( 
.A(n_616),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_555),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_638),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_498),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_537),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_538),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_542),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_539),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_545),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_549),
.Y(n_852)
);

NOR2xp67_ASAP7_75t_L g853 ( 
.A(n_693),
.B(n_1),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_553),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_551),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_561),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_501),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_569),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_560),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_576),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_555),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_579),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_528),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_562),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_580),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_563),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_536),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_544),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_555),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_602),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_555),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_606),
.Y(n_872)
);

INVx1_ASAP7_75t_SL g873 ( 
.A(n_684),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_530),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_546),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_607),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_547),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_608),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_631),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_634),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_552),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_554),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_635),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_565),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_643),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_663),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_671),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_680),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_697),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_582),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_583),
.Y(n_891)
);

INVxp67_ASAP7_75t_SL g892 ( 
.A(n_550),
.Y(n_892)
);

CKINVDCx20_ASAP7_75t_R g893 ( 
.A(n_532),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_708),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_564),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_711),
.Y(n_896)
);

CKINVDCx20_ASAP7_75t_R g897 ( 
.A(n_599),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_584),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_566),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_721),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_724),
.Y(n_901)
);

CKINVDCx20_ASAP7_75t_R g902 ( 
.A(n_611),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_725),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_730),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_589),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_733),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_590),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_746),
.Y(n_908)
);

CKINVDCx20_ASAP7_75t_R g909 ( 
.A(n_618),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_596),
.Y(n_910)
);

INVx1_ASAP7_75t_SL g911 ( 
.A(n_649),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_550),
.B(n_556),
.Y(n_912)
);

CKINVDCx6p67_ASAP7_75t_R g913 ( 
.A(n_548),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_753),
.Y(n_914)
);

CKINVDCx16_ASAP7_75t_R g915 ( 
.A(n_567),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_759),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_780),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_598),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_556),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_615),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_615),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_718),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_600),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_473),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_604),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_610),
.Y(n_926)
);

CKINVDCx16_ASAP7_75t_R g927 ( 
.A(n_667),
.Y(n_927)
);

NOR2xp67_ASAP7_75t_L g928 ( 
.A(n_714),
.B(n_2),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_617),
.Y(n_929)
);

INVx1_ASAP7_75t_SL g930 ( 
.A(n_683),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_718),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_623),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_625),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_799),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_799),
.Y(n_935)
);

CKINVDCx14_ASAP7_75t_R g936 ( 
.A(n_496),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_507),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_508),
.Y(n_938)
);

BUFx2_ASAP7_75t_L g939 ( 
.A(n_473),
.Y(n_939)
);

INVx1_ASAP7_75t_SL g940 ( 
.A(n_763),
.Y(n_940)
);

CKINVDCx20_ASAP7_75t_R g941 ( 
.A(n_784),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_511),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_517),
.Y(n_943)
);

INVx1_ASAP7_75t_SL g944 ( 
.A(n_667),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_626),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_518),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_519),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_521),
.Y(n_948)
);

BUFx10_ASAP7_75t_L g949 ( 
.A(n_659),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_627),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_572),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_630),
.Y(n_952)
);

CKINVDCx16_ASAP7_75t_R g953 ( 
.A(n_667),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_555),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_525),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_535),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_555),
.Y(n_957)
);

CKINVDCx16_ASAP7_75t_R g958 ( 
.A(n_696),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_543),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_568),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_570),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_571),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_474),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_574),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_573),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_575),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_585),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_587),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_578),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_632),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_641),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_645),
.Y(n_972)
);

CKINVDCx20_ASAP7_75t_R g973 ( 
.A(n_474),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_581),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_646),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_652),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_555),
.Y(n_977)
);

BUFx5_ASAP7_75t_L g978 ( 
.A(n_586),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_597),
.Y(n_979)
);

CKINVDCx16_ASAP7_75t_R g980 ( 
.A(n_696),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_619),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_656),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_479),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_658),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_664),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_665),
.Y(n_986)
);

CKINVDCx14_ASAP7_75t_R g987 ( 
.A(n_496),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_620),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_621),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_670),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_622),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_673),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_676),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_629),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_637),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_677),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_487),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_678),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_479),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_679),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_650),
.Y(n_1001)
);

BUFx10_ASAP7_75t_L g1002 ( 
.A(n_659),
.Y(n_1002)
);

CKINVDCx20_ASAP7_75t_R g1003 ( 
.A(n_481),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_685),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_653),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_674),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_686),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_692),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_691),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_700),
.Y(n_1010)
);

INVxp67_ASAP7_75t_SL g1011 ( 
.A(n_717),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_722),
.Y(n_1012)
);

CKINVDCx16_ASAP7_75t_R g1013 ( 
.A(n_696),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_481),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_735),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_736),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_750),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_751),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_773),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_695),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_493),
.Y(n_1021)
);

CKINVDCx16_ASAP7_75t_R g1022 ( 
.A(n_495),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_774),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_779),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_701),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_487),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_675),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_706),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_712),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_713),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_720),
.Y(n_1031)
);

INVxp67_ASAP7_75t_L g1032 ( 
.A(n_493),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_793),
.Y(n_1033)
);

CKINVDCx20_ASAP7_75t_R g1034 ( 
.A(n_503),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_796),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_797),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_727),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_500),
.Y(n_1038)
);

INVx1_ASAP7_75t_SL g1039 ( 
.A(n_492),
.Y(n_1039)
);

INVx1_ASAP7_75t_SL g1040 ( 
.A(n_502),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_729),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_500),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_522),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_732),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_734),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_522),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_533),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_741),
.Y(n_1048)
);

BUFx8_ASAP7_75t_SL g1049 ( 
.A(n_804),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_742),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_700),
.Y(n_1051)
);

CKINVDCx20_ASAP7_75t_R g1052 ( 
.A(n_503),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_700),
.Y(n_1053)
);

NOR2xp67_ASAP7_75t_L g1054 ( 
.A(n_682),
.B(n_2),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_744),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_745),
.Y(n_1056)
);

CKINVDCx20_ASAP7_75t_R g1057 ( 
.A(n_509),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_747),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_533),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_749),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_612),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_612),
.Y(n_1062)
);

INVx1_ASAP7_75t_SL g1063 ( 
.A(n_504),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_757),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_687),
.Y(n_1065)
);

BUFx10_ASAP7_75t_L g1066 ( 
.A(n_788),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_761),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_687),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_675),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_509),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_512),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_688),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_688),
.Y(n_1073)
);

CKINVDCx16_ASAP7_75t_R g1074 ( 
.A(n_499),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_700),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_588),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_710),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_710),
.Y(n_1078)
);

INVxp33_ASAP7_75t_L g1079 ( 
.A(n_739),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_739),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_788),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_591),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_512),
.Y(n_1083)
);

CKINVDCx20_ASAP7_75t_R g1084 ( 
.A(n_513),
.Y(n_1084)
);

BUFx10_ASAP7_75t_L g1085 ( 
.A(n_682),
.Y(n_1085)
);

INVxp67_ASAP7_75t_L g1086 ( 
.A(n_513),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_592),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_700),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_593),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_786),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_786),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_594),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_595),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_777),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_777),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_601),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_603),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_609),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_777),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_613),
.Y(n_1100)
);

CKINVDCx20_ASAP7_75t_R g1101 ( 
.A(n_515),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_614),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_496),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_624),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_633),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_639),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_642),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_644),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_647),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_648),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_651),
.Y(n_1111)
);

CKINVDCx20_ASAP7_75t_R g1112 ( 
.A(n_515),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_777),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_654),
.Y(n_1114)
);

INVxp67_ASAP7_75t_L g1115 ( 
.A(n_804),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_516),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_660),
.Y(n_1117)
);

CKINVDCx16_ASAP7_75t_R g1118 ( 
.A(n_540),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_661),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_662),
.Y(n_1120)
);

CKINVDCx20_ASAP7_75t_R g1121 ( 
.A(n_516),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_520),
.Y(n_1122)
);

CKINVDCx20_ASAP7_75t_R g1123 ( 
.A(n_520),
.Y(n_1123)
);

CKINVDCx16_ASAP7_75t_R g1124 ( 
.A(n_541),
.Y(n_1124)
);

CKINVDCx14_ASAP7_75t_R g1125 ( 
.A(n_655),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_557),
.Y(n_1126)
);

INVx1_ASAP7_75t_SL g1127 ( 
.A(n_707),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_666),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_777),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_669),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_655),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_672),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_636),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_689),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_681),
.Y(n_1135)
);

INVx1_ASAP7_75t_SL g1136 ( 
.A(n_690),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_699),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_655),
.Y(n_1138)
);

CKINVDCx20_ASAP7_75t_R g1139 ( 
.A(n_527),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_702),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_758),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_703),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_704),
.Y(n_1143)
);

INVxp67_ASAP7_75t_L g1144 ( 
.A(n_527),
.Y(n_1144)
);

CKINVDCx20_ASAP7_75t_R g1145 ( 
.A(n_529),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_705),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_709),
.Y(n_1147)
);

INVxp67_ASAP7_75t_L g1148 ( 
.A(n_529),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_715),
.Y(n_1149)
);

INVxp67_ASAP7_75t_L g1150 ( 
.A(n_762),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_716),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_719),
.Y(n_1152)
);

NOR2xp67_ASAP7_75t_L g1153 ( 
.A(n_723),
.B(n_3),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_668),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_668),
.Y(n_1155)
);

INVxp67_ASAP7_75t_L g1156 ( 
.A(n_762),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_726),
.Y(n_1157)
);

INVxp67_ASAP7_75t_L g1158 ( 
.A(n_764),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_728),
.Y(n_1159)
);

INVxp67_ASAP7_75t_SL g1160 ( 
.A(n_559),
.Y(n_1160)
);

CKINVDCx20_ASAP7_75t_R g1161 ( 
.A(n_764),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_731),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_668),
.Y(n_1163)
);

CKINVDCx16_ASAP7_75t_R g1164 ( 
.A(n_698),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_738),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_740),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_743),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_748),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_824),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_822),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_829),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_826),
.Y(n_1172)
);

CKINVDCx20_ASAP7_75t_R g1173 ( 
.A(n_817),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_828),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_1039),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_824),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_1040),
.Y(n_1177)
);

INVxp33_ASAP7_75t_SL g1178 ( 
.A(n_832),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_867),
.Y(n_1179)
);

AND2x6_ASAP7_75t_L g1180 ( 
.A(n_912),
.B(n_785),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_830),
.Y(n_1181)
);

HB1xp67_ASAP7_75t_L g1182 ( 
.A(n_1063),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_868),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_973),
.Y(n_1184)
);

CKINVDCx20_ASAP7_75t_R g1185 ( 
.A(n_817),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_833),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_1127),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_833),
.Y(n_1188)
);

INVxp67_ASAP7_75t_SL g1189 ( 
.A(n_1138),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_875),
.Y(n_1190)
);

CKINVDCx20_ASAP7_75t_R g1191 ( 
.A(n_821),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_834),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_877),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_834),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1088),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_881),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_811),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_937),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_882),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1088),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_884),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_938),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_942),
.Y(n_1203)
);

INVxp67_ASAP7_75t_SL g1204 ( 
.A(n_1138),
.Y(n_1204)
);

INVxp67_ASAP7_75t_L g1205 ( 
.A(n_924),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_943),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_890),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_946),
.Y(n_1208)
);

INVxp33_ASAP7_75t_L g1209 ( 
.A(n_939),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_947),
.Y(n_1210)
);

CKINVDCx20_ASAP7_75t_R g1211 ( 
.A(n_821),
.Y(n_1211)
);

CKINVDCx20_ASAP7_75t_R g1212 ( 
.A(n_863),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_948),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_955),
.Y(n_1214)
);

CKINVDCx20_ASAP7_75t_R g1215 ( 
.A(n_863),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_1126),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_1133),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_956),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_959),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_960),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_961),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1160),
.B(n_800),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_962),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_964),
.Y(n_1224)
);

INVxp67_ASAP7_75t_SL g1225 ( 
.A(n_1138),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_891),
.Y(n_1226)
);

INVxp67_ASAP7_75t_SL g1227 ( 
.A(n_1138),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1094),
.Y(n_1228)
);

CKINVDCx20_ASAP7_75t_R g1229 ( 
.A(n_874),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1136),
.B(n_476),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_966),
.Y(n_1231)
);

CKINVDCx20_ASAP7_75t_R g1232 ( 
.A(n_874),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_1164),
.B(n_476),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_969),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_898),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_905),
.Y(n_1236)
);

CKINVDCx20_ASAP7_75t_R g1237 ( 
.A(n_893),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1163),
.B(n_477),
.Y(n_1238)
);

HB1xp67_ASAP7_75t_L g1239 ( 
.A(n_1142),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1163),
.B(n_477),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_907),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_974),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1094),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_910),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1095),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_918),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1163),
.B(n_1146),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_SL g1248 ( 
.A(n_1103),
.Y(n_1248)
);

HB1xp67_ASAP7_75t_L g1249 ( 
.A(n_1147),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_979),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_981),
.Y(n_1251)
);

INVxp67_ASAP7_75t_SL g1252 ( 
.A(n_1163),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_988),
.Y(n_1253)
);

CKINVDCx20_ASAP7_75t_R g1254 ( 
.A(n_893),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_989),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_991),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_994),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_923),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_995),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_897),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_1149),
.Y(n_1261)
);

CKINVDCx20_ASAP7_75t_R g1262 ( 
.A(n_897),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1151),
.Y(n_1263)
);

INVxp67_ASAP7_75t_SL g1264 ( 
.A(n_857),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_925),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1001),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_926),
.Y(n_1267)
);

INVxp67_ASAP7_75t_L g1268 ( 
.A(n_963),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1095),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_929),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_902),
.Y(n_1271)
);

CKINVDCx20_ASAP7_75t_R g1272 ( 
.A(n_902),
.Y(n_1272)
);

CKINVDCx20_ASAP7_75t_R g1273 ( 
.A(n_909),
.Y(n_1273)
);

NOR2xp67_ASAP7_75t_L g1274 ( 
.A(n_1032),
.B(n_480),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1005),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_909),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_857),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1006),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1007),
.Y(n_1279)
);

INVxp67_ASAP7_75t_L g1280 ( 
.A(n_999),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1009),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_932),
.Y(n_1282)
);

INVxp67_ASAP7_75t_SL g1283 ( 
.A(n_892),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1157),
.B(n_480),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1012),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1015),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1016),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1017),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_933),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1159),
.Y(n_1290)
);

INVxp67_ASAP7_75t_L g1291 ( 
.A(n_1014),
.Y(n_1291)
);

INVxp33_ASAP7_75t_SL g1292 ( 
.A(n_832),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1018),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_1167),
.B(n_482),
.Y(n_1294)
);

CKINVDCx16_ASAP7_75t_R g1295 ( 
.A(n_1022),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1019),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_945),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1023),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_950),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_952),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_941),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1024),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_973),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1033),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1035),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1036),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_835),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_837),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_970),
.B(n_482),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_971),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_972),
.B(n_975),
.Y(n_1311)
);

CKINVDCx20_ASAP7_75t_R g1312 ( 
.A(n_941),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_838),
.Y(n_1313)
);

INVxp33_ASAP7_75t_SL g1314 ( 
.A(n_976),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_841),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_982),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_984),
.Y(n_1317)
);

OR2x2_ASAP7_75t_L g1318 ( 
.A(n_843),
.B(n_752),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_985),
.B(n_485),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_846),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1099),
.Y(n_1321)
);

BUFx2_ASAP7_75t_SL g1322 ( 
.A(n_983),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_986),
.B(n_485),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_990),
.B(n_488),
.Y(n_1324)
);

INVxp67_ASAP7_75t_L g1325 ( 
.A(n_1071),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1099),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_847),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_848),
.Y(n_1328)
);

CKINVDCx20_ASAP7_75t_R g1329 ( 
.A(n_1049),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_992),
.B(n_488),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_849),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_993),
.Y(n_1332)
);

CKINVDCx20_ASAP7_75t_R g1333 ( 
.A(n_1049),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_852),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_855),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_996),
.Y(n_1336)
);

INVxp67_ASAP7_75t_SL g1337 ( 
.A(n_823),
.Y(n_1337)
);

NOR2xp67_ASAP7_75t_L g1338 ( 
.A(n_1086),
.B(n_489),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_856),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_850),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_998),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_825),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_1000),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_858),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1004),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_1074),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_860),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_862),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_865),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_870),
.Y(n_1350)
);

INVx2_ASAP7_75t_SL g1351 ( 
.A(n_1085),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_983),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1008),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_SL g1354 ( 
.A(n_1103),
.Y(n_1354)
);

INVxp67_ASAP7_75t_L g1355 ( 
.A(n_1122),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1020),
.B(n_489),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_872),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_876),
.Y(n_1358)
);

INVxp33_ASAP7_75t_L g1359 ( 
.A(n_1093),
.Y(n_1359)
);

CKINVDCx14_ASAP7_75t_R g1360 ( 
.A(n_936),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_878),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_1025),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_879),
.Y(n_1363)
);

INVx3_ASAP7_75t_L g1364 ( 
.A(n_811),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_1118),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_880),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_883),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_885),
.Y(n_1368)
);

INVxp33_ASAP7_75t_SL g1369 ( 
.A(n_1028),
.Y(n_1369)
);

CKINVDCx20_ASAP7_75t_R g1370 ( 
.A(n_1124),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_886),
.Y(n_1371)
);

CKINVDCx14_ASAP7_75t_R g1372 ( 
.A(n_936),
.Y(n_1372)
);

NOR2xp67_ASAP7_75t_L g1373 ( 
.A(n_1115),
.B(n_491),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_1029),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1030),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_887),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1031),
.Y(n_1377)
);

NOR2xp67_ASAP7_75t_L g1378 ( 
.A(n_1144),
.B(n_491),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_888),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1037),
.B(n_494),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_987),
.B(n_494),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1041),
.Y(n_1382)
);

CKINVDCx20_ASAP7_75t_R g1383 ( 
.A(n_1003),
.Y(n_1383)
);

CKINVDCx14_ASAP7_75t_R g1384 ( 
.A(n_987),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1044),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_850),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_889),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_894),
.Y(n_1388)
);

INVxp67_ASAP7_75t_L g1389 ( 
.A(n_944),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_1045),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_1048),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_896),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_900),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_901),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_1134),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1113),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_903),
.Y(n_1397)
);

CKINVDCx20_ASAP7_75t_R g1398 ( 
.A(n_1003),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_904),
.Y(n_1399)
);

CKINVDCx20_ASAP7_75t_R g1400 ( 
.A(n_1021),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_1021),
.Y(n_1401)
);

INVxp67_ASAP7_75t_SL g1402 ( 
.A(n_1097),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_1034),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_1034),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_906),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_908),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_914),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_916),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_917),
.Y(n_1409)
);

CKINVDCx16_ASAP7_75t_R g1410 ( 
.A(n_1125),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_1052),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_805),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_806),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1141),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_913),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_919),
.Y(n_1416)
);

INVxp67_ASAP7_75t_SL g1417 ( 
.A(n_1104),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_913),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_807),
.Y(n_1419)
);

INVxp67_ASAP7_75t_SL g1420 ( 
.A(n_1107),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_808),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_851),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_1052),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_812),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_814),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_818),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1090),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_1050),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1091),
.Y(n_1429)
);

CKINVDCx20_ASAP7_75t_R g1430 ( 
.A(n_1057),
.Y(n_1430)
);

CKINVDCx20_ASAP7_75t_R g1431 ( 
.A(n_1057),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_1070),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_1055),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1056),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_851),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1011),
.B(n_803),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1070),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1038),
.Y(n_1438)
);

CKINVDCx20_ASAP7_75t_R g1439 ( 
.A(n_1083),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1113),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1042),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1043),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1046),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_1058),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1047),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1059),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1125),
.B(n_1148),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1060),
.Y(n_1448)
);

INVxp33_ASAP7_75t_SL g1449 ( 
.A(n_1064),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1067),
.B(n_505),
.Y(n_1450)
);

CKINVDCx20_ASAP7_75t_R g1451 ( 
.A(n_1083),
.Y(n_1451)
);

CKINVDCx16_ASAP7_75t_R g1452 ( 
.A(n_927),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_854),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1061),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1062),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1065),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_1084),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1068),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_920),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_854),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_921),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_859),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_811),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_859),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_922),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_864),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_864),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_931),
.Y(n_1468)
);

CKINVDCx20_ASAP7_75t_R g1469 ( 
.A(n_1084),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_934),
.Y(n_1470)
);

CKINVDCx20_ASAP7_75t_R g1471 ( 
.A(n_1101),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_935),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1081),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_866),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1175),
.B(n_873),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1195),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1307),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1169),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1169),
.B(n_997),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_1177),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1337),
.B(n_819),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1189),
.B(n_1204),
.Y(n_1482)
);

AND2x6_ASAP7_75t_L g1483 ( 
.A(n_1381),
.B(n_1131),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_SL g1484 ( 
.A(n_1182),
.B(n_915),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1195),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1200),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1359),
.A2(n_815),
.B1(n_810),
.B2(n_1150),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_1176),
.Y(n_1488)
);

BUFx6f_ASAP7_75t_L g1489 ( 
.A(n_1463),
.Y(n_1489)
);

BUFx3_ASAP7_75t_L g1490 ( 
.A(n_1176),
.Y(n_1490)
);

INVx2_ASAP7_75t_SL g1491 ( 
.A(n_1187),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1389),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1308),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_SL g1494 ( 
.A1(n_1342),
.A2(n_1112),
.B1(n_1116),
.B2(n_1101),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1200),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1313),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1228),
.Y(n_1497)
);

INVx6_ASAP7_75t_L g1498 ( 
.A(n_1277),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1228),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1225),
.B(n_819),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1227),
.B(n_1252),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1315),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1463),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1243),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1243),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1320),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1277),
.B(n_997),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1342),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1245),
.Y(n_1509)
);

OA21x2_ASAP7_75t_L g1510 ( 
.A1(n_1412),
.A2(n_1129),
.B(n_820),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1230),
.B(n_1156),
.Y(n_1511)
);

OA21x2_ASAP7_75t_L g1512 ( 
.A1(n_1413),
.A2(n_1129),
.B(n_820),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1283),
.B(n_1238),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1327),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1328),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1331),
.Y(n_1516)
);

OA21x2_ASAP7_75t_L g1517 ( 
.A1(n_1419),
.A2(n_844),
.B(n_840),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1416),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1334),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1351),
.B(n_1222),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1335),
.Y(n_1521)
);

BUFx6f_ASAP7_75t_L g1522 ( 
.A(n_1463),
.Y(n_1522)
);

BUFx6f_ASAP7_75t_L g1523 ( 
.A(n_1463),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_1245),
.Y(n_1524)
);

AND2x4_ASAP7_75t_L g1525 ( 
.A(n_1264),
.B(n_1026),
.Y(n_1525)
);

BUFx6f_ASAP7_75t_L g1526 ( 
.A(n_1197),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_1197),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1339),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_1197),
.Y(n_1529)
);

CKINVDCx11_ASAP7_75t_R g1530 ( 
.A(n_1329),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1240),
.B(n_819),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1344),
.Y(n_1532)
);

BUFx6f_ASAP7_75t_L g1533 ( 
.A(n_1364),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1347),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1348),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1349),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1350),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1357),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1346),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1416),
.B(n_1468),
.Y(n_1540)
);

XNOR2xp5_ASAP7_75t_L g1541 ( 
.A(n_1346),
.B(n_911),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1351),
.B(n_1158),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1318),
.Y(n_1543)
);

AOI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1180),
.A2(n_866),
.B1(n_965),
.B2(n_899),
.Y(n_1544)
);

AOI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1180),
.A2(n_899),
.B1(n_967),
.B2(n_965),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1269),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_1216),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1269),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1321),
.Y(n_1549)
);

BUFx6f_ASAP7_75t_L g1550 ( 
.A(n_1364),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1360),
.B(n_816),
.Y(n_1551)
);

OA21x2_ASAP7_75t_L g1552 ( 
.A1(n_1421),
.A2(n_844),
.B(n_840),
.Y(n_1552)
);

BUFx6f_ASAP7_75t_L g1553 ( 
.A(n_1364),
.Y(n_1553)
);

BUFx6f_ASAP7_75t_L g1554 ( 
.A(n_1321),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1326),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1358),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1436),
.Y(n_1557)
);

AOI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1180),
.A2(n_967),
.B1(n_1076),
.B2(n_968),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1326),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1459),
.B(n_1026),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1361),
.Y(n_1561)
);

OA21x2_ASAP7_75t_L g1562 ( 
.A1(n_1424),
.A2(n_1426),
.B(n_1425),
.Y(n_1562)
);

BUFx6f_ASAP7_75t_L g1563 ( 
.A(n_1396),
.Y(n_1563)
);

BUFx6f_ASAP7_75t_L g1564 ( 
.A(n_1396),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_SL g1565 ( 
.A1(n_1365),
.A2(n_1116),
.B1(n_1121),
.B2(n_1112),
.Y(n_1565)
);

INVx3_ASAP7_75t_L g1566 ( 
.A(n_1440),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1363),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1366),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_SL g1569 ( 
.A(n_1410),
.B(n_839),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1367),
.Y(n_1570)
);

BUFx6f_ASAP7_75t_L g1571 ( 
.A(n_1440),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1372),
.B(n_1384),
.Y(n_1572)
);

OA21x2_ASAP7_75t_L g1573 ( 
.A1(n_1170),
.A2(n_869),
.B(n_861),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1359),
.B(n_1402),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1186),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1188),
.Y(n_1576)
);

CKINVDCx8_ASAP7_75t_R g1577 ( 
.A(n_1322),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1368),
.Y(n_1578)
);

CKINVDCx11_ASAP7_75t_R g1579 ( 
.A(n_1329),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1436),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1192),
.Y(n_1581)
);

OA21x2_ASAP7_75t_L g1582 ( 
.A1(n_1171),
.A2(n_869),
.B(n_861),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1371),
.Y(n_1583)
);

XNOR2xp5_ASAP7_75t_L g1584 ( 
.A(n_1365),
.B(n_930),
.Y(n_1584)
);

BUFx6f_ASAP7_75t_L g1585 ( 
.A(n_1198),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1376),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1436),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1461),
.B(n_1027),
.Y(n_1588)
);

INVxp67_ASAP7_75t_L g1589 ( 
.A(n_1233),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1379),
.Y(n_1590)
);

INVx4_ASAP7_75t_L g1591 ( 
.A(n_1180),
.Y(n_1591)
);

INVx6_ASAP7_75t_L g1592 ( 
.A(n_1447),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1194),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_SL g1594 ( 
.A1(n_1370),
.A2(n_1121),
.B1(n_1139),
.B2(n_1123),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1181),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1438),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1465),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1387),
.Y(n_1598)
);

INVx3_ASAP7_75t_L g1599 ( 
.A(n_1441),
.Y(n_1599)
);

BUFx6f_ASAP7_75t_L g1600 ( 
.A(n_1202),
.Y(n_1600)
);

INVx6_ASAP7_75t_L g1601 ( 
.A(n_1295),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1388),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1417),
.B(n_819),
.Y(n_1603)
);

INVx5_ASAP7_75t_L g1604 ( 
.A(n_1180),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1392),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1442),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1209),
.B(n_1205),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1393),
.Y(n_1608)
);

CKINVDCx20_ASAP7_75t_R g1609 ( 
.A(n_1173),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1394),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1397),
.Y(n_1611)
);

INVx3_ASAP7_75t_L g1612 ( 
.A(n_1443),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1420),
.B(n_819),
.Y(n_1613)
);

AOI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1180),
.A2(n_968),
.B1(n_1082),
.B2(n_1076),
.Y(n_1614)
);

INVx3_ASAP7_75t_L g1615 ( 
.A(n_1445),
.Y(n_1615)
);

INVx6_ASAP7_75t_L g1616 ( 
.A(n_1452),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1399),
.Y(n_1617)
);

BUFx8_ASAP7_75t_L g1618 ( 
.A(n_1248),
.Y(n_1618)
);

AOI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1268),
.A2(n_1082),
.B1(n_1089),
.B2(n_1087),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1470),
.B(n_1027),
.Y(n_1620)
);

INVx3_ASAP7_75t_L g1621 ( 
.A(n_1446),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1405),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1454),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1455),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1406),
.Y(n_1625)
);

AOI22x1_ASAP7_75t_SL g1626 ( 
.A1(n_1333),
.A2(n_768),
.B1(n_770),
.B2(n_767),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1323),
.A2(n_809),
.B1(n_853),
.B2(n_827),
.Y(n_1627)
);

AOI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1280),
.A2(n_1089),
.B1(n_1092),
.B2(n_1087),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1407),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1247),
.B(n_819),
.Y(n_1630)
);

BUFx6f_ASAP7_75t_L g1631 ( 
.A(n_1203),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1274),
.Y(n_1632)
);

AND2x4_ASAP7_75t_L g1633 ( 
.A(n_1472),
.B(n_1069),
.Y(n_1633)
);

AND2x6_ASAP7_75t_L g1634 ( 
.A(n_1311),
.B(n_1131),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1206),
.B(n_1072),
.Y(n_1635)
);

AND2x2_ASAP7_75t_SL g1636 ( 
.A(n_1309),
.B(n_1154),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1408),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1456),
.Y(n_1638)
);

BUFx6f_ASAP7_75t_L g1639 ( 
.A(n_1208),
.Y(n_1639)
);

INVx3_ASAP7_75t_L g1640 ( 
.A(n_1458),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1210),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1213),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1216),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1409),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1214),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1218),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1291),
.A2(n_928),
.B1(n_1096),
.B2(n_1092),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1219),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1220),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1370),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1284),
.B(n_1096),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1221),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1319),
.B(n_819),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1223),
.B(n_1073),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1224),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1231),
.Y(n_1656)
);

INVx2_ASAP7_75t_SL g1657 ( 
.A(n_1340),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1324),
.B(n_978),
.Y(n_1658)
);

BUFx8_ASAP7_75t_L g1659 ( 
.A(n_1248),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1234),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1242),
.Y(n_1661)
);

OA21x2_ASAP7_75t_L g1662 ( 
.A1(n_1250),
.A2(n_1253),
.B(n_1251),
.Y(n_1662)
);

OA21x2_ASAP7_75t_L g1663 ( 
.A1(n_1255),
.A2(n_954),
.B(n_871),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1256),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1257),
.B(n_1259),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1266),
.Y(n_1666)
);

NOR2x1_ASAP7_75t_L g1667 ( 
.A(n_1330),
.B(n_1108),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1275),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1209),
.B(n_816),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1278),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1279),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1281),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1338),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1217),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1356),
.B(n_978),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1294),
.B(n_836),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1285),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1286),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1325),
.B(n_836),
.Y(n_1679)
);

AND2x4_ASAP7_75t_L g1680 ( 
.A(n_1287),
.B(n_1077),
.Y(n_1680)
);

INVx4_ASAP7_75t_L g1681 ( 
.A(n_1172),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1288),
.B(n_1078),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1293),
.Y(n_1683)
);

BUFx6f_ASAP7_75t_L g1684 ( 
.A(n_1296),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1380),
.B(n_978),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1298),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1450),
.B(n_1373),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1302),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1304),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1355),
.A2(n_1100),
.B1(n_1102),
.B2(n_1098),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1305),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1306),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1473),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1427),
.Y(n_1694)
);

BUFx3_ASAP7_75t_L g1695 ( 
.A(n_1429),
.Y(n_1695)
);

AOI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1314),
.A2(n_1100),
.B1(n_1102),
.B2(n_1098),
.Y(n_1696)
);

INVx2_ASAP7_75t_SL g1697 ( 
.A(n_1386),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1378),
.B(n_1080),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1248),
.Y(n_1699)
);

BUFx6f_ASAP7_75t_L g1700 ( 
.A(n_1174),
.Y(n_1700)
);

INVx3_ASAP7_75t_L g1701 ( 
.A(n_1354),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1354),
.Y(n_1702)
);

INVx5_ASAP7_75t_L g1703 ( 
.A(n_1354),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1239),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1179),
.B(n_978),
.Y(n_1705)
);

INVx5_ASAP7_75t_L g1706 ( 
.A(n_1314),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1249),
.Y(n_1707)
);

AND2x4_ASAP7_75t_L g1708 ( 
.A(n_1261),
.B(n_1054),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1263),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1290),
.B(n_1111),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1422),
.Y(n_1711)
);

INVx3_ASAP7_75t_L g1712 ( 
.A(n_1183),
.Y(n_1712)
);

NOR2x1_ASAP7_75t_L g1713 ( 
.A(n_1184),
.B(n_1114),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1435),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1369),
.B(n_1105),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1190),
.B(n_978),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1193),
.Y(n_1717)
);

BUFx12f_ASAP7_75t_L g1718 ( 
.A(n_1415),
.Y(n_1718)
);

AOI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1369),
.A2(n_1449),
.B1(n_1199),
.B2(n_1201),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1449),
.A2(n_1106),
.B1(n_1109),
.B2(n_1105),
.Y(n_1720)
);

INVx4_ASAP7_75t_L g1721 ( 
.A(n_1196),
.Y(n_1721)
);

AOI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1207),
.A2(n_1109),
.B1(n_1110),
.B2(n_1106),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1226),
.B(n_1117),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1235),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1236),
.B(n_978),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1241),
.Y(n_1726)
);

BUFx3_ASAP7_75t_L g1727 ( 
.A(n_1453),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1244),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1246),
.Y(n_1729)
);

BUFx6f_ASAP7_75t_L g1730 ( 
.A(n_1258),
.Y(n_1730)
);

OA21x2_ASAP7_75t_L g1731 ( 
.A1(n_1265),
.A2(n_954),
.B(n_871),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1267),
.A2(n_1110),
.B1(n_1120),
.B2(n_1119),
.Y(n_1732)
);

INVx3_ASAP7_75t_L g1733 ( 
.A(n_1270),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1282),
.Y(n_1734)
);

BUFx6f_ASAP7_75t_L g1735 ( 
.A(n_1289),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1297),
.B(n_895),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1299),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1300),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1310),
.B(n_895),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_SL g1740 ( 
.A(n_1316),
.B(n_953),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1317),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1332),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1336),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1341),
.B(n_978),
.Y(n_1744)
);

BUFx2_ASAP7_75t_L g1745 ( 
.A(n_1217),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1343),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1345),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1353),
.B(n_1128),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_1362),
.Y(n_1749)
);

INVx3_ASAP7_75t_L g1750 ( 
.A(n_1374),
.Y(n_1750)
);

BUFx6f_ASAP7_75t_L g1751 ( 
.A(n_1375),
.Y(n_1751)
);

BUFx8_ASAP7_75t_L g1752 ( 
.A(n_1303),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1377),
.B(n_1130),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1382),
.B(n_1132),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1385),
.Y(n_1755)
);

INVx3_ASAP7_75t_L g1756 ( 
.A(n_1390),
.Y(n_1756)
);

BUFx6f_ASAP7_75t_L g1757 ( 
.A(n_1391),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1428),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1433),
.Y(n_1759)
);

INVx4_ASAP7_75t_L g1760 ( 
.A(n_1434),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1444),
.Y(n_1761)
);

INVx3_ASAP7_75t_L g1762 ( 
.A(n_1448),
.Y(n_1762)
);

INVx3_ASAP7_75t_L g1763 ( 
.A(n_1460),
.Y(n_1763)
);

OAI22xp5_ASAP7_75t_SL g1764 ( 
.A1(n_1494),
.A2(n_1398),
.B1(n_1400),
.B2(n_1383),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1665),
.B(n_1135),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_SL g1766 ( 
.A(n_1604),
.B(n_1462),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1510),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1513),
.B(n_1137),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1574),
.B(n_1464),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1475),
.B(n_1140),
.Y(n_1770)
);

BUFx8_ASAP7_75t_L g1771 ( 
.A(n_1508),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1479),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1479),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1510),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1479),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1557),
.B(n_1143),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1507),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1507),
.Y(n_1778)
);

AND2x6_ASAP7_75t_L g1779 ( 
.A(n_1701),
.B(n_1154),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1510),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1507),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1641),
.Y(n_1782)
);

BUFx6f_ASAP7_75t_L g1783 ( 
.A(n_1663),
.Y(n_1783)
);

INVxp67_ASAP7_75t_L g1784 ( 
.A(n_1492),
.Y(n_1784)
);

INVxp67_ASAP7_75t_L g1785 ( 
.A(n_1492),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1512),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1641),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1574),
.B(n_1152),
.Y(n_1788)
);

HB1xp67_ASAP7_75t_L g1789 ( 
.A(n_1491),
.Y(n_1789)
);

BUFx6f_ASAP7_75t_L g1790 ( 
.A(n_1663),
.Y(n_1790)
);

BUFx3_ASAP7_75t_L g1791 ( 
.A(n_1498),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1512),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1642),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1642),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1656),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1520),
.B(n_1162),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1557),
.B(n_1165),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_L g1798 ( 
.A(n_1589),
.B(n_1466),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1656),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1512),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1660),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1573),
.Y(n_1802)
);

OAI21x1_ASAP7_75t_L g1803 ( 
.A1(n_1531),
.A2(n_977),
.B(n_957),
.Y(n_1803)
);

INVxp67_ASAP7_75t_L g1804 ( 
.A(n_1491),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1660),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1668),
.Y(n_1806)
);

BUFx6f_ASAP7_75t_L g1807 ( 
.A(n_1663),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1573),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1668),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1580),
.B(n_1166),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1481),
.B(n_1168),
.Y(n_1811)
);

HB1xp67_ASAP7_75t_L g1812 ( 
.A(n_1480),
.Y(n_1812)
);

BUFx2_ASAP7_75t_L g1813 ( 
.A(n_1480),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1573),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1670),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_SL g1816 ( 
.A(n_1604),
.B(n_1467),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_SL g1817 ( 
.A(n_1604),
.B(n_1591),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_L g1818 ( 
.A(n_1511),
.B(n_1474),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1670),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1677),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1677),
.Y(n_1821)
);

AND2x4_ASAP7_75t_L g1822 ( 
.A(n_1665),
.B(n_1518),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1582),
.Y(n_1823)
);

BUFx6f_ASAP7_75t_L g1824 ( 
.A(n_1585),
.Y(n_1824)
);

AND2x6_ASAP7_75t_L g1825 ( 
.A(n_1701),
.B(n_1155),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1678),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1678),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1634),
.B(n_1155),
.Y(n_1828)
);

INVx3_ASAP7_75t_L g1829 ( 
.A(n_1582),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1582),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1580),
.B(n_1079),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1683),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1665),
.B(n_1153),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1683),
.Y(n_1834)
);

BUFx6f_ASAP7_75t_L g1835 ( 
.A(n_1585),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1686),
.Y(n_1836)
);

BUFx8_ASAP7_75t_L g1837 ( 
.A(n_1539),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_SL g1838 ( 
.A(n_1681),
.B(n_1415),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1517),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1634),
.B(n_949),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1686),
.Y(n_1841)
);

BUFx6f_ASAP7_75t_L g1842 ( 
.A(n_1585),
.Y(n_1842)
);

AND2x4_ASAP7_75t_L g1843 ( 
.A(n_1518),
.B(n_234),
.Y(n_1843)
);

CKINVDCx16_ASAP7_75t_R g1844 ( 
.A(n_1609),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1688),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1517),
.Y(n_1846)
);

AND2x4_ASAP7_75t_L g1847 ( 
.A(n_1525),
.B(n_239),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1517),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1688),
.Y(n_1849)
);

BUFx6f_ASAP7_75t_L g1850 ( 
.A(n_1585),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1552),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_SL g1852 ( 
.A(n_1604),
.B(n_1178),
.Y(n_1852)
);

BUFx3_ASAP7_75t_L g1853 ( 
.A(n_1498),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1634),
.B(n_949),
.Y(n_1854)
);

BUFx2_ASAP7_75t_L g1855 ( 
.A(n_1609),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1689),
.Y(n_1856)
);

INVx3_ASAP7_75t_L g1857 ( 
.A(n_1552),
.Y(n_1857)
);

BUFx6f_ASAP7_75t_L g1858 ( 
.A(n_1600),
.Y(n_1858)
);

INVx3_ASAP7_75t_L g1859 ( 
.A(n_1552),
.Y(n_1859)
);

HB1xp67_ASAP7_75t_L g1860 ( 
.A(n_1669),
.Y(n_1860)
);

BUFx6f_ASAP7_75t_L g1861 ( 
.A(n_1600),
.Y(n_1861)
);

BUFx6f_ASAP7_75t_L g1862 ( 
.A(n_1600),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1691),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1476),
.Y(n_1864)
);

INVxp67_ASAP7_75t_L g1865 ( 
.A(n_1607),
.Y(n_1865)
);

INVx1_ASAP7_75t_SL g1866 ( 
.A(n_1679),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1476),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1587),
.Y(n_1868)
);

INVx1_ASAP7_75t_SL g1869 ( 
.A(n_1736),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1691),
.Y(n_1870)
);

HB1xp67_ASAP7_75t_L g1871 ( 
.A(n_1587),
.Y(n_1871)
);

INVx3_ASAP7_75t_L g1872 ( 
.A(n_1731),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1692),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1485),
.Y(n_1874)
);

INVx3_ASAP7_75t_L g1875 ( 
.A(n_1731),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1485),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_SL g1877 ( 
.A(n_1591),
.B(n_1178),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1662),
.B(n_1079),
.Y(n_1878)
);

INVx3_ASAP7_75t_L g1879 ( 
.A(n_1731),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1692),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1694),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1634),
.B(n_949),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1694),
.Y(n_1883)
);

BUFx6f_ASAP7_75t_L g1884 ( 
.A(n_1600),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1635),
.Y(n_1885)
);

AND2x4_ASAP7_75t_L g1886 ( 
.A(n_1525),
.B(n_240),
.Y(n_1886)
);

OAI21x1_ASAP7_75t_L g1887 ( 
.A1(n_1603),
.A2(n_977),
.B(n_957),
.Y(n_1887)
);

OA21x2_ASAP7_75t_L g1888 ( 
.A1(n_1613),
.A2(n_506),
.B(n_505),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1635),
.Y(n_1889)
);

BUFx6f_ASAP7_75t_L g1890 ( 
.A(n_1631),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1486),
.Y(n_1891)
);

BUFx6f_ASAP7_75t_L g1892 ( 
.A(n_1631),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1635),
.Y(n_1893)
);

OAI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1591),
.A2(n_1687),
.B1(n_1636),
.B2(n_1592),
.Y(n_1894)
);

AND2x4_ASAP7_75t_L g1895 ( 
.A(n_1525),
.B(n_241),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1478),
.B(n_242),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1634),
.B(n_1002),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1654),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1654),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1654),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_SL g1901 ( 
.A(n_1636),
.B(n_1292),
.Y(n_1901)
);

NAND2xp33_ASAP7_75t_L g1902 ( 
.A(n_1483),
.B(n_506),
.Y(n_1902)
);

INVx3_ASAP7_75t_L g1903 ( 
.A(n_1554),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1680),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1486),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1680),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1662),
.B(n_940),
.Y(n_1907)
);

BUFx2_ASAP7_75t_L g1908 ( 
.A(n_1650),
.Y(n_1908)
);

INVx3_ASAP7_75t_L g1909 ( 
.A(n_1554),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1680),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1682),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1682),
.Y(n_1912)
);

HB1xp67_ASAP7_75t_L g1913 ( 
.A(n_1542),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1495),
.Y(n_1914)
);

INVx3_ASAP7_75t_L g1915 ( 
.A(n_1554),
.Y(n_1915)
);

INVx3_ASAP7_75t_L g1916 ( 
.A(n_1554),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1682),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1633),
.Y(n_1918)
);

BUFx6f_ASAP7_75t_L g1919 ( 
.A(n_1631),
.Y(n_1919)
);

INVxp67_ASAP7_75t_L g1920 ( 
.A(n_1543),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_SL g1921 ( 
.A(n_1676),
.B(n_1292),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1705),
.B(n_1002),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1633),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1633),
.Y(n_1924)
);

INVx3_ASAP7_75t_L g1925 ( 
.A(n_1563),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1495),
.Y(n_1926)
);

OAI21x1_ASAP7_75t_L g1927 ( 
.A1(n_1500),
.A2(n_1630),
.B(n_1653),
.Y(n_1927)
);

INVxp67_ASAP7_75t_L g1928 ( 
.A(n_1543),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1478),
.B(n_244),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1477),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1493),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1662),
.B(n_1085),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1496),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1716),
.B(n_1002),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1497),
.Y(n_1935)
);

BUFx6f_ASAP7_75t_L g1936 ( 
.A(n_1631),
.Y(n_1936)
);

BUFx2_ASAP7_75t_L g1937 ( 
.A(n_1711),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1502),
.Y(n_1938)
);

HB1xp67_ASAP7_75t_L g1939 ( 
.A(n_1711),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1506),
.Y(n_1940)
);

NAND3xp33_ASAP7_75t_L g1941 ( 
.A(n_1732),
.B(n_1414),
.C(n_1395),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1514),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1515),
.Y(n_1943)
);

INVxp67_ASAP7_75t_L g1944 ( 
.A(n_1484),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1497),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1739),
.B(n_1085),
.Y(n_1946)
);

INVxp67_ASAP7_75t_L g1947 ( 
.A(n_1715),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1499),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1516),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1519),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1499),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1521),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1725),
.B(n_1066),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1698),
.B(n_958),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1698),
.B(n_980),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1528),
.Y(n_1956)
);

AND2x6_ASAP7_75t_L g1957 ( 
.A(n_1699),
.B(n_811),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1744),
.B(n_1066),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1621),
.B(n_1623),
.Y(n_1959)
);

NAND2xp33_ASAP7_75t_SL g1960 ( 
.A(n_1632),
.B(n_1123),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1532),
.Y(n_1961)
);

INVx3_ASAP7_75t_L g1962 ( 
.A(n_1563),
.Y(n_1962)
);

BUFx12f_ASAP7_75t_L g1963 ( 
.A(n_1618),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1534),
.Y(n_1964)
);

OAI22xp5_ASAP7_75t_SL g1965 ( 
.A1(n_1565),
.A2(n_1398),
.B1(n_1400),
.B2(n_1383),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1504),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1535),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1536),
.Y(n_1968)
);

BUFx6f_ASAP7_75t_L g1969 ( 
.A(n_1639),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1537),
.Y(n_1970)
);

NOR2xp33_ASAP7_75t_SL g1971 ( 
.A(n_1681),
.B(n_1418),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1538),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1621),
.B(n_1066),
.Y(n_1973)
);

BUFx6f_ASAP7_75t_L g1974 ( 
.A(n_1639),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1556),
.Y(n_1975)
);

NAND2x1_ASAP7_75t_L g1976 ( 
.A(n_1503),
.B(n_1524),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1561),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1567),
.Y(n_1978)
);

BUFx3_ASAP7_75t_L g1979 ( 
.A(n_1498),
.Y(n_1979)
);

AND2x4_ASAP7_75t_L g1980 ( 
.A(n_1488),
.B(n_1490),
.Y(n_1980)
);

AND2x4_ASAP7_75t_L g1981 ( 
.A(n_1488),
.B(n_246),
.Y(n_1981)
);

BUFx6f_ASAP7_75t_L g1982 ( 
.A(n_1639),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1568),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1570),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1578),
.Y(n_1985)
);

OAI21x1_ASAP7_75t_L g1986 ( 
.A1(n_1658),
.A2(n_514),
.B(n_510),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1504),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1583),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1586),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1590),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1598),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1602),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1505),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1505),
.Y(n_1994)
);

HB1xp67_ASAP7_75t_L g1995 ( 
.A(n_1708),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1509),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1605),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1608),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1610),
.Y(n_1999)
);

HB1xp67_ASAP7_75t_L g2000 ( 
.A(n_1708),
.Y(n_2000)
);

BUFx6f_ASAP7_75t_L g2001 ( 
.A(n_1639),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1698),
.B(n_1013),
.Y(n_2002)
);

HB1xp67_ASAP7_75t_L g2003 ( 
.A(n_1708),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1611),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_1530),
.Y(n_2005)
);

BUFx2_ASAP7_75t_L g2006 ( 
.A(n_1541),
.Y(n_2006)
);

CKINVDCx5p33_ASAP7_75t_R g2007 ( 
.A(n_1530),
.Y(n_2007)
);

BUFx2_ASAP7_75t_L g2008 ( 
.A(n_1584),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1509),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1546),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1546),
.Y(n_2011)
);

AND2x4_ASAP7_75t_L g2012 ( 
.A(n_1490),
.B(n_247),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1617),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1548),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1622),
.Y(n_2015)
);

INVx3_ASAP7_75t_L g2016 ( 
.A(n_1563),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1548),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1549),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1625),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_SL g2020 ( 
.A(n_1675),
.B(n_1685),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1632),
.B(n_1395),
.Y(n_2021)
);

INVxp67_ASAP7_75t_L g2022 ( 
.A(n_1715),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1629),
.Y(n_2023)
);

BUFx2_ASAP7_75t_L g2024 ( 
.A(n_1657),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1621),
.B(n_510),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1549),
.Y(n_2026)
);

AND2x6_ASAP7_75t_L g2027 ( 
.A(n_1667),
.B(n_813),
.Y(n_2027)
);

HB1xp67_ASAP7_75t_L g2028 ( 
.A(n_1657),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1637),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1555),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1644),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1555),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1645),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1576),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1646),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1576),
.Y(n_2036)
);

INVx4_ASAP7_75t_L g2037 ( 
.A(n_1526),
.Y(n_2037)
);

BUFx6f_ASAP7_75t_L g2038 ( 
.A(n_1684),
.Y(n_2038)
);

INVx3_ASAP7_75t_L g2039 ( 
.A(n_1563),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1673),
.B(n_1414),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1581),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_SL g2042 ( 
.A(n_1684),
.B(n_1418),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1581),
.Y(n_2043)
);

AND2x2_ASAP7_75t_SL g2044 ( 
.A(n_1651),
.B(n_1352),
.Y(n_2044)
);

INVx1_ASAP7_75t_SL g2045 ( 
.A(n_1745),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1648),
.Y(n_2046)
);

NAND2xp33_ASAP7_75t_SL g2047 ( 
.A(n_1673),
.B(n_1139),
.Y(n_2047)
);

BUFx6f_ASAP7_75t_L g2048 ( 
.A(n_1684),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1593),
.Y(n_2049)
);

BUFx2_ASAP7_75t_L g2050 ( 
.A(n_1697),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1593),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1649),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_SL g2053 ( 
.A(n_1684),
.B(n_514),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1652),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1655),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1524),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1524),
.Y(n_2057)
);

INVx3_ASAP7_75t_L g2058 ( 
.A(n_1564),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1661),
.Y(n_2059)
);

NAND2xp33_ASAP7_75t_SL g2060 ( 
.A(n_1627),
.B(n_1145),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_1697),
.B(n_839),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1664),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1768),
.B(n_1651),
.Y(n_2063)
);

INVx4_ASAP7_75t_L g2064 ( 
.A(n_1824),
.Y(n_2064)
);

NOR2xp33_ASAP7_75t_L g2065 ( 
.A(n_1947),
.B(n_2022),
.Y(n_2065)
);

AND2x4_ASAP7_75t_L g2066 ( 
.A(n_1980),
.B(n_1540),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1788),
.B(n_1811),
.Y(n_2067)
);

NAND2xp33_ASAP7_75t_L g2068 ( 
.A(n_1779),
.B(n_1483),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1772),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1864),
.Y(n_2070)
);

AOI22xp33_ASAP7_75t_L g2071 ( 
.A1(n_1878),
.A2(n_1562),
.B1(n_1483),
.B2(n_1487),
.Y(n_2071)
);

BUFx6f_ASAP7_75t_L g2072 ( 
.A(n_1824),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_1831),
.B(n_1704),
.Y(n_2073)
);

NOR2xp33_ASAP7_75t_L g2074 ( 
.A(n_1769),
.B(n_1712),
.Y(n_2074)
);

INVx3_ASAP7_75t_L g2075 ( 
.A(n_1824),
.Y(n_2075)
);

AND2x2_ASAP7_75t_SL g2076 ( 
.A(n_2044),
.B(n_1700),
.Y(n_2076)
);

AOI22xp5_ASAP7_75t_L g2077 ( 
.A1(n_1894),
.A2(n_1483),
.B1(n_1592),
.B2(n_1754),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1773),
.Y(n_2078)
);

INVx3_ASAP7_75t_L g2079 ( 
.A(n_1824),
.Y(n_2079)
);

INVx3_ASAP7_75t_L g2080 ( 
.A(n_1835),
.Y(n_2080)
);

NOR2xp33_ASAP7_75t_L g2081 ( 
.A(n_1769),
.B(n_1798),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_1864),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1775),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1777),
.Y(n_2084)
);

INVx4_ASAP7_75t_L g2085 ( 
.A(n_1835),
.Y(n_2085)
);

NOR3xp33_ASAP7_75t_L g2086 ( 
.A(n_1901),
.B(n_1647),
.C(n_1754),
.Y(n_2086)
);

INVx3_ASAP7_75t_L g2087 ( 
.A(n_1835),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_1831),
.B(n_1704),
.Y(n_2088)
);

AND2x4_ASAP7_75t_L g2089 ( 
.A(n_1980),
.B(n_1540),
.Y(n_2089)
);

AND2x4_ASAP7_75t_L g2090 ( 
.A(n_1980),
.B(n_1540),
.Y(n_2090)
);

AND2x4_ASAP7_75t_L g2091 ( 
.A(n_1791),
.B(n_1695),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_1770),
.B(n_1763),
.Y(n_2092)
);

CKINVDCx20_ASAP7_75t_R g2093 ( 
.A(n_1844),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1778),
.Y(n_2094)
);

INVx3_ASAP7_75t_L g2095 ( 
.A(n_1835),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_1867),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1781),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_1770),
.B(n_1866),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1878),
.B(n_1623),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_SL g2100 ( 
.A(n_1847),
.B(n_1706),
.Y(n_2100)
);

INVx2_ASAP7_75t_SL g2101 ( 
.A(n_1789),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_1946),
.B(n_1763),
.Y(n_2102)
);

NOR2x1p5_ASAP7_75t_L g2103 ( 
.A(n_1963),
.B(n_1762),
.Y(n_2103)
);

AND2x4_ASAP7_75t_L g2104 ( 
.A(n_1791),
.B(n_1695),
.Y(n_2104)
);

INVx2_ASAP7_75t_SL g2105 ( 
.A(n_2028),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2034),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1907),
.B(n_1623),
.Y(n_2107)
);

NAND2xp33_ASAP7_75t_L g2108 ( 
.A(n_1779),
.B(n_1700),
.Y(n_2108)
);

BUFx2_ASAP7_75t_L g2109 ( 
.A(n_1908),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2034),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2036),
.Y(n_2111)
);

NOR2xp33_ASAP7_75t_L g2112 ( 
.A(n_1798),
.B(n_1712),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1907),
.B(n_1640),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_SL g2114 ( 
.A(n_1847),
.B(n_1706),
.Y(n_2114)
);

INVxp67_ASAP7_75t_L g2115 ( 
.A(n_2024),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_SL g2116 ( 
.A(n_1847),
.B(n_1706),
.Y(n_2116)
);

INVx3_ASAP7_75t_L g2117 ( 
.A(n_1842),
.Y(n_2117)
);

INVx3_ASAP7_75t_L g2118 ( 
.A(n_1842),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2036),
.Y(n_2119)
);

AND2x4_ASAP7_75t_L g2120 ( 
.A(n_1853),
.B(n_1699),
.Y(n_2120)
);

INVx5_ASAP7_75t_L g2121 ( 
.A(n_1783),
.Y(n_2121)
);

INVx2_ASAP7_75t_SL g2122 ( 
.A(n_2050),
.Y(n_2122)
);

INVxp33_ASAP7_75t_L g2123 ( 
.A(n_1812),
.Y(n_2123)
);

NAND2xp33_ASAP7_75t_L g2124 ( 
.A(n_1779),
.B(n_1483),
.Y(n_2124)
);

BUFx6f_ASAP7_75t_SL g2125 ( 
.A(n_2044),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1796),
.B(n_1640),
.Y(n_2126)
);

INVxp67_ASAP7_75t_L g2127 ( 
.A(n_1937),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1886),
.B(n_1640),
.Y(n_2128)
);

INVx3_ASAP7_75t_L g2129 ( 
.A(n_1842),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_1886),
.B(n_1599),
.Y(n_2130)
);

CKINVDCx20_ASAP7_75t_R g2131 ( 
.A(n_1764),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1867),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_1886),
.B(n_1599),
.Y(n_2133)
);

NAND2x1p5_ASAP7_75t_L g2134 ( 
.A(n_1895),
.B(n_1700),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2041),
.Y(n_2135)
);

AND3x4_ASAP7_75t_L g2136 ( 
.A(n_1765),
.B(n_1713),
.C(n_1710),
.Y(n_2136)
);

INVx3_ASAP7_75t_L g2137 ( 
.A(n_1842),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1874),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1874),
.Y(n_2139)
);

INVx1_ASAP7_75t_SL g2140 ( 
.A(n_2045),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_1895),
.B(n_1612),
.Y(n_2141)
);

NOR2xp33_ASAP7_75t_L g2142 ( 
.A(n_1865),
.B(n_1869),
.Y(n_2142)
);

NAND2xp33_ASAP7_75t_L g2143 ( 
.A(n_1779),
.B(n_1700),
.Y(n_2143)
);

AOI22xp33_ASAP7_75t_L g2144 ( 
.A1(n_1932),
.A2(n_1895),
.B1(n_1875),
.B2(n_1879),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_1876),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_1932),
.B(n_1612),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_1946),
.B(n_1762),
.Y(n_2147)
);

BUFx4f_ASAP7_75t_L g2148 ( 
.A(n_1963),
.Y(n_2148)
);

BUFx8_ASAP7_75t_SL g2149 ( 
.A(n_2005),
.Y(n_2149)
);

INVx3_ASAP7_75t_L g2150 ( 
.A(n_1850),
.Y(n_2150)
);

BUFx10_ASAP7_75t_L g2151 ( 
.A(n_1818),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2041),
.Y(n_2152)
);

INVx3_ASAP7_75t_L g2153 ( 
.A(n_1850),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2043),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_SL g2155 ( 
.A(n_1850),
.B(n_1706),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2043),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2049),
.Y(n_2157)
);

INVx3_ASAP7_75t_L g2158 ( 
.A(n_1850),
.Y(n_2158)
);

NOR2xp33_ASAP7_75t_L g2159 ( 
.A(n_1818),
.B(n_1712),
.Y(n_2159)
);

AND2x6_ASAP7_75t_L g2160 ( 
.A(n_1802),
.B(n_1702),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1922),
.B(n_1615),
.Y(n_2161)
);

BUFx2_ASAP7_75t_L g2162 ( 
.A(n_1855),
.Y(n_2162)
);

INVx3_ASAP7_75t_L g2163 ( 
.A(n_1858),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_1876),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1891),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2049),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2051),
.Y(n_2167)
);

INVx4_ASAP7_75t_L g2168 ( 
.A(n_1858),
.Y(n_2168)
);

INVx5_ASAP7_75t_L g2169 ( 
.A(n_1783),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_SL g2170 ( 
.A(n_1858),
.B(n_1730),
.Y(n_2170)
);

NOR2xp33_ASAP7_75t_L g2171 ( 
.A(n_1913),
.B(n_1733),
.Y(n_2171)
);

INVx2_ASAP7_75t_SL g2172 ( 
.A(n_1939),
.Y(n_2172)
);

INVxp67_ASAP7_75t_L g2173 ( 
.A(n_1813),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2051),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_SL g2175 ( 
.A(n_1858),
.B(n_1730),
.Y(n_2175)
);

OR2x6_ASAP7_75t_L g2176 ( 
.A(n_1804),
.B(n_1601),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1782),
.Y(n_2177)
);

INVx4_ASAP7_75t_L g2178 ( 
.A(n_1861),
.Y(n_2178)
);

BUFx3_ASAP7_75t_L g2179 ( 
.A(n_1853),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1787),
.Y(n_2180)
);

BUFx3_ASAP7_75t_L g2181 ( 
.A(n_1979),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1793),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1794),
.Y(n_2183)
);

NOR2xp33_ASAP7_75t_L g2184 ( 
.A(n_1860),
.B(n_1733),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_1934),
.B(n_1615),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_1953),
.B(n_1482),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2061),
.B(n_1733),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1795),
.Y(n_2188)
);

INVx3_ASAP7_75t_L g2189 ( 
.A(n_1861),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1799),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1801),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_SL g2192 ( 
.A(n_1861),
.B(n_1730),
.Y(n_2192)
);

BUFx5_ASAP7_75t_L g2193 ( 
.A(n_1779),
.Y(n_2193)
);

INVx5_ASAP7_75t_L g2194 ( 
.A(n_1783),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1805),
.Y(n_2195)
);

AND2x6_ASAP7_75t_L g2196 ( 
.A(n_1802),
.B(n_1808),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1806),
.Y(n_2197)
);

INVx3_ASAP7_75t_L g2198 ( 
.A(n_1861),
.Y(n_2198)
);

BUFx10_ASAP7_75t_L g2199 ( 
.A(n_1765),
.Y(n_2199)
);

XNOR2xp5_ASAP7_75t_L g2200 ( 
.A(n_2006),
.B(n_1173),
.Y(n_2200)
);

NOR2xp33_ASAP7_75t_L g2201 ( 
.A(n_1784),
.B(n_1749),
.Y(n_2201)
);

INVxp67_ASAP7_75t_SL g2202 ( 
.A(n_1783),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_1958),
.B(n_1501),
.Y(n_2203)
);

INVx3_ASAP7_75t_L g2204 ( 
.A(n_1862),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_1776),
.B(n_1748),
.Y(n_2205)
);

INVx3_ASAP7_75t_L g2206 ( 
.A(n_1862),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_1891),
.Y(n_2207)
);

AOI22xp5_ASAP7_75t_L g2208 ( 
.A1(n_1828),
.A2(n_1592),
.B1(n_1710),
.B2(n_1723),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_1776),
.B(n_1666),
.Y(n_2209)
);

OAI22xp5_ASAP7_75t_L g2210 ( 
.A1(n_1959),
.A2(n_1734),
.B1(n_1742),
.B2(n_1726),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_1905),
.Y(n_2211)
);

NOR2xp33_ASAP7_75t_L g2212 ( 
.A(n_1785),
.B(n_1749),
.Y(n_2212)
);

INVx3_ASAP7_75t_L g2213 ( 
.A(n_1862),
.Y(n_2213)
);

CKINVDCx5p33_ASAP7_75t_R g2214 ( 
.A(n_2005),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_1797),
.B(n_1671),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_1905),
.Y(n_2216)
);

AND2x4_ASAP7_75t_L g2217 ( 
.A(n_1979),
.B(n_1702),
.Y(n_2217)
);

AOI22xp33_ASAP7_75t_L g2218 ( 
.A1(n_1872),
.A2(n_1562),
.B1(n_1606),
.B2(n_1596),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1809),
.Y(n_2219)
);

CKINVDCx5p33_ASAP7_75t_R g2220 ( 
.A(n_2007),
.Y(n_2220)
);

AOI22xp33_ASAP7_75t_L g2221 ( 
.A1(n_1872),
.A2(n_1562),
.B1(n_1606),
.B2(n_1596),
.Y(n_2221)
);

NOR2x1p5_ASAP7_75t_L g2222 ( 
.A(n_1941),
.B(n_1749),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1815),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1819),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_1797),
.B(n_1672),
.Y(n_2225)
);

OAI22x1_ASAP7_75t_SL g2226 ( 
.A1(n_2007),
.A2(n_1333),
.B1(n_1191),
.B2(n_1211),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1820),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_SL g2228 ( 
.A(n_1862),
.B(n_1730),
.Y(n_2228)
);

INVx5_ASAP7_75t_L g2229 ( 
.A(n_1790),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1821),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_1810),
.B(n_1726),
.Y(n_2231)
);

INVx5_ASAP7_75t_L g2232 ( 
.A(n_1790),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_1810),
.B(n_1734),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_1826),
.B(n_1742),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1827),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_1914),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_1914),
.Y(n_2237)
);

NOR2xp33_ASAP7_75t_L g2238 ( 
.A(n_1901),
.B(n_1750),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_SL g2239 ( 
.A(n_1884),
.B(n_1735),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1832),
.Y(n_2240)
);

NOR2x1p5_ASAP7_75t_L g2241 ( 
.A(n_1954),
.B(n_1750),
.Y(n_2241)
);

INVx5_ASAP7_75t_L g2242 ( 
.A(n_1790),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_1834),
.B(n_1758),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_SL g2244 ( 
.A(n_1884),
.B(n_1735),
.Y(n_2244)
);

AOI22xp33_ASAP7_75t_L g2245 ( 
.A1(n_1872),
.A2(n_1638),
.B1(n_1624),
.B2(n_1588),
.Y(n_2245)
);

AOI21x1_ASAP7_75t_L g2246 ( 
.A1(n_1976),
.A2(n_1595),
.B(n_1624),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_1836),
.B(n_1758),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2061),
.B(n_2021),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_1926),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1841),
.Y(n_2250)
);

NOR2x1p5_ASAP7_75t_L g2251 ( 
.A(n_1954),
.B(n_1750),
.Y(n_2251)
);

INVx3_ASAP7_75t_L g2252 ( 
.A(n_1884),
.Y(n_2252)
);

CKINVDCx5p33_ASAP7_75t_R g2253 ( 
.A(n_1771),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_1926),
.Y(n_2254)
);

NAND3xp33_ASAP7_75t_L g2255 ( 
.A(n_1920),
.B(n_1628),
.C(n_1619),
.Y(n_2255)
);

INVx3_ASAP7_75t_L g2256 ( 
.A(n_1884),
.Y(n_2256)
);

INVx3_ASAP7_75t_L g2257 ( 
.A(n_1890),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_1845),
.B(n_1710),
.Y(n_2258)
);

BUFx3_ASAP7_75t_L g2259 ( 
.A(n_1822),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_1849),
.B(n_1595),
.Y(n_2260)
);

NAND2xp33_ASAP7_75t_L g2261 ( 
.A(n_1779),
.B(n_1735),
.Y(n_2261)
);

AND3x2_ASAP7_75t_L g2262 ( 
.A(n_1838),
.B(n_1437),
.C(n_1569),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_1935),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_2021),
.B(n_1756),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1935),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1856),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1945),
.Y(n_2267)
);

NAND2xp33_ASAP7_75t_L g2268 ( 
.A(n_1825),
.B(n_1735),
.Y(n_2268)
);

INVx1_ASAP7_75t_SL g2269 ( 
.A(n_2040),
.Y(n_2269)
);

BUFx3_ASAP7_75t_L g2270 ( 
.A(n_1822),
.Y(n_2270)
);

AOI22xp33_ASAP7_75t_L g2271 ( 
.A1(n_1875),
.A2(n_1638),
.B1(n_1588),
.B2(n_1620),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_1863),
.B(n_1723),
.Y(n_2272)
);

AOI22xp33_ASAP7_75t_L g2273 ( 
.A1(n_1875),
.A2(n_1588),
.B1(n_1620),
.B2(n_1560),
.Y(n_2273)
);

NAND2x1p5_ASAP7_75t_L g2274 ( 
.A(n_1890),
.B(n_1751),
.Y(n_2274)
);

INVx2_ASAP7_75t_SL g2275 ( 
.A(n_1765),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1870),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_SL g2277 ( 
.A(n_1890),
.B(n_1751),
.Y(n_2277)
);

INVx2_ASAP7_75t_SL g2278 ( 
.A(n_1833),
.Y(n_2278)
);

INVx5_ASAP7_75t_L g2279 ( 
.A(n_1790),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_1873),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_1880),
.Y(n_2281)
);

OR2x6_ASAP7_75t_L g2282 ( 
.A(n_1965),
.B(n_1601),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1881),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_2040),
.B(n_1955),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_1883),
.B(n_1723),
.Y(n_2285)
);

AND2x2_ASAP7_75t_L g2286 ( 
.A(n_1955),
.B(n_1756),
.Y(n_2286)
);

BUFx8_ASAP7_75t_SL g2287 ( 
.A(n_2008),
.Y(n_2287)
);

INVx1_ASAP7_75t_SL g2288 ( 
.A(n_2002),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_1945),
.Y(n_2289)
);

BUFx3_ASAP7_75t_L g2290 ( 
.A(n_1822),
.Y(n_2290)
);

OR2x2_ASAP7_75t_L g2291 ( 
.A(n_1928),
.B(n_1714),
.Y(n_2291)
);

INVx4_ASAP7_75t_L g2292 ( 
.A(n_1890),
.Y(n_2292)
);

AOI22xp33_ASAP7_75t_L g2293 ( 
.A1(n_1879),
.A2(n_1620),
.B1(n_1560),
.B2(n_1575),
.Y(n_2293)
);

NOR2xp33_ASAP7_75t_L g2294 ( 
.A(n_1921),
.B(n_1756),
.Y(n_2294)
);

CKINVDCx20_ASAP7_75t_R g2295 ( 
.A(n_1771),
.Y(n_2295)
);

OAI22xp33_ASAP7_75t_L g2296 ( 
.A1(n_1885),
.A2(n_1757),
.B1(n_1751),
.B2(n_1545),
.Y(n_2296)
);

NOR2xp33_ASAP7_75t_L g2297 ( 
.A(n_1921),
.B(n_1868),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_SL g2298 ( 
.A(n_1892),
.B(n_1751),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_1948),
.Y(n_2299)
);

INVx3_ASAP7_75t_L g2300 ( 
.A(n_1892),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_1930),
.B(n_1753),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_1948),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_2002),
.B(n_1757),
.Y(n_2303)
);

INVxp67_ASAP7_75t_SL g2304 ( 
.A(n_1807),
.Y(n_2304)
);

BUFx2_ASAP7_75t_L g2305 ( 
.A(n_1771),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_1951),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_1951),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_1966),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_1931),
.B(n_1753),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_1966),
.Y(n_2310)
);

INVx5_ASAP7_75t_L g2311 ( 
.A(n_1807),
.Y(n_2311)
);

AND2x2_ASAP7_75t_SL g2312 ( 
.A(n_1902),
.B(n_1757),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_1933),
.B(n_1753),
.Y(n_2313)
);

OR2x2_ASAP7_75t_L g2314 ( 
.A(n_1871),
.B(n_1690),
.Y(n_2314)
);

INVx4_ASAP7_75t_L g2315 ( 
.A(n_1892),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_1938),
.B(n_1693),
.Y(n_2316)
);

NOR2xp33_ASAP7_75t_SL g2317 ( 
.A(n_1971),
.B(n_1547),
.Y(n_2317)
);

NOR2xp33_ASAP7_75t_L g2318 ( 
.A(n_1944),
.B(n_1681),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_1987),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_1987),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_1940),
.B(n_1597),
.Y(n_2321)
);

NAND3xp33_ASAP7_75t_L g2322 ( 
.A(n_2060),
.B(n_1722),
.C(n_1720),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_1942),
.B(n_1597),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_1993),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_1943),
.B(n_1717),
.Y(n_2325)
);

INVxp33_ASAP7_75t_L g2326 ( 
.A(n_1995),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_1949),
.B(n_1724),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_1950),
.B(n_1952),
.Y(n_2328)
);

BUFx3_ASAP7_75t_L g2329 ( 
.A(n_1896),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2000),
.B(n_1757),
.Y(n_2330)
);

INVx3_ASAP7_75t_L g2331 ( 
.A(n_1892),
.Y(n_2331)
);

INVx4_ASAP7_75t_L g2332 ( 
.A(n_1919),
.Y(n_2332)
);

NOR2xp33_ASAP7_75t_L g2333 ( 
.A(n_2003),
.B(n_1721),
.Y(n_2333)
);

INVx3_ASAP7_75t_L g2334 ( 
.A(n_1919),
.Y(n_2334)
);

INVx2_ASAP7_75t_SL g2335 ( 
.A(n_1833),
.Y(n_2335)
);

BUFx2_ASAP7_75t_L g2336 ( 
.A(n_1837),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_SL g2337 ( 
.A(n_1919),
.B(n_1721),
.Y(n_2337)
);

BUFx10_ASAP7_75t_L g2338 ( 
.A(n_1833),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2042),
.B(n_1727),
.Y(n_2339)
);

OAI22xp33_ASAP7_75t_L g2340 ( 
.A1(n_1889),
.A2(n_1558),
.B1(n_1614),
.B2(n_1544),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_1993),
.Y(n_2341)
);

AOI22xp33_ASAP7_75t_L g2342 ( 
.A1(n_1879),
.A2(n_1560),
.B1(n_1575),
.B2(n_1161),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_1994),
.Y(n_2343)
);

INVx4_ASAP7_75t_L g2344 ( 
.A(n_1919),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_1994),
.Y(n_2345)
);

BUFx10_ASAP7_75t_L g2346 ( 
.A(n_1896),
.Y(n_2346)
);

INVx3_ASAP7_75t_L g2347 ( 
.A(n_1936),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_1996),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_1996),
.Y(n_2349)
);

AOI22xp33_ASAP7_75t_L g2350 ( 
.A1(n_1808),
.A2(n_1575),
.B1(n_1161),
.B2(n_1145),
.Y(n_2350)
);

AO22x2_ASAP7_75t_L g2351 ( 
.A1(n_1877),
.A2(n_1729),
.B1(n_1737),
.B2(n_1728),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2009),
.Y(n_2352)
);

NOR2xp33_ASAP7_75t_L g2353 ( 
.A(n_1956),
.B(n_1721),
.Y(n_2353)
);

BUFx3_ASAP7_75t_L g2354 ( 
.A(n_1896),
.Y(n_2354)
);

INVx2_ASAP7_75t_SL g2355 ( 
.A(n_1961),
.Y(n_2355)
);

NAND2xp33_ASAP7_75t_SL g2356 ( 
.A(n_1843),
.B(n_1760),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2009),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_2010),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_1964),
.B(n_1738),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_2010),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_1967),
.B(n_1741),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_2011),
.Y(n_2362)
);

INVx3_ASAP7_75t_L g2363 ( 
.A(n_1936),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2011),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2014),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_1968),
.B(n_1743),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2070),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2106),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2110),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_SL g2370 ( 
.A(n_2159),
.B(n_2112),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2063),
.B(n_1843),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2070),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_2082),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2082),
.Y(n_2374)
);

NOR2xp33_ASAP7_75t_L g2375 ( 
.A(n_2081),
.B(n_1547),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2111),
.Y(n_2376)
);

INVxp67_ASAP7_75t_L g2377 ( 
.A(n_2109),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2119),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2135),
.Y(n_2379)
);

OAI21xp33_ASAP7_75t_L g2380 ( 
.A1(n_2081),
.A2(n_1696),
.B(n_1674),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_SL g2381 ( 
.A(n_2112),
.B(n_1760),
.Y(n_2381)
);

AND2x2_ASAP7_75t_L g2382 ( 
.A(n_2098),
.B(n_2073),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2067),
.B(n_1829),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2152),
.Y(n_2384)
);

NOR2xp33_ASAP7_75t_L g2385 ( 
.A(n_2065),
.B(n_1643),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2074),
.B(n_1829),
.Y(n_2386)
);

CKINVDCx5p33_ASAP7_75t_R g2387 ( 
.A(n_2149),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2074),
.B(n_1829),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2202),
.B(n_1857),
.Y(n_2389)
);

BUFx6f_ASAP7_75t_L g2390 ( 
.A(n_2072),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_2096),
.Y(n_2391)
);

NAND3xp33_ASAP7_75t_L g2392 ( 
.A(n_2086),
.B(n_1972),
.C(n_1970),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2154),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2156),
.Y(n_2394)
);

NOR2xp33_ASAP7_75t_L g2395 ( 
.A(n_2065),
.B(n_2205),
.Y(n_2395)
);

OR2x2_ASAP7_75t_L g2396 ( 
.A(n_2269),
.B(n_1643),
.Y(n_2396)
);

NAND2xp33_ASAP7_75t_L g2397 ( 
.A(n_2134),
.B(n_1825),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_SL g2398 ( 
.A(n_2092),
.B(n_1727),
.Y(n_2398)
);

BUFx6f_ASAP7_75t_SL g2399 ( 
.A(n_2176),
.Y(n_2399)
);

AO221x1_ASAP7_75t_L g2400 ( 
.A1(n_2296),
.A2(n_1594),
.B1(n_1755),
.B2(n_1747),
.C(n_1746),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2157),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2166),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_SL g2403 ( 
.A(n_2147),
.B(n_1719),
.Y(n_2403)
);

NOR2xp33_ASAP7_75t_L g2404 ( 
.A(n_2231),
.B(n_1674),
.Y(n_2404)
);

NAND3xp33_ASAP7_75t_SL g2405 ( 
.A(n_2086),
.B(n_1403),
.C(n_1401),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_2233),
.B(n_1843),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2167),
.Y(n_2407)
);

NOR2xp33_ASAP7_75t_L g2408 ( 
.A(n_2318),
.B(n_1759),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2174),
.Y(n_2409)
);

BUFx5_ASAP7_75t_L g2410 ( 
.A(n_2196),
.Y(n_2410)
);

NOR2xp33_ASAP7_75t_L g2411 ( 
.A(n_2318),
.B(n_1761),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2096),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_2186),
.B(n_1929),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2069),
.Y(n_2414)
);

NOR2xp33_ASAP7_75t_L g2415 ( 
.A(n_2142),
.B(n_1401),
.Y(n_2415)
);

NOR3xp33_ASAP7_75t_L g2416 ( 
.A(n_2322),
.B(n_1740),
.C(n_1960),
.Y(n_2416)
);

NOR3xp33_ASAP7_75t_L g2417 ( 
.A(n_2255),
.B(n_1740),
.C(n_1960),
.Y(n_2417)
);

NOR2xp33_ASAP7_75t_L g2418 ( 
.A(n_2142),
.B(n_1403),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2078),
.Y(n_2419)
);

AND2x6_ASAP7_75t_L g2420 ( 
.A(n_2329),
.B(n_1814),
.Y(n_2420)
);

BUFx6f_ASAP7_75t_L g2421 ( 
.A(n_2072),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2203),
.B(n_1929),
.Y(n_2422)
);

NOR2xp33_ASAP7_75t_L g2423 ( 
.A(n_2140),
.B(n_1404),
.Y(n_2423)
);

NOR2xp33_ASAP7_75t_L g2424 ( 
.A(n_2127),
.B(n_1404),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_SL g2425 ( 
.A(n_2102),
.B(n_1577),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2132),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2083),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2084),
.Y(n_2428)
);

BUFx6f_ASAP7_75t_L g2429 ( 
.A(n_2072),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2094),
.Y(n_2430)
);

OR2x6_ASAP7_75t_L g2431 ( 
.A(n_2176),
.B(n_1601),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2097),
.Y(n_2432)
);

BUFx6f_ASAP7_75t_L g2433 ( 
.A(n_2072),
.Y(n_2433)
);

NOR2xp33_ASAP7_75t_L g2434 ( 
.A(n_2115),
.B(n_1411),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2306),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2132),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2209),
.B(n_1929),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_SL g2438 ( 
.A(n_2076),
.B(n_1577),
.Y(n_2438)
);

AO221x1_ASAP7_75t_L g2439 ( 
.A1(n_2296),
.A2(n_1709),
.B1(n_1707),
.B2(n_1969),
.C(n_1936),
.Y(n_2439)
);

INVx2_ASAP7_75t_SL g2440 ( 
.A(n_2122),
.Y(n_2440)
);

NOR2xp33_ASAP7_75t_L g2441 ( 
.A(n_2123),
.B(n_1411),
.Y(n_2441)
);

NAND2xp33_ASAP7_75t_L g2442 ( 
.A(n_2134),
.B(n_1825),
.Y(n_2442)
);

NOR2xp33_ASAP7_75t_L g2443 ( 
.A(n_2123),
.B(n_1423),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_2138),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2138),
.Y(n_2445)
);

NOR2xp33_ASAP7_75t_L g2446 ( 
.A(n_2288),
.B(n_1423),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2215),
.B(n_1981),
.Y(n_2447)
);

INVxp67_ASAP7_75t_L g2448 ( 
.A(n_2291),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2225),
.B(n_1981),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2310),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2088),
.B(n_1981),
.Y(n_2451)
);

NAND3xp33_ASAP7_75t_L g2452 ( 
.A(n_2238),
.B(n_1977),
.C(n_1975),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_SL g2453 ( 
.A(n_2076),
.B(n_1973),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2126),
.B(n_2012),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2238),
.B(n_2012),
.Y(n_2455)
);

INVx2_ASAP7_75t_SL g2456 ( 
.A(n_2101),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2187),
.B(n_2012),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_SL g2458 ( 
.A(n_2264),
.B(n_1703),
.Y(n_2458)
);

BUFx5_ASAP7_75t_L g2459 ( 
.A(n_2196),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2324),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_2202),
.B(n_1857),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_2353),
.B(n_1978),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_SL g2463 ( 
.A(n_2294),
.B(n_1703),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2341),
.Y(n_2464)
);

AND2x2_ASAP7_75t_L g2465 ( 
.A(n_2248),
.B(n_1551),
.Y(n_2465)
);

NOR2xp67_ASAP7_75t_L g2466 ( 
.A(n_2173),
.B(n_1703),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_SL g2467 ( 
.A(n_2294),
.B(n_1703),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_2139),
.Y(n_2468)
);

BUFx8_ASAP7_75t_L g2469 ( 
.A(n_2305),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_SL g2470 ( 
.A(n_2353),
.B(n_2047),
.Y(n_2470)
);

HB1xp67_ASAP7_75t_L g2471 ( 
.A(n_2172),
.Y(n_2471)
);

BUFx3_ASAP7_75t_L g2472 ( 
.A(n_2162),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2348),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_L g2474 ( 
.A(n_2329),
.B(n_1983),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2139),
.Y(n_2475)
);

NOR3xp33_ASAP7_75t_L g2476 ( 
.A(n_2333),
.B(n_2047),
.C(n_2060),
.Y(n_2476)
);

NOR3xp33_ASAP7_75t_L g2477 ( 
.A(n_2333),
.B(n_2042),
.C(n_1579),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2304),
.B(n_1857),
.Y(n_2478)
);

NAND2xp33_ASAP7_75t_L g2479 ( 
.A(n_2356),
.B(n_1825),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_SL g2480 ( 
.A(n_2317),
.B(n_1840),
.Y(n_2480)
);

NOR2xp33_ASAP7_75t_L g2481 ( 
.A(n_2201),
.B(n_1430),
.Y(n_2481)
);

NOR2xp33_ASAP7_75t_L g2482 ( 
.A(n_2201),
.B(n_1430),
.Y(n_2482)
);

INVxp67_ASAP7_75t_L g2483 ( 
.A(n_2284),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_SL g2484 ( 
.A(n_2171),
.B(n_1854),
.Y(n_2484)
);

XOR2xp5_ASAP7_75t_L g2485 ( 
.A(n_2200),
.B(n_1185),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_SL g2486 ( 
.A(n_2171),
.B(n_1882),
.Y(n_2486)
);

AND2x2_ASAP7_75t_L g2487 ( 
.A(n_2303),
.B(n_1893),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2145),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2145),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2304),
.B(n_1859),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_SL g2491 ( 
.A(n_2184),
.B(n_1897),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2164),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2144),
.B(n_1859),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2352),
.Y(n_2494)
);

INVxp67_ASAP7_75t_L g2495 ( 
.A(n_2105),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2164),
.Y(n_2496)
);

AND2x6_ASAP7_75t_SL g2497 ( 
.A(n_2282),
.B(n_1572),
.Y(n_2497)
);

BUFx8_ASAP7_75t_L g2498 ( 
.A(n_2336),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_SL g2499 ( 
.A(n_2184),
.B(n_1936),
.Y(n_2499)
);

INVx2_ASAP7_75t_L g2500 ( 
.A(n_2165),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2144),
.B(n_1859),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2357),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2165),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_SL g2504 ( 
.A(n_2301),
.B(n_1969),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2354),
.B(n_1984),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2364),
.Y(n_2506)
);

INVxp67_ASAP7_75t_SL g2507 ( 
.A(n_2354),
.Y(n_2507)
);

INVxp33_ASAP7_75t_L g2508 ( 
.A(n_2287),
.Y(n_2508)
);

INVx8_ASAP7_75t_L g2509 ( 
.A(n_2176),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2207),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2099),
.B(n_1814),
.Y(n_2511)
);

NOR2xp67_ASAP7_75t_L g2512 ( 
.A(n_2214),
.B(n_1718),
.Y(n_2512)
);

NOR2xp67_ASAP7_75t_L g2513 ( 
.A(n_2220),
.B(n_1718),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2107),
.B(n_1823),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_2113),
.B(n_1823),
.Y(n_2515)
);

AO221x1_ASAP7_75t_L g2516 ( 
.A1(n_2340),
.A2(n_2351),
.B1(n_2210),
.B2(n_2080),
.C(n_2087),
.Y(n_2516)
);

CKINVDCx20_ASAP7_75t_R g2517 ( 
.A(n_2093),
.Y(n_2517)
);

BUFx6f_ASAP7_75t_L g2518 ( 
.A(n_2259),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2207),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_SL g2520 ( 
.A(n_2309),
.B(n_1969),
.Y(n_2520)
);

BUFx6f_ASAP7_75t_L g2521 ( 
.A(n_2259),
.Y(n_2521)
);

NOR2xp33_ASAP7_75t_L g2522 ( 
.A(n_2212),
.B(n_1431),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_SL g2523 ( 
.A(n_2313),
.B(n_1969),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_SL g2524 ( 
.A(n_2286),
.B(n_1974),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_SL g2525 ( 
.A(n_2325),
.B(n_1974),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2151),
.B(n_1898),
.Y(n_2526)
);

NOR2xp33_ASAP7_75t_L g2527 ( 
.A(n_2212),
.B(n_1431),
.Y(n_2527)
);

NOR2xp33_ASAP7_75t_L g2528 ( 
.A(n_2314),
.B(n_1432),
.Y(n_2528)
);

NOR2xp33_ASAP7_75t_L g2529 ( 
.A(n_2151),
.B(n_1432),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_SL g2530 ( 
.A(n_2327),
.B(n_1974),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2211),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_SL g2532 ( 
.A(n_2359),
.B(n_1974),
.Y(n_2532)
);

NOR2xp33_ASAP7_75t_L g2533 ( 
.A(n_2297),
.B(n_1439),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2211),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_2161),
.B(n_1985),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2185),
.B(n_1988),
.Y(n_2536)
);

BUFx5_ASAP7_75t_L g2537 ( 
.A(n_2196),
.Y(n_2537)
);

BUFx6f_ASAP7_75t_SL g2538 ( 
.A(n_2282),
.Y(n_2538)
);

NOR2xp33_ASAP7_75t_L g2539 ( 
.A(n_2297),
.B(n_1439),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2234),
.B(n_1989),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2196),
.B(n_1830),
.Y(n_2541)
);

NAND3xp33_ASAP7_75t_L g2542 ( 
.A(n_2077),
.B(n_2208),
.C(n_2361),
.Y(n_2542)
);

BUFx3_ASAP7_75t_L g2543 ( 
.A(n_2093),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2196),
.B(n_1830),
.Y(n_2544)
);

NOR2xp67_ASAP7_75t_L g2545 ( 
.A(n_2355),
.B(n_1990),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2216),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2216),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2236),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_SL g2549 ( 
.A(n_2366),
.B(n_1982),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2146),
.B(n_1839),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2236),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2237),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2243),
.B(n_1991),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2247),
.B(n_1992),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2237),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_SL g2556 ( 
.A(n_2066),
.B(n_1982),
.Y(n_2556)
);

BUFx6f_ASAP7_75t_L g2557 ( 
.A(n_2270),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2249),
.Y(n_2558)
);

NOR3xp33_ASAP7_75t_L g2559 ( 
.A(n_2330),
.B(n_1579),
.C(n_1877),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2249),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2254),
.Y(n_2561)
);

AND2x4_ASAP7_75t_L g2562 ( 
.A(n_2270),
.B(n_1899),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2254),
.Y(n_2563)
);

AOI21xp5_ASAP7_75t_L g2564 ( 
.A1(n_2121),
.A2(n_1817),
.B(n_2020),
.Y(n_2564)
);

AND2x2_ASAP7_75t_L g2565 ( 
.A(n_2339),
.B(n_1900),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_L g2566 ( 
.A(n_2328),
.B(n_1997),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2258),
.B(n_1998),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2272),
.B(n_1999),
.Y(n_2568)
);

NOR2xp33_ASAP7_75t_L g2569 ( 
.A(n_2326),
.B(n_1451),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2285),
.B(n_2004),
.Y(n_2570)
);

BUFx3_ASAP7_75t_L g2571 ( 
.A(n_2287),
.Y(n_2571)
);

INVx3_ASAP7_75t_L g2572 ( 
.A(n_2064),
.Y(n_2572)
);

NOR2xp67_ASAP7_75t_L g2573 ( 
.A(n_2278),
.B(n_2013),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2263),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2263),
.Y(n_2575)
);

NOR2xp33_ASAP7_75t_L g2576 ( 
.A(n_2326),
.B(n_1451),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_2316),
.B(n_2015),
.Y(n_2577)
);

INVxp67_ASAP7_75t_L g2578 ( 
.A(n_2179),
.Y(n_2578)
);

INVx1_ASAP7_75t_SL g2579 ( 
.A(n_2066),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_L g2580 ( 
.A(n_2321),
.B(n_2019),
.Y(n_2580)
);

NOR3xp33_ASAP7_75t_L g2581 ( 
.A(n_2340),
.B(n_1906),
.C(n_1904),
.Y(n_2581)
);

NOR3xp33_ASAP7_75t_L g2582 ( 
.A(n_2275),
.B(n_1911),
.C(n_1910),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_2121),
.B(n_1839),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2265),
.Y(n_2584)
);

NOR2xp33_ASAP7_75t_L g2585 ( 
.A(n_2323),
.B(n_1457),
.Y(n_2585)
);

AND2x2_ASAP7_75t_L g2586 ( 
.A(n_2350),
.B(n_1912),
.Y(n_2586)
);

NOR2xp67_ASAP7_75t_L g2587 ( 
.A(n_2335),
.B(n_2023),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2265),
.Y(n_2588)
);

INVx2_ASAP7_75t_L g2589 ( 
.A(n_2267),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2267),
.Y(n_2590)
);

AND2x2_ASAP7_75t_L g2591 ( 
.A(n_2350),
.B(n_1917),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_2121),
.B(n_1846),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2289),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_2289),
.Y(n_2594)
);

INVxp67_ASAP7_75t_SL g2595 ( 
.A(n_2128),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2299),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2121),
.B(n_1846),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_L g2598 ( 
.A(n_2169),
.B(n_1848),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2299),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_2302),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2169),
.B(n_1848),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_SL g2602 ( 
.A(n_2089),
.B(n_1982),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_2302),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2307),
.Y(n_2604)
);

NOR3xp33_ASAP7_75t_L g2605 ( 
.A(n_2100),
.B(n_1923),
.C(n_1918),
.Y(n_2605)
);

NOR2xp33_ASAP7_75t_L g2606 ( 
.A(n_2125),
.B(n_1457),
.Y(n_2606)
);

NOR2xp33_ASAP7_75t_SL g2607 ( 
.A(n_2125),
.B(n_2312),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2307),
.Y(n_2608)
);

NAND2xp33_ASAP7_75t_L g2609 ( 
.A(n_2356),
.B(n_2193),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2308),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_SL g2611 ( 
.A(n_2089),
.B(n_2090),
.Y(n_2611)
);

AND2x2_ASAP7_75t_L g2612 ( 
.A(n_2382),
.B(n_2090),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2395),
.B(n_2091),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2414),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2375),
.B(n_2091),
.Y(n_2615)
);

INVxp67_ASAP7_75t_L g2616 ( 
.A(n_2471),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2367),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2419),
.Y(n_2618)
);

NOR2xp33_ASAP7_75t_L g2619 ( 
.A(n_2385),
.B(n_2136),
.Y(n_2619)
);

INVx2_ASAP7_75t_L g2620 ( 
.A(n_2372),
.Y(n_2620)
);

A2O1A1Ixp33_ASAP7_75t_L g2621 ( 
.A1(n_2413),
.A2(n_2312),
.B(n_2222),
.C(n_2133),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2427),
.Y(n_2622)
);

NAND2x1_ASAP7_75t_L g2623 ( 
.A(n_2420),
.B(n_2064),
.Y(n_2623)
);

NOR2x2_ASAP7_75t_L g2624 ( 
.A(n_2431),
.B(n_2282),
.Y(n_2624)
);

OAI22xp5_ASAP7_75t_SL g2625 ( 
.A1(n_2533),
.A2(n_2131),
.B1(n_1471),
.B2(n_1469),
.Y(n_2625)
);

AOI21xp5_ASAP7_75t_L g2626 ( 
.A1(n_2422),
.A2(n_2261),
.B(n_2143),
.Y(n_2626)
);

BUFx3_ASAP7_75t_L g2627 ( 
.A(n_2472),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_L g2628 ( 
.A(n_2371),
.B(n_2104),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_L g2629 ( 
.A(n_2408),
.B(n_2104),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2428),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_SL g2631 ( 
.A(n_2404),
.B(n_2199),
.Y(n_2631)
);

BUFx6f_ASAP7_75t_L g2632 ( 
.A(n_2390),
.Y(n_2632)
);

OAI22xp5_ASAP7_75t_L g2633 ( 
.A1(n_2437),
.A2(n_2342),
.B1(n_2141),
.B2(n_2130),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2411),
.B(n_2342),
.Y(n_2634)
);

OAI22xp5_ASAP7_75t_L g2635 ( 
.A1(n_2447),
.A2(n_2071),
.B1(n_2114),
.B2(n_2100),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2577),
.B(n_2290),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2430),
.Y(n_2637)
);

BUFx3_ASAP7_75t_L g2638 ( 
.A(n_2509),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2432),
.Y(n_2639)
);

A2O1A1Ixp33_ASAP7_75t_L g2640 ( 
.A1(n_2380),
.A2(n_2416),
.B(n_2417),
.C(n_2455),
.Y(n_2640)
);

NOR2xp33_ASAP7_75t_L g2641 ( 
.A(n_2415),
.B(n_2136),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2373),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_2374),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2368),
.Y(n_2644)
);

AOI22xp5_ASAP7_75t_L g2645 ( 
.A1(n_2418),
.A2(n_1471),
.B1(n_1469),
.B2(n_2241),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2369),
.Y(n_2646)
);

INVx4_ASAP7_75t_L g2647 ( 
.A(n_2509),
.Y(n_2647)
);

AOI22xp5_ASAP7_75t_L g2648 ( 
.A1(n_2528),
.A2(n_2539),
.B1(n_2585),
.B2(n_2482),
.Y(n_2648)
);

INVx2_ASAP7_75t_L g2649 ( 
.A(n_2391),
.Y(n_2649)
);

AOI22xp5_ASAP7_75t_L g2650 ( 
.A1(n_2481),
.A2(n_2251),
.B1(n_1185),
.B2(n_1211),
.Y(n_2650)
);

AND2x2_ASAP7_75t_L g2651 ( 
.A(n_2465),
.B(n_2483),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2376),
.Y(n_2652)
);

HB1xp67_ASAP7_75t_L g2653 ( 
.A(n_2487),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2566),
.B(n_2290),
.Y(n_2654)
);

OR2x2_ASAP7_75t_L g2655 ( 
.A(n_2396),
.B(n_2179),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2412),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_L g2657 ( 
.A(n_2370),
.B(n_2120),
.Y(n_2657)
);

INVx2_ASAP7_75t_L g2658 ( 
.A(n_2426),
.Y(n_2658)
);

NOR2xp33_ASAP7_75t_L g2659 ( 
.A(n_2522),
.B(n_1191),
.Y(n_2659)
);

AND2x2_ASAP7_75t_L g2660 ( 
.A(n_2565),
.B(n_2120),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_L g2661 ( 
.A(n_2449),
.B(n_2217),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2462),
.B(n_2217),
.Y(n_2662)
);

OR2x2_ASAP7_75t_L g2663 ( 
.A(n_2446),
.B(n_2448),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2378),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2436),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_2540),
.B(n_2553),
.Y(n_2666)
);

HB1xp67_ASAP7_75t_L g2667 ( 
.A(n_2451),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_2554),
.B(n_2346),
.Y(n_2668)
);

AND2x6_ASAP7_75t_SL g2669 ( 
.A(n_2606),
.B(n_2226),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2568),
.B(n_2346),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2379),
.Y(n_2671)
);

AND2x2_ASAP7_75t_L g2672 ( 
.A(n_2527),
.B(n_2181),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2384),
.Y(n_2673)
);

OR2x2_ASAP7_75t_L g2674 ( 
.A(n_2405),
.B(n_2181),
.Y(n_2674)
);

HB1xp67_ASAP7_75t_L g2675 ( 
.A(n_2377),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2393),
.Y(n_2676)
);

INVx2_ASAP7_75t_L g2677 ( 
.A(n_2444),
.Y(n_2677)
);

BUFx6f_ASAP7_75t_L g2678 ( 
.A(n_2390),
.Y(n_2678)
);

AND2x4_ASAP7_75t_L g2679 ( 
.A(n_2518),
.B(n_1924),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2394),
.Y(n_2680)
);

NAND3xp33_ASAP7_75t_L g2681 ( 
.A(n_2476),
.B(n_845),
.C(n_1752),
.Y(n_2681)
);

AOI22xp33_ASAP7_75t_L g2682 ( 
.A1(n_2400),
.A2(n_2351),
.B1(n_2071),
.B2(n_2180),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2401),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2570),
.B(n_2029),
.Y(n_2684)
);

AOI21xp5_ASAP7_75t_L g2685 ( 
.A1(n_2609),
.A2(n_2261),
.B(n_2108),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2402),
.Y(n_2686)
);

BUFx3_ASAP7_75t_L g2687 ( 
.A(n_2509),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2567),
.B(n_2031),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_SL g2689 ( 
.A(n_2545),
.B(n_2199),
.Y(n_2689)
);

OR2x2_ASAP7_75t_L g2690 ( 
.A(n_2423),
.B(n_2033),
.Y(n_2690)
);

NAND3xp33_ASAP7_75t_L g2691 ( 
.A(n_2470),
.B(n_845),
.C(n_1752),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2580),
.B(n_2035),
.Y(n_2692)
);

OAI221xp5_ASAP7_75t_L g2693 ( 
.A1(n_2403),
.A2(n_2046),
.B1(n_2055),
.B2(n_2054),
.C(n_2052),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2407),
.Y(n_2694)
);

INVx3_ASAP7_75t_L g2695 ( 
.A(n_2420),
.Y(n_2695)
);

BUFx3_ASAP7_75t_L g2696 ( 
.A(n_2440),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2409),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_SL g2698 ( 
.A(n_2406),
.B(n_2169),
.Y(n_2698)
);

XOR2xp5_ASAP7_75t_L g2699 ( 
.A(n_2485),
.B(n_1212),
.Y(n_2699)
);

INVx2_ASAP7_75t_L g2700 ( 
.A(n_2445),
.Y(n_2700)
);

AND2x2_ASAP7_75t_L g2701 ( 
.A(n_2569),
.B(n_2576),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_2535),
.B(n_2536),
.Y(n_2702)
);

AOI21xp5_ASAP7_75t_L g2703 ( 
.A1(n_2454),
.A2(n_2194),
.B(n_2169),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_SL g2704 ( 
.A(n_2542),
.B(n_2194),
.Y(n_2704)
);

INVx2_ASAP7_75t_SL g2705 ( 
.A(n_2456),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2586),
.B(n_2059),
.Y(n_2706)
);

NOR2xp33_ASAP7_75t_L g2707 ( 
.A(n_2424),
.B(n_1212),
.Y(n_2707)
);

BUFx8_ASAP7_75t_L g2708 ( 
.A(n_2399),
.Y(n_2708)
);

BUFx12f_ASAP7_75t_L g2709 ( 
.A(n_2469),
.Y(n_2709)
);

OAI22xp5_ASAP7_75t_L g2710 ( 
.A1(n_2457),
.A2(n_2114),
.B1(n_2116),
.B2(n_2274),
.Y(n_2710)
);

OR2x6_ASAP7_75t_L g2711 ( 
.A(n_2431),
.B(n_2274),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2468),
.Y(n_2712)
);

BUFx3_ASAP7_75t_L g2713 ( 
.A(n_2469),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2591),
.B(n_2062),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2526),
.B(n_2177),
.Y(n_2715)
);

INVx3_ASAP7_75t_L g2716 ( 
.A(n_2420),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2475),
.Y(n_2717)
);

OAI22xp33_ASAP7_75t_L g2718 ( 
.A1(n_2607),
.A2(n_2182),
.B1(n_2188),
.B2(n_2183),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2579),
.B(n_2190),
.Y(n_2719)
);

NOR2xp33_ASAP7_75t_L g2720 ( 
.A(n_2434),
.B(n_1215),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2435),
.Y(n_2721)
);

AOI21xp5_ASAP7_75t_L g2722 ( 
.A1(n_2479),
.A2(n_2229),
.B(n_2194),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_L g2723 ( 
.A(n_2579),
.B(n_2191),
.Y(n_2723)
);

NOR2xp67_ASAP7_75t_L g2724 ( 
.A(n_2495),
.B(n_2253),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2488),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_SL g2726 ( 
.A(n_2441),
.B(n_2338),
.Y(n_2726)
);

CKINVDCx20_ASAP7_75t_R g2727 ( 
.A(n_2517),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2595),
.B(n_2195),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_L g2729 ( 
.A(n_2383),
.B(n_2197),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_SL g2730 ( 
.A(n_2542),
.B(n_2194),
.Y(n_2730)
);

AND2x2_ASAP7_75t_L g2731 ( 
.A(n_2443),
.B(n_2338),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_SL g2732 ( 
.A(n_2453),
.B(n_2229),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2383),
.B(n_2219),
.Y(n_2733)
);

NOR2xp33_ASAP7_75t_L g2734 ( 
.A(n_2438),
.B(n_2607),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_2392),
.B(n_2223),
.Y(n_2735)
);

INVx3_ASAP7_75t_L g2736 ( 
.A(n_2420),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2392),
.B(n_2224),
.Y(n_2737)
);

AND2x2_ASAP7_75t_L g2738 ( 
.A(n_2477),
.B(n_2227),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2474),
.B(n_2230),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2505),
.B(n_2235),
.Y(n_2740)
);

INVx8_ASAP7_75t_L g2741 ( 
.A(n_2431),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2450),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2489),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2562),
.B(n_2240),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2562),
.B(n_2250),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_SL g2746 ( 
.A(n_2512),
.B(n_2148),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_SL g2747 ( 
.A(n_2452),
.B(n_2229),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2398),
.B(n_2266),
.Y(n_2748)
);

OAI22xp5_ASAP7_75t_SL g2749 ( 
.A1(n_2529),
.A2(n_2131),
.B1(n_1229),
.B2(n_1232),
.Y(n_2749)
);

INVx3_ASAP7_75t_L g2750 ( 
.A(n_2572),
.Y(n_2750)
);

NOR3xp33_ASAP7_75t_L g2751 ( 
.A(n_2425),
.B(n_2116),
.C(n_2053),
.Y(n_2751)
);

INVx2_ASAP7_75t_L g2752 ( 
.A(n_2492),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2460),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_2496),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_SL g2755 ( 
.A(n_2513),
.B(n_2148),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2464),
.Y(n_2756)
);

NOR2xp33_ASAP7_75t_L g2757 ( 
.A(n_2452),
.B(n_1215),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_SL g2758 ( 
.A(n_2573),
.B(n_2229),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_SL g2759 ( 
.A(n_2587),
.B(n_2232),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_SL g2760 ( 
.A(n_2381),
.B(n_2232),
.Y(n_2760)
);

NOR2xp33_ASAP7_75t_SL g2761 ( 
.A(n_2387),
.B(n_2149),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2484),
.B(n_2276),
.Y(n_2762)
);

OR2x2_ASAP7_75t_L g2763 ( 
.A(n_2543),
.B(n_2280),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2486),
.B(n_2281),
.Y(n_2764)
);

INVx2_ASAP7_75t_SL g2765 ( 
.A(n_2498),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_2491),
.B(n_2283),
.Y(n_2766)
);

CKINVDCx5p33_ASAP7_75t_R g2767 ( 
.A(n_2399),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_2581),
.B(n_2262),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_SL g2769 ( 
.A(n_2518),
.B(n_2232),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_SL g2770 ( 
.A(n_2518),
.B(n_2232),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2500),
.Y(n_2771)
);

INVx3_ASAP7_75t_L g2772 ( 
.A(n_2572),
.Y(n_2772)
);

AND2x6_ASAP7_75t_SL g2773 ( 
.A(n_2508),
.B(n_1229),
.Y(n_2773)
);

NAND2xp5_ASAP7_75t_L g2774 ( 
.A(n_2507),
.B(n_2262),
.Y(n_2774)
);

AOI22xp33_ASAP7_75t_L g2775 ( 
.A1(n_2516),
.A2(n_2351),
.B1(n_2260),
.B2(n_1902),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_L g2776 ( 
.A(n_2611),
.B(n_2245),
.Y(n_2776)
);

NOR2xp33_ASAP7_75t_L g2777 ( 
.A(n_2578),
.B(n_1232),
.Y(n_2777)
);

NAND2xp33_ASAP7_75t_L g2778 ( 
.A(n_2410),
.B(n_2193),
.Y(n_2778)
);

NAND2xp5_ASAP7_75t_L g2779 ( 
.A(n_2521),
.B(n_2245),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_L g2780 ( 
.A(n_2521),
.B(n_2271),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_L g2781 ( 
.A(n_2521),
.B(n_2271),
.Y(n_2781)
);

INVxp67_ASAP7_75t_SL g2782 ( 
.A(n_2389),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_SL g2783 ( 
.A(n_2410),
.B(n_2242),
.Y(n_2783)
);

AOI22xp33_ASAP7_75t_L g2784 ( 
.A1(n_2439),
.A2(n_2337),
.B1(n_2053),
.B2(n_1888),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_L g2785 ( 
.A(n_2557),
.B(n_2273),
.Y(n_2785)
);

O2A1O1Ixp5_ASAP7_75t_L g2786 ( 
.A1(n_2480),
.A2(n_2020),
.B(n_2337),
.C(n_2175),
.Y(n_2786)
);

CKINVDCx11_ASAP7_75t_R g2787 ( 
.A(n_2571),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2557),
.B(n_2514),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_SL g2789 ( 
.A(n_2557),
.B(n_2242),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2514),
.B(n_2273),
.Y(n_2790)
);

AOI22xp33_ASAP7_75t_L g2791 ( 
.A1(n_2605),
.A2(n_1888),
.B1(n_2175),
.B2(n_2170),
.Y(n_2791)
);

AND2x2_ASAP7_75t_L g2792 ( 
.A(n_2559),
.B(n_1888),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2473),
.Y(n_2793)
);

NOR2xp33_ASAP7_75t_L g2794 ( 
.A(n_2494),
.B(n_1237),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2502),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2506),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_2515),
.B(n_2293),
.Y(n_2797)
);

INVx2_ASAP7_75t_L g2798 ( 
.A(n_2503),
.Y(n_2798)
);

NAND2xp33_ASAP7_75t_L g2799 ( 
.A(n_2410),
.B(n_2193),
.Y(n_2799)
);

CKINVDCx5p33_ASAP7_75t_R g2800 ( 
.A(n_2498),
.Y(n_2800)
);

AOI21x1_ASAP7_75t_L g2801 ( 
.A1(n_2463),
.A2(n_2155),
.B(n_2170),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_SL g2802 ( 
.A(n_2582),
.B(n_2242),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2510),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2548),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_SL g2805 ( 
.A(n_2466),
.B(n_2242),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2551),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_SL g2807 ( 
.A(n_2410),
.B(n_2279),
.Y(n_2807)
);

AOI21xp33_ASAP7_75t_L g2808 ( 
.A1(n_2634),
.A2(n_2458),
.B(n_2467),
.Y(n_2808)
);

AND2x2_ASAP7_75t_L g2809 ( 
.A(n_2651),
.B(n_2555),
.Y(n_2809)
);

NOR2xp33_ASAP7_75t_L g2810 ( 
.A(n_2648),
.B(n_1237),
.Y(n_2810)
);

AOI21xp5_ASAP7_75t_L g2811 ( 
.A1(n_2685),
.A2(n_2268),
.B(n_2397),
.Y(n_2811)
);

AOI21xp5_ASAP7_75t_L g2812 ( 
.A1(n_2685),
.A2(n_2442),
.B(n_2311),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_2702),
.B(n_2560),
.Y(n_2813)
);

AOI21xp5_ASAP7_75t_L g2814 ( 
.A1(n_2778),
.A2(n_2311),
.B(n_2279),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2614),
.Y(n_2815)
);

A2O1A1Ixp33_ASAP7_75t_L g2816 ( 
.A1(n_2619),
.A2(n_2228),
.B(n_2239),
.C(n_2192),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_L g2817 ( 
.A(n_2666),
.B(n_2589),
.Y(n_2817)
);

AOI21xp5_ASAP7_75t_L g2818 ( 
.A1(n_2799),
.A2(n_2311),
.B(n_2279),
.Y(n_2818)
);

A2O1A1Ixp33_ASAP7_75t_L g2819 ( 
.A1(n_2619),
.A2(n_2228),
.B(n_2239),
.C(n_2192),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2613),
.B(n_2590),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_L g2821 ( 
.A(n_2629),
.B(n_2594),
.Y(n_2821)
);

AND2x2_ASAP7_75t_L g2822 ( 
.A(n_2701),
.B(n_2600),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_L g2823 ( 
.A(n_2692),
.B(n_2603),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2684),
.B(n_2604),
.Y(n_2824)
);

CKINVDCx5p33_ASAP7_75t_R g2825 ( 
.A(n_2727),
.Y(n_2825)
);

BUFx6f_ASAP7_75t_L g2826 ( 
.A(n_2632),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_L g2827 ( 
.A(n_2688),
.B(n_2519),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2615),
.B(n_2531),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_2653),
.B(n_2534),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2653),
.B(n_2546),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2612),
.B(n_2547),
.Y(n_2831)
);

HB1xp67_ASAP7_75t_L g2832 ( 
.A(n_2675),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_2660),
.B(n_2552),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_SL g2834 ( 
.A(n_2690),
.B(n_1254),
.Y(n_2834)
);

AOI21xp33_ASAP7_75t_L g2835 ( 
.A1(n_2757),
.A2(n_2520),
.B(n_2504),
.Y(n_2835)
);

O2A1O1Ixp33_ASAP7_75t_L g2836 ( 
.A1(n_2640),
.A2(n_2277),
.B(n_2298),
.C(n_2244),
.Y(n_2836)
);

NOR2xp33_ASAP7_75t_L g2837 ( 
.A(n_2659),
.B(n_1254),
.Y(n_2837)
);

NOR2xp33_ASAP7_75t_L g2838 ( 
.A(n_2659),
.B(n_1260),
.Y(n_2838)
);

AOI21xp5_ASAP7_75t_L g2839 ( 
.A1(n_2626),
.A2(n_2124),
.B(n_2068),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_SL g2840 ( 
.A(n_2670),
.B(n_2641),
.Y(n_2840)
);

BUFx2_ASAP7_75t_L g2841 ( 
.A(n_2627),
.Y(n_2841)
);

BUFx3_ASAP7_75t_L g2842 ( 
.A(n_2696),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2617),
.Y(n_2843)
);

BUFx4f_ASAP7_75t_L g2844 ( 
.A(n_2709),
.Y(n_2844)
);

OAI22xp5_ASAP7_75t_L g2845 ( 
.A1(n_2734),
.A2(n_2650),
.B1(n_2645),
.B2(n_2757),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2667),
.B(n_2558),
.Y(n_2846)
);

AOI22xp5_ASAP7_75t_L g2847 ( 
.A1(n_2641),
.A2(n_1262),
.B1(n_1271),
.B2(n_1260),
.Y(n_2847)
);

AOI22xp5_ASAP7_75t_L g2848 ( 
.A1(n_2707),
.A2(n_1271),
.B1(n_1272),
.B2(n_1262),
.Y(n_2848)
);

NAND2xp33_ASAP7_75t_L g2849 ( 
.A(n_2751),
.B(n_2410),
.Y(n_2849)
);

O2A1O1Ixp33_ASAP7_75t_L g2850 ( 
.A1(n_2768),
.A2(n_2277),
.B(n_2298),
.C(n_2244),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_SL g2851 ( 
.A(n_2668),
.B(n_1272),
.Y(n_2851)
);

AOI21xp5_ASAP7_75t_L g2852 ( 
.A1(n_2722),
.A2(n_1817),
.B(n_2389),
.Y(n_2852)
);

AOI21xp5_ASAP7_75t_L g2853 ( 
.A1(n_2782),
.A2(n_2478),
.B(n_2461),
.Y(n_2853)
);

OAI22xp5_ASAP7_75t_L g2854 ( 
.A1(n_2734),
.A2(n_2538),
.B1(n_1276),
.B2(n_1301),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_2667),
.B(n_2561),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2672),
.B(n_2563),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_2663),
.B(n_2574),
.Y(n_2857)
);

AOI21xp5_ASAP7_75t_L g2858 ( 
.A1(n_2782),
.A2(n_2478),
.B(n_2461),
.Y(n_2858)
);

AOI21xp5_ASAP7_75t_L g2859 ( 
.A1(n_2704),
.A2(n_2490),
.B(n_2388),
.Y(n_2859)
);

A2O1A1Ixp33_ASAP7_75t_L g2860 ( 
.A1(n_2751),
.A2(n_2530),
.B(n_2532),
.C(n_2525),
.Y(n_2860)
);

O2A1O1Ixp33_ASAP7_75t_L g2861 ( 
.A1(n_2718),
.A2(n_2549),
.B(n_2499),
.C(n_2523),
.Y(n_2861)
);

BUFx4f_ASAP7_75t_L g2862 ( 
.A(n_2741),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_2628),
.B(n_2575),
.Y(n_2863)
);

INVx3_ASAP7_75t_L g2864 ( 
.A(n_2695),
.Y(n_2864)
);

NOR2xp33_ASAP7_75t_L g2865 ( 
.A(n_2707),
.B(n_1273),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2739),
.B(n_2584),
.Y(n_2866)
);

AND2x2_ASAP7_75t_L g2867 ( 
.A(n_2794),
.B(n_2731),
.Y(n_2867)
);

AOI21xp5_ASAP7_75t_L g2868 ( 
.A1(n_2704),
.A2(n_2490),
.B(n_2388),
.Y(n_2868)
);

NAND2x1_ASAP7_75t_L g2869 ( 
.A(n_2695),
.B(n_2085),
.Y(n_2869)
);

HB1xp67_ASAP7_75t_L g2870 ( 
.A(n_2675),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2618),
.Y(n_2871)
);

AOI21xp5_ASAP7_75t_L g2872 ( 
.A1(n_2730),
.A2(n_2386),
.B(n_2564),
.Y(n_2872)
);

AOI22xp33_ASAP7_75t_L g2873 ( 
.A1(n_2720),
.A2(n_2538),
.B1(n_1276),
.B2(n_1301),
.Y(n_2873)
);

AOI21xp5_ASAP7_75t_L g2874 ( 
.A1(n_2730),
.A2(n_2386),
.B(n_2221),
.Y(n_2874)
);

AOI21xp5_ASAP7_75t_L g2875 ( 
.A1(n_2635),
.A2(n_2221),
.B(n_2218),
.Y(n_2875)
);

OAI21xp33_ASAP7_75t_L g2876 ( 
.A1(n_2794),
.A2(n_1312),
.B(n_1273),
.Y(n_2876)
);

NAND2xp33_ASAP7_75t_L g2877 ( 
.A(n_2741),
.B(n_2774),
.Y(n_2877)
);

AOI21xp5_ASAP7_75t_L g2878 ( 
.A1(n_2703),
.A2(n_2218),
.B(n_2583),
.Y(n_2878)
);

OAI21xp5_ASAP7_75t_L g2879 ( 
.A1(n_2786),
.A2(n_1986),
.B(n_2493),
.Y(n_2879)
);

OAI21xp5_ASAP7_75t_L g2880 ( 
.A1(n_2786),
.A2(n_1986),
.B(n_2493),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2620),
.Y(n_2881)
);

AOI21xp5_ASAP7_75t_L g2882 ( 
.A1(n_2703),
.A2(n_2592),
.B(n_2583),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_SL g2883 ( 
.A(n_2738),
.B(n_2636),
.Y(n_2883)
);

AOI21xp5_ASAP7_75t_L g2884 ( 
.A1(n_2621),
.A2(n_2597),
.B(n_2592),
.Y(n_2884)
);

AO21x1_ASAP7_75t_L g2885 ( 
.A1(n_2718),
.A2(n_2524),
.B(n_2155),
.Y(n_2885)
);

AOI21x1_ASAP7_75t_L g2886 ( 
.A1(n_2747),
.A2(n_2550),
.B(n_1803),
.Y(n_2886)
);

CKINVDCx5p33_ASAP7_75t_R g2887 ( 
.A(n_2787),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2622),
.Y(n_2888)
);

AOI21xp5_ASAP7_75t_L g2889 ( 
.A1(n_2729),
.A2(n_2598),
.B(n_2597),
.Y(n_2889)
);

O2A1O1Ixp33_ASAP7_75t_L g2890 ( 
.A1(n_2631),
.A2(n_1766),
.B(n_1816),
.C(n_1852),
.Y(n_2890)
);

BUFx6f_ASAP7_75t_L g2891 ( 
.A(n_2632),
.Y(n_2891)
);

OAI22xp5_ASAP7_75t_L g2892 ( 
.A1(n_2720),
.A2(n_1312),
.B1(n_1616),
.B2(n_2295),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_2740),
.B(n_2588),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2630),
.Y(n_2894)
);

HB1xp67_ASAP7_75t_L g2895 ( 
.A(n_2616),
.Y(n_2895)
);

OAI21xp5_ASAP7_75t_L g2896 ( 
.A1(n_2633),
.A2(n_2775),
.B(n_2790),
.Y(n_2896)
);

AOI21xp5_ASAP7_75t_L g2897 ( 
.A1(n_2733),
.A2(n_2747),
.B(n_2797),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2654),
.B(n_2593),
.Y(n_2898)
);

OAI21xp5_ASAP7_75t_L g2899 ( 
.A1(n_2775),
.A2(n_2501),
.B(n_1927),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_SL g2900 ( 
.A(n_2715),
.B(n_1752),
.Y(n_2900)
);

OR2x2_ASAP7_75t_L g2901 ( 
.A(n_2763),
.B(n_2596),
.Y(n_2901)
);

OAI21xp5_ASAP7_75t_L g2902 ( 
.A1(n_2776),
.A2(n_2501),
.B(n_1927),
.Y(n_2902)
);

NOR2xp33_ASAP7_75t_SL g2903 ( 
.A(n_2647),
.B(n_2295),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2706),
.B(n_2599),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2637),
.Y(n_2905)
);

NOR2xp33_ASAP7_75t_L g2906 ( 
.A(n_2699),
.B(n_1616),
.Y(n_2906)
);

INVx2_ASAP7_75t_L g2907 ( 
.A(n_2642),
.Y(n_2907)
);

INVx2_ASAP7_75t_L g2908 ( 
.A(n_2643),
.Y(n_2908)
);

OAI21xp5_ASAP7_75t_L g2909 ( 
.A1(n_2784),
.A2(n_2550),
.B(n_2515),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_L g2910 ( 
.A(n_2714),
.B(n_2608),
.Y(n_2910)
);

INVxp67_ASAP7_75t_L g2911 ( 
.A(n_2777),
.Y(n_2911)
);

AND2x2_ASAP7_75t_L g2912 ( 
.A(n_2777),
.B(n_2610),
.Y(n_2912)
);

O2A1O1Ixp33_ASAP7_75t_L g2913 ( 
.A1(n_2693),
.A2(n_1816),
.B(n_1766),
.C(n_1852),
.Y(n_2913)
);

AOI21xp5_ASAP7_75t_L g2914 ( 
.A1(n_2760),
.A2(n_2601),
.B(n_2598),
.Y(n_2914)
);

A2O1A1Ixp33_ASAP7_75t_L g2915 ( 
.A1(n_2691),
.A2(n_2025),
.B(n_2602),
.C(n_2556),
.Y(n_2915)
);

NOR2xp33_ASAP7_75t_L g2916 ( 
.A(n_2625),
.B(n_1616),
.Y(n_2916)
);

NOR2xp33_ASAP7_75t_L g2917 ( 
.A(n_2749),
.B(n_1626),
.Y(n_2917)
);

OAI22xp5_ASAP7_75t_L g2918 ( 
.A1(n_2674),
.A2(n_2293),
.B1(n_2103),
.B2(n_2168),
.Y(n_2918)
);

AOI21xp5_ASAP7_75t_L g2919 ( 
.A1(n_2760),
.A2(n_2601),
.B(n_2511),
.Y(n_2919)
);

AOI21xp5_ASAP7_75t_L g2920 ( 
.A1(n_2698),
.A2(n_2511),
.B(n_2541),
.Y(n_2920)
);

NOR2x1p5_ASAP7_75t_SL g2921 ( 
.A(n_2801),
.B(n_2193),
.Y(n_2921)
);

AOI21x1_ASAP7_75t_L g2922 ( 
.A1(n_2792),
.A2(n_1803),
.B(n_2246),
.Y(n_2922)
);

AOI22xp5_ASAP7_75t_L g2923 ( 
.A1(n_2726),
.A2(n_1837),
.B1(n_1825),
.B2(n_1659),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2662),
.B(n_2497),
.Y(n_2924)
);

NAND2xp5_ASAP7_75t_SL g2925 ( 
.A(n_2728),
.B(n_1837),
.Y(n_2925)
);

CKINVDCx8_ASAP7_75t_R g2926 ( 
.A(n_2773),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_SL g2927 ( 
.A(n_2744),
.B(n_2745),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2657),
.B(n_2308),
.Y(n_2928)
);

AND2x2_ASAP7_75t_L g2929 ( 
.A(n_2655),
.B(n_523),
.Y(n_2929)
);

CKINVDCx8_ASAP7_75t_R g2930 ( 
.A(n_2669),
.Y(n_2930)
);

AOI21xp5_ASAP7_75t_L g2931 ( 
.A1(n_2698),
.A2(n_2544),
.B(n_2541),
.Y(n_2931)
);

NAND2xp5_ASAP7_75t_L g2932 ( 
.A(n_2719),
.B(n_2723),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2639),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_SL g2934 ( 
.A(n_2661),
.B(n_2459),
.Y(n_2934)
);

OAI21xp5_ASAP7_75t_L g2935 ( 
.A1(n_2784),
.A2(n_2544),
.B(n_1887),
.Y(n_2935)
);

AOI21xp5_ASAP7_75t_L g2936 ( 
.A1(n_2783),
.A2(n_2807),
.B(n_2737),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2644),
.Y(n_2937)
);

AND2x2_ASAP7_75t_L g2938 ( 
.A(n_2679),
.B(n_523),
.Y(n_2938)
);

AOI21xp5_ASAP7_75t_L g2939 ( 
.A1(n_2783),
.A2(n_2807),
.B(n_2735),
.Y(n_2939)
);

AOI21xp5_ASAP7_75t_L g2940 ( 
.A1(n_2710),
.A2(n_2001),
.B(n_1982),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2646),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_2788),
.B(n_2319),
.Y(n_2942)
);

INVx3_ASAP7_75t_L g2943 ( 
.A(n_2716),
.Y(n_2943)
);

AOI22xp5_ASAP7_75t_L g2944 ( 
.A1(n_2681),
.A2(n_1659),
.B1(n_1618),
.B2(n_2027),
.Y(n_2944)
);

NOR3xp33_ASAP7_75t_L g2945 ( 
.A(n_2746),
.B(n_768),
.C(n_767),
.Y(n_2945)
);

AOI21x1_ASAP7_75t_L g2946 ( 
.A1(n_2732),
.A2(n_1887),
.B(n_2014),
.Y(n_2946)
);

AOI22xp33_ASAP7_75t_L g2947 ( 
.A1(n_2682),
.A2(n_2027),
.B1(n_2160),
.B2(n_1659),
.Y(n_2947)
);

NOR2xp33_ASAP7_75t_L g2948 ( 
.A(n_2616),
.B(n_1618),
.Y(n_2948)
);

AOI21xp5_ASAP7_75t_L g2949 ( 
.A1(n_2623),
.A2(n_2038),
.B(n_2001),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_L g2950 ( 
.A(n_2762),
.B(n_2319),
.Y(n_2950)
);

NOR2xp33_ASAP7_75t_L g2951 ( 
.A(n_2705),
.B(n_524),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2652),
.Y(n_2952)
);

A2O1A1Ixp33_ASAP7_75t_L g2953 ( 
.A1(n_2682),
.A2(n_2079),
.B(n_2080),
.C(n_2075),
.Y(n_2953)
);

INVx3_ASAP7_75t_L g2954 ( 
.A(n_2736),
.Y(n_2954)
);

BUFx2_ASAP7_75t_L g2955 ( 
.A(n_2638),
.Y(n_2955)
);

OAI21xp5_ASAP7_75t_L g2956 ( 
.A1(n_2764),
.A2(n_2027),
.B(n_2160),
.Y(n_2956)
);

AOI21xp5_ASAP7_75t_L g2957 ( 
.A1(n_2766),
.A2(n_2038),
.B(n_2001),
.Y(n_2957)
);

OAI21xp5_ASAP7_75t_L g2958 ( 
.A1(n_2791),
.A2(n_2027),
.B(n_2160),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2664),
.Y(n_2959)
);

AOI21xp5_ASAP7_75t_L g2960 ( 
.A1(n_2779),
.A2(n_2048),
.B(n_2038),
.Y(n_2960)
);

AOI22xp5_ASAP7_75t_L g2961 ( 
.A1(n_2755),
.A2(n_2027),
.B1(n_2160),
.B2(n_755),
.Y(n_2961)
);

OAI21xp5_ASAP7_75t_L g2962 ( 
.A1(n_2791),
.A2(n_2343),
.B(n_2320),
.Y(n_2962)
);

AND2x4_ASAP7_75t_L g2963 ( 
.A(n_2647),
.B(n_2390),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2649),
.Y(n_2964)
);

BUFx6f_ASAP7_75t_L g2965 ( 
.A(n_2632),
.Y(n_2965)
);

AOI21xp5_ASAP7_75t_L g2966 ( 
.A1(n_2732),
.A2(n_2802),
.B(n_2781),
.Y(n_2966)
);

O2A1O1Ixp33_ASAP7_75t_L g2967 ( 
.A1(n_2689),
.A2(n_2343),
.B(n_2345),
.C(n_2320),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_L g2968 ( 
.A(n_2748),
.B(n_2345),
.Y(n_2968)
);

OAI321xp33_ASAP7_75t_L g2969 ( 
.A1(n_2785),
.A2(n_2362),
.A3(n_2358),
.B1(n_2365),
.B2(n_2360),
.C(n_2349),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2671),
.Y(n_2970)
);

AND2x2_ASAP7_75t_L g2971 ( 
.A(n_2679),
.B(n_524),
.Y(n_2971)
);

CKINVDCx5p33_ASAP7_75t_R g2972 ( 
.A(n_2800),
.Y(n_2972)
);

AOI21x1_ASAP7_75t_L g2973 ( 
.A1(n_2758),
.A2(n_2759),
.B(n_2769),
.Y(n_2973)
);

AOI21xp5_ASAP7_75t_L g2974 ( 
.A1(n_2780),
.A2(n_2048),
.B(n_2085),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2673),
.Y(n_2975)
);

INVx2_ASAP7_75t_SL g2976 ( 
.A(n_2708),
.Y(n_2976)
);

HB1xp67_ASAP7_75t_L g2977 ( 
.A(n_2676),
.Y(n_2977)
);

AND2x2_ASAP7_75t_L g2978 ( 
.A(n_2656),
.B(n_526),
.Y(n_2978)
);

AND2x4_ASAP7_75t_L g2979 ( 
.A(n_2687),
.B(n_2421),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_SL g2980 ( 
.A(n_2724),
.B(n_2459),
.Y(n_2980)
);

AOI21xp5_ASAP7_75t_L g2981 ( 
.A1(n_2805),
.A2(n_2048),
.B(n_2168),
.Y(n_2981)
);

AOI22xp33_ASAP7_75t_L g2982 ( 
.A1(n_2741),
.A2(n_2160),
.B1(n_1957),
.B2(n_2459),
.Y(n_2982)
);

NOR2xp33_ASAP7_75t_SL g2983 ( 
.A(n_2708),
.B(n_2459),
.Y(n_2983)
);

AND2x2_ASAP7_75t_L g2984 ( 
.A(n_2658),
.B(n_526),
.Y(n_2984)
);

AOI21xp5_ASAP7_75t_L g2985 ( 
.A1(n_2770),
.A2(n_2048),
.B(n_2178),
.Y(n_2985)
);

NOR2x1_ASAP7_75t_L g2986 ( 
.A(n_2711),
.B(n_2178),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2680),
.Y(n_2987)
);

A2O1A1Ixp33_ASAP7_75t_L g2988 ( 
.A1(n_2683),
.A2(n_2079),
.B(n_2087),
.C(n_2075),
.Y(n_2988)
);

AOI21xp5_ASAP7_75t_L g2989 ( 
.A1(n_2789),
.A2(n_2736),
.B(n_2711),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2686),
.B(n_2349),
.Y(n_2990)
);

AOI21xp5_ASAP7_75t_L g2991 ( 
.A1(n_2711),
.A2(n_2315),
.B(n_2292),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2694),
.B(n_2358),
.Y(n_2992)
);

OAI21xp33_ASAP7_75t_L g2993 ( 
.A1(n_2697),
.A2(n_2742),
.B(n_2721),
.Y(n_2993)
);

AOI21xp5_ASAP7_75t_L g2994 ( 
.A1(n_2750),
.A2(n_2315),
.B(n_2292),
.Y(n_2994)
);

INVx2_ASAP7_75t_L g2995 ( 
.A(n_2665),
.Y(n_2995)
);

NOR2xp33_ASAP7_75t_L g2996 ( 
.A(n_2767),
.B(n_765),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2977),
.Y(n_2997)
);

AOI22xp5_ASAP7_75t_L g2998 ( 
.A1(n_2810),
.A2(n_2765),
.B1(n_2756),
.B2(n_2753),
.Y(n_2998)
);

INVx4_ASAP7_75t_L g2999 ( 
.A(n_2862),
.Y(n_2999)
);

INVxp67_ASAP7_75t_SL g3000 ( 
.A(n_2832),
.Y(n_3000)
);

INVx3_ASAP7_75t_L g3001 ( 
.A(n_2862),
.Y(n_3001)
);

AOI22xp5_ASAP7_75t_L g3002 ( 
.A1(n_2845),
.A2(n_2795),
.B1(n_2796),
.B2(n_2793),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2815),
.Y(n_3003)
);

BUFx12f_ASAP7_75t_L g3004 ( 
.A(n_2887),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_2897),
.B(n_2932),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_2843),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2871),
.Y(n_3007)
);

INVx5_ASAP7_75t_L g3008 ( 
.A(n_2826),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2888),
.Y(n_3009)
);

INVx2_ASAP7_75t_L g3010 ( 
.A(n_2881),
.Y(n_3010)
);

BUFx3_ASAP7_75t_L g3011 ( 
.A(n_2841),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_L g3012 ( 
.A(n_2883),
.B(n_2803),
.Y(n_3012)
);

BUFx6f_ASAP7_75t_L g3013 ( 
.A(n_2842),
.Y(n_3013)
);

INVx2_ASAP7_75t_SL g3014 ( 
.A(n_2844),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_SL g3015 ( 
.A(n_2840),
.B(n_2750),
.Y(n_3015)
);

INVx4_ASAP7_75t_L g3016 ( 
.A(n_2826),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2904),
.B(n_2677),
.Y(n_3017)
);

BUFx3_ASAP7_75t_L g3018 ( 
.A(n_2955),
.Y(n_3018)
);

INVx2_ASAP7_75t_L g3019 ( 
.A(n_2907),
.Y(n_3019)
);

BUFx2_ASAP7_75t_L g3020 ( 
.A(n_2870),
.Y(n_3020)
);

NOR2xp33_ASAP7_75t_L g3021 ( 
.A(n_2837),
.B(n_2761),
.Y(n_3021)
);

NOR2xp33_ASAP7_75t_R g3022 ( 
.A(n_2825),
.B(n_2713),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_SL g3023 ( 
.A(n_2924),
.B(n_2772),
.Y(n_3023)
);

INVx3_ASAP7_75t_L g3024 ( 
.A(n_2826),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2894),
.Y(n_3025)
);

BUFx6f_ASAP7_75t_L g3026 ( 
.A(n_2891),
.Y(n_3026)
);

O2A1O1Ixp33_ASAP7_75t_L g3027 ( 
.A1(n_2925),
.A2(n_2712),
.B(n_2717),
.C(n_2700),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2905),
.Y(n_3028)
);

HB1xp67_ASAP7_75t_SL g3029 ( 
.A(n_2926),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2933),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_SL g3031 ( 
.A(n_2867),
.B(n_2772),
.Y(n_3031)
);

INVx2_ASAP7_75t_L g3032 ( 
.A(n_2908),
.Y(n_3032)
);

INVx2_ASAP7_75t_L g3033 ( 
.A(n_2964),
.Y(n_3033)
);

NOR2xp33_ASAP7_75t_L g3034 ( 
.A(n_2838),
.B(n_2725),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2927),
.B(n_2743),
.Y(n_3035)
);

BUFx6f_ASAP7_75t_L g3036 ( 
.A(n_2891),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_SL g3037 ( 
.A(n_2923),
.B(n_2900),
.Y(n_3037)
);

INVx2_ASAP7_75t_L g3038 ( 
.A(n_2995),
.Y(n_3038)
);

AND2x4_ASAP7_75t_L g3039 ( 
.A(n_2989),
.B(n_2632),
.Y(n_3039)
);

OAI22xp5_ASAP7_75t_L g3040 ( 
.A1(n_2911),
.A2(n_771),
.B1(n_772),
.B2(n_770),
.Y(n_3040)
);

CKINVDCx5p33_ASAP7_75t_R g3041 ( 
.A(n_2972),
.Y(n_3041)
);

BUFx4f_ASAP7_75t_SL g3042 ( 
.A(n_2976),
.Y(n_3042)
);

INVx3_ASAP7_75t_L g3043 ( 
.A(n_2891),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_L g3044 ( 
.A(n_2828),
.B(n_2806),
.Y(n_3044)
);

CKINVDCx5p33_ASAP7_75t_R g3045 ( 
.A(n_2844),
.Y(n_3045)
);

INVx2_ASAP7_75t_L g3046 ( 
.A(n_2937),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_SL g3047 ( 
.A(n_2944),
.B(n_2752),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_2822),
.B(n_2804),
.Y(n_3048)
);

INVx2_ASAP7_75t_L g3049 ( 
.A(n_2941),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_SL g3050 ( 
.A(n_2856),
.B(n_2754),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_2910),
.B(n_2771),
.Y(n_3051)
);

INVx2_ASAP7_75t_L g3052 ( 
.A(n_2952),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_2966),
.B(n_2798),
.Y(n_3053)
);

INVx2_ASAP7_75t_L g3054 ( 
.A(n_2959),
.Y(n_3054)
);

AND2x2_ASAP7_75t_L g3055 ( 
.A(n_2912),
.B(n_2678),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_2821),
.B(n_2678),
.Y(n_3056)
);

INVx2_ASAP7_75t_L g3057 ( 
.A(n_2970),
.Y(n_3057)
);

AO22x1_ASAP7_75t_L g3058 ( 
.A1(n_2916),
.A2(n_772),
.B1(n_775),
.B2(n_771),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2975),
.Y(n_3059)
);

INVxp67_ASAP7_75t_L g3060 ( 
.A(n_2895),
.Y(n_3060)
);

NOR2xp67_ASAP7_75t_L g3061 ( 
.A(n_2974),
.B(n_2678),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2987),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_SL g3063 ( 
.A(n_2890),
.B(n_2459),
.Y(n_3063)
);

INVx2_ASAP7_75t_L g3064 ( 
.A(n_2809),
.Y(n_3064)
);

BUFx6f_ASAP7_75t_L g3065 ( 
.A(n_2965),
.Y(n_3065)
);

AND2x6_ASAP7_75t_L g3066 ( 
.A(n_2986),
.B(n_2678),
.Y(n_3066)
);

A2O1A1Ixp33_ASAP7_75t_L g3067 ( 
.A1(n_2913),
.A2(n_766),
.B(n_778),
.C(n_765),
.Y(n_3067)
);

INVx1_ASAP7_75t_SL g3068 ( 
.A(n_2901),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2993),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2831),
.Y(n_3070)
);

AND2x4_ASAP7_75t_L g3071 ( 
.A(n_2963),
.B(n_2421),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_SL g3072 ( 
.A(n_2918),
.B(n_2537),
.Y(n_3072)
);

INVx3_ASAP7_75t_L g3073 ( 
.A(n_2965),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_L g3074 ( 
.A(n_2820),
.B(n_754),
.Y(n_3074)
);

AOI22xp5_ASAP7_75t_L g3075 ( 
.A1(n_2876),
.A2(n_776),
.B1(n_781),
.B2(n_775),
.Y(n_3075)
);

OAI221xp5_ASAP7_75t_L g3076 ( 
.A1(n_2873),
.A2(n_776),
.B1(n_787),
.B2(n_782),
.C(n_781),
.Y(n_3076)
);

INVx2_ASAP7_75t_L g3077 ( 
.A(n_2833),
.Y(n_3077)
);

NOR2xp67_ASAP7_75t_L g3078 ( 
.A(n_2936),
.B(n_2360),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_SL g3079 ( 
.A(n_2854),
.B(n_2537),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_SL g3080 ( 
.A(n_2903),
.B(n_2537),
.Y(n_3080)
);

INVx2_ASAP7_75t_L g3081 ( 
.A(n_2829),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2830),
.Y(n_3082)
);

INVx3_ASAP7_75t_L g3083 ( 
.A(n_2965),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_L g3084 ( 
.A(n_2857),
.B(n_756),
.Y(n_3084)
);

BUFx6f_ASAP7_75t_L g3085 ( 
.A(n_2979),
.Y(n_3085)
);

INVx2_ASAP7_75t_L g3086 ( 
.A(n_2990),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_L g3087 ( 
.A(n_2813),
.B(n_760),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2817),
.B(n_2362),
.Y(n_3088)
);

INVx2_ASAP7_75t_L g3089 ( 
.A(n_2992),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2846),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_L g3091 ( 
.A(n_2827),
.B(n_2863),
.Y(n_3091)
);

BUFx2_ASAP7_75t_R g3092 ( 
.A(n_2930),
.Y(n_3092)
);

AOI22xp33_ASAP7_75t_L g3093 ( 
.A1(n_2865),
.A2(n_787),
.B1(n_789),
.B2(n_782),
.Y(n_3093)
);

INVx3_ASAP7_75t_L g3094 ( 
.A(n_2963),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2823),
.B(n_2824),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_2866),
.B(n_2365),
.Y(n_3096)
);

BUFx6f_ASAP7_75t_L g3097 ( 
.A(n_2979),
.Y(n_3097)
);

OAI21xp5_ASAP7_75t_L g3098 ( 
.A1(n_2884),
.A2(n_2057),
.B(n_2056),
.Y(n_3098)
);

AND2x4_ASAP7_75t_L g3099 ( 
.A(n_2864),
.B(n_2421),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_2893),
.B(n_789),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2855),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_L g3102 ( 
.A(n_2898),
.B(n_790),
.Y(n_3102)
);

AND2x4_ASAP7_75t_L g3103 ( 
.A(n_2864),
.B(n_2429),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2942),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_2950),
.Y(n_3105)
);

OAI22xp33_ASAP7_75t_L g3106 ( 
.A1(n_2903),
.A2(n_791),
.B1(n_792),
.B2(n_790),
.Y(n_3106)
);

AOI21xp5_ASAP7_75t_L g3107 ( 
.A1(n_2853),
.A2(n_2344),
.B(n_2332),
.Y(n_3107)
);

HB1xp67_ASAP7_75t_L g3108 ( 
.A(n_2928),
.Y(n_3108)
);

NOR2xp33_ASAP7_75t_L g3109 ( 
.A(n_2848),
.B(n_766),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_2896),
.B(n_2537),
.Y(n_3110)
);

NOR2xp67_ASAP7_75t_L g3111 ( 
.A(n_2939),
.B(n_2095),
.Y(n_3111)
);

INVx2_ASAP7_75t_SL g3112 ( 
.A(n_2929),
.Y(n_3112)
);

INVx3_ASAP7_75t_L g3113 ( 
.A(n_2943),
.Y(n_3113)
);

AOI22xp33_ASAP7_75t_L g3114 ( 
.A1(n_2834),
.A2(n_792),
.B1(n_795),
.B2(n_791),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_L g3115 ( 
.A(n_2851),
.B(n_795),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2968),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_2943),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_2896),
.B(n_2537),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_L g3119 ( 
.A(n_2877),
.B(n_798),
.Y(n_3119)
);

NOR2xp33_ASAP7_75t_L g3120 ( 
.A(n_2892),
.B(n_778),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2885),
.Y(n_3121)
);

INVx2_ASAP7_75t_SL g3122 ( 
.A(n_2938),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_2849),
.Y(n_3123)
);

CKINVDCx8_ASAP7_75t_R g3124 ( 
.A(n_2906),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_2858),
.Y(n_3125)
);

INVxp67_ASAP7_75t_L g3126 ( 
.A(n_2951),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2978),
.B(n_798),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_2984),
.B(n_801),
.Y(n_3128)
);

AND2x2_ASAP7_75t_SL g3129 ( 
.A(n_2983),
.B(n_2624),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_2973),
.Y(n_3130)
);

INVx2_ASAP7_75t_L g3131 ( 
.A(n_2954),
.Y(n_3131)
);

CKINVDCx8_ASAP7_75t_R g3132 ( 
.A(n_2996),
.Y(n_3132)
);

INVx2_ASAP7_75t_SL g3133 ( 
.A(n_2971),
.Y(n_3133)
);

INVx3_ASAP7_75t_L g3134 ( 
.A(n_2954),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_SL g3135 ( 
.A(n_2835),
.B(n_2945),
.Y(n_3135)
);

INVx3_ASAP7_75t_L g3136 ( 
.A(n_2869),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_L g3137 ( 
.A(n_2847),
.B(n_801),
.Y(n_3137)
);

INVx2_ASAP7_75t_L g3138 ( 
.A(n_2886),
.Y(n_3138)
);

BUFx6f_ASAP7_75t_L g3139 ( 
.A(n_2980),
.Y(n_3139)
);

INVxp67_ASAP7_75t_SL g3140 ( 
.A(n_2889),
.Y(n_3140)
);

OR2x2_ASAP7_75t_L g3141 ( 
.A(n_2902),
.B(n_2934),
.Y(n_3141)
);

INVxp67_ASAP7_75t_L g3142 ( 
.A(n_2948),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_2816),
.B(n_802),
.Y(n_3143)
);

BUFx2_ASAP7_75t_L g3144 ( 
.A(n_2819),
.Y(n_3144)
);

BUFx6f_ASAP7_75t_L g3145 ( 
.A(n_2917),
.Y(n_3145)
);

INVx2_ASAP7_75t_L g3146 ( 
.A(n_2946),
.Y(n_3146)
);

BUFx6f_ASAP7_75t_L g3147 ( 
.A(n_2922),
.Y(n_3147)
);

NOR2xp67_ASAP7_75t_L g3148 ( 
.A(n_2882),
.B(n_2095),
.Y(n_3148)
);

AND2x2_ASAP7_75t_L g3149 ( 
.A(n_2808),
.B(n_783),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_SL g3150 ( 
.A(n_2983),
.B(n_2429),
.Y(n_3150)
);

OR2x6_ASAP7_75t_L g3151 ( 
.A(n_2811),
.B(n_2429),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2859),
.Y(n_3152)
);

BUFx2_ASAP7_75t_L g3153 ( 
.A(n_2988),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_2868),
.B(n_2433),
.Y(n_3154)
);

INVx4_ASAP7_75t_L g3155 ( 
.A(n_2991),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_2931),
.Y(n_3156)
);

BUFx2_ASAP7_75t_L g3157 ( 
.A(n_2956),
.Y(n_3157)
);

NAND2xp5_ASAP7_75t_L g3158 ( 
.A(n_2874),
.B(n_2433),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_SL g3159 ( 
.A(n_2915),
.B(n_2433),
.Y(n_3159)
);

INVxp33_ASAP7_75t_SL g3160 ( 
.A(n_2961),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2902),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2861),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_2962),
.Y(n_3163)
);

AOI221x1_ASAP7_75t_L g3164 ( 
.A1(n_2879),
.A2(n_2129),
.B1(n_2137),
.B2(n_2118),
.C(n_2117),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_2920),
.B(n_2117),
.Y(n_3165)
);

BUFx2_ASAP7_75t_L g3166 ( 
.A(n_2860),
.Y(n_3166)
);

BUFx4f_ASAP7_75t_L g3167 ( 
.A(n_2850),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_SL g3168 ( 
.A(n_2836),
.B(n_2332),
.Y(n_3168)
);

INVx4_ASAP7_75t_L g3169 ( 
.A(n_2994),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2962),
.Y(n_3170)
);

INVx4_ASAP7_75t_L g3171 ( 
.A(n_2967),
.Y(n_3171)
);

BUFx6f_ASAP7_75t_L g3172 ( 
.A(n_2921),
.Y(n_3172)
);

CKINVDCx5p33_ASAP7_75t_R g3173 ( 
.A(n_2914),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_SL g3174 ( 
.A(n_2947),
.B(n_2344),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2919),
.Y(n_3175)
);

INVxp67_ASAP7_75t_L g3176 ( 
.A(n_2899),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_SL g3177 ( 
.A(n_2953),
.B(n_2118),
.Y(n_3177)
);

INVx2_ASAP7_75t_L g3178 ( 
.A(n_2879),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_2880),
.Y(n_3179)
);

AND2x2_ASAP7_75t_L g3180 ( 
.A(n_2880),
.B(n_783),
.Y(n_3180)
);

HB1xp67_ASAP7_75t_L g3181 ( 
.A(n_2899),
.Y(n_3181)
);

NOR2xp33_ASAP7_75t_L g3182 ( 
.A(n_2872),
.B(n_794),
.Y(n_3182)
);

BUFx8_ASAP7_75t_SL g3183 ( 
.A(n_2982),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2909),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_L g3185 ( 
.A(n_2909),
.B(n_802),
.Y(n_3185)
);

INVx2_ASAP7_75t_SL g3186 ( 
.A(n_2985),
.Y(n_3186)
);

AND2x2_ASAP7_75t_L g3187 ( 
.A(n_2935),
.B(n_794),
.Y(n_3187)
);

AOI21xp5_ASAP7_75t_L g3188 ( 
.A1(n_2814),
.A2(n_1851),
.B(n_1807),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2957),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_L g3190 ( 
.A(n_2875),
.B(n_803),
.Y(n_3190)
);

NAND2xp5_ASAP7_75t_L g3191 ( 
.A(n_2878),
.B(n_2017),
.Y(n_3191)
);

INVx4_ASAP7_75t_L g3192 ( 
.A(n_2981),
.Y(n_3192)
);

BUFx6f_ASAP7_75t_L g3193 ( 
.A(n_2949),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_L g3194 ( 
.A(n_2852),
.B(n_2017),
.Y(n_3194)
);

INVx2_ASAP7_75t_L g3195 ( 
.A(n_2935),
.Y(n_3195)
);

BUFx10_ASAP7_75t_L g3196 ( 
.A(n_2940),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_SL g3197 ( 
.A(n_2818),
.B(n_2129),
.Y(n_3197)
);

INVx3_ASAP7_75t_L g3198 ( 
.A(n_3139),
.Y(n_3198)
);

HB1xp67_ASAP7_75t_L g3199 ( 
.A(n_3020),
.Y(n_3199)
);

AOI22xp5_ASAP7_75t_L g3200 ( 
.A1(n_3160),
.A2(n_2839),
.B1(n_2958),
.B2(n_2812),
.Y(n_3200)
);

BUFx12f_ASAP7_75t_L g3201 ( 
.A(n_3045),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_3003),
.Y(n_3202)
);

BUFx3_ASAP7_75t_L g3203 ( 
.A(n_3013),
.Y(n_3203)
);

NOR2xp33_ASAP7_75t_L g3204 ( 
.A(n_3126),
.B(n_4),
.Y(n_3204)
);

INVx1_ASAP7_75t_SL g3205 ( 
.A(n_3011),
.Y(n_3205)
);

AND2x2_ASAP7_75t_L g3206 ( 
.A(n_3055),
.B(n_3068),
.Y(n_3206)
);

AND2x4_ASAP7_75t_L g3207 ( 
.A(n_3000),
.B(n_2960),
.Y(n_3207)
);

BUFx6f_ASAP7_75t_L g3208 ( 
.A(n_3013),
.Y(n_3208)
);

AOI21xp5_ASAP7_75t_L g3209 ( 
.A1(n_3140),
.A2(n_2969),
.B(n_1851),
.Y(n_3209)
);

INVx3_ASAP7_75t_SL g3210 ( 
.A(n_3041),
.Y(n_3210)
);

BUFx8_ASAP7_75t_L g3211 ( 
.A(n_3004),
.Y(n_3211)
);

AOI22xp33_ASAP7_75t_SL g3212 ( 
.A1(n_3166),
.A2(n_2193),
.B1(n_1957),
.B2(n_2969),
.Y(n_3212)
);

O2A1O1Ixp33_ASAP7_75t_L g3213 ( 
.A1(n_3135),
.A2(n_2026),
.B(n_2030),
.C(n_2018),
.Y(n_3213)
);

AND2x2_ASAP7_75t_L g3214 ( 
.A(n_3068),
.B(n_4),
.Y(n_3214)
);

O2A1O1Ixp33_ASAP7_75t_L g3215 ( 
.A1(n_3185),
.A2(n_2026),
.B(n_2030),
.C(n_2018),
.Y(n_3215)
);

OAI22xp5_ASAP7_75t_L g3216 ( 
.A1(n_2998),
.A2(n_2363),
.B1(n_2150),
.B2(n_2153),
.Y(n_3216)
);

BUFx2_ASAP7_75t_L g3217 ( 
.A(n_3018),
.Y(n_3217)
);

INVx1_ASAP7_75t_L g3218 ( 
.A(n_2997),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_L g3219 ( 
.A(n_3090),
.B(n_5),
.Y(n_3219)
);

INVx2_ASAP7_75t_L g3220 ( 
.A(n_3046),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_3007),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_SL g3222 ( 
.A(n_3173),
.B(n_2137),
.Y(n_3222)
);

NOR2xp67_ASAP7_75t_L g3223 ( 
.A(n_3142),
.B(n_3112),
.Y(n_3223)
);

AND2x2_ASAP7_75t_SL g3224 ( 
.A(n_3167),
.B(n_3129),
.Y(n_3224)
);

HB1xp67_ASAP7_75t_L g3225 ( 
.A(n_3069),
.Y(n_3225)
);

INVx2_ASAP7_75t_L g3226 ( 
.A(n_3049),
.Y(n_3226)
);

NOR2xp33_ASAP7_75t_L g3227 ( 
.A(n_3132),
.B(n_3124),
.Y(n_3227)
);

NOR2xp33_ASAP7_75t_L g3228 ( 
.A(n_3034),
.B(n_5),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_3009),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_3101),
.B(n_6),
.Y(n_3230)
);

HB1xp67_ASAP7_75t_L g3231 ( 
.A(n_3108),
.Y(n_3231)
);

AOI21xp5_ASAP7_75t_L g3232 ( 
.A1(n_3005),
.A2(n_1807),
.B(n_2193),
.Y(n_3232)
);

HB1xp67_ASAP7_75t_L g3233 ( 
.A(n_3081),
.Y(n_3233)
);

AOI22xp5_ASAP7_75t_L g3234 ( 
.A1(n_3037),
.A2(n_1957),
.B1(n_2163),
.B2(n_2158),
.Y(n_3234)
);

INVx2_ASAP7_75t_L g3235 ( 
.A(n_3052),
.Y(n_3235)
);

AOI22xp33_ASAP7_75t_L g3236 ( 
.A1(n_3144),
.A2(n_1957),
.B1(n_2189),
.B2(n_2163),
.Y(n_3236)
);

AOI21xp5_ASAP7_75t_L g3237 ( 
.A1(n_3005),
.A2(n_1774),
.B(n_1767),
.Y(n_3237)
);

OAI22xp33_ASAP7_75t_L g3238 ( 
.A1(n_3143),
.A2(n_2198),
.B1(n_2204),
.B2(n_2189),
.Y(n_3238)
);

INVx2_ASAP7_75t_L g3239 ( 
.A(n_3054),
.Y(n_3239)
);

INVx2_ASAP7_75t_L g3240 ( 
.A(n_3057),
.Y(n_3240)
);

INVx2_ASAP7_75t_L g3241 ( 
.A(n_3025),
.Y(n_3241)
);

AOI221xp5_ASAP7_75t_L g3242 ( 
.A1(n_3120),
.A2(n_2032),
.B1(n_842),
.B2(n_951),
.C(n_831),
.Y(n_3242)
);

INVx2_ASAP7_75t_L g3243 ( 
.A(n_3028),
.Y(n_3243)
);

BUFx2_ASAP7_75t_L g3244 ( 
.A(n_3060),
.Y(n_3244)
);

AO21x1_ASAP7_75t_L g3245 ( 
.A1(n_3182),
.A2(n_9),
.B(n_11),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_3030),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_3059),
.Y(n_3247)
);

AOI21xp5_ASAP7_75t_L g3248 ( 
.A1(n_3125),
.A2(n_1774),
.B(n_1767),
.Y(n_3248)
);

NOR2x1_ASAP7_75t_L g3249 ( 
.A(n_3130),
.B(n_2198),
.Y(n_3249)
);

AOI21xp5_ASAP7_75t_L g3250 ( 
.A1(n_3067),
.A2(n_1786),
.B(n_1780),
.Y(n_3250)
);

AND2x4_ASAP7_75t_L g3251 ( 
.A(n_3039),
.B(n_3062),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_3082),
.Y(n_3252)
);

BUFx2_ASAP7_75t_SL g3253 ( 
.A(n_3013),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_3152),
.Y(n_3254)
);

NOR2xp33_ASAP7_75t_L g3255 ( 
.A(n_3021),
.B(n_9),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_3012),
.Y(n_3256)
);

AOI22xp33_ASAP7_75t_L g3257 ( 
.A1(n_3109),
.A2(n_1957),
.B1(n_2206),
.B2(n_2204),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_3012),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_3006),
.Y(n_3259)
);

INVx2_ASAP7_75t_L g3260 ( 
.A(n_3010),
.Y(n_3260)
);

AND2x4_ASAP7_75t_L g3261 ( 
.A(n_3039),
.B(n_2206),
.Y(n_3261)
);

AOI22xp33_ASAP7_75t_L g3262 ( 
.A1(n_3187),
.A2(n_1957),
.B1(n_2252),
.B2(n_2213),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_3175),
.Y(n_3263)
);

INVx3_ASAP7_75t_L g3264 ( 
.A(n_3139),
.Y(n_3264)
);

OAI22xp5_ASAP7_75t_L g3265 ( 
.A1(n_3137),
.A2(n_2363),
.B1(n_2252),
.B2(n_2256),
.Y(n_3265)
);

INVx2_ASAP7_75t_SL g3266 ( 
.A(n_3026),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_3091),
.B(n_12),
.Y(n_3267)
);

AOI21xp5_ASAP7_75t_L g3268 ( 
.A1(n_3148),
.A2(n_1786),
.B(n_1780),
.Y(n_3268)
);

INVx3_ASAP7_75t_L g3269 ( 
.A(n_3139),
.Y(n_3269)
);

INVx2_ASAP7_75t_L g3270 ( 
.A(n_3019),
.Y(n_3270)
);

AOI21xp5_ASAP7_75t_L g3271 ( 
.A1(n_3148),
.A2(n_1800),
.B(n_1792),
.Y(n_3271)
);

O2A1O1Ixp33_ASAP7_75t_L g3272 ( 
.A1(n_3106),
.A2(n_2032),
.B(n_2256),
.C(n_2213),
.Y(n_3272)
);

NAND2xp5_ASAP7_75t_SL g3273 ( 
.A(n_3162),
.B(n_2257),
.Y(n_3273)
);

BUFx2_ASAP7_75t_L g3274 ( 
.A(n_3070),
.Y(n_3274)
);

BUFx3_ASAP7_75t_L g3275 ( 
.A(n_3042),
.Y(n_3275)
);

O2A1O1Ixp33_ASAP7_75t_L g3276 ( 
.A1(n_3190),
.A2(n_2300),
.B(n_2331),
.C(n_2257),
.Y(n_3276)
);

INVx2_ASAP7_75t_SL g3277 ( 
.A(n_3026),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_3156),
.Y(n_3278)
);

INVx5_ASAP7_75t_L g3279 ( 
.A(n_3147),
.Y(n_3279)
);

INVx4_ASAP7_75t_L g3280 ( 
.A(n_3008),
.Y(n_3280)
);

AO21x2_ASAP7_75t_L g3281 ( 
.A1(n_3191),
.A2(n_1800),
.B(n_1792),
.Y(n_3281)
);

OAI221xp5_ASAP7_75t_L g3282 ( 
.A1(n_3076),
.A2(n_2334),
.B1(n_2347),
.B2(n_2331),
.C(n_2300),
.Y(n_3282)
);

A2O1A1Ixp33_ASAP7_75t_L g3283 ( 
.A1(n_3180),
.A2(n_2347),
.B(n_2334),
.C(n_1909),
.Y(n_3283)
);

INVx2_ASAP7_75t_L g3284 ( 
.A(n_3032),
.Y(n_3284)
);

AND2x4_ASAP7_75t_L g3285 ( 
.A(n_3094),
.B(n_1903),
.Y(n_3285)
);

BUFx6f_ASAP7_75t_L g3286 ( 
.A(n_3085),
.Y(n_3286)
);

AOI22xp33_ASAP7_75t_L g3287 ( 
.A1(n_3079),
.A2(n_1909),
.B1(n_1915),
.B2(n_1903),
.Y(n_3287)
);

INVx2_ASAP7_75t_L g3288 ( 
.A(n_3033),
.Y(n_3288)
);

BUFx6f_ASAP7_75t_L g3289 ( 
.A(n_3085),
.Y(n_3289)
);

NOR2x1_ASAP7_75t_L g3290 ( 
.A(n_3053),
.B(n_1903),
.Y(n_3290)
);

INVx2_ASAP7_75t_L g3291 ( 
.A(n_3038),
.Y(n_3291)
);

NOR2xp33_ASAP7_75t_L g3292 ( 
.A(n_3122),
.B(n_13),
.Y(n_3292)
);

AND2x4_ASAP7_75t_L g3293 ( 
.A(n_3094),
.B(n_1909),
.Y(n_3293)
);

A2O1A1Ixp33_ASAP7_75t_L g3294 ( 
.A1(n_3176),
.A2(n_1916),
.B(n_1925),
.C(n_1915),
.Y(n_3294)
);

BUFx3_ASAP7_75t_L g3295 ( 
.A(n_3014),
.Y(n_3295)
);

HB1xp67_ASAP7_75t_L g3296 ( 
.A(n_3158),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_SL g3297 ( 
.A(n_3077),
.B(n_3002),
.Y(n_3297)
);

INVxp67_ASAP7_75t_SL g3298 ( 
.A(n_3158),
.Y(n_3298)
);

AOI21xp5_ASAP7_75t_L g3299 ( 
.A1(n_3063),
.A2(n_3168),
.B(n_3107),
.Y(n_3299)
);

BUFx6f_ASAP7_75t_L g3300 ( 
.A(n_3085),
.Y(n_3300)
);

BUFx12f_ASAP7_75t_L g3301 ( 
.A(n_3133),
.Y(n_3301)
);

AND2x2_ASAP7_75t_L g3302 ( 
.A(n_3064),
.B(n_14),
.Y(n_3302)
);

BUFx6f_ASAP7_75t_L g3303 ( 
.A(n_3097),
.Y(n_3303)
);

AND2x2_ASAP7_75t_L g3304 ( 
.A(n_3157),
.B(n_14),
.Y(n_3304)
);

O2A1O1Ixp33_ASAP7_75t_L g3305 ( 
.A1(n_3119),
.A2(n_2057),
.B(n_2056),
.C(n_1915),
.Y(n_3305)
);

AOI222xp33_ASAP7_75t_L g3306 ( 
.A1(n_3093),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.C1(n_19),
.C2(n_20),
.Y(n_3306)
);

INVx6_ASAP7_75t_L g3307 ( 
.A(n_3097),
.Y(n_3307)
);

NOR2x1_ASAP7_75t_L g3308 ( 
.A(n_3053),
.B(n_1916),
.Y(n_3308)
);

AOI21xp5_ASAP7_75t_L g3309 ( 
.A1(n_3188),
.A2(n_1925),
.B(n_1916),
.Y(n_3309)
);

INVx4_ASAP7_75t_L g3310 ( 
.A(n_3008),
.Y(n_3310)
);

INVx5_ASAP7_75t_L g3311 ( 
.A(n_3147),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_SL g3312 ( 
.A(n_3002),
.B(n_1925),
.Y(n_3312)
);

AOI21xp5_ASAP7_75t_L g3313 ( 
.A1(n_3111),
.A2(n_2016),
.B(n_1962),
.Y(n_3313)
);

BUFx6f_ASAP7_75t_L g3314 ( 
.A(n_3097),
.Y(n_3314)
);

AND2x4_ASAP7_75t_L g3315 ( 
.A(n_2999),
.B(n_1962),
.Y(n_3315)
);

INVx2_ASAP7_75t_SL g3316 ( 
.A(n_3026),
.Y(n_3316)
);

INVx2_ASAP7_75t_L g3317 ( 
.A(n_3117),
.Y(n_3317)
);

AOI33xp33_ASAP7_75t_L g3318 ( 
.A1(n_3114),
.A2(n_16),
.A3(n_17),
.B1(n_18),
.B2(n_21),
.B3(n_22),
.Y(n_3318)
);

AOI21xp5_ASAP7_75t_L g3319 ( 
.A1(n_3111),
.A2(n_2016),
.B(n_1962),
.Y(n_3319)
);

NAND2xp5_ASAP7_75t_L g3320 ( 
.A(n_3095),
.B(n_21),
.Y(n_3320)
);

AOI21xp33_ASAP7_75t_L g3321 ( 
.A1(n_3149),
.A2(n_2039),
.B(n_2016),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_3131),
.Y(n_3322)
);

NOR2xp33_ASAP7_75t_L g3323 ( 
.A(n_3092),
.B(n_22),
.Y(n_3323)
);

INVx1_ASAP7_75t_SL g3324 ( 
.A(n_3022),
.Y(n_3324)
);

AOI21xp5_ASAP7_75t_L g3325 ( 
.A1(n_3194),
.A2(n_2058),
.B(n_2039),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_3184),
.Y(n_3326)
);

INVxp67_ASAP7_75t_L g3327 ( 
.A(n_3048),
.Y(n_3327)
);

INVx2_ASAP7_75t_L g3328 ( 
.A(n_3056),
.Y(n_3328)
);

BUFx6f_ASAP7_75t_L g3329 ( 
.A(n_3036),
.Y(n_3329)
);

AOI21xp5_ASAP7_75t_L g3330 ( 
.A1(n_3165),
.A2(n_2058),
.B(n_2039),
.Y(n_3330)
);

NOR2xp67_ASAP7_75t_L g3331 ( 
.A(n_2999),
.B(n_23),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_3104),
.B(n_24),
.Y(n_3332)
);

INVxp67_ASAP7_75t_L g3333 ( 
.A(n_3127),
.Y(n_3333)
);

O2A1O1Ixp33_ASAP7_75t_L g3334 ( 
.A1(n_3047),
.A2(n_2058),
.B(n_1503),
.C(n_1566),
.Y(n_3334)
);

INVx2_ASAP7_75t_L g3335 ( 
.A(n_3086),
.Y(n_3335)
);

AND2x4_ASAP7_75t_L g3336 ( 
.A(n_3001),
.B(n_253),
.Y(n_3336)
);

OAI22xp5_ASAP7_75t_L g3337 ( 
.A1(n_3075),
.A2(n_3145),
.B1(n_3023),
.B2(n_3029),
.Y(n_3337)
);

INVx3_ASAP7_75t_L g3338 ( 
.A(n_3016),
.Y(n_3338)
);

O2A1O1Ixp5_ASAP7_75t_L g3339 ( 
.A1(n_3072),
.A2(n_2037),
.B(n_1503),
.C(n_1566),
.Y(n_3339)
);

A2O1A1Ixp33_ASAP7_75t_SL g3340 ( 
.A1(n_3121),
.A2(n_1559),
.B(n_26),
.C(n_24),
.Y(n_3340)
);

INVx4_ASAP7_75t_L g3341 ( 
.A(n_3008),
.Y(n_3341)
);

O2A1O1Ixp33_ASAP7_75t_L g3342 ( 
.A1(n_3040),
.A2(n_1559),
.B(n_27),
.C(n_25),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_3141),
.Y(n_3343)
);

AND2x4_ASAP7_75t_L g3344 ( 
.A(n_3001),
.B(n_255),
.Y(n_3344)
);

INVx3_ASAP7_75t_L g3345 ( 
.A(n_3016),
.Y(n_3345)
);

INVx2_ASAP7_75t_L g3346 ( 
.A(n_3089),
.Y(n_3346)
);

NOR2xp67_ASAP7_75t_L g3347 ( 
.A(n_3084),
.B(n_26),
.Y(n_3347)
);

INVx2_ASAP7_75t_L g3348 ( 
.A(n_3113),
.Y(n_3348)
);

AOI21xp5_ASAP7_75t_L g3349 ( 
.A1(n_3165),
.A2(n_2037),
.B(n_1571),
.Y(n_3349)
);

CKINVDCx20_ASAP7_75t_R g3350 ( 
.A(n_3031),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3154),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3154),
.Y(n_3352)
);

AND2x4_ASAP7_75t_L g3353 ( 
.A(n_3113),
.B(n_258),
.Y(n_3353)
);

NAND2x1p5_ASAP7_75t_L g3354 ( 
.A(n_3150),
.B(n_2037),
.Y(n_3354)
);

BUFx6f_ASAP7_75t_L g3355 ( 
.A(n_3036),
.Y(n_3355)
);

AND2x2_ASAP7_75t_L g3356 ( 
.A(n_3181),
.B(n_27),
.Y(n_3356)
);

BUFx6f_ASAP7_75t_L g3357 ( 
.A(n_3036),
.Y(n_3357)
);

NOR2xp33_ASAP7_75t_L g3358 ( 
.A(n_3074),
.B(n_29),
.Y(n_3358)
);

NAND3xp33_ASAP7_75t_L g3359 ( 
.A(n_3075),
.B(n_831),
.C(n_813),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3123),
.Y(n_3360)
);

NOR2xp33_ASAP7_75t_L g3361 ( 
.A(n_3087),
.B(n_29),
.Y(n_3361)
);

O2A1O1Ixp33_ASAP7_75t_SL g3362 ( 
.A1(n_3015),
.A2(n_33),
.B(n_31),
.C(n_32),
.Y(n_3362)
);

HB1xp67_ASAP7_75t_L g3363 ( 
.A(n_3105),
.Y(n_3363)
);

INVx2_ASAP7_75t_SL g3364 ( 
.A(n_3065),
.Y(n_3364)
);

AOI22xp33_ASAP7_75t_L g3365 ( 
.A1(n_3153),
.A2(n_1571),
.B1(n_1564),
.B2(n_1527),
.Y(n_3365)
);

AND2x4_ASAP7_75t_L g3366 ( 
.A(n_3134),
.B(n_259),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_3163),
.Y(n_3367)
);

AND2x4_ASAP7_75t_L g3368 ( 
.A(n_3134),
.B(n_260),
.Y(n_3368)
);

INVx1_ASAP7_75t_L g3369 ( 
.A(n_3170),
.Y(n_3369)
);

A2O1A1Ixp33_ASAP7_75t_L g3370 ( 
.A1(n_3115),
.A2(n_34),
.B(n_31),
.C(n_33),
.Y(n_3370)
);

BUFx2_ASAP7_75t_L g3371 ( 
.A(n_3024),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_L g3372 ( 
.A(n_3116),
.B(n_35),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_3050),
.B(n_35),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_3035),
.Y(n_3374)
);

AOI21xp5_ASAP7_75t_L g3375 ( 
.A1(n_3078),
.A2(n_1571),
.B(n_1564),
.Y(n_3375)
);

AND2x2_ASAP7_75t_L g3376 ( 
.A(n_3110),
.B(n_3118),
.Y(n_3376)
);

INVx1_ASAP7_75t_SL g3377 ( 
.A(n_3065),
.Y(n_3377)
);

INVx3_ASAP7_75t_L g3378 ( 
.A(n_3065),
.Y(n_3378)
);

AND2x2_ASAP7_75t_L g3379 ( 
.A(n_3110),
.B(n_36),
.Y(n_3379)
);

AND2x4_ASAP7_75t_L g3380 ( 
.A(n_3080),
.B(n_263),
.Y(n_3380)
);

AOI22xp33_ASAP7_75t_L g3381 ( 
.A1(n_3174),
.A2(n_1571),
.B1(n_1564),
.B2(n_1527),
.Y(n_3381)
);

AND2x4_ASAP7_75t_L g3382 ( 
.A(n_3155),
.B(n_264),
.Y(n_3382)
);

INVx2_ASAP7_75t_SL g3383 ( 
.A(n_3024),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_3161),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_3044),
.B(n_37),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_3189),
.Y(n_3386)
);

INVx2_ASAP7_75t_L g3387 ( 
.A(n_3043),
.Y(n_3387)
);

OAI22xp5_ASAP7_75t_L g3388 ( 
.A1(n_3145),
.A2(n_831),
.B1(n_842),
.B2(n_813),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_3179),
.Y(n_3389)
);

INVx2_ASAP7_75t_L g3390 ( 
.A(n_3043),
.Y(n_3390)
);

OR2x6_ASAP7_75t_L g3391 ( 
.A(n_3151),
.B(n_813),
.Y(n_3391)
);

BUFx6f_ASAP7_75t_L g3392 ( 
.A(n_3071),
.Y(n_3392)
);

HB1xp67_ASAP7_75t_L g3393 ( 
.A(n_3151),
.Y(n_3393)
);

BUFx6f_ASAP7_75t_L g3394 ( 
.A(n_3071),
.Y(n_3394)
);

O2A1O1Ixp33_ASAP7_75t_SL g3395 ( 
.A1(n_3159),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_3395)
);

O2A1O1Ixp33_ASAP7_75t_L g3396 ( 
.A1(n_3040),
.A2(n_42),
.B(n_39),
.C(n_41),
.Y(n_3396)
);

AND2x2_ASAP7_75t_L g3397 ( 
.A(n_3118),
.B(n_43),
.Y(n_3397)
);

OAI22xp33_ASAP7_75t_L g3398 ( 
.A1(n_3171),
.A2(n_3102),
.B1(n_3100),
.B2(n_3128),
.Y(n_3398)
);

AOI22xp5_ASAP7_75t_L g3399 ( 
.A1(n_3058),
.A2(n_1553),
.B1(n_1527),
.B2(n_1529),
.Y(n_3399)
);

AOI21xp5_ASAP7_75t_L g3400 ( 
.A1(n_3164),
.A2(n_1522),
.B(n_1489),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_3017),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_3017),
.Y(n_3402)
);

INVx2_ASAP7_75t_L g3403 ( 
.A(n_3073),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_3051),
.Y(n_3404)
);

INVx2_ASAP7_75t_SL g3405 ( 
.A(n_3073),
.Y(n_3405)
);

BUFx6f_ASAP7_75t_L g3406 ( 
.A(n_3208),
.Y(n_3406)
);

INVx3_ASAP7_75t_L g3407 ( 
.A(n_3251),
.Y(n_3407)
);

INVx2_ASAP7_75t_L g3408 ( 
.A(n_3241),
.Y(n_3408)
);

AOI21xp5_ASAP7_75t_L g3409 ( 
.A1(n_3299),
.A2(n_3197),
.B(n_3177),
.Y(n_3409)
);

INVx2_ASAP7_75t_L g3410 ( 
.A(n_3243),
.Y(n_3410)
);

NAND2xp5_ASAP7_75t_L g3411 ( 
.A(n_3231),
.B(n_3178),
.Y(n_3411)
);

INVx1_ASAP7_75t_SL g3412 ( 
.A(n_3205),
.Y(n_3412)
);

OAI22xp5_ASAP7_75t_L g3413 ( 
.A1(n_3224),
.A2(n_3171),
.B1(n_3151),
.B2(n_3155),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_3202),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3343),
.B(n_3195),
.Y(n_3415)
);

HB1xp67_ASAP7_75t_L g3416 ( 
.A(n_3296),
.Y(n_3416)
);

AND2x4_ASAP7_75t_L g3417 ( 
.A(n_3251),
.B(n_3061),
.Y(n_3417)
);

AND2x2_ASAP7_75t_L g3418 ( 
.A(n_3206),
.B(n_3147),
.Y(n_3418)
);

INVx3_ASAP7_75t_L g3419 ( 
.A(n_3198),
.Y(n_3419)
);

OR2x6_ASAP7_75t_L g3420 ( 
.A(n_3253),
.B(n_3186),
.Y(n_3420)
);

BUFx6f_ASAP7_75t_L g3421 ( 
.A(n_3208),
.Y(n_3421)
);

INVx3_ASAP7_75t_L g3422 ( 
.A(n_3198),
.Y(n_3422)
);

AO22x1_ASAP7_75t_L g3423 ( 
.A1(n_3298),
.A2(n_3066),
.B1(n_3136),
.B2(n_3193),
.Y(n_3423)
);

BUFx2_ASAP7_75t_L g3424 ( 
.A(n_3199),
.Y(n_3424)
);

BUFx3_ASAP7_75t_L g3425 ( 
.A(n_3275),
.Y(n_3425)
);

AOI21xp5_ASAP7_75t_L g3426 ( 
.A1(n_3359),
.A2(n_3098),
.B(n_3027),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_L g3427 ( 
.A(n_3328),
.B(n_3138),
.Y(n_3427)
);

CKINVDCx5p33_ASAP7_75t_R g3428 ( 
.A(n_3210),
.Y(n_3428)
);

INVx2_ASAP7_75t_L g3429 ( 
.A(n_3220),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_L g3430 ( 
.A(n_3401),
.B(n_3402),
.Y(n_3430)
);

NOR2xp33_ASAP7_75t_L g3431 ( 
.A(n_3398),
.B(n_3083),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3202),
.Y(n_3432)
);

BUFx4f_ASAP7_75t_SL g3433 ( 
.A(n_3201),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_3351),
.Y(n_3434)
);

CKINVDCx5p33_ASAP7_75t_R g3435 ( 
.A(n_3211),
.Y(n_3435)
);

AND2x4_ASAP7_75t_L g3436 ( 
.A(n_3393),
.B(n_3061),
.Y(n_3436)
);

BUFx4_ASAP7_75t_SL g3437 ( 
.A(n_3295),
.Y(n_3437)
);

INVx1_ASAP7_75t_L g3438 ( 
.A(n_3221),
.Y(n_3438)
);

AOI22xp33_ASAP7_75t_L g3439 ( 
.A1(n_3245),
.A2(n_3183),
.B1(n_3172),
.B2(n_3192),
.Y(n_3439)
);

INVx3_ASAP7_75t_L g3440 ( 
.A(n_3264),
.Y(n_3440)
);

AOI21xp5_ASAP7_75t_L g3441 ( 
.A1(n_3312),
.A2(n_3098),
.B(n_3169),
.Y(n_3441)
);

NOR2x1_ASAP7_75t_SL g3442 ( 
.A(n_3297),
.B(n_3278),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_3229),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_3404),
.B(n_3172),
.Y(n_3444)
);

INVx5_ASAP7_75t_L g3445 ( 
.A(n_3208),
.Y(n_3445)
);

NOR2xp33_ASAP7_75t_L g3446 ( 
.A(n_3333),
.B(n_3255),
.Y(n_3446)
);

BUFx6f_ASAP7_75t_L g3447 ( 
.A(n_3203),
.Y(n_3447)
);

AOI22xp5_ASAP7_75t_L g3448 ( 
.A1(n_3337),
.A2(n_3066),
.B1(n_3192),
.B2(n_3196),
.Y(n_3448)
);

OAI22xp5_ASAP7_75t_L g3449 ( 
.A1(n_3370),
.A2(n_3096),
.B1(n_3136),
.B2(n_3193),
.Y(n_3449)
);

A2O1A1Ixp33_ASAP7_75t_SL g3450 ( 
.A1(n_3396),
.A2(n_3146),
.B(n_3088),
.C(n_3196),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_3246),
.Y(n_3451)
);

INVx2_ASAP7_75t_L g3452 ( 
.A(n_3226),
.Y(n_3452)
);

AOI22xp5_ASAP7_75t_L g3453 ( 
.A1(n_3306),
.A2(n_3066),
.B1(n_3172),
.B2(n_3193),
.Y(n_3453)
);

INVx2_ASAP7_75t_L g3454 ( 
.A(n_3235),
.Y(n_3454)
);

OR2x6_ASAP7_75t_L g3455 ( 
.A(n_3223),
.B(n_3099),
.Y(n_3455)
);

INVx3_ASAP7_75t_L g3456 ( 
.A(n_3264),
.Y(n_3456)
);

NAND2x1p5_ASAP7_75t_L g3457 ( 
.A(n_3280),
.B(n_3099),
.Y(n_3457)
);

OR2x2_ASAP7_75t_L g3458 ( 
.A(n_3376),
.B(n_3103),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_3352),
.Y(n_3459)
);

BUFx6f_ASAP7_75t_L g3460 ( 
.A(n_3329),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_L g3461 ( 
.A(n_3233),
.B(n_3066),
.Y(n_3461)
);

INVx2_ASAP7_75t_L g3462 ( 
.A(n_3239),
.Y(n_3462)
);

HB1xp67_ASAP7_75t_L g3463 ( 
.A(n_3225),
.Y(n_3463)
);

BUFx3_ASAP7_75t_L g3464 ( 
.A(n_3211),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_3240),
.Y(n_3465)
);

AOI22xp33_ASAP7_75t_L g3466 ( 
.A1(n_3358),
.A2(n_1527),
.B1(n_1529),
.B2(n_1526),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_L g3467 ( 
.A(n_3256),
.B(n_43),
.Y(n_3467)
);

INVx2_ASAP7_75t_L g3468 ( 
.A(n_3247),
.Y(n_3468)
);

INVx5_ASAP7_75t_L g3469 ( 
.A(n_3280),
.Y(n_3469)
);

AOI21xp5_ASAP7_75t_L g3470 ( 
.A1(n_3334),
.A2(n_1522),
.B(n_1489),
.Y(n_3470)
);

INVx1_ASAP7_75t_SL g3471 ( 
.A(n_3217),
.Y(n_3471)
);

INVx1_ASAP7_75t_SL g3472 ( 
.A(n_3301),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_L g3473 ( 
.A(n_3258),
.B(n_44),
.Y(n_3473)
);

INVx3_ASAP7_75t_L g3474 ( 
.A(n_3269),
.Y(n_3474)
);

INVx4_ASAP7_75t_L g3475 ( 
.A(n_3310),
.Y(n_3475)
);

AND2x4_ASAP7_75t_L g3476 ( 
.A(n_3207),
.B(n_44),
.Y(n_3476)
);

INVx2_ASAP7_75t_L g3477 ( 
.A(n_3252),
.Y(n_3477)
);

BUFx6f_ASAP7_75t_L g3478 ( 
.A(n_3329),
.Y(n_3478)
);

HB1xp67_ASAP7_75t_L g3479 ( 
.A(n_3363),
.Y(n_3479)
);

INVx3_ASAP7_75t_L g3480 ( 
.A(n_3269),
.Y(n_3480)
);

NAND3xp33_ASAP7_75t_L g3481 ( 
.A(n_3318),
.B(n_842),
.C(n_831),
.Y(n_3481)
);

INVx2_ASAP7_75t_L g3482 ( 
.A(n_3218),
.Y(n_3482)
);

AND2x4_ASAP7_75t_L g3483 ( 
.A(n_3207),
.B(n_45),
.Y(n_3483)
);

INVx2_ASAP7_75t_SL g3484 ( 
.A(n_3307),
.Y(n_3484)
);

AOI22xp33_ASAP7_75t_L g3485 ( 
.A1(n_3361),
.A2(n_1529),
.B1(n_1533),
.B2(n_1526),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3254),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3263),
.Y(n_3487)
);

BUFx3_ASAP7_75t_L g3488 ( 
.A(n_3244),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_L g3489 ( 
.A(n_3374),
.B(n_46),
.Y(n_3489)
);

AO32x2_ASAP7_75t_L g3490 ( 
.A1(n_3383),
.A2(n_46),
.A3(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_3490)
);

INVx2_ASAP7_75t_L g3491 ( 
.A(n_3274),
.Y(n_3491)
);

CKINVDCx6p67_ASAP7_75t_R g3492 ( 
.A(n_3324),
.Y(n_3492)
);

BUFx12f_ASAP7_75t_L g3493 ( 
.A(n_3214),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3278),
.Y(n_3494)
);

AOI22xp5_ASAP7_75t_L g3495 ( 
.A1(n_3200),
.A2(n_1529),
.B1(n_1533),
.B2(n_1526),
.Y(n_3495)
);

INVx2_ASAP7_75t_SL g3496 ( 
.A(n_3307),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3327),
.B(n_47),
.Y(n_3497)
);

INVx2_ASAP7_75t_L g3498 ( 
.A(n_3360),
.Y(n_3498)
);

AO21x1_ASAP7_75t_L g3499 ( 
.A1(n_3228),
.A2(n_53),
.B(n_56),
.Y(n_3499)
);

AO21x2_ASAP7_75t_L g3500 ( 
.A1(n_3349),
.A2(n_53),
.B(n_56),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3386),
.Y(n_3501)
);

INVx3_ASAP7_75t_L g3502 ( 
.A(n_3387),
.Y(n_3502)
);

AOI22xp33_ASAP7_75t_L g3503 ( 
.A1(n_3347),
.A2(n_1550),
.B1(n_1553),
.B2(n_1533),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_3335),
.B(n_57),
.Y(n_3504)
);

BUFx4_ASAP7_75t_SL g3505 ( 
.A(n_3350),
.Y(n_3505)
);

INVx3_ASAP7_75t_L g3506 ( 
.A(n_3390),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3386),
.Y(n_3507)
);

HB1xp67_ASAP7_75t_L g3508 ( 
.A(n_3326),
.Y(n_3508)
);

O2A1O1Ixp33_ASAP7_75t_L g3509 ( 
.A1(n_3342),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_3509)
);

OAI22xp5_ASAP7_75t_L g3510 ( 
.A1(n_3222),
.A2(n_3399),
.B1(n_3257),
.B2(n_3234),
.Y(n_3510)
);

OR2x6_ASAP7_75t_L g3511 ( 
.A(n_3310),
.B(n_3341),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_L g3512 ( 
.A(n_3346),
.B(n_58),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_L g3513 ( 
.A(n_3379),
.B(n_59),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3384),
.Y(n_3514)
);

NOR2xp33_ASAP7_75t_L g3515 ( 
.A(n_3227),
.B(n_60),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3384),
.Y(n_3516)
);

INVx2_ASAP7_75t_L g3517 ( 
.A(n_3317),
.Y(n_3517)
);

BUFx6f_ASAP7_75t_L g3518 ( 
.A(n_3329),
.Y(n_3518)
);

INVx1_ASAP7_75t_L g3519 ( 
.A(n_3389),
.Y(n_3519)
);

HB1xp67_ASAP7_75t_L g3520 ( 
.A(n_3326),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_3389),
.Y(n_3521)
);

OAI22xp5_ASAP7_75t_L g3522 ( 
.A1(n_3282),
.A2(n_951),
.B1(n_1010),
.B2(n_842),
.Y(n_3522)
);

INVx4_ASAP7_75t_L g3523 ( 
.A(n_3341),
.Y(n_3523)
);

INVx2_ASAP7_75t_SL g3524 ( 
.A(n_3355),
.Y(n_3524)
);

AND2x2_ASAP7_75t_L g3525 ( 
.A(n_3371),
.B(n_60),
.Y(n_3525)
);

AND2x4_ASAP7_75t_L g3526 ( 
.A(n_3348),
.B(n_61),
.Y(n_3526)
);

OR2x2_ASAP7_75t_L g3527 ( 
.A(n_3367),
.B(n_62),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_3397),
.B(n_62),
.Y(n_3528)
);

O2A1O1Ixp33_ASAP7_75t_SL g3529 ( 
.A1(n_3323),
.A2(n_65),
.B(n_63),
.C(n_64),
.Y(n_3529)
);

BUFx6f_ASAP7_75t_L g3530 ( 
.A(n_3355),
.Y(n_3530)
);

NOR2xp33_ASAP7_75t_L g3531 ( 
.A(n_3320),
.B(n_65),
.Y(n_3531)
);

AOI21xp5_ASAP7_75t_L g3532 ( 
.A1(n_3209),
.A2(n_1523),
.B(n_1489),
.Y(n_3532)
);

BUFx3_ASAP7_75t_L g3533 ( 
.A(n_3355),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_L g3534 ( 
.A(n_3259),
.B(n_66),
.Y(n_3534)
);

INVx1_ASAP7_75t_SL g3535 ( 
.A(n_3377),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3367),
.Y(n_3536)
);

INVx2_ASAP7_75t_SL g3537 ( 
.A(n_3357),
.Y(n_3537)
);

INVx3_ASAP7_75t_L g3538 ( 
.A(n_3403),
.Y(n_3538)
);

AOI22xp33_ASAP7_75t_L g3539 ( 
.A1(n_3380),
.A2(n_1550),
.B1(n_1553),
.B2(n_1533),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_3369),
.Y(n_3540)
);

BUFx6f_ASAP7_75t_L g3541 ( 
.A(n_3357),
.Y(n_3541)
);

BUFx6f_ASAP7_75t_L g3542 ( 
.A(n_3357),
.Y(n_3542)
);

INVx4_ASAP7_75t_L g3543 ( 
.A(n_3338),
.Y(n_3543)
);

INVx2_ASAP7_75t_SL g3544 ( 
.A(n_3286),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3369),
.Y(n_3545)
);

INVx4_ASAP7_75t_L g3546 ( 
.A(n_3338),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3260),
.Y(n_3547)
);

AND2x2_ASAP7_75t_L g3548 ( 
.A(n_3322),
.B(n_66),
.Y(n_3548)
);

NOR2x1_ASAP7_75t_L g3549 ( 
.A(n_3249),
.B(n_951),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_3270),
.B(n_67),
.Y(n_3550)
);

BUFx6f_ASAP7_75t_L g3551 ( 
.A(n_3286),
.Y(n_3551)
);

BUFx2_ASAP7_75t_L g3552 ( 
.A(n_3286),
.Y(n_3552)
);

INVx2_ASAP7_75t_L g3553 ( 
.A(n_3284),
.Y(n_3553)
);

NOR2xp33_ASAP7_75t_L g3554 ( 
.A(n_3267),
.B(n_67),
.Y(n_3554)
);

INVx1_ASAP7_75t_L g3555 ( 
.A(n_3288),
.Y(n_3555)
);

CKINVDCx5p33_ASAP7_75t_R g3556 ( 
.A(n_3289),
.Y(n_3556)
);

INVx2_ASAP7_75t_SL g3557 ( 
.A(n_3289),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_3291),
.B(n_68),
.Y(n_3558)
);

AOI22xp5_ASAP7_75t_L g3559 ( 
.A1(n_3331),
.A2(n_1553),
.B1(n_1550),
.B2(n_1010),
.Y(n_3559)
);

INVx2_ASAP7_75t_L g3560 ( 
.A(n_3405),
.Y(n_3560)
);

AOI21xp5_ASAP7_75t_L g3561 ( 
.A1(n_3340),
.A2(n_1523),
.B(n_1550),
.Y(n_3561)
);

INVx2_ASAP7_75t_SL g3562 ( 
.A(n_3289),
.Y(n_3562)
);

INVx2_ASAP7_75t_L g3563 ( 
.A(n_3378),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_3356),
.B(n_68),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3219),
.Y(n_3565)
);

AOI222xp33_ASAP7_75t_L g3566 ( 
.A1(n_3204),
.A2(n_70),
.B1(n_72),
.B2(n_74),
.C1(n_75),
.C2(n_76),
.Y(n_3566)
);

OR2x6_ASAP7_75t_L g3567 ( 
.A(n_3391),
.B(n_951),
.Y(n_3567)
);

AND2x2_ASAP7_75t_L g3568 ( 
.A(n_3392),
.B(n_70),
.Y(n_3568)
);

BUFx2_ASAP7_75t_L g3569 ( 
.A(n_3300),
.Y(n_3569)
);

INVx2_ASAP7_75t_SL g3570 ( 
.A(n_3300),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3230),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3290),
.Y(n_3572)
);

AOI222xp33_ASAP7_75t_L g3573 ( 
.A1(n_3304),
.A2(n_72),
.B1(n_78),
.B2(n_79),
.C1(n_80),
.C2(n_82),
.Y(n_3573)
);

BUFx4f_ASAP7_75t_L g3574 ( 
.A(n_3492),
.Y(n_3574)
);

OAI21x1_ASAP7_75t_L g3575 ( 
.A1(n_3409),
.A2(n_3232),
.B(n_3308),
.Y(n_3575)
);

O2A1O1Ixp33_ASAP7_75t_SL g3576 ( 
.A1(n_3471),
.A2(n_3372),
.B(n_3332),
.C(n_3292),
.Y(n_3576)
);

OR2x2_ASAP7_75t_L g3577 ( 
.A(n_3416),
.B(n_3385),
.Y(n_3577)
);

HB1xp67_ASAP7_75t_L g3578 ( 
.A(n_3463),
.Y(n_3578)
);

OA21x2_ASAP7_75t_L g3579 ( 
.A1(n_3494),
.A2(n_3375),
.B(n_3273),
.Y(n_3579)
);

AOI22xp5_ASAP7_75t_L g3580 ( 
.A1(n_3413),
.A2(n_3238),
.B1(n_3380),
.B2(n_3382),
.Y(n_3580)
);

OR2x2_ASAP7_75t_L g3581 ( 
.A(n_3491),
.B(n_3373),
.Y(n_3581)
);

NAND2x1p5_ASAP7_75t_L g3582 ( 
.A(n_3445),
.B(n_3279),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3494),
.Y(n_3583)
);

OAI21x1_ASAP7_75t_L g3584 ( 
.A1(n_3549),
.A2(n_3237),
.B(n_3330),
.Y(n_3584)
);

OAI22x1_ASAP7_75t_L g3585 ( 
.A1(n_3424),
.A2(n_3302),
.B1(n_3277),
.B2(n_3266),
.Y(n_3585)
);

NOR2x1_ASAP7_75t_SL g3586 ( 
.A(n_3420),
.B(n_3391),
.Y(n_3586)
);

OR2x2_ASAP7_75t_L g3587 ( 
.A(n_3479),
.B(n_3281),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3508),
.Y(n_3588)
);

OAI21x1_ASAP7_75t_L g3589 ( 
.A1(n_3441),
.A2(n_3248),
.B(n_3268),
.Y(n_3589)
);

HB1xp67_ASAP7_75t_L g3590 ( 
.A(n_3520),
.Y(n_3590)
);

INVx1_ASAP7_75t_L g3591 ( 
.A(n_3414),
.Y(n_3591)
);

AOI211xp5_ASAP7_75t_L g3592 ( 
.A1(n_3499),
.A2(n_3395),
.B(n_3362),
.C(n_3321),
.Y(n_3592)
);

INVx6_ASAP7_75t_L g3593 ( 
.A(n_3447),
.Y(n_3593)
);

OA21x2_ASAP7_75t_L g3594 ( 
.A1(n_3501),
.A2(n_3294),
.B(n_3271),
.Y(n_3594)
);

NOR2xp33_ASAP7_75t_L g3595 ( 
.A(n_3428),
.B(n_3392),
.Y(n_3595)
);

INVx1_ASAP7_75t_L g3596 ( 
.A(n_3432),
.Y(n_3596)
);

AOI22xp33_ASAP7_75t_L g3597 ( 
.A1(n_3566),
.A2(n_3382),
.B1(n_3261),
.B2(n_3265),
.Y(n_3597)
);

O2A1O1Ixp33_ASAP7_75t_L g3598 ( 
.A1(n_3529),
.A2(n_3283),
.B(n_3216),
.C(n_3276),
.Y(n_3598)
);

OAI21x1_ASAP7_75t_SL g3599 ( 
.A1(n_3442),
.A2(n_3364),
.B(n_3316),
.Y(n_3599)
);

OAI21x1_ASAP7_75t_L g3600 ( 
.A1(n_3532),
.A2(n_3572),
.B(n_3426),
.Y(n_3600)
);

INVx5_ASAP7_75t_L g3601 ( 
.A(n_3511),
.Y(n_3601)
);

OAI21xp5_ASAP7_75t_L g3602 ( 
.A1(n_3509),
.A2(n_3554),
.B(n_3531),
.Y(n_3602)
);

OAI21x1_ASAP7_75t_L g3603 ( 
.A1(n_3448),
.A2(n_3325),
.B(n_3400),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_L g3604 ( 
.A(n_3434),
.B(n_3261),
.Y(n_3604)
);

INVx1_ASAP7_75t_L g3605 ( 
.A(n_3514),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3516),
.Y(n_3606)
);

AND2x2_ASAP7_75t_L g3607 ( 
.A(n_3407),
.B(n_3394),
.Y(n_3607)
);

OAI21x1_ASAP7_75t_L g3608 ( 
.A1(n_3457),
.A2(n_3339),
.B(n_3345),
.Y(n_3608)
);

INVxp67_ASAP7_75t_SL g3609 ( 
.A(n_3442),
.Y(n_3609)
);

NAND2x1p5_ASAP7_75t_L g3610 ( 
.A(n_3445),
.B(n_3279),
.Y(n_3610)
);

BUFx3_ASAP7_75t_L g3611 ( 
.A(n_3464),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3519),
.Y(n_3612)
);

OAI21xp5_ASAP7_75t_L g3613 ( 
.A1(n_3481),
.A2(n_3305),
.B(n_3353),
.Y(n_3613)
);

NOR2xp67_ASAP7_75t_L g3614 ( 
.A(n_3469),
.B(n_3279),
.Y(n_3614)
);

OAI21x1_ASAP7_75t_L g3615 ( 
.A1(n_3444),
.A2(n_3345),
.B(n_3319),
.Y(n_3615)
);

AND2x4_ASAP7_75t_L g3616 ( 
.A(n_3436),
.B(n_3311),
.Y(n_3616)
);

OAI21xp5_ASAP7_75t_L g3617 ( 
.A1(n_3431),
.A2(n_3366),
.B(n_3353),
.Y(n_3617)
);

CKINVDCx5p33_ASAP7_75t_R g3618 ( 
.A(n_3435),
.Y(n_3618)
);

HB1xp67_ASAP7_75t_L g3619 ( 
.A(n_3411),
.Y(n_3619)
);

INVxp67_ASAP7_75t_L g3620 ( 
.A(n_3565),
.Y(n_3620)
);

CKINVDCx16_ASAP7_75t_R g3621 ( 
.A(n_3493),
.Y(n_3621)
);

OA21x2_ASAP7_75t_L g3622 ( 
.A1(n_3507),
.A2(n_3313),
.B(n_3309),
.Y(n_3622)
);

NOR2xp33_ASAP7_75t_SL g3623 ( 
.A(n_3433),
.B(n_3336),
.Y(n_3623)
);

INVx2_ASAP7_75t_L g3624 ( 
.A(n_3459),
.Y(n_3624)
);

NAND2x1p5_ASAP7_75t_L g3625 ( 
.A(n_3445),
.B(n_3311),
.Y(n_3625)
);

INVx1_ASAP7_75t_L g3626 ( 
.A(n_3521),
.Y(n_3626)
);

AND2x4_ASAP7_75t_L g3627 ( 
.A(n_3436),
.B(n_3311),
.Y(n_3627)
);

OAI221xp5_ASAP7_75t_L g3628 ( 
.A1(n_3439),
.A2(n_3262),
.B1(n_3394),
.B2(n_3392),
.C(n_3287),
.Y(n_3628)
);

AOI21xp5_ASAP7_75t_L g3629 ( 
.A1(n_3450),
.A2(n_3215),
.B(n_3272),
.Y(n_3629)
);

BUFx4f_ASAP7_75t_L g3630 ( 
.A(n_3447),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3536),
.Y(n_3631)
);

OAI21x1_ASAP7_75t_L g3632 ( 
.A1(n_3427),
.A2(n_3354),
.B(n_3378),
.Y(n_3632)
);

AND2x4_ASAP7_75t_L g3633 ( 
.A(n_3407),
.B(n_3303),
.Y(n_3633)
);

AOI21xp5_ASAP7_75t_L g3634 ( 
.A1(n_3423),
.A2(n_3242),
.B(n_3250),
.Y(n_3634)
);

OAI21xp5_ASAP7_75t_L g3635 ( 
.A1(n_3446),
.A2(n_3368),
.B(n_3366),
.Y(n_3635)
);

INVx2_ASAP7_75t_SL g3636 ( 
.A(n_3437),
.Y(n_3636)
);

OAI21x1_ASAP7_75t_L g3637 ( 
.A1(n_3470),
.A2(n_3388),
.B(n_3381),
.Y(n_3637)
);

INVx1_ASAP7_75t_L g3638 ( 
.A(n_3540),
.Y(n_3638)
);

NOR2xp33_ASAP7_75t_L g3639 ( 
.A(n_3472),
.B(n_3394),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3545),
.Y(n_3640)
);

BUFx2_ASAP7_75t_R g3641 ( 
.A(n_3425),
.Y(n_3641)
);

OAI222xp33_ASAP7_75t_L g3642 ( 
.A1(n_3449),
.A2(n_3212),
.B1(n_3368),
.B2(n_3344),
.C1(n_3336),
.C2(n_3365),
.Y(n_3642)
);

OAI21x1_ASAP7_75t_L g3643 ( 
.A1(n_3415),
.A2(n_3213),
.B(n_3236),
.Y(n_3643)
);

OAI21x1_ASAP7_75t_L g3644 ( 
.A1(n_3461),
.A2(n_3314),
.B(n_3303),
.Y(n_3644)
);

OAI21x1_ASAP7_75t_L g3645 ( 
.A1(n_3419),
.A2(n_3440),
.B(n_3422),
.Y(n_3645)
);

OA21x2_ASAP7_75t_L g3646 ( 
.A1(n_3486),
.A2(n_3293),
.B(n_3285),
.Y(n_3646)
);

OAI22xp5_ASAP7_75t_SL g3647 ( 
.A1(n_3515),
.A2(n_3344),
.B1(n_3314),
.B2(n_3303),
.Y(n_3647)
);

AO31x2_ASAP7_75t_L g3648 ( 
.A1(n_3475),
.A2(n_82),
.A3(n_79),
.B(n_80),
.Y(n_3648)
);

OAI22xp33_ASAP7_75t_L g3649 ( 
.A1(n_3453),
.A2(n_3314),
.B1(n_3293),
.B2(n_3285),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3438),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_3438),
.Y(n_3651)
);

OAI22xp5_ASAP7_75t_SL g3652 ( 
.A1(n_3455),
.A2(n_3315),
.B1(n_85),
.B2(n_83),
.Y(n_3652)
);

INVx2_ASAP7_75t_SL g3653 ( 
.A(n_3488),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_L g3654 ( 
.A(n_3430),
.B(n_3315),
.Y(n_3654)
);

AOI22xp5_ASAP7_75t_L g3655 ( 
.A1(n_3510),
.A2(n_1051),
.B1(n_1053),
.B2(n_1010),
.Y(n_3655)
);

OAI22xp5_ASAP7_75t_L g3656 ( 
.A1(n_3466),
.A2(n_1051),
.B1(n_1053),
.B2(n_1010),
.Y(n_3656)
);

AND2x4_ASAP7_75t_L g3657 ( 
.A(n_3417),
.B(n_84),
.Y(n_3657)
);

AND2x2_ASAP7_75t_L g3658 ( 
.A(n_3418),
.B(n_84),
.Y(n_3658)
);

AO21x2_ASAP7_75t_L g3659 ( 
.A1(n_3467),
.A2(n_85),
.B(n_87),
.Y(n_3659)
);

BUFx10_ASAP7_75t_L g3660 ( 
.A(n_3526),
.Y(n_3660)
);

OAI21x1_ASAP7_75t_L g3661 ( 
.A1(n_3419),
.A2(n_87),
.B(n_88),
.Y(n_3661)
);

OAI21x1_ASAP7_75t_L g3662 ( 
.A1(n_3422),
.A2(n_3456),
.B(n_3440),
.Y(n_3662)
);

OAI21x1_ASAP7_75t_SL g3663 ( 
.A1(n_3473),
.A2(n_88),
.B(n_89),
.Y(n_3663)
);

OAI21x1_ASAP7_75t_L g3664 ( 
.A1(n_3456),
.A2(n_89),
.B(n_90),
.Y(n_3664)
);

INVx2_ASAP7_75t_SL g3665 ( 
.A(n_3447),
.Y(n_3665)
);

OAI21x1_ASAP7_75t_SL g3666 ( 
.A1(n_3475),
.A2(n_94),
.B(n_95),
.Y(n_3666)
);

NOR2xp33_ASAP7_75t_L g3667 ( 
.A(n_3571),
.B(n_94),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3547),
.B(n_95),
.Y(n_3668)
);

AOI21xp5_ASAP7_75t_L g3669 ( 
.A1(n_3423),
.A2(n_1053),
.B(n_1051),
.Y(n_3669)
);

OAI21xp5_ASAP7_75t_L g3670 ( 
.A1(n_3573),
.A2(n_98),
.B(n_99),
.Y(n_3670)
);

BUFx3_ASAP7_75t_L g3671 ( 
.A(n_3556),
.Y(n_3671)
);

AND2x4_ASAP7_75t_L g3672 ( 
.A(n_3417),
.B(n_98),
.Y(n_3672)
);

NOR2xp33_ASAP7_75t_L g3673 ( 
.A(n_3412),
.B(n_3513),
.Y(n_3673)
);

OAI21x1_ASAP7_75t_L g3674 ( 
.A1(n_3474),
.A2(n_100),
.B(n_101),
.Y(n_3674)
);

BUFx6f_ASAP7_75t_L g3675 ( 
.A(n_3406),
.Y(n_3675)
);

AO21x2_ASAP7_75t_L g3676 ( 
.A1(n_3489),
.A2(n_100),
.B(n_102),
.Y(n_3676)
);

INVx2_ASAP7_75t_L g3677 ( 
.A(n_3502),
.Y(n_3677)
);

INVx2_ASAP7_75t_L g3678 ( 
.A(n_3502),
.Y(n_3678)
);

OAI21x1_ASAP7_75t_L g3679 ( 
.A1(n_3474),
.A2(n_102),
.B(n_103),
.Y(n_3679)
);

CKINVDCx5p33_ASAP7_75t_R g3680 ( 
.A(n_3505),
.Y(n_3680)
);

OAI21xp5_ASAP7_75t_L g3681 ( 
.A1(n_3497),
.A2(n_103),
.B(n_105),
.Y(n_3681)
);

INVx1_ASAP7_75t_SL g3682 ( 
.A(n_3535),
.Y(n_3682)
);

OR3x4_ASAP7_75t_SL g3683 ( 
.A(n_3490),
.B(n_106),
.C(n_107),
.Y(n_3683)
);

INVx1_ASAP7_75t_L g3684 ( 
.A(n_3443),
.Y(n_3684)
);

NAND2x1p5_ASAP7_75t_L g3685 ( 
.A(n_3469),
.B(n_1051),
.Y(n_3685)
);

OAI21x1_ASAP7_75t_L g3686 ( 
.A1(n_3480),
.A2(n_107),
.B(n_108),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_3443),
.Y(n_3687)
);

AOI21x1_ASAP7_75t_L g3688 ( 
.A1(n_3511),
.A2(n_109),
.B(n_110),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_3451),
.Y(n_3689)
);

INVx2_ASAP7_75t_L g3690 ( 
.A(n_3506),
.Y(n_3690)
);

BUFx6f_ASAP7_75t_L g3691 ( 
.A(n_3406),
.Y(n_3691)
);

NAND2x1p5_ASAP7_75t_L g3692 ( 
.A(n_3469),
.B(n_1053),
.Y(n_3692)
);

INVx2_ASAP7_75t_SL g3693 ( 
.A(n_3406),
.Y(n_3693)
);

NOR2xp33_ASAP7_75t_L g3694 ( 
.A(n_3528),
.B(n_3564),
.Y(n_3694)
);

AO21x2_ASAP7_75t_L g3695 ( 
.A1(n_3451),
.A2(n_109),
.B(n_110),
.Y(n_3695)
);

INVx2_ASAP7_75t_L g3696 ( 
.A(n_3506),
.Y(n_3696)
);

OAI21x1_ASAP7_75t_L g3697 ( 
.A1(n_3480),
.A2(n_111),
.B(n_112),
.Y(n_3697)
);

AOI22xp33_ASAP7_75t_L g3698 ( 
.A1(n_3476),
.A2(n_1075),
.B1(n_1523),
.B2(n_116),
.Y(n_3698)
);

AND2x2_ASAP7_75t_L g3699 ( 
.A(n_3458),
.B(n_112),
.Y(n_3699)
);

O2A1O1Ixp33_ASAP7_75t_SL g3700 ( 
.A1(n_3527),
.A2(n_114),
.B(n_117),
.C(n_119),
.Y(n_3700)
);

OAI21x1_ASAP7_75t_L g3701 ( 
.A1(n_3487),
.A2(n_114),
.B(n_117),
.Y(n_3701)
);

OR2x2_ASAP7_75t_L g3702 ( 
.A(n_3482),
.B(n_120),
.Y(n_3702)
);

AOI22xp33_ASAP7_75t_L g3703 ( 
.A1(n_3476),
.A2(n_1075),
.B1(n_1523),
.B2(n_123),
.Y(n_3703)
);

NAND2xp5_ASAP7_75t_SL g3704 ( 
.A(n_3483),
.B(n_1075),
.Y(n_3704)
);

A2O1A1Ixp33_ASAP7_75t_L g3705 ( 
.A1(n_3503),
.A2(n_120),
.B(n_121),
.C(n_123),
.Y(n_3705)
);

OAI21x1_ASAP7_75t_L g3706 ( 
.A1(n_3498),
.A2(n_124),
.B(n_125),
.Y(n_3706)
);

INVx2_ASAP7_75t_SL g3707 ( 
.A(n_3421),
.Y(n_3707)
);

OR2x6_ASAP7_75t_L g3708 ( 
.A(n_3420),
.B(n_1075),
.Y(n_3708)
);

AND2x2_ASAP7_75t_L g3709 ( 
.A(n_3607),
.B(n_3552),
.Y(n_3709)
);

INVxp67_ASAP7_75t_SL g3710 ( 
.A(n_3590),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3650),
.Y(n_3711)
);

OAI21xp5_ASAP7_75t_L g3712 ( 
.A1(n_3602),
.A2(n_3681),
.B(n_3670),
.Y(n_3712)
);

BUFx2_ASAP7_75t_L g3713 ( 
.A(n_3616),
.Y(n_3713)
);

AOI22xp33_ASAP7_75t_L g3714 ( 
.A1(n_3667),
.A2(n_3500),
.B1(n_3483),
.B2(n_3485),
.Y(n_3714)
);

INVx1_ASAP7_75t_L g3715 ( 
.A(n_3650),
.Y(n_3715)
);

AO21x1_ASAP7_75t_SL g3716 ( 
.A1(n_3642),
.A2(n_3495),
.B(n_3555),
.Y(n_3716)
);

BUFx6f_ASAP7_75t_L g3717 ( 
.A(n_3611),
.Y(n_3717)
);

HB1xp67_ASAP7_75t_L g3718 ( 
.A(n_3583),
.Y(n_3718)
);

AOI21x1_ASAP7_75t_L g3719 ( 
.A1(n_3614),
.A2(n_3512),
.B(n_3504),
.Y(n_3719)
);

INVx2_ASAP7_75t_SL g3720 ( 
.A(n_3593),
.Y(n_3720)
);

INVx2_ASAP7_75t_L g3721 ( 
.A(n_3651),
.Y(n_3721)
);

HB1xp67_ASAP7_75t_L g3722 ( 
.A(n_3583),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_3651),
.Y(n_3723)
);

INVx1_ASAP7_75t_SL g3724 ( 
.A(n_3641),
.Y(n_3724)
);

BUFx2_ASAP7_75t_R g3725 ( 
.A(n_3680),
.Y(n_3725)
);

AO21x2_ASAP7_75t_L g3726 ( 
.A1(n_3599),
.A2(n_3550),
.B(n_3534),
.Y(n_3726)
);

BUFx6f_ASAP7_75t_L g3727 ( 
.A(n_3688),
.Y(n_3727)
);

INVx2_ASAP7_75t_L g3728 ( 
.A(n_3684),
.Y(n_3728)
);

AND2x2_ASAP7_75t_L g3729 ( 
.A(n_3616),
.B(n_3569),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_3684),
.Y(n_3730)
);

AOI22xp33_ASAP7_75t_L g3731 ( 
.A1(n_3663),
.A2(n_3526),
.B1(n_3522),
.B2(n_3525),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3687),
.Y(n_3732)
);

BUFx2_ASAP7_75t_L g3733 ( 
.A(n_3627),
.Y(n_3733)
);

INVx2_ASAP7_75t_L g3734 ( 
.A(n_3689),
.Y(n_3734)
);

INVx3_ASAP7_75t_L g3735 ( 
.A(n_3627),
.Y(n_3735)
);

AOI22xp33_ASAP7_75t_SL g3736 ( 
.A1(n_3683),
.A2(n_3490),
.B1(n_3455),
.B2(n_3568),
.Y(n_3736)
);

CKINVDCx11_ASAP7_75t_R g3737 ( 
.A(n_3621),
.Y(n_3737)
);

OAI21x1_ASAP7_75t_L g3738 ( 
.A1(n_3645),
.A2(n_3538),
.B(n_3468),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3596),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3596),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3605),
.Y(n_3741)
);

AOI22xp33_ASAP7_75t_L g3742 ( 
.A1(n_3676),
.A2(n_3548),
.B1(n_3558),
.B2(n_3539),
.Y(n_3742)
);

OAI22xp33_ASAP7_75t_L g3743 ( 
.A1(n_3580),
.A2(n_3490),
.B1(n_3559),
.B2(n_3523),
.Y(n_3743)
);

AND2x2_ASAP7_75t_L g3744 ( 
.A(n_3653),
.B(n_3560),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3605),
.Y(n_3745)
);

INVxp33_ASAP7_75t_L g3746 ( 
.A(n_3586),
.Y(n_3746)
);

OAI22xp5_ASAP7_75t_L g3747 ( 
.A1(n_3597),
.A2(n_3496),
.B1(n_3484),
.B2(n_3567),
.Y(n_3747)
);

AO21x1_ASAP7_75t_L g3748 ( 
.A1(n_3609),
.A2(n_3523),
.B(n_3543),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3606),
.Y(n_3749)
);

AOI22xp33_ASAP7_75t_L g3750 ( 
.A1(n_3659),
.A2(n_3477),
.B1(n_3452),
.B2(n_3454),
.Y(n_3750)
);

CKINVDCx11_ASAP7_75t_R g3751 ( 
.A(n_3660),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3606),
.Y(n_3752)
);

AND2x4_ASAP7_75t_L g3753 ( 
.A(n_3601),
.B(n_3543),
.Y(n_3753)
);

AND2x4_ASAP7_75t_SL g3754 ( 
.A(n_3708),
.B(n_3546),
.Y(n_3754)
);

AND2x4_ASAP7_75t_L g3755 ( 
.A(n_3601),
.B(n_3546),
.Y(n_3755)
);

AOI22xp33_ASAP7_75t_L g3756 ( 
.A1(n_3652),
.A2(n_3462),
.B1(n_3465),
.B2(n_3429),
.Y(n_3756)
);

INVx2_ASAP7_75t_L g3757 ( 
.A(n_3612),
.Y(n_3757)
);

AND2x2_ASAP7_75t_L g3758 ( 
.A(n_3619),
.B(n_3538),
.Y(n_3758)
);

INVx3_ASAP7_75t_L g3759 ( 
.A(n_3662),
.Y(n_3759)
);

AOI22xp33_ASAP7_75t_SL g3760 ( 
.A1(n_3695),
.A2(n_3421),
.B1(n_3551),
.B2(n_3478),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3612),
.Y(n_3761)
);

AND2x2_ASAP7_75t_L g3762 ( 
.A(n_3633),
.B(n_3578),
.Y(n_3762)
);

AND2x2_ASAP7_75t_L g3763 ( 
.A(n_3633),
.B(n_3563),
.Y(n_3763)
);

NAND2xp5_ASAP7_75t_L g3764 ( 
.A(n_3620),
.B(n_3555),
.Y(n_3764)
);

INVx1_ASAP7_75t_SL g3765 ( 
.A(n_3593),
.Y(n_3765)
);

AND2x2_ASAP7_75t_L g3766 ( 
.A(n_3682),
.B(n_3553),
.Y(n_3766)
);

HB1xp67_ASAP7_75t_L g3767 ( 
.A(n_3646),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3626),
.Y(n_3768)
);

INVx2_ASAP7_75t_L g3769 ( 
.A(n_3646),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_3626),
.Y(n_3770)
);

INVx4_ASAP7_75t_L g3771 ( 
.A(n_3618),
.Y(n_3771)
);

INVx2_ASAP7_75t_L g3772 ( 
.A(n_3631),
.Y(n_3772)
);

INVx2_ASAP7_75t_L g3773 ( 
.A(n_3631),
.Y(n_3773)
);

AOI22xp33_ASAP7_75t_SL g3774 ( 
.A1(n_3647),
.A2(n_3421),
.B1(n_3551),
.B2(n_3460),
.Y(n_3774)
);

BUFx6f_ASAP7_75t_L g3775 ( 
.A(n_3708),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3638),
.Y(n_3776)
);

NAND2x1p5_ASAP7_75t_L g3777 ( 
.A(n_3601),
.B(n_3551),
.Y(n_3777)
);

INVx1_ASAP7_75t_SL g3778 ( 
.A(n_3671),
.Y(n_3778)
);

INVx1_ASAP7_75t_L g3779 ( 
.A(n_3638),
.Y(n_3779)
);

OAI21xp5_ASAP7_75t_L g3780 ( 
.A1(n_3629),
.A2(n_3410),
.B(n_3408),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3640),
.Y(n_3781)
);

INVx2_ASAP7_75t_L g3782 ( 
.A(n_3640),
.Y(n_3782)
);

BUFx2_ASAP7_75t_SL g3783 ( 
.A(n_3636),
.Y(n_3783)
);

AOI22xp33_ASAP7_75t_L g3784 ( 
.A1(n_3694),
.A2(n_3517),
.B1(n_3567),
.B2(n_3561),
.Y(n_3784)
);

HB1xp67_ASAP7_75t_L g3785 ( 
.A(n_3588),
.Y(n_3785)
);

INVx2_ASAP7_75t_L g3786 ( 
.A(n_3644),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3588),
.Y(n_3787)
);

AOI21x1_ASAP7_75t_L g3788 ( 
.A1(n_3669),
.A2(n_3537),
.B(n_3524),
.Y(n_3788)
);

OAI21x1_ASAP7_75t_L g3789 ( 
.A1(n_3615),
.A2(n_3557),
.B(n_3544),
.Y(n_3789)
);

INVx2_ASAP7_75t_L g3790 ( 
.A(n_3591),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_3624),
.Y(n_3791)
);

NAND2x1p5_ASAP7_75t_L g3792 ( 
.A(n_3579),
.B(n_3533),
.Y(n_3792)
);

AO21x2_ASAP7_75t_L g3793 ( 
.A1(n_3668),
.A2(n_3570),
.B(n_3562),
.Y(n_3793)
);

BUFx3_ASAP7_75t_L g3794 ( 
.A(n_3574),
.Y(n_3794)
);

INVx2_ASAP7_75t_L g3795 ( 
.A(n_3587),
.Y(n_3795)
);

NOR2xp33_ASAP7_75t_L g3796 ( 
.A(n_3576),
.B(n_3542),
.Y(n_3796)
);

INVx1_ASAP7_75t_SL g3797 ( 
.A(n_3577),
.Y(n_3797)
);

OAI22xp5_ASAP7_75t_L g3798 ( 
.A1(n_3592),
.A2(n_3541),
.B1(n_3530),
.B2(n_3518),
.Y(n_3798)
);

INVx2_ASAP7_75t_L g3799 ( 
.A(n_3581),
.Y(n_3799)
);

BUFx4_ASAP7_75t_SL g3800 ( 
.A(n_3702),
.Y(n_3800)
);

AO21x1_ASAP7_75t_SL g3801 ( 
.A1(n_3617),
.A2(n_3478),
.B(n_3460),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3604),
.Y(n_3802)
);

INVx1_ASAP7_75t_L g3803 ( 
.A(n_3654),
.Y(n_3803)
);

INVx2_ASAP7_75t_L g3804 ( 
.A(n_3632),
.Y(n_3804)
);

OAI21x1_ASAP7_75t_L g3805 ( 
.A1(n_3600),
.A2(n_3478),
.B(n_3460),
.Y(n_3805)
);

INVx5_ASAP7_75t_L g3806 ( 
.A(n_3675),
.Y(n_3806)
);

OA21x2_ASAP7_75t_L g3807 ( 
.A1(n_3575),
.A2(n_3542),
.B(n_3530),
.Y(n_3807)
);

INVx1_ASAP7_75t_L g3808 ( 
.A(n_3677),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_3678),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3690),
.Y(n_3810)
);

INVx2_ASAP7_75t_L g3811 ( 
.A(n_3696),
.Y(n_3811)
);

INVx2_ASAP7_75t_L g3812 ( 
.A(n_3648),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3585),
.Y(n_3813)
);

INVx2_ASAP7_75t_SL g3814 ( 
.A(n_3574),
.Y(n_3814)
);

AO21x1_ASAP7_75t_L g3815 ( 
.A1(n_3673),
.A2(n_124),
.B(n_125),
.Y(n_3815)
);

INVx1_ASAP7_75t_L g3816 ( 
.A(n_3693),
.Y(n_3816)
);

OAI21x1_ASAP7_75t_L g3817 ( 
.A1(n_3603),
.A2(n_3530),
.B(n_3518),
.Y(n_3817)
);

AO21x1_ASAP7_75t_L g3818 ( 
.A1(n_3657),
.A2(n_126),
.B(n_128),
.Y(n_3818)
);

OAI21x1_ASAP7_75t_L g3819 ( 
.A1(n_3582),
.A2(n_3541),
.B(n_3518),
.Y(n_3819)
);

INVx2_ASAP7_75t_L g3820 ( 
.A(n_3648),
.Y(n_3820)
);

INVx2_ASAP7_75t_L g3821 ( 
.A(n_3675),
.Y(n_3821)
);

OA21x2_ASAP7_75t_L g3822 ( 
.A1(n_3608),
.A2(n_3542),
.B(n_3541),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3707),
.Y(n_3823)
);

BUFx12f_ASAP7_75t_L g3824 ( 
.A(n_3657),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_3648),
.Y(n_3825)
);

AOI22xp5_ASAP7_75t_L g3826 ( 
.A1(n_3649),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_3826)
);

AND2x2_ASAP7_75t_L g3827 ( 
.A(n_3665),
.B(n_130),
.Y(n_3827)
);

AOI22xp33_ASAP7_75t_L g3828 ( 
.A1(n_3666),
.A2(n_131),
.B1(n_132),
.B2(n_134),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_3675),
.Y(n_3829)
);

AOI22xp33_ASAP7_75t_L g3830 ( 
.A1(n_3613),
.A2(n_131),
.B1(n_135),
.B2(n_136),
.Y(n_3830)
);

INVx1_ASAP7_75t_L g3831 ( 
.A(n_3691),
.Y(n_3831)
);

AOI22xp33_ASAP7_75t_SL g3832 ( 
.A1(n_3623),
.A2(n_135),
.B1(n_138),
.B2(n_139),
.Y(n_3832)
);

OAI22xp5_ASAP7_75t_L g3833 ( 
.A1(n_3698),
.A2(n_138),
.B1(n_140),
.B2(n_141),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3718),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3718),
.Y(n_3835)
);

INVx1_ASAP7_75t_L g3836 ( 
.A(n_3722),
.Y(n_3836)
);

INVx1_ASAP7_75t_L g3837 ( 
.A(n_3722),
.Y(n_3837)
);

INVx2_ASAP7_75t_L g3838 ( 
.A(n_3769),
.Y(n_3838)
);

INVx3_ASAP7_75t_L g3839 ( 
.A(n_3777),
.Y(n_3839)
);

OA21x2_ASAP7_75t_L g3840 ( 
.A1(n_3789),
.A2(n_3701),
.B(n_3664),
.Y(n_3840)
);

INVx1_ASAP7_75t_L g3841 ( 
.A(n_3739),
.Y(n_3841)
);

AND2x2_ASAP7_75t_L g3842 ( 
.A(n_3735),
.B(n_3746),
.Y(n_3842)
);

INVx2_ASAP7_75t_L g3843 ( 
.A(n_3769),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3740),
.Y(n_3844)
);

OR2x6_ASAP7_75t_L g3845 ( 
.A(n_3777),
.B(n_3634),
.Y(n_3845)
);

INVx3_ASAP7_75t_L g3846 ( 
.A(n_3792),
.Y(n_3846)
);

AOI22xp5_ASAP7_75t_L g3847 ( 
.A1(n_3743),
.A2(n_3672),
.B1(n_3655),
.B2(n_3704),
.Y(n_3847)
);

OA21x2_ASAP7_75t_L g3848 ( 
.A1(n_3805),
.A2(n_3674),
.B(n_3661),
.Y(n_3848)
);

AND2x2_ASAP7_75t_L g3849 ( 
.A(n_3735),
.B(n_3586),
.Y(n_3849)
);

NOR2x1p5_ASAP7_75t_L g3850 ( 
.A(n_3794),
.B(n_3672),
.Y(n_3850)
);

INVx1_ASAP7_75t_L g3851 ( 
.A(n_3741),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_L g3852 ( 
.A(n_3797),
.B(n_3699),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_3745),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3772),
.Y(n_3854)
);

INVx1_ASAP7_75t_L g3855 ( 
.A(n_3749),
.Y(n_3855)
);

INVx6_ASAP7_75t_L g3856 ( 
.A(n_3806),
.Y(n_3856)
);

AND2x2_ASAP7_75t_L g3857 ( 
.A(n_3746),
.B(n_3610),
.Y(n_3857)
);

BUFx3_ASAP7_75t_L g3858 ( 
.A(n_3737),
.Y(n_3858)
);

INVx2_ASAP7_75t_L g3859 ( 
.A(n_3728),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_3752),
.Y(n_3860)
);

OAI21x1_ASAP7_75t_L g3861 ( 
.A1(n_3792),
.A2(n_3738),
.B(n_3759),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_3761),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3772),
.Y(n_3863)
);

AND2x2_ASAP7_75t_L g3864 ( 
.A(n_3713),
.B(n_3625),
.Y(n_3864)
);

INVx1_ASAP7_75t_L g3865 ( 
.A(n_3773),
.Y(n_3865)
);

AND2x2_ASAP7_75t_L g3866 ( 
.A(n_3733),
.B(n_3639),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3773),
.Y(n_3867)
);

NAND2x1p5_ASAP7_75t_L g3868 ( 
.A(n_3807),
.B(n_3579),
.Y(n_3868)
);

INVx1_ASAP7_75t_L g3869 ( 
.A(n_3782),
.Y(n_3869)
);

INVx2_ASAP7_75t_L g3870 ( 
.A(n_3782),
.Y(n_3870)
);

INVx2_ASAP7_75t_L g3871 ( 
.A(n_3767),
.Y(n_3871)
);

INVx2_ASAP7_75t_L g3872 ( 
.A(n_3767),
.Y(n_3872)
);

INVx2_ASAP7_75t_L g3873 ( 
.A(n_3721),
.Y(n_3873)
);

BUFx6f_ASAP7_75t_L g3874 ( 
.A(n_3794),
.Y(n_3874)
);

AO21x2_ASAP7_75t_L g3875 ( 
.A1(n_3812),
.A2(n_3700),
.B(n_3686),
.Y(n_3875)
);

NOR2x1_ASAP7_75t_R g3876 ( 
.A(n_3737),
.B(n_3658),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3711),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3715),
.Y(n_3878)
);

BUFx6f_ASAP7_75t_L g3879 ( 
.A(n_3806),
.Y(n_3879)
);

OAI21x1_ASAP7_75t_L g3880 ( 
.A1(n_3759),
.A2(n_3622),
.B(n_3589),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3768),
.Y(n_3881)
);

OAI22xp5_ASAP7_75t_L g3882 ( 
.A1(n_3736),
.A2(n_3630),
.B1(n_3703),
.B2(n_3628),
.Y(n_3882)
);

INVx2_ASAP7_75t_L g3883 ( 
.A(n_3734),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_3770),
.Y(n_3884)
);

INVx2_ASAP7_75t_L g3885 ( 
.A(n_3757),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3776),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3779),
.Y(n_3887)
);

HB1xp67_ASAP7_75t_L g3888 ( 
.A(n_3812),
.Y(n_3888)
);

AND2x4_ASAP7_75t_L g3889 ( 
.A(n_3753),
.B(n_3635),
.Y(n_3889)
);

AO21x2_ASAP7_75t_L g3890 ( 
.A1(n_3820),
.A2(n_3697),
.B(n_3679),
.Y(n_3890)
);

INVx3_ASAP7_75t_L g3891 ( 
.A(n_3753),
.Y(n_3891)
);

INVx3_ASAP7_75t_L g3892 ( 
.A(n_3755),
.Y(n_3892)
);

INVx2_ASAP7_75t_L g3893 ( 
.A(n_3790),
.Y(n_3893)
);

AOI22xp33_ASAP7_75t_L g3894 ( 
.A1(n_3712),
.A2(n_3643),
.B1(n_3594),
.B2(n_3660),
.Y(n_3894)
);

INVx1_ASAP7_75t_L g3895 ( 
.A(n_3781),
.Y(n_3895)
);

INVx2_ASAP7_75t_L g3896 ( 
.A(n_3790),
.Y(n_3896)
);

HB1xp67_ASAP7_75t_L g3897 ( 
.A(n_3820),
.Y(n_3897)
);

INVx1_ASAP7_75t_L g3898 ( 
.A(n_3723),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_3730),
.Y(n_3899)
);

INVx2_ASAP7_75t_L g3900 ( 
.A(n_3732),
.Y(n_3900)
);

INVx3_ASAP7_75t_L g3901 ( 
.A(n_3755),
.Y(n_3901)
);

INVx3_ASAP7_75t_L g3902 ( 
.A(n_3822),
.Y(n_3902)
);

INVx2_ASAP7_75t_L g3903 ( 
.A(n_3811),
.Y(n_3903)
);

INVx1_ASAP7_75t_L g3904 ( 
.A(n_3785),
.Y(n_3904)
);

BUFx2_ASAP7_75t_L g3905 ( 
.A(n_3793),
.Y(n_3905)
);

INVx1_ASAP7_75t_L g3906 ( 
.A(n_3785),
.Y(n_3906)
);

INVx1_ASAP7_75t_L g3907 ( 
.A(n_3787),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3764),
.Y(n_3908)
);

INVx3_ASAP7_75t_L g3909 ( 
.A(n_3822),
.Y(n_3909)
);

AO21x2_ASAP7_75t_L g3910 ( 
.A1(n_3743),
.A2(n_3706),
.B(n_3705),
.Y(n_3910)
);

AND2x2_ASAP7_75t_L g3911 ( 
.A(n_3729),
.B(n_3691),
.Y(n_3911)
);

INVx1_ASAP7_75t_L g3912 ( 
.A(n_3799),
.Y(n_3912)
);

INVx2_ASAP7_75t_L g3913 ( 
.A(n_3811),
.Y(n_3913)
);

INVx3_ASAP7_75t_L g3914 ( 
.A(n_3822),
.Y(n_3914)
);

INVx2_ASAP7_75t_SL g3915 ( 
.A(n_3806),
.Y(n_3915)
);

INVx2_ASAP7_75t_L g3916 ( 
.A(n_3793),
.Y(n_3916)
);

BUFx3_ASAP7_75t_L g3917 ( 
.A(n_3717),
.Y(n_3917)
);

INVx2_ASAP7_75t_L g3918 ( 
.A(n_3799),
.Y(n_3918)
);

OAI22xp5_ASAP7_75t_L g3919 ( 
.A1(n_3736),
.A2(n_3630),
.B1(n_3598),
.B2(n_3685),
.Y(n_3919)
);

INVx2_ASAP7_75t_L g3920 ( 
.A(n_3795),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_3791),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_3825),
.Y(n_3922)
);

INVx2_ASAP7_75t_L g3923 ( 
.A(n_3795),
.Y(n_3923)
);

INVx3_ASAP7_75t_L g3924 ( 
.A(n_3807),
.Y(n_3924)
);

OR2x2_ASAP7_75t_L g3925 ( 
.A(n_3710),
.B(n_3594),
.Y(n_3925)
);

INVx2_ASAP7_75t_L g3926 ( 
.A(n_3758),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3710),
.Y(n_3927)
);

AND2x4_ASAP7_75t_L g3928 ( 
.A(n_3817),
.B(n_3691),
.Y(n_3928)
);

AND2x2_ASAP7_75t_L g3929 ( 
.A(n_3801),
.B(n_3595),
.Y(n_3929)
);

BUFx2_ASAP7_75t_SL g3930 ( 
.A(n_3806),
.Y(n_3930)
);

BUFx2_ASAP7_75t_L g3931 ( 
.A(n_3726),
.Y(n_3931)
);

INVx2_ASAP7_75t_SL g3932 ( 
.A(n_3717),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_3802),
.Y(n_3933)
);

BUFx2_ASAP7_75t_L g3934 ( 
.A(n_3726),
.Y(n_3934)
);

BUFx3_ASAP7_75t_L g3935 ( 
.A(n_3717),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3803),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3829),
.Y(n_3937)
);

INVx1_ASAP7_75t_L g3938 ( 
.A(n_3831),
.Y(n_3938)
);

INVx5_ASAP7_75t_L g3939 ( 
.A(n_3727),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3808),
.Y(n_3940)
);

HB1xp67_ASAP7_75t_L g3941 ( 
.A(n_3800),
.Y(n_3941)
);

AO21x2_ASAP7_75t_L g3942 ( 
.A1(n_3815),
.A2(n_3584),
.B(n_3637),
.Y(n_3942)
);

AND2x2_ASAP7_75t_L g3943 ( 
.A(n_3813),
.B(n_3762),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3809),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3810),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3804),
.Y(n_3946)
);

BUFx3_ASAP7_75t_L g3947 ( 
.A(n_3717),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3804),
.Y(n_3948)
);

INVx1_ASAP7_75t_L g3949 ( 
.A(n_3807),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3786),
.Y(n_3950)
);

BUFx3_ASAP7_75t_L g3951 ( 
.A(n_3751),
.Y(n_3951)
);

INVx1_ASAP7_75t_L g3952 ( 
.A(n_3922),
.Y(n_3952)
);

AOI22xp33_ASAP7_75t_L g3953 ( 
.A1(n_3910),
.A2(n_3716),
.B1(n_3727),
.B2(n_3830),
.Y(n_3953)
);

NAND3xp33_ASAP7_75t_L g3954 ( 
.A(n_3939),
.B(n_3830),
.C(n_3828),
.Y(n_3954)
);

A2O1A1Ixp33_ASAP7_75t_L g3955 ( 
.A1(n_3919),
.A2(n_3796),
.B(n_3724),
.C(n_3826),
.Y(n_3955)
);

AOI222xp33_ASAP7_75t_L g3956 ( 
.A1(n_3882),
.A2(n_3833),
.B1(n_3828),
.B2(n_3747),
.C1(n_3756),
.C2(n_3742),
.Y(n_3956)
);

OAI22xp5_ASAP7_75t_L g3957 ( 
.A1(n_3847),
.A2(n_3774),
.B1(n_3760),
.B2(n_3756),
.Y(n_3957)
);

OAI22xp5_ASAP7_75t_L g3958 ( 
.A1(n_3894),
.A2(n_3774),
.B1(n_3760),
.B2(n_3714),
.Y(n_3958)
);

INVx1_ASAP7_75t_L g3959 ( 
.A(n_3877),
.Y(n_3959)
);

AOI21x1_ASAP7_75t_L g3960 ( 
.A1(n_3931),
.A2(n_3934),
.B(n_3941),
.Y(n_3960)
);

OAI211xp5_ASAP7_75t_L g3961 ( 
.A1(n_3931),
.A2(n_3832),
.B(n_3731),
.C(n_3742),
.Y(n_3961)
);

AOI221xp5_ASAP7_75t_L g3962 ( 
.A1(n_3934),
.A2(n_3780),
.B1(n_3750),
.B2(n_3818),
.C(n_3727),
.Y(n_3962)
);

NAND2xp5_ASAP7_75t_L g3963 ( 
.A(n_3937),
.B(n_3938),
.Y(n_3963)
);

OAI22xp5_ASAP7_75t_L g3964 ( 
.A1(n_3845),
.A2(n_3714),
.B1(n_3727),
.B2(n_3796),
.Y(n_3964)
);

BUFx12f_ASAP7_75t_L g3965 ( 
.A(n_3858),
.Y(n_3965)
);

AND2x2_ASAP7_75t_L g3966 ( 
.A(n_3911),
.B(n_3783),
.Y(n_3966)
);

AOI22xp33_ASAP7_75t_L g3967 ( 
.A1(n_3910),
.A2(n_3832),
.B1(n_3824),
.B2(n_3751),
.Y(n_3967)
);

AND2x4_ASAP7_75t_L g3968 ( 
.A(n_3951),
.B(n_3814),
.Y(n_3968)
);

AOI22xp33_ASAP7_75t_L g3969 ( 
.A1(n_3910),
.A2(n_3775),
.B1(n_3784),
.B2(n_3748),
.Y(n_3969)
);

NAND3xp33_ASAP7_75t_L g3970 ( 
.A(n_3939),
.B(n_3750),
.C(n_3731),
.Y(n_3970)
);

OR2x2_ASAP7_75t_L g3971 ( 
.A(n_3908),
.B(n_3821),
.Y(n_3971)
);

INVx1_ASAP7_75t_L g3972 ( 
.A(n_3877),
.Y(n_3972)
);

OAI22xp5_ASAP7_75t_L g3973 ( 
.A1(n_3845),
.A2(n_3784),
.B1(n_3765),
.B2(n_3720),
.Y(n_3973)
);

OAI211xp5_ASAP7_75t_L g3974 ( 
.A1(n_3939),
.A2(n_3719),
.B(n_3827),
.C(n_3775),
.Y(n_3974)
);

AOI22xp33_ASAP7_75t_L g3975 ( 
.A1(n_3889),
.A2(n_3845),
.B1(n_3874),
.B2(n_3942),
.Y(n_3975)
);

AOI22xp33_ASAP7_75t_L g3976 ( 
.A1(n_3889),
.A2(n_3775),
.B1(n_3766),
.B2(n_3778),
.Y(n_3976)
);

AND2x2_ASAP7_75t_L g3977 ( 
.A(n_3911),
.B(n_3763),
.Y(n_3977)
);

OAI22xp5_ASAP7_75t_L g3978 ( 
.A1(n_3845),
.A2(n_3775),
.B1(n_3754),
.B2(n_3798),
.Y(n_3978)
);

OAI21xp5_ASAP7_75t_L g3979 ( 
.A1(n_3939),
.A2(n_3819),
.B(n_3788),
.Y(n_3979)
);

OAI222xp33_ASAP7_75t_L g3980 ( 
.A1(n_3939),
.A2(n_3823),
.B1(n_3816),
.B2(n_3744),
.C1(n_3800),
.C2(n_3709),
.Y(n_3980)
);

AOI22xp33_ASAP7_75t_L g3981 ( 
.A1(n_3889),
.A2(n_3771),
.B1(n_3754),
.B2(n_3692),
.Y(n_3981)
);

AO21x1_ASAP7_75t_SL g3982 ( 
.A1(n_3927),
.A2(n_3725),
.B(n_3771),
.Y(n_3982)
);

OA21x2_ASAP7_75t_L g3983 ( 
.A1(n_3861),
.A2(n_3656),
.B(n_140),
.Y(n_3983)
);

INVx1_ASAP7_75t_L g3984 ( 
.A(n_3878),
.Y(n_3984)
);

OAI22xp5_ASAP7_75t_L g3985 ( 
.A1(n_3951),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_3985)
);

AOI222xp33_ASAP7_75t_L g3986 ( 
.A1(n_3876),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.C1(n_146),
.C2(n_147),
.Y(n_3986)
);

AOI22xp33_ASAP7_75t_L g3987 ( 
.A1(n_3874),
.A2(n_3942),
.B1(n_3858),
.B2(n_3943),
.Y(n_3987)
);

OAI211xp5_ASAP7_75t_L g3988 ( 
.A1(n_3905),
.A2(n_3925),
.B(n_3842),
.C(n_3846),
.Y(n_3988)
);

OAI21x1_ASAP7_75t_L g3989 ( 
.A1(n_3861),
.A2(n_147),
.B(n_148),
.Y(n_3989)
);

AOI22xp33_ASAP7_75t_L g3990 ( 
.A1(n_3874),
.A2(n_149),
.B1(n_151),
.B2(n_152),
.Y(n_3990)
);

AND2x2_ASAP7_75t_L g3991 ( 
.A(n_3929),
.B(n_149),
.Y(n_3991)
);

AOI22xp33_ASAP7_75t_L g3992 ( 
.A1(n_3874),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_3992)
);

HB1xp67_ASAP7_75t_L g3993 ( 
.A(n_3875),
.Y(n_3993)
);

AOI222xp33_ASAP7_75t_L g3994 ( 
.A1(n_3874),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.C1(n_157),
.C2(n_159),
.Y(n_3994)
);

INVx2_ASAP7_75t_L g3995 ( 
.A(n_3891),
.Y(n_3995)
);

AND2x2_ASAP7_75t_L g3996 ( 
.A(n_3929),
.B(n_156),
.Y(n_3996)
);

AOI22xp33_ASAP7_75t_L g3997 ( 
.A1(n_3942),
.A2(n_3943),
.B1(n_3926),
.B2(n_3864),
.Y(n_3997)
);

INVxp33_ASAP7_75t_L g3998 ( 
.A(n_3866),
.Y(n_3998)
);

AOI221xp5_ASAP7_75t_L g3999 ( 
.A1(n_3933),
.A2(n_3905),
.B1(n_3912),
.B2(n_3936),
.C(n_3918),
.Y(n_3999)
);

AOI22xp33_ASAP7_75t_SL g4000 ( 
.A1(n_3930),
.A2(n_159),
.B1(n_162),
.B2(n_163),
.Y(n_4000)
);

AOI22xp33_ASAP7_75t_L g4001 ( 
.A1(n_3926),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_4001)
);

AOI22xp33_ASAP7_75t_L g4002 ( 
.A1(n_3864),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_4002)
);

AOI22xp33_ASAP7_75t_SL g4003 ( 
.A1(n_3930),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_4003)
);

OAI22xp5_ASAP7_75t_L g4004 ( 
.A1(n_3850),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_4004)
);

AOI22xp33_ASAP7_75t_L g4005 ( 
.A1(n_3857),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_4005)
);

AND2x6_ASAP7_75t_L g4006 ( 
.A(n_3917),
.B(n_172),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3878),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_3841),
.Y(n_4008)
);

INVx1_ASAP7_75t_L g4009 ( 
.A(n_3844),
.Y(n_4009)
);

AND2x4_ASAP7_75t_L g4010 ( 
.A(n_3891),
.B(n_172),
.Y(n_4010)
);

OAI211xp5_ASAP7_75t_L g4011 ( 
.A1(n_3925),
.A2(n_173),
.B(n_174),
.C(n_175),
.Y(n_4011)
);

A2O1A1Ixp33_ASAP7_75t_L g4012 ( 
.A1(n_3846),
.A2(n_173),
.B(n_174),
.C(n_175),
.Y(n_4012)
);

BUFx4f_ASAP7_75t_SL g4013 ( 
.A(n_3917),
.Y(n_4013)
);

AOI221xp5_ASAP7_75t_L g4014 ( 
.A1(n_3918),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.C(n_180),
.Y(n_4014)
);

OR2x6_ASAP7_75t_L g4015 ( 
.A(n_3856),
.B(n_178),
.Y(n_4015)
);

OAI22xp5_ASAP7_75t_L g4016 ( 
.A1(n_3932),
.A2(n_180),
.B1(n_181),
.B2(n_183),
.Y(n_4016)
);

OAI221xp5_ASAP7_75t_L g4017 ( 
.A1(n_3891),
.A2(n_181),
.B1(n_183),
.B2(n_185),
.C(n_188),
.Y(n_4017)
);

OAI221xp5_ASAP7_75t_SL g4018 ( 
.A1(n_3842),
.A2(n_185),
.B1(n_189),
.B2(n_190),
.C(n_191),
.Y(n_4018)
);

AOI22xp33_ASAP7_75t_L g4019 ( 
.A1(n_3857),
.A2(n_189),
.B1(n_190),
.B2(n_192),
.Y(n_4019)
);

A2O1A1Ixp33_ASAP7_75t_L g4020 ( 
.A1(n_3846),
.A2(n_192),
.B(n_193),
.C(n_195),
.Y(n_4020)
);

AOI22xp33_ASAP7_75t_L g4021 ( 
.A1(n_3892),
.A2(n_3901),
.B1(n_3866),
.B2(n_3875),
.Y(n_4021)
);

AOI22xp33_ASAP7_75t_L g4022 ( 
.A1(n_3892),
.A2(n_193),
.B1(n_197),
.B2(n_198),
.Y(n_4022)
);

AOI22xp33_ASAP7_75t_L g4023 ( 
.A1(n_3892),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_4023)
);

NAND3xp33_ASAP7_75t_L g4024 ( 
.A(n_3904),
.B(n_200),
.C(n_202),
.Y(n_4024)
);

INVx2_ASAP7_75t_L g4025 ( 
.A(n_3901),
.Y(n_4025)
);

AOI22xp33_ASAP7_75t_L g4026 ( 
.A1(n_3901),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_4026)
);

AOI21xp5_ASAP7_75t_L g4027 ( 
.A1(n_3875),
.A2(n_205),
.B(n_206),
.Y(n_4027)
);

AOI22xp33_ASAP7_75t_L g4028 ( 
.A1(n_3856),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_4028)
);

INVx2_ASAP7_75t_L g4029 ( 
.A(n_3879),
.Y(n_4029)
);

OAI22xp5_ASAP7_75t_L g4030 ( 
.A1(n_3932),
.A2(n_208),
.B1(n_210),
.B2(n_211),
.Y(n_4030)
);

AND2x4_ASAP7_75t_SL g4031 ( 
.A(n_3849),
.B(n_210),
.Y(n_4031)
);

AOI211xp5_ASAP7_75t_L g4032 ( 
.A1(n_3879),
.A2(n_211),
.B(n_212),
.C(n_213),
.Y(n_4032)
);

AOI22xp33_ASAP7_75t_L g4033 ( 
.A1(n_3856),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_4033)
);

AOI22xp33_ASAP7_75t_L g4034 ( 
.A1(n_3856),
.A2(n_214),
.B1(n_216),
.B2(n_217),
.Y(n_4034)
);

INVx2_ASAP7_75t_L g4035 ( 
.A(n_3879),
.Y(n_4035)
);

NOR3xp33_ASAP7_75t_L g4036 ( 
.A(n_3915),
.B(n_218),
.C(n_219),
.Y(n_4036)
);

AND2x2_ASAP7_75t_L g4037 ( 
.A(n_3935),
.B(n_3947),
.Y(n_4037)
);

INVxp67_ASAP7_75t_SL g4038 ( 
.A(n_3935),
.Y(n_4038)
);

AND2x4_ASAP7_75t_L g4039 ( 
.A(n_3947),
.B(n_3915),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_L g4040 ( 
.A(n_3852),
.B(n_218),
.Y(n_4040)
);

AND2x2_ASAP7_75t_L g4041 ( 
.A(n_3849),
.B(n_219),
.Y(n_4041)
);

INVxp67_ASAP7_75t_L g4042 ( 
.A(n_3890),
.Y(n_4042)
);

NAND4xp25_ASAP7_75t_L g4043 ( 
.A(n_3906),
.B(n_220),
.C(n_223),
.D(n_225),
.Y(n_4043)
);

OAI221xp5_ASAP7_75t_L g4044 ( 
.A1(n_3839),
.A2(n_223),
.B1(n_226),
.B2(n_229),
.C(n_265),
.Y(n_4044)
);

AO31x2_ASAP7_75t_L g4045 ( 
.A1(n_3871),
.A2(n_267),
.A3(n_269),
.B(n_272),
.Y(n_4045)
);

AOI22xp33_ASAP7_75t_L g4046 ( 
.A1(n_3879),
.A2(n_274),
.B1(n_276),
.B2(n_279),
.Y(n_4046)
);

INVx1_ASAP7_75t_L g4047 ( 
.A(n_3851),
.Y(n_4047)
);

AOI221xp5_ASAP7_75t_L g4048 ( 
.A1(n_3950),
.A2(n_280),
.B1(n_290),
.B2(n_294),
.C(n_300),
.Y(n_4048)
);

AOI21xp5_ASAP7_75t_L g4049 ( 
.A1(n_3840),
.A2(n_302),
.B(n_303),
.Y(n_4049)
);

BUFx3_ASAP7_75t_L g4050 ( 
.A(n_3879),
.Y(n_4050)
);

INVxp33_ASAP7_75t_L g4051 ( 
.A(n_3840),
.Y(n_4051)
);

OAI22xp5_ASAP7_75t_L g4052 ( 
.A1(n_3839),
.A2(n_305),
.B1(n_307),
.B2(n_309),
.Y(n_4052)
);

OAI221xp5_ASAP7_75t_SL g4053 ( 
.A1(n_3916),
.A2(n_3872),
.B1(n_3871),
.B2(n_3839),
.C(n_3949),
.Y(n_4053)
);

AOI22xp33_ASAP7_75t_L g4054 ( 
.A1(n_3840),
.A2(n_310),
.B1(n_314),
.B2(n_316),
.Y(n_4054)
);

INVx1_ASAP7_75t_L g4055 ( 
.A(n_3853),
.Y(n_4055)
);

OAI22xp5_ASAP7_75t_L g4056 ( 
.A1(n_3868),
.A2(n_318),
.B1(n_320),
.B2(n_322),
.Y(n_4056)
);

OAI22xp5_ASAP7_75t_L g4057 ( 
.A1(n_3868),
.A2(n_324),
.B1(n_327),
.B2(n_329),
.Y(n_4057)
);

NOR2xp33_ASAP7_75t_L g4058 ( 
.A(n_3940),
.B(n_330),
.Y(n_4058)
);

NAND2x1p5_ASAP7_75t_L g4059 ( 
.A(n_3928),
.B(n_333),
.Y(n_4059)
);

OAI211xp5_ASAP7_75t_SL g4060 ( 
.A1(n_3946),
.A2(n_336),
.B(n_338),
.C(n_340),
.Y(n_4060)
);

NAND3xp33_ASAP7_75t_L g4061 ( 
.A(n_3872),
.B(n_341),
.C(n_344),
.Y(n_4061)
);

AOI21xp5_ASAP7_75t_L g4062 ( 
.A1(n_3890),
.A2(n_3848),
.B(n_3928),
.Y(n_4062)
);

NAND2xp5_ASAP7_75t_L g4063 ( 
.A(n_3907),
.B(n_472),
.Y(n_4063)
);

AOI22xp33_ASAP7_75t_SL g4064 ( 
.A1(n_3848),
.A2(n_345),
.B1(n_346),
.B2(n_347),
.Y(n_4064)
);

AOI22xp33_ASAP7_75t_L g4065 ( 
.A1(n_3890),
.A2(n_350),
.B1(n_351),
.B2(n_353),
.Y(n_4065)
);

NOR2xp33_ASAP7_75t_SL g4066 ( 
.A(n_3928),
.B(n_3868),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_3921),
.B(n_3944),
.Y(n_4067)
);

INVx2_ASAP7_75t_L g4068 ( 
.A(n_3838),
.Y(n_4068)
);

OAI22xp5_ASAP7_75t_L g4069 ( 
.A1(n_3848),
.A2(n_354),
.B1(n_356),
.B2(n_358),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_3855),
.Y(n_4070)
);

AND2x2_ASAP7_75t_L g4071 ( 
.A(n_3982),
.B(n_3920),
.Y(n_4071)
);

BUFx3_ASAP7_75t_L g4072 ( 
.A(n_3965),
.Y(n_4072)
);

BUFx3_ASAP7_75t_L g4073 ( 
.A(n_4006),
.Y(n_4073)
);

INVx2_ASAP7_75t_L g4074 ( 
.A(n_4039),
.Y(n_4074)
);

INVx1_ASAP7_75t_L g4075 ( 
.A(n_3959),
.Y(n_4075)
);

BUFx2_ASAP7_75t_L g4076 ( 
.A(n_4039),
.Y(n_4076)
);

INVx2_ASAP7_75t_L g4077 ( 
.A(n_4050),
.Y(n_4077)
);

INVx2_ASAP7_75t_L g4078 ( 
.A(n_4015),
.Y(n_4078)
);

AND2x2_ASAP7_75t_L g4079 ( 
.A(n_3966),
.B(n_3920),
.Y(n_4079)
);

AND2x4_ASAP7_75t_L g4080 ( 
.A(n_3995),
.B(n_3834),
.Y(n_4080)
);

AND2x2_ASAP7_75t_L g4081 ( 
.A(n_4037),
.B(n_3923),
.Y(n_4081)
);

INVx1_ASAP7_75t_L g4082 ( 
.A(n_3972),
.Y(n_4082)
);

AND2x2_ASAP7_75t_L g4083 ( 
.A(n_4038),
.B(n_3923),
.Y(n_4083)
);

BUFx2_ASAP7_75t_L g4084 ( 
.A(n_4013),
.Y(n_4084)
);

AND2x2_ASAP7_75t_L g4085 ( 
.A(n_3998),
.B(n_3885),
.Y(n_4085)
);

INVx2_ASAP7_75t_L g4086 ( 
.A(n_4015),
.Y(n_4086)
);

INVx2_ASAP7_75t_L g4087 ( 
.A(n_4015),
.Y(n_4087)
);

INVx1_ASAP7_75t_L g4088 ( 
.A(n_3984),
.Y(n_4088)
);

AND2x4_ASAP7_75t_L g4089 ( 
.A(n_4025),
.B(n_3835),
.Y(n_4089)
);

AND2x2_ASAP7_75t_L g4090 ( 
.A(n_3977),
.B(n_3885),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_4007),
.Y(n_4091)
);

INVx1_ASAP7_75t_L g4092 ( 
.A(n_4067),
.Y(n_4092)
);

HB1xp67_ASAP7_75t_L g4093 ( 
.A(n_3960),
.Y(n_4093)
);

HB1xp67_ASAP7_75t_L g4094 ( 
.A(n_3993),
.Y(n_4094)
);

INVx1_ASAP7_75t_L g4095 ( 
.A(n_3952),
.Y(n_4095)
);

AND2x2_ASAP7_75t_L g4096 ( 
.A(n_3968),
.B(n_3903),
.Y(n_4096)
);

HB1xp67_ASAP7_75t_L g4097 ( 
.A(n_4041),
.Y(n_4097)
);

INVx1_ASAP7_75t_L g4098 ( 
.A(n_4008),
.Y(n_4098)
);

NAND2xp5_ASAP7_75t_L g4099 ( 
.A(n_3991),
.B(n_3921),
.Y(n_4099)
);

INVx4_ASAP7_75t_SL g4100 ( 
.A(n_4006),
.Y(n_4100)
);

AND2x4_ASAP7_75t_L g4101 ( 
.A(n_4029),
.B(n_3836),
.Y(n_4101)
);

BUFx2_ASAP7_75t_SL g4102 ( 
.A(n_4006),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_4009),
.Y(n_4103)
);

BUFx4f_ASAP7_75t_SL g4104 ( 
.A(n_3968),
.Y(n_4104)
);

BUFx3_ASAP7_75t_L g4105 ( 
.A(n_4006),
.Y(n_4105)
);

BUFx2_ASAP7_75t_L g4106 ( 
.A(n_4035),
.Y(n_4106)
);

HB1xp67_ASAP7_75t_L g4107 ( 
.A(n_4010),
.Y(n_4107)
);

INVx2_ASAP7_75t_L g4108 ( 
.A(n_3989),
.Y(n_4108)
);

BUFx2_ASAP7_75t_L g4109 ( 
.A(n_3979),
.Y(n_4109)
);

INVx1_ASAP7_75t_L g4110 ( 
.A(n_4047),
.Y(n_4110)
);

INVx1_ASAP7_75t_L g4111 ( 
.A(n_4055),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_4070),
.Y(n_4112)
);

INVx1_ASAP7_75t_L g4113 ( 
.A(n_4068),
.Y(n_4113)
);

AND2x2_ASAP7_75t_L g4114 ( 
.A(n_3976),
.B(n_3903),
.Y(n_4114)
);

INVx1_ASAP7_75t_L g4115 ( 
.A(n_3963),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_3971),
.Y(n_4116)
);

BUFx12f_ASAP7_75t_L g4117 ( 
.A(n_4010),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_3996),
.Y(n_4118)
);

BUFx6f_ASAP7_75t_L g4119 ( 
.A(n_4061),
.Y(n_4119)
);

BUFx3_ASAP7_75t_L g4120 ( 
.A(n_4031),
.Y(n_4120)
);

NAND2xp5_ASAP7_75t_L g4121 ( 
.A(n_3956),
.B(n_3860),
.Y(n_4121)
);

AND2x4_ASAP7_75t_L g4122 ( 
.A(n_3970),
.B(n_3837),
.Y(n_4122)
);

AND2x2_ASAP7_75t_L g4123 ( 
.A(n_3975),
.B(n_3913),
.Y(n_4123)
);

HB1xp67_ASAP7_75t_L g4124 ( 
.A(n_3970),
.Y(n_4124)
);

INVx2_ASAP7_75t_L g4125 ( 
.A(n_3983),
.Y(n_4125)
);

HB1xp67_ASAP7_75t_L g4126 ( 
.A(n_3988),
.Y(n_4126)
);

AND2x2_ASAP7_75t_L g4127 ( 
.A(n_3987),
.B(n_3913),
.Y(n_4127)
);

INVx2_ASAP7_75t_L g4128 ( 
.A(n_3983),
.Y(n_4128)
);

CKINVDCx11_ASAP7_75t_R g4129 ( 
.A(n_4004),
.Y(n_4129)
);

HB1xp67_ASAP7_75t_L g4130 ( 
.A(n_4042),
.Y(n_4130)
);

AOI22xp33_ASAP7_75t_L g4131 ( 
.A1(n_3967),
.A2(n_3958),
.B1(n_3953),
.B2(n_3954),
.Y(n_4131)
);

BUFx2_ASAP7_75t_L g4132 ( 
.A(n_3962),
.Y(n_4132)
);

INVxp67_ASAP7_75t_SL g4133 ( 
.A(n_4066),
.Y(n_4133)
);

AND2x4_ASAP7_75t_L g4134 ( 
.A(n_3954),
.B(n_3900),
.Y(n_4134)
);

BUFx3_ASAP7_75t_L g4135 ( 
.A(n_4059),
.Y(n_4135)
);

AND2x4_ASAP7_75t_L g4136 ( 
.A(n_4027),
.B(n_3900),
.Y(n_4136)
);

INVxp67_ASAP7_75t_SL g4137 ( 
.A(n_3978),
.Y(n_4137)
);

AND2x2_ASAP7_75t_L g4138 ( 
.A(n_3969),
.B(n_3873),
.Y(n_4138)
);

INVx1_ASAP7_75t_L g4139 ( 
.A(n_4063),
.Y(n_4139)
);

INVx1_ASAP7_75t_L g4140 ( 
.A(n_4040),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_4011),
.Y(n_4141)
);

INVx1_ASAP7_75t_L g4142 ( 
.A(n_4024),
.Y(n_4142)
);

BUFx2_ASAP7_75t_L g4143 ( 
.A(n_3957),
.Y(n_4143)
);

BUFx3_ASAP7_75t_L g4144 ( 
.A(n_4058),
.Y(n_4144)
);

AND2x4_ASAP7_75t_L g4145 ( 
.A(n_3981),
.B(n_3916),
.Y(n_4145)
);

AND2x2_ASAP7_75t_L g4146 ( 
.A(n_3997),
.B(n_3873),
.Y(n_4146)
);

AND2x2_ASAP7_75t_L g4147 ( 
.A(n_4021),
.B(n_3883),
.Y(n_4147)
);

INVx1_ASAP7_75t_L g4148 ( 
.A(n_3961),
.Y(n_4148)
);

NAND2xp5_ASAP7_75t_L g4149 ( 
.A(n_3955),
.B(n_3986),
.Y(n_4149)
);

INVx2_ASAP7_75t_L g4150 ( 
.A(n_4045),
.Y(n_4150)
);

AND2x2_ASAP7_75t_L g4151 ( 
.A(n_3974),
.B(n_3883),
.Y(n_4151)
);

AND2x4_ASAP7_75t_L g4152 ( 
.A(n_4036),
.B(n_3893),
.Y(n_4152)
);

INVx3_ASAP7_75t_L g4153 ( 
.A(n_4045),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_4051),
.Y(n_4154)
);

INVx2_ASAP7_75t_L g4155 ( 
.A(n_4045),
.Y(n_4155)
);

BUFx3_ASAP7_75t_L g4156 ( 
.A(n_4017),
.Y(n_4156)
);

BUFx6f_ASAP7_75t_L g4157 ( 
.A(n_4061),
.Y(n_4157)
);

INVx2_ASAP7_75t_L g4158 ( 
.A(n_3973),
.Y(n_4158)
);

OR2x2_ASAP7_75t_L g4159 ( 
.A(n_4053),
.B(n_3944),
.Y(n_4159)
);

INVxp67_ASAP7_75t_L g4160 ( 
.A(n_3964),
.Y(n_4160)
);

AND2x2_ASAP7_75t_L g4161 ( 
.A(n_3999),
.B(n_3893),
.Y(n_4161)
);

INVx3_ASAP7_75t_L g4162 ( 
.A(n_3980),
.Y(n_4162)
);

AND2x4_ASAP7_75t_L g4163 ( 
.A(n_4062),
.B(n_3896),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_4076),
.Y(n_4164)
);

NAND2xp33_ASAP7_75t_R g4165 ( 
.A(n_4132),
.B(n_4143),
.Y(n_4165)
);

AND2x2_ASAP7_75t_L g4166 ( 
.A(n_4084),
.B(n_3945),
.Y(n_4166)
);

INVx2_ASAP7_75t_L g4167 ( 
.A(n_4076),
.Y(n_4167)
);

OR2x2_ASAP7_75t_L g4168 ( 
.A(n_4118),
.B(n_4043),
.Y(n_4168)
);

OR2x2_ASAP7_75t_L g4169 ( 
.A(n_4118),
.B(n_4012),
.Y(n_4169)
);

BUFx2_ASAP7_75t_L g4170 ( 
.A(n_4117),
.Y(n_4170)
);

AND2x4_ASAP7_75t_L g4171 ( 
.A(n_4100),
.B(n_3902),
.Y(n_4171)
);

AND2x2_ASAP7_75t_L g4172 ( 
.A(n_4084),
.B(n_3945),
.Y(n_4172)
);

AND2x2_ASAP7_75t_L g4173 ( 
.A(n_4072),
.B(n_3862),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_4106),
.Y(n_4174)
);

OR2x2_ASAP7_75t_L g4175 ( 
.A(n_4097),
.B(n_4020),
.Y(n_4175)
);

INVxp67_ASAP7_75t_SL g4176 ( 
.A(n_4119),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_4106),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_4094),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_4075),
.Y(n_4179)
);

AND2x2_ASAP7_75t_L g4180 ( 
.A(n_4072),
.B(n_4120),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_4075),
.Y(n_4181)
);

OAI22xp5_ASAP7_75t_L g4182 ( 
.A1(n_4162),
.A2(n_4018),
.B1(n_4032),
.B2(n_4000),
.Y(n_4182)
);

BUFx2_ASAP7_75t_L g4183 ( 
.A(n_4117),
.Y(n_4183)
);

INVx1_ASAP7_75t_L g4184 ( 
.A(n_4082),
.Y(n_4184)
);

INVx2_ASAP7_75t_L g4185 ( 
.A(n_4100),
.Y(n_4185)
);

BUFx2_ASAP7_75t_L g4186 ( 
.A(n_4104),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_4082),
.Y(n_4187)
);

NAND2xp5_ASAP7_75t_L g4188 ( 
.A(n_4107),
.B(n_4032),
.Y(n_4188)
);

INVx1_ASAP7_75t_SL g4189 ( 
.A(n_4102),
.Y(n_4189)
);

AND2x2_ASAP7_75t_SL g4190 ( 
.A(n_4132),
.B(n_4014),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_L g4191 ( 
.A(n_4141),
.B(n_3994),
.Y(n_4191)
);

NAND2xp5_ASAP7_75t_L g4192 ( 
.A(n_4141),
.B(n_4126),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_4088),
.Y(n_4193)
);

AND2x2_ASAP7_75t_L g4194 ( 
.A(n_4120),
.B(n_3881),
.Y(n_4194)
);

HB1xp67_ASAP7_75t_L g4195 ( 
.A(n_4093),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_4088),
.Y(n_4196)
);

INVx1_ASAP7_75t_L g4197 ( 
.A(n_4091),
.Y(n_4197)
);

AOI22x1_ASAP7_75t_L g4198 ( 
.A1(n_4124),
.A2(n_4049),
.B1(n_3909),
.B2(n_3902),
.Y(n_4198)
);

INVx1_ASAP7_75t_L g4199 ( 
.A(n_4091),
.Y(n_4199)
);

AND2x2_ASAP7_75t_L g4200 ( 
.A(n_4079),
.B(n_3884),
.Y(n_4200)
);

AND2x2_ASAP7_75t_L g4201 ( 
.A(n_4079),
.B(n_3886),
.Y(n_4201)
);

NAND2xp5_ASAP7_75t_L g4202 ( 
.A(n_4078),
.B(n_4003),
.Y(n_4202)
);

INVx2_ASAP7_75t_L g4203 ( 
.A(n_4100),
.Y(n_4203)
);

NAND2xp5_ASAP7_75t_L g4204 ( 
.A(n_4078),
.B(n_3985),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_4083),
.Y(n_4205)
);

NAND2x1p5_ASAP7_75t_L g4206 ( 
.A(n_4119),
.B(n_3902),
.Y(n_4206)
);

OR2x2_ASAP7_75t_L g4207 ( 
.A(n_4086),
.B(n_4016),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_L g4208 ( 
.A(n_4086),
.B(n_4002),
.Y(n_4208)
);

AND2x4_ASAP7_75t_L g4209 ( 
.A(n_4100),
.B(n_3909),
.Y(n_4209)
);

AND2x4_ASAP7_75t_L g4210 ( 
.A(n_4074),
.B(n_4073),
.Y(n_4210)
);

NAND2xp5_ASAP7_75t_L g4211 ( 
.A(n_4087),
.B(n_4143),
.Y(n_4211)
);

AOI22xp33_ASAP7_75t_L g4212 ( 
.A1(n_4162),
.A2(n_4149),
.B1(n_4131),
.B2(n_4119),
.Y(n_4212)
);

INVx2_ASAP7_75t_SL g4213 ( 
.A(n_4074),
.Y(n_4213)
);

INVx2_ASAP7_75t_L g4214 ( 
.A(n_4119),
.Y(n_4214)
);

INVxp67_ASAP7_75t_SL g4215 ( 
.A(n_4119),
.Y(n_4215)
);

INVx1_ASAP7_75t_L g4216 ( 
.A(n_4083),
.Y(n_4216)
);

AND2x4_ASAP7_75t_L g4217 ( 
.A(n_4073),
.B(n_3909),
.Y(n_4217)
);

NAND2xp5_ASAP7_75t_L g4218 ( 
.A(n_4210),
.B(n_4087),
.Y(n_4218)
);

HB1xp67_ASAP7_75t_L g4219 ( 
.A(n_4167),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_L g4220 ( 
.A(n_4210),
.B(n_4077),
.Y(n_4220)
);

AND2x4_ASAP7_75t_L g4221 ( 
.A(n_4167),
.B(n_4105),
.Y(n_4221)
);

AND2x2_ASAP7_75t_L g4222 ( 
.A(n_4180),
.B(n_4102),
.Y(n_4222)
);

BUFx3_ASAP7_75t_L g4223 ( 
.A(n_4170),
.Y(n_4223)
);

AO21x2_ASAP7_75t_L g4224 ( 
.A1(n_4176),
.A2(n_4148),
.B(n_4154),
.Y(n_4224)
);

INVx2_ASAP7_75t_L g4225 ( 
.A(n_4206),
.Y(n_4225)
);

HB1xp67_ASAP7_75t_L g4226 ( 
.A(n_4206),
.Y(n_4226)
);

OR2x2_ASAP7_75t_L g4227 ( 
.A(n_4176),
.B(n_4148),
.Y(n_4227)
);

NAND2xp5_ASAP7_75t_L g4228 ( 
.A(n_4210),
.B(n_4077),
.Y(n_4228)
);

BUFx2_ASAP7_75t_SL g4229 ( 
.A(n_4215),
.Y(n_4229)
);

AOI22xp33_ASAP7_75t_L g4230 ( 
.A1(n_4190),
.A2(n_4162),
.B1(n_4157),
.B2(n_4158),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_4195),
.Y(n_4231)
);

INVx3_ASAP7_75t_L g4232 ( 
.A(n_4171),
.Y(n_4232)
);

INVxp67_ASAP7_75t_SL g4233 ( 
.A(n_4165),
.Y(n_4233)
);

OR2x2_ASAP7_75t_L g4234 ( 
.A(n_4215),
.B(n_4125),
.Y(n_4234)
);

INVx1_ASAP7_75t_L g4235 ( 
.A(n_4195),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_4174),
.Y(n_4236)
);

AND2x2_ASAP7_75t_L g4237 ( 
.A(n_4186),
.B(n_4071),
.Y(n_4237)
);

INVx2_ASAP7_75t_L g4238 ( 
.A(n_4171),
.Y(n_4238)
);

AND2x2_ASAP7_75t_L g4239 ( 
.A(n_4183),
.B(n_4071),
.Y(n_4239)
);

INVx5_ASAP7_75t_SL g4240 ( 
.A(n_4171),
.Y(n_4240)
);

AND2x2_ASAP7_75t_L g4241 ( 
.A(n_4189),
.B(n_4096),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_4177),
.Y(n_4242)
);

AO21x2_ASAP7_75t_L g4243 ( 
.A1(n_4214),
.A2(n_4154),
.B(n_4128),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_L g4244 ( 
.A(n_4182),
.B(n_4156),
.Y(n_4244)
);

AND2x2_ASAP7_75t_L g4245 ( 
.A(n_4164),
.B(n_4096),
.Y(n_4245)
);

INVx2_ASAP7_75t_L g4246 ( 
.A(n_4198),
.Y(n_4246)
);

INVx2_ASAP7_75t_SL g4247 ( 
.A(n_4209),
.Y(n_4247)
);

AND2x2_ASAP7_75t_L g4248 ( 
.A(n_4166),
.B(n_4105),
.Y(n_4248)
);

BUFx2_ASAP7_75t_L g4249 ( 
.A(n_4209),
.Y(n_4249)
);

NAND2xp5_ASAP7_75t_L g4250 ( 
.A(n_4212),
.B(n_4156),
.Y(n_4250)
);

INVx1_ASAP7_75t_L g4251 ( 
.A(n_4213),
.Y(n_4251)
);

OR2x2_ASAP7_75t_L g4252 ( 
.A(n_4192),
.B(n_4125),
.Y(n_4252)
);

AND2x2_ASAP7_75t_L g4253 ( 
.A(n_4172),
.B(n_4081),
.Y(n_4253)
);

INVx2_ASAP7_75t_L g4254 ( 
.A(n_4214),
.Y(n_4254)
);

HB1xp67_ASAP7_75t_L g4255 ( 
.A(n_4213),
.Y(n_4255)
);

AND2x2_ASAP7_75t_L g4256 ( 
.A(n_4205),
.B(n_4081),
.Y(n_4256)
);

OR2x2_ASAP7_75t_L g4257 ( 
.A(n_4211),
.B(n_4128),
.Y(n_4257)
);

INVx1_ASAP7_75t_L g4258 ( 
.A(n_4216),
.Y(n_4258)
);

INVx2_ASAP7_75t_L g4259 ( 
.A(n_4190),
.Y(n_4259)
);

AND2x2_ASAP7_75t_L g4260 ( 
.A(n_4194),
.B(n_4151),
.Y(n_4260)
);

INVx1_ASAP7_75t_L g4261 ( 
.A(n_4178),
.Y(n_4261)
);

INVx3_ASAP7_75t_L g4262 ( 
.A(n_4209),
.Y(n_4262)
);

INVxp67_ASAP7_75t_L g4263 ( 
.A(n_4165),
.Y(n_4263)
);

HB1xp67_ASAP7_75t_L g4264 ( 
.A(n_4217),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_4179),
.Y(n_4265)
);

INVx1_ASAP7_75t_L g4266 ( 
.A(n_4181),
.Y(n_4266)
);

NAND2xp5_ASAP7_75t_L g4267 ( 
.A(n_4212),
.B(n_4137),
.Y(n_4267)
);

INVx2_ASAP7_75t_L g4268 ( 
.A(n_4217),
.Y(n_4268)
);

HB1xp67_ASAP7_75t_L g4269 ( 
.A(n_4217),
.Y(n_4269)
);

AND2x2_ASAP7_75t_L g4270 ( 
.A(n_4237),
.B(n_4185),
.Y(n_4270)
);

AND2x2_ASAP7_75t_L g4271 ( 
.A(n_4237),
.B(n_4185),
.Y(n_4271)
);

AND2x2_ASAP7_75t_L g4272 ( 
.A(n_4239),
.B(n_4222),
.Y(n_4272)
);

INVx2_ASAP7_75t_L g4273 ( 
.A(n_4243),
.Y(n_4273)
);

INVx2_ASAP7_75t_L g4274 ( 
.A(n_4243),
.Y(n_4274)
);

OR2x2_ASAP7_75t_L g4275 ( 
.A(n_4233),
.B(n_4188),
.Y(n_4275)
);

AND2x2_ASAP7_75t_L g4276 ( 
.A(n_4239),
.B(n_4203),
.Y(n_4276)
);

OR2x2_ASAP7_75t_L g4277 ( 
.A(n_4224),
.B(n_4191),
.Y(n_4277)
);

INVxp67_ASAP7_75t_L g4278 ( 
.A(n_4229),
.Y(n_4278)
);

INVx2_ASAP7_75t_L g4279 ( 
.A(n_4243),
.Y(n_4279)
);

INVx2_ASAP7_75t_L g4280 ( 
.A(n_4224),
.Y(n_4280)
);

AND2x4_ASAP7_75t_L g4281 ( 
.A(n_4249),
.B(n_4203),
.Y(n_4281)
);

AND2x2_ASAP7_75t_L g4282 ( 
.A(n_4222),
.B(n_4173),
.Y(n_4282)
);

OR2x2_ASAP7_75t_L g4283 ( 
.A(n_4224),
.B(n_4168),
.Y(n_4283)
);

HB1xp67_ASAP7_75t_L g4284 ( 
.A(n_4249),
.Y(n_4284)
);

INVx2_ASAP7_75t_L g4285 ( 
.A(n_4259),
.Y(n_4285)
);

AND2x2_ASAP7_75t_L g4286 ( 
.A(n_4241),
.B(n_4134),
.Y(n_4286)
);

AND2x2_ASAP7_75t_L g4287 ( 
.A(n_4241),
.B(n_4134),
.Y(n_4287)
);

INVx5_ASAP7_75t_L g4288 ( 
.A(n_4232),
.Y(n_4288)
);

OR2x2_ASAP7_75t_L g4289 ( 
.A(n_4259),
.B(n_4159),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_4229),
.Y(n_4290)
);

OR2x2_ASAP7_75t_L g4291 ( 
.A(n_4259),
.B(n_4263),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_4255),
.Y(n_4292)
);

NAND2xp5_ASAP7_75t_L g4293 ( 
.A(n_4221),
.B(n_4142),
.Y(n_4293)
);

INVx2_ASAP7_75t_L g4294 ( 
.A(n_4232),
.Y(n_4294)
);

AND2x2_ASAP7_75t_L g4295 ( 
.A(n_4260),
.B(n_4253),
.Y(n_4295)
);

INVx2_ASAP7_75t_L g4296 ( 
.A(n_4232),
.Y(n_4296)
);

AND2x2_ASAP7_75t_L g4297 ( 
.A(n_4260),
.B(n_4134),
.Y(n_4297)
);

NAND2xp5_ASAP7_75t_L g4298 ( 
.A(n_4221),
.B(n_4142),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_4219),
.Y(n_4299)
);

INVx2_ASAP7_75t_SL g4300 ( 
.A(n_4232),
.Y(n_4300)
);

NAND2xp5_ASAP7_75t_L g4301 ( 
.A(n_4221),
.B(n_4160),
.Y(n_4301)
);

AND2x4_ASAP7_75t_L g4302 ( 
.A(n_4262),
.B(n_4122),
.Y(n_4302)
);

AND2x2_ASAP7_75t_L g4303 ( 
.A(n_4253),
.B(n_4114),
.Y(n_4303)
);

AND2x2_ASAP7_75t_L g4304 ( 
.A(n_4248),
.B(n_4223),
.Y(n_4304)
);

AND2x2_ASAP7_75t_L g4305 ( 
.A(n_4248),
.B(n_4114),
.Y(n_4305)
);

AND2x2_ASAP7_75t_L g4306 ( 
.A(n_4223),
.B(n_4200),
.Y(n_4306)
);

OR2x2_ASAP7_75t_L g4307 ( 
.A(n_4227),
.B(n_4159),
.Y(n_4307)
);

HB1xp67_ASAP7_75t_L g4308 ( 
.A(n_4262),
.Y(n_4308)
);

AND2x2_ASAP7_75t_L g4309 ( 
.A(n_4272),
.B(n_4223),
.Y(n_4309)
);

NAND2xp5_ASAP7_75t_L g4310 ( 
.A(n_4272),
.B(n_4304),
.Y(n_4310)
);

NOR2xp33_ASAP7_75t_L g4311 ( 
.A(n_4277),
.B(n_4218),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_4308),
.Y(n_4312)
);

AND2x2_ASAP7_75t_L g4313 ( 
.A(n_4305),
.B(n_4245),
.Y(n_4313)
);

INVx1_ASAP7_75t_L g4314 ( 
.A(n_4284),
.Y(n_4314)
);

NAND2xp5_ASAP7_75t_L g4315 ( 
.A(n_4304),
.B(n_4221),
.Y(n_4315)
);

AND2x2_ASAP7_75t_L g4316 ( 
.A(n_4270),
.B(n_4245),
.Y(n_4316)
);

AND2x2_ASAP7_75t_L g4317 ( 
.A(n_4270),
.B(n_4256),
.Y(n_4317)
);

AND2x2_ASAP7_75t_SL g4318 ( 
.A(n_4277),
.B(n_4250),
.Y(n_4318)
);

NAND2xp5_ASAP7_75t_L g4319 ( 
.A(n_4271),
.B(n_4230),
.Y(n_4319)
);

NOR2xp33_ASAP7_75t_L g4320 ( 
.A(n_4283),
.B(n_4267),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_4294),
.Y(n_4321)
);

AND2x2_ASAP7_75t_SL g4322 ( 
.A(n_4283),
.B(n_4244),
.Y(n_4322)
);

OR2x2_ASAP7_75t_L g4323 ( 
.A(n_4307),
.B(n_4227),
.Y(n_4323)
);

BUFx2_ASAP7_75t_L g4324 ( 
.A(n_4302),
.Y(n_4324)
);

HB1xp67_ASAP7_75t_L g4325 ( 
.A(n_4280),
.Y(n_4325)
);

AND2x2_ASAP7_75t_L g4326 ( 
.A(n_4305),
.B(n_4256),
.Y(n_4326)
);

OR2x2_ASAP7_75t_L g4327 ( 
.A(n_4307),
.B(n_4202),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_4294),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_4294),
.Y(n_4329)
);

NOR2x1_ASAP7_75t_L g4330 ( 
.A(n_4280),
.B(n_4262),
.Y(n_4330)
);

INVx2_ASAP7_75t_L g4331 ( 
.A(n_4280),
.Y(n_4331)
);

NAND2xp5_ASAP7_75t_L g4332 ( 
.A(n_4271),
.B(n_4264),
.Y(n_4332)
);

NAND2xp5_ASAP7_75t_L g4333 ( 
.A(n_4276),
.B(n_4269),
.Y(n_4333)
);

AND2x2_ASAP7_75t_L g4334 ( 
.A(n_4295),
.B(n_4240),
.Y(n_4334)
);

INVx1_ASAP7_75t_L g4335 ( 
.A(n_4324),
.Y(n_4335)
);

AND2x4_ASAP7_75t_L g4336 ( 
.A(n_4309),
.B(n_4281),
.Y(n_4336)
);

AND3x2_ASAP7_75t_L g4337 ( 
.A(n_4320),
.B(n_4279),
.C(n_4273),
.Y(n_4337)
);

AND2x2_ASAP7_75t_L g4338 ( 
.A(n_4313),
.B(n_4295),
.Y(n_4338)
);

INVx2_ASAP7_75t_SL g4339 ( 
.A(n_4309),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_SL g4340 ( 
.A(n_4318),
.B(n_4157),
.Y(n_4340)
);

AND2x2_ASAP7_75t_L g4341 ( 
.A(n_4326),
.B(n_4282),
.Y(n_4341)
);

AND2x2_ASAP7_75t_L g4342 ( 
.A(n_4316),
.B(n_4282),
.Y(n_4342)
);

OR2x2_ASAP7_75t_L g4343 ( 
.A(n_4310),
.B(n_4289),
.Y(n_4343)
);

INVx6_ASAP7_75t_L g4344 ( 
.A(n_4334),
.Y(n_4344)
);

AND2x2_ASAP7_75t_L g4345 ( 
.A(n_4316),
.B(n_4303),
.Y(n_4345)
);

AND2x2_ASAP7_75t_L g4346 ( 
.A(n_4317),
.B(n_4303),
.Y(n_4346)
);

AOI22xp5_ASAP7_75t_L g4347 ( 
.A1(n_4322),
.A2(n_4157),
.B1(n_4246),
.B2(n_4286),
.Y(n_4347)
);

OR2x2_ASAP7_75t_L g4348 ( 
.A(n_4323),
.B(n_4289),
.Y(n_4348)
);

OR2x2_ASAP7_75t_L g4349 ( 
.A(n_4332),
.B(n_4275),
.Y(n_4349)
);

INVx2_ASAP7_75t_L g4350 ( 
.A(n_4317),
.Y(n_4350)
);

AND2x2_ASAP7_75t_L g4351 ( 
.A(n_4314),
.B(n_4286),
.Y(n_4351)
);

AND2x2_ASAP7_75t_L g4352 ( 
.A(n_4333),
.B(n_4287),
.Y(n_4352)
);

NAND2xp5_ASAP7_75t_L g4353 ( 
.A(n_4318),
.B(n_4300),
.Y(n_4353)
);

AND2x2_ASAP7_75t_L g4354 ( 
.A(n_4315),
.B(n_4287),
.Y(n_4354)
);

NAND2xp67_ASAP7_75t_SL g4355 ( 
.A(n_4345),
.B(n_4276),
.Y(n_4355)
);

OAI322xp33_ASAP7_75t_L g4356 ( 
.A1(n_4340),
.A2(n_4320),
.A3(n_4275),
.B1(n_4252),
.B2(n_4246),
.C1(n_4322),
.C2(n_4311),
.Y(n_4356)
);

INVx1_ASAP7_75t_L g4357 ( 
.A(n_4336),
.Y(n_4357)
);

INVx3_ASAP7_75t_L g4358 ( 
.A(n_4336),
.Y(n_4358)
);

INVx2_ASAP7_75t_L g4359 ( 
.A(n_4348),
.Y(n_4359)
);

INVx2_ASAP7_75t_L g4360 ( 
.A(n_4344),
.Y(n_4360)
);

OR2x2_ASAP7_75t_L g4361 ( 
.A(n_4339),
.B(n_4293),
.Y(n_4361)
);

AND2x4_ASAP7_75t_L g4362 ( 
.A(n_4342),
.B(n_4306),
.Y(n_4362)
);

INVx2_ASAP7_75t_L g4363 ( 
.A(n_4344),
.Y(n_4363)
);

INVx1_ASAP7_75t_L g4364 ( 
.A(n_4353),
.Y(n_4364)
);

NAND2x1_ASAP7_75t_L g4365 ( 
.A(n_4346),
.B(n_4302),
.Y(n_4365)
);

INVx3_ASAP7_75t_L g4366 ( 
.A(n_4344),
.Y(n_4366)
);

INVx1_ASAP7_75t_L g4367 ( 
.A(n_4353),
.Y(n_4367)
);

NAND2xp5_ASAP7_75t_L g4368 ( 
.A(n_4338),
.B(n_4297),
.Y(n_4368)
);

AOI22xp33_ASAP7_75t_L g4369 ( 
.A1(n_4340),
.A2(n_4109),
.B1(n_4158),
.B2(n_4122),
.Y(n_4369)
);

OAI22xp33_ASAP7_75t_SL g4370 ( 
.A1(n_4335),
.A2(n_4246),
.B1(n_4234),
.B2(n_4278),
.Y(n_4370)
);

AOI22xp5_ASAP7_75t_L g4371 ( 
.A1(n_4341),
.A2(n_4157),
.B1(n_4122),
.B2(n_4354),
.Y(n_4371)
);

HB1xp67_ASAP7_75t_L g4372 ( 
.A(n_4365),
.Y(n_4372)
);

AND2x2_ASAP7_75t_L g4373 ( 
.A(n_4362),
.B(n_4351),
.Y(n_4373)
);

AND2x2_ASAP7_75t_L g4374 ( 
.A(n_4362),
.B(n_4352),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_4358),
.Y(n_4375)
);

NAND2xp5_ASAP7_75t_L g4376 ( 
.A(n_4358),
.B(n_4337),
.Y(n_4376)
);

AND2x2_ASAP7_75t_L g4377 ( 
.A(n_4366),
.B(n_4306),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_4365),
.Y(n_4378)
);

NAND2x1p5_ASAP7_75t_L g4379 ( 
.A(n_4360),
.B(n_4288),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_4368),
.Y(n_4380)
);

NAND2xp5_ASAP7_75t_L g4381 ( 
.A(n_4357),
.B(n_4337),
.Y(n_4381)
);

AND2x2_ASAP7_75t_L g4382 ( 
.A(n_4359),
.B(n_4350),
.Y(n_4382)
);

BUFx2_ASAP7_75t_L g4383 ( 
.A(n_4355),
.Y(n_4383)
);

INVx1_ASAP7_75t_SL g4384 ( 
.A(n_4373),
.Y(n_4384)
);

AOI22xp33_ASAP7_75t_L g4385 ( 
.A1(n_4374),
.A2(n_4109),
.B1(n_4157),
.B2(n_4363),
.Y(n_4385)
);

INVxp67_ASAP7_75t_L g4386 ( 
.A(n_4372),
.Y(n_4386)
);

INVx1_ASAP7_75t_SL g4387 ( 
.A(n_4377),
.Y(n_4387)
);

OR2x2_ASAP7_75t_L g4388 ( 
.A(n_4375),
.B(n_4327),
.Y(n_4388)
);

AOI22xp33_ASAP7_75t_L g4389 ( 
.A1(n_4382),
.A2(n_4133),
.B1(n_4297),
.B2(n_4302),
.Y(n_4389)
);

INVx1_ASAP7_75t_SL g4390 ( 
.A(n_4376),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_4378),
.Y(n_4391)
);

OAI22xp5_ASAP7_75t_L g4392 ( 
.A1(n_4389),
.A2(n_4369),
.B1(n_4371),
.B2(n_4347),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_4388),
.Y(n_4393)
);

OR2x2_ASAP7_75t_L g4394 ( 
.A(n_4384),
.B(n_4220),
.Y(n_4394)
);

OAI221xp5_ASAP7_75t_L g4395 ( 
.A1(n_4385),
.A2(n_4347),
.B1(n_4319),
.B2(n_4298),
.C(n_4290),
.Y(n_4395)
);

AND2x2_ASAP7_75t_L g4396 ( 
.A(n_4387),
.B(n_4281),
.Y(n_4396)
);

INVxp67_ASAP7_75t_L g4397 ( 
.A(n_4391),
.Y(n_4397)
);

NAND2xp5_ASAP7_75t_L g4398 ( 
.A(n_4386),
.B(n_4281),
.Y(n_4398)
);

O2A1O1Ixp33_ASAP7_75t_L g4399 ( 
.A1(n_4390),
.A2(n_4356),
.B(n_4370),
.C(n_4311),
.Y(n_4399)
);

OAI221xp5_ASAP7_75t_L g4400 ( 
.A1(n_4389),
.A2(n_4290),
.B1(n_4301),
.B2(n_4291),
.C(n_4257),
.Y(n_4400)
);

AOI21xp5_ASAP7_75t_SL g4401 ( 
.A1(n_4388),
.A2(n_4349),
.B(n_4376),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_4388),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_4388),
.Y(n_4403)
);

AOI21xp5_ASAP7_75t_L g4404 ( 
.A1(n_4384),
.A2(n_4381),
.B(n_4343),
.Y(n_4404)
);

AOI22xp5_ASAP7_75t_L g4405 ( 
.A1(n_4396),
.A2(n_4247),
.B1(n_4302),
.B2(n_4228),
.Y(n_4405)
);

INVxp67_ASAP7_75t_L g4406 ( 
.A(n_4398),
.Y(n_4406)
);

OAI21xp5_ASAP7_75t_L g4407 ( 
.A1(n_4404),
.A2(n_4291),
.B(n_4299),
.Y(n_4407)
);

AOI31xp33_ASAP7_75t_L g4408 ( 
.A1(n_4394),
.A2(n_4361),
.A3(n_4379),
.B(n_4381),
.Y(n_4408)
);

NAND2xp5_ASAP7_75t_L g4409 ( 
.A(n_4393),
.B(n_4281),
.Y(n_4409)
);

AOI21xp33_ASAP7_75t_L g4410 ( 
.A1(n_4399),
.A2(n_4367),
.B(n_4364),
.Y(n_4410)
);

AOI22xp33_ASAP7_75t_SL g4411 ( 
.A1(n_4400),
.A2(n_4240),
.B1(n_4247),
.B2(n_4262),
.Y(n_4411)
);

NAND2xp5_ASAP7_75t_L g4412 ( 
.A(n_4402),
.B(n_4299),
.Y(n_4412)
);

NOR2x1_ASAP7_75t_L g4413 ( 
.A(n_4401),
.B(n_4330),
.Y(n_4413)
);

AOI22xp33_ASAP7_75t_L g4414 ( 
.A1(n_4403),
.A2(n_4292),
.B1(n_4238),
.B2(n_4268),
.Y(n_4414)
);

AOI21xp33_ASAP7_75t_SL g4415 ( 
.A1(n_4395),
.A2(n_4312),
.B(n_4285),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_4392),
.Y(n_4416)
);

AOI22xp5_ASAP7_75t_L g4417 ( 
.A1(n_4397),
.A2(n_4292),
.B1(n_4251),
.B2(n_4380),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_4396),
.Y(n_4418)
);

INVx1_ASAP7_75t_L g4419 ( 
.A(n_4396),
.Y(n_4419)
);

OAI22xp5_ASAP7_75t_L g4420 ( 
.A1(n_4400),
.A2(n_4240),
.B1(n_4257),
.B2(n_4252),
.Y(n_4420)
);

NAND2xp5_ASAP7_75t_L g4421 ( 
.A(n_4396),
.B(n_4285),
.Y(n_4421)
);

AOI21xp5_ASAP7_75t_L g4422 ( 
.A1(n_4401),
.A2(n_4383),
.B(n_4279),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_4396),
.Y(n_4423)
);

OAI31xp33_ASAP7_75t_L g4424 ( 
.A1(n_4400),
.A2(n_4231),
.A3(n_4235),
.B(n_4234),
.Y(n_4424)
);

OAI211xp5_ASAP7_75t_L g4425 ( 
.A1(n_4399),
.A2(n_4285),
.B(n_4288),
.C(n_4328),
.Y(n_4425)
);

NAND2x1_ASAP7_75t_L g4426 ( 
.A(n_4401),
.B(n_4300),
.Y(n_4426)
);

NAND2xp5_ASAP7_75t_L g4427 ( 
.A(n_4405),
.B(n_4236),
.Y(n_4427)
);

NAND2xp5_ASAP7_75t_L g4428 ( 
.A(n_4411),
.B(n_4236),
.Y(n_4428)
);

AOI21xp33_ASAP7_75t_L g4429 ( 
.A1(n_4426),
.A2(n_4329),
.B(n_4321),
.Y(n_4429)
);

NAND2xp5_ASAP7_75t_L g4430 ( 
.A(n_4414),
.B(n_4242),
.Y(n_4430)
);

NOR2xp33_ASAP7_75t_L g4431 ( 
.A(n_4409),
.B(n_4261),
.Y(n_4431)
);

INVx1_ASAP7_75t_SL g4432 ( 
.A(n_4413),
.Y(n_4432)
);

HB1xp67_ASAP7_75t_L g4433 ( 
.A(n_4407),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_L g4434 ( 
.A(n_4424),
.B(n_4242),
.Y(n_4434)
);

AOI221x1_ASAP7_75t_SL g4435 ( 
.A1(n_4420),
.A2(n_4235),
.B1(n_4231),
.B2(n_4296),
.C(n_4331),
.Y(n_4435)
);

NOR2x1_ASAP7_75t_L g4436 ( 
.A(n_4421),
.B(n_4331),
.Y(n_4436)
);

INVxp67_ASAP7_75t_L g4437 ( 
.A(n_4412),
.Y(n_4437)
);

NAND2xp5_ASAP7_75t_L g4438 ( 
.A(n_4415),
.B(n_4261),
.Y(n_4438)
);

NAND2xp5_ASAP7_75t_L g4439 ( 
.A(n_4418),
.B(n_4258),
.Y(n_4439)
);

OAI22xp5_ASAP7_75t_L g4440 ( 
.A1(n_4417),
.A2(n_4240),
.B1(n_4251),
.B2(n_4238),
.Y(n_4440)
);

INVx1_ASAP7_75t_L g4441 ( 
.A(n_4419),
.Y(n_4441)
);

INVx1_ASAP7_75t_L g4442 ( 
.A(n_4423),
.Y(n_4442)
);

INVxp67_ASAP7_75t_L g4443 ( 
.A(n_4408),
.Y(n_4443)
);

INVx1_ASAP7_75t_SL g4444 ( 
.A(n_4422),
.Y(n_4444)
);

AND2x2_ASAP7_75t_L g4445 ( 
.A(n_4416),
.B(n_4296),
.Y(n_4445)
);

NAND2xp33_ASAP7_75t_L g4446 ( 
.A(n_4425),
.B(n_4288),
.Y(n_4446)
);

NAND2xp5_ASAP7_75t_L g4447 ( 
.A(n_4406),
.B(n_4258),
.Y(n_4447)
);

AND2x2_ASAP7_75t_SL g4448 ( 
.A(n_4410),
.B(n_4325),
.Y(n_4448)
);

INVx1_ASAP7_75t_L g4449 ( 
.A(n_4413),
.Y(n_4449)
);

NAND2xp5_ASAP7_75t_L g4450 ( 
.A(n_4405),
.B(n_4288),
.Y(n_4450)
);

NAND2xp33_ASAP7_75t_SL g4451 ( 
.A(n_4426),
.B(n_4254),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_L g4452 ( 
.A(n_4405),
.B(n_4288),
.Y(n_4452)
);

OAI21xp5_ASAP7_75t_L g4453 ( 
.A1(n_4443),
.A2(n_4288),
.B(n_4254),
.Y(n_4453)
);

AND2x2_ASAP7_75t_L g4454 ( 
.A(n_4445),
.B(n_4441),
.Y(n_4454)
);

INVx1_ASAP7_75t_L g4455 ( 
.A(n_4440),
.Y(n_4455)
);

INVx1_ASAP7_75t_L g4456 ( 
.A(n_4436),
.Y(n_4456)
);

AO21x2_ASAP7_75t_L g4457 ( 
.A1(n_4449),
.A2(n_4325),
.B(n_4279),
.Y(n_4457)
);

XOR2xp5_ASAP7_75t_L g4458 ( 
.A(n_4433),
.B(n_4254),
.Y(n_4458)
);

INVx1_ASAP7_75t_L g4459 ( 
.A(n_4430),
.Y(n_4459)
);

INVx1_ASAP7_75t_L g4460 ( 
.A(n_4451),
.Y(n_4460)
);

INVx1_ASAP7_75t_L g4461 ( 
.A(n_4450),
.Y(n_4461)
);

NOR4xp25_ASAP7_75t_SL g4462 ( 
.A(n_4429),
.B(n_4442),
.C(n_4435),
.D(n_4266),
.Y(n_4462)
);

INVx1_ASAP7_75t_L g4463 ( 
.A(n_4452),
.Y(n_4463)
);

INVx1_ASAP7_75t_L g4464 ( 
.A(n_4427),
.Y(n_4464)
);

OAI22xp33_ASAP7_75t_L g4465 ( 
.A1(n_4428),
.A2(n_4268),
.B1(n_4226),
.B2(n_4225),
.Y(n_4465)
);

INVx1_ASAP7_75t_SL g4466 ( 
.A(n_4448),
.Y(n_4466)
);

INVx1_ASAP7_75t_L g4467 ( 
.A(n_4434),
.Y(n_4467)
);

INVx1_ASAP7_75t_L g4468 ( 
.A(n_4438),
.Y(n_4468)
);

NAND2xp5_ASAP7_75t_L g4469 ( 
.A(n_4432),
.B(n_4240),
.Y(n_4469)
);

NAND2xp5_ASAP7_75t_L g4470 ( 
.A(n_4431),
.B(n_4265),
.Y(n_4470)
);

INVx1_ASAP7_75t_L g4471 ( 
.A(n_4439),
.Y(n_4471)
);

NAND2xp5_ASAP7_75t_L g4472 ( 
.A(n_4444),
.B(n_4265),
.Y(n_4472)
);

INVx1_ASAP7_75t_L g4473 ( 
.A(n_4446),
.Y(n_4473)
);

NAND3x1_ASAP7_75t_L g4474 ( 
.A(n_4447),
.B(n_4266),
.C(n_4204),
.Y(n_4474)
);

NAND2xp5_ASAP7_75t_SL g4475 ( 
.A(n_4437),
.B(n_4225),
.Y(n_4475)
);

AND2x2_ASAP7_75t_L g4476 ( 
.A(n_4445),
.B(n_4207),
.Y(n_4476)
);

INVxp67_ASAP7_75t_L g4477 ( 
.A(n_4458),
.Y(n_4477)
);

AOI21xp5_ASAP7_75t_L g4478 ( 
.A1(n_4469),
.A2(n_4273),
.B(n_4274),
.Y(n_4478)
);

AO22x2_ASAP7_75t_L g4479 ( 
.A1(n_4456),
.A2(n_4273),
.B1(n_4274),
.B2(n_4225),
.Y(n_4479)
);

OA22x2_ASAP7_75t_L g4480 ( 
.A1(n_4453),
.A2(n_4476),
.B1(n_4473),
.B2(n_4466),
.Y(n_4480)
);

NAND3xp33_ASAP7_75t_SL g4481 ( 
.A(n_4462),
.B(n_4187),
.C(n_4184),
.Y(n_4481)
);

OAI21xp5_ASAP7_75t_L g4482 ( 
.A1(n_4474),
.A2(n_4196),
.B(n_4193),
.Y(n_4482)
);

NAND2xp5_ASAP7_75t_L g4483 ( 
.A(n_4465),
.B(n_4208),
.Y(n_4483)
);

NAND2xp5_ASAP7_75t_SL g4484 ( 
.A(n_4455),
.B(n_4197),
.Y(n_4484)
);

NAND4xp25_ASAP7_75t_L g4485 ( 
.A(n_4454),
.B(n_4199),
.C(n_4121),
.D(n_4169),
.Y(n_4485)
);

AOI21xp5_ASAP7_75t_L g4486 ( 
.A1(n_4475),
.A2(n_4460),
.B(n_4472),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_4457),
.Y(n_4487)
);

AOI21xp5_ASAP7_75t_L g4488 ( 
.A1(n_4470),
.A2(n_4175),
.B(n_4140),
.Y(n_4488)
);

AOI21xp5_ASAP7_75t_L g4489 ( 
.A1(n_4467),
.A2(n_4459),
.B(n_4461),
.Y(n_4489)
);

NOR2x1_ASAP7_75t_SL g4490 ( 
.A(n_4457),
.B(n_4095),
.Y(n_4490)
);

OAI21xp5_ASAP7_75t_L g4491 ( 
.A1(n_4463),
.A2(n_4130),
.B(n_4127),
.Y(n_4491)
);

NOR3xp33_ASAP7_75t_L g4492 ( 
.A(n_4464),
.B(n_4129),
.C(n_4140),
.Y(n_4492)
);

NOR2xp33_ASAP7_75t_L g4493 ( 
.A(n_4468),
.B(n_4115),
.Y(n_4493)
);

OAI222xp33_ASAP7_75t_L g4494 ( 
.A1(n_4480),
.A2(n_4471),
.B1(n_4092),
.B2(n_4112),
.C1(n_4103),
.C2(n_4095),
.Y(n_4494)
);

INVx1_ASAP7_75t_L g4495 ( 
.A(n_4479),
.Y(n_4495)
);

INVxp67_ASAP7_75t_L g4496 ( 
.A(n_4483),
.Y(n_4496)
);

OAI221xp5_ASAP7_75t_L g4497 ( 
.A1(n_4492),
.A2(n_4092),
.B1(n_4110),
.B2(n_4098),
.C(n_4103),
.Y(n_4497)
);

NOR3xp33_ASAP7_75t_L g4498 ( 
.A(n_4477),
.B(n_4127),
.C(n_4123),
.Y(n_4498)
);

OR2x2_ASAP7_75t_L g4499 ( 
.A(n_4485),
.B(n_4098),
.Y(n_4499)
);

NOR4xp25_ASAP7_75t_L g4500 ( 
.A(n_4484),
.B(n_4110),
.C(n_4112),
.D(n_4111),
.Y(n_4500)
);

OAI221xp5_ASAP7_75t_L g4501 ( 
.A1(n_4491),
.A2(n_4111),
.B1(n_4138),
.B2(n_4123),
.C(n_4113),
.Y(n_4501)
);

AOI211xp5_ASAP7_75t_L g4502 ( 
.A1(n_4481),
.A2(n_4138),
.B(n_4161),
.C(n_4145),
.Y(n_4502)
);

INVx1_ASAP7_75t_L g4503 ( 
.A(n_4479),
.Y(n_4503)
);

OAI21xp5_ASAP7_75t_L g4504 ( 
.A1(n_4488),
.A2(n_4145),
.B(n_4151),
.Y(n_4504)
);

AND2x2_ASAP7_75t_L g4505 ( 
.A(n_4493),
.B(n_4201),
.Y(n_4505)
);

NAND2xp5_ASAP7_75t_SL g4506 ( 
.A(n_4486),
.B(n_4145),
.Y(n_4506)
);

AOI22xp5_ASAP7_75t_L g4507 ( 
.A1(n_4489),
.A2(n_4161),
.B1(n_4147),
.B2(n_4146),
.Y(n_4507)
);

INVx1_ASAP7_75t_L g4508 ( 
.A(n_4490),
.Y(n_4508)
);

OAI211xp5_ASAP7_75t_SL g4509 ( 
.A1(n_4506),
.A2(n_4478),
.B(n_4487),
.C(n_4482),
.Y(n_4509)
);

AOI21xp5_ASAP7_75t_L g4510 ( 
.A1(n_4508),
.A2(n_4147),
.B(n_4163),
.Y(n_4510)
);

NAND3xp33_ASAP7_75t_SL g4511 ( 
.A(n_4502),
.B(n_4108),
.C(n_4146),
.Y(n_4511)
);

AOI221xp5_ASAP7_75t_L g4512 ( 
.A1(n_4498),
.A2(n_4494),
.B1(n_4504),
.B2(n_4500),
.C(n_4501),
.Y(n_4512)
);

OAI321xp33_ASAP7_75t_L g4513 ( 
.A1(n_4507),
.A2(n_4113),
.A3(n_4116),
.B1(n_4030),
.B2(n_4085),
.C(n_4155),
.Y(n_4513)
);

OAI211xp5_ASAP7_75t_SL g4514 ( 
.A1(n_4496),
.A2(n_4139),
.B(n_4108),
.C(n_4153),
.Y(n_4514)
);

XNOR2x1_ASAP7_75t_L g4515 ( 
.A(n_4499),
.B(n_4144),
.Y(n_4515)
);

INVx1_ASAP7_75t_SL g4516 ( 
.A(n_4505),
.Y(n_4516)
);

NOR3xp33_ASAP7_75t_L g4517 ( 
.A(n_4495),
.B(n_4139),
.C(n_4153),
.Y(n_4517)
);

INVx2_ASAP7_75t_L g4518 ( 
.A(n_4503),
.Y(n_4518)
);

OAI22xp5_ASAP7_75t_L g4519 ( 
.A1(n_4497),
.A2(n_4101),
.B1(n_4163),
.B2(n_4089),
.Y(n_4519)
);

AOI211x1_ASAP7_75t_SL g4520 ( 
.A1(n_4506),
.A2(n_4155),
.B(n_4150),
.C(n_4099),
.Y(n_4520)
);

AOI322xp5_ASAP7_75t_L g4521 ( 
.A1(n_4498),
.A2(n_4163),
.A3(n_4101),
.B1(n_4085),
.B2(n_4080),
.C1(n_4089),
.C2(n_4153),
.Y(n_4521)
);

INVx1_ASAP7_75t_L g4522 ( 
.A(n_4506),
.Y(n_4522)
);

AOI321xp33_ASAP7_75t_L g4523 ( 
.A1(n_4506),
.A2(n_4101),
.A3(n_4044),
.B1(n_3990),
.B2(n_3992),
.C(n_4034),
.Y(n_4523)
);

NOR2xp33_ASAP7_75t_L g4524 ( 
.A(n_4506),
.B(n_4144),
.Y(n_4524)
);

NOR3xp33_ASAP7_75t_L g4525 ( 
.A(n_4496),
.B(n_4150),
.C(n_4135),
.Y(n_4525)
);

NOR3xp33_ASAP7_75t_L g4526 ( 
.A(n_4496),
.B(n_4135),
.C(n_4152),
.Y(n_4526)
);

INVx1_ASAP7_75t_L g4527 ( 
.A(n_4526),
.Y(n_4527)
);

NAND4xp75_ASAP7_75t_L g4528 ( 
.A(n_4512),
.B(n_4522),
.C(n_4518),
.D(n_4524),
.Y(n_4528)
);

INVx1_ASAP7_75t_L g4529 ( 
.A(n_4515),
.Y(n_4529)
);

NOR3xp33_ASAP7_75t_L g4530 ( 
.A(n_4509),
.B(n_4152),
.C(n_4069),
.Y(n_4530)
);

NOR2xp33_ASAP7_75t_L g4531 ( 
.A(n_4511),
.B(n_4080),
.Y(n_4531)
);

INVx2_ASAP7_75t_L g4532 ( 
.A(n_4516),
.Y(n_4532)
);

NAND4xp75_ASAP7_75t_L g4533 ( 
.A(n_4510),
.B(n_4090),
.C(n_3949),
.D(n_3948),
.Y(n_4533)
);

NAND4xp75_ASAP7_75t_L g4534 ( 
.A(n_4520),
.B(n_4090),
.C(n_3946),
.D(n_3948),
.Y(n_4534)
);

NOR4xp75_ASAP7_75t_L g4535 ( 
.A(n_4519),
.B(n_4057),
.C(n_4056),
.D(n_4052),
.Y(n_4535)
);

NAND3xp33_ASAP7_75t_SL g4536 ( 
.A(n_4525),
.B(n_4033),
.C(n_4028),
.Y(n_4536)
);

NOR2x1_ASAP7_75t_L g4537 ( 
.A(n_4514),
.B(n_4136),
.Y(n_4537)
);

OR2x2_ASAP7_75t_L g4538 ( 
.A(n_4517),
.B(n_4080),
.Y(n_4538)
);

NAND2xp5_ASAP7_75t_L g4539 ( 
.A(n_4521),
.B(n_4136),
.Y(n_4539)
);

NAND3xp33_ASAP7_75t_L g4540 ( 
.A(n_4523),
.B(n_4089),
.C(n_4136),
.Y(n_4540)
);

NAND2xp5_ASAP7_75t_L g4541 ( 
.A(n_4513),
.B(n_4152),
.Y(n_4541)
);

NAND2xp33_ASAP7_75t_L g4542 ( 
.A(n_4525),
.B(n_3838),
.Y(n_4542)
);

OA22x2_ASAP7_75t_L g4543 ( 
.A1(n_4516),
.A2(n_3914),
.B1(n_3924),
.B2(n_3897),
.Y(n_4543)
);

NAND3xp33_ASAP7_75t_SL g4544 ( 
.A(n_4532),
.B(n_4026),
.C(n_4022),
.Y(n_4544)
);

AOI221x1_ASAP7_75t_L g4545 ( 
.A1(n_4527),
.A2(n_3924),
.B1(n_3914),
.B2(n_3843),
.C(n_3950),
.Y(n_4545)
);

AOI21xp5_ASAP7_75t_L g4546 ( 
.A1(n_4539),
.A2(n_3843),
.B(n_3914),
.Y(n_4546)
);

OAI211xp5_ASAP7_75t_L g4547 ( 
.A1(n_4529),
.A2(n_4005),
.B(n_4019),
.C(n_4023),
.Y(n_4547)
);

AOI211xp5_ASAP7_75t_L g4548 ( 
.A1(n_4531),
.A2(n_3888),
.B(n_3924),
.C(n_4048),
.Y(n_4548)
);

NOR3xp33_ASAP7_75t_L g4549 ( 
.A(n_4528),
.B(n_4541),
.C(n_4540),
.Y(n_4549)
);

NAND2xp5_ASAP7_75t_L g4550 ( 
.A(n_4530),
.B(n_4001),
.Y(n_4550)
);

O2A1O1Ixp5_ASAP7_75t_L g4551 ( 
.A1(n_4538),
.A2(n_3896),
.B(n_3870),
.C(n_3859),
.Y(n_4551)
);

AOI221xp5_ASAP7_75t_L g4552 ( 
.A1(n_4542),
.A2(n_3869),
.B1(n_3863),
.B2(n_3865),
.C(n_3867),
.Y(n_4552)
);

AOI21xp33_ASAP7_75t_SL g4553 ( 
.A1(n_4543),
.A2(n_359),
.B(n_361),
.Y(n_4553)
);

AND2x2_ASAP7_75t_L g4554 ( 
.A(n_4537),
.B(n_3887),
.Y(n_4554)
);

INVx1_ASAP7_75t_L g4555 ( 
.A(n_4554),
.Y(n_4555)
);

INVx1_ASAP7_75t_SL g4556 ( 
.A(n_4550),
.Y(n_4556)
);

INVx2_ASAP7_75t_L g4557 ( 
.A(n_4551),
.Y(n_4557)
);

NAND2xp5_ASAP7_75t_L g4558 ( 
.A(n_4546),
.B(n_4533),
.Y(n_4558)
);

NOR2x1_ASAP7_75t_L g4559 ( 
.A(n_4544),
.B(n_4536),
.Y(n_4559)
);

AND2x4_ASAP7_75t_L g4560 ( 
.A(n_4549),
.B(n_4535),
.Y(n_4560)
);

NAND4xp75_ASAP7_75t_L g4561 ( 
.A(n_4559),
.B(n_4545),
.C(n_4553),
.D(n_4552),
.Y(n_4561)
);

NOR5xp2_ASAP7_75t_L g4562 ( 
.A(n_4555),
.B(n_4547),
.C(n_4534),
.D(n_4548),
.E(n_3854),
.Y(n_4562)
);

OAI211xp5_ASAP7_75t_L g4563 ( 
.A1(n_4558),
.A2(n_4064),
.B(n_4046),
.C(n_4054),
.Y(n_4563)
);

HB1xp67_ASAP7_75t_L g4564 ( 
.A(n_4561),
.Y(n_4564)
);

INVx2_ASAP7_75t_L g4565 ( 
.A(n_4562),
.Y(n_4565)
);

INVx2_ASAP7_75t_L g4566 ( 
.A(n_4565),
.Y(n_4566)
);

OAI22x1_ASAP7_75t_L g4567 ( 
.A1(n_4566),
.A2(n_4560),
.B1(n_4564),
.B2(n_4557),
.Y(n_4567)
);

INVx1_ASAP7_75t_L g4568 ( 
.A(n_4567),
.Y(n_4568)
);

NAND4xp25_ASAP7_75t_SL g4569 ( 
.A(n_4568),
.B(n_4556),
.C(n_4563),
.D(n_4065),
.Y(n_4569)
);

AOI22xp5_ASAP7_75t_L g4570 ( 
.A1(n_4569),
.A2(n_3895),
.B1(n_3899),
.B2(n_3898),
.Y(n_4570)
);

OAI221xp5_ASAP7_75t_L g4571 ( 
.A1(n_4570),
.A2(n_4060),
.B1(n_363),
.B2(n_364),
.C(n_366),
.Y(n_4571)
);

OAI22xp33_ASAP7_75t_SL g4572 ( 
.A1(n_4571),
.A2(n_362),
.B1(n_367),
.B2(n_372),
.Y(n_4572)
);

AOI22xp5_ASAP7_75t_L g4573 ( 
.A1(n_4572),
.A2(n_3870),
.B1(n_3869),
.B2(n_3863),
.Y(n_4573)
);

XNOR2xp5_ASAP7_75t_L g4574 ( 
.A(n_4573),
.B(n_374),
.Y(n_4574)
);

AOI21xp5_ASAP7_75t_L g4575 ( 
.A1(n_4574),
.A2(n_376),
.B(n_378),
.Y(n_4575)
);

NAND2xp5_ASAP7_75t_L g4576 ( 
.A(n_4574),
.B(n_386),
.Y(n_4576)
);

HB1xp67_ASAP7_75t_L g4577 ( 
.A(n_4576),
.Y(n_4577)
);

XNOR2xp5_ASAP7_75t_L g4578 ( 
.A(n_4575),
.B(n_393),
.Y(n_4578)
);

OA21x2_ASAP7_75t_L g4579 ( 
.A1(n_4577),
.A2(n_3880),
.B(n_3867),
.Y(n_4579)
);

XNOR2xp5_ASAP7_75t_L g4580 ( 
.A(n_4578),
.B(n_394),
.Y(n_4580)
);

OAI221xp5_ASAP7_75t_R g4581 ( 
.A1(n_4580),
.A2(n_398),
.B1(n_403),
.B2(n_405),
.C(n_416),
.Y(n_4581)
);

OAI221xp5_ASAP7_75t_R g4582 ( 
.A1(n_4579),
.A2(n_418),
.B1(n_421),
.B2(n_427),
.C(n_432),
.Y(n_4582)
);

AOI22xp5_ASAP7_75t_L g4583 ( 
.A1(n_4582),
.A2(n_4581),
.B1(n_3854),
.B2(n_3865),
.Y(n_4583)
);

AOI211xp5_ASAP7_75t_L g4584 ( 
.A1(n_4583),
.A2(n_434),
.B(n_435),
.C(n_436),
.Y(n_4584)
);


endmodule