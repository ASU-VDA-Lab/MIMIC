module real_aes_7121_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_505;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g259 ( .A1(n_0), .A2(n_260), .B(n_261), .C(n_264), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_1), .B(n_248), .Y(n_265) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_2), .B(n_107), .C(n_108), .Y(n_106) );
INVx1_ASAP7_75t_L g455 ( .A(n_2), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_3), .B(n_176), .Y(n_175) );
A2O1A1Ixp33_ASAP7_75t_L g539 ( .A1(n_4), .A2(n_137), .B(n_140), .C(n_540), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_5), .A2(n_132), .B(n_564), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_6), .A2(n_132), .B(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_7), .B(n_248), .Y(n_570) );
AO21x2_ASAP7_75t_L g203 ( .A1(n_8), .A2(n_167), .B(n_204), .Y(n_203) );
AND2x6_ASAP7_75t_L g137 ( .A(n_9), .B(n_138), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_10), .A2(n_137), .B(n_140), .C(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g508 ( .A(n_11), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_12), .B(n_105), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_12), .B(n_41), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_13), .B(n_224), .Y(n_542) );
INVx1_ASAP7_75t_L g158 ( .A(n_14), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_15), .B(n_176), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_16), .A2(n_177), .B(n_526), .C(n_528), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_17), .B(n_248), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_18), .B(n_152), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g139 ( .A1(n_19), .A2(n_140), .B(n_143), .C(n_151), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_20), .A2(n_212), .B(n_263), .C(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_21), .B(n_224), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_22), .A2(n_102), .B1(n_111), .B2(n_752), .Y(n_101) );
AOI22xp5_ASAP7_75t_L g118 ( .A1(n_23), .A2(n_119), .B1(n_120), .B2(n_448), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_23), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_24), .B(n_224), .Y(n_481) );
CKINVDCx16_ASAP7_75t_R g555 ( .A(n_25), .Y(n_555) );
INVx1_ASAP7_75t_L g480 ( .A(n_26), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_27), .A2(n_140), .B(n_151), .C(n_207), .Y(n_206) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_28), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_29), .Y(n_538) );
INVx1_ASAP7_75t_L g496 ( .A(n_30), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_31), .B(n_458), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_32), .A2(n_132), .B(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g135 ( .A(n_33), .Y(n_135) );
A2O1A1Ixp33_ASAP7_75t_L g188 ( .A1(n_34), .A2(n_180), .B(n_189), .C(n_191), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_35), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g566 ( .A1(n_36), .A2(n_263), .B(n_567), .C(n_569), .Y(n_566) );
INVxp67_ASAP7_75t_L g497 ( .A(n_37), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_38), .B(n_209), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_39), .A2(n_140), .B(n_151), .C(n_479), .Y(n_478) );
CKINVDCx14_ASAP7_75t_R g565 ( .A(n_40), .Y(n_565) );
INVx1_ASAP7_75t_L g105 ( .A(n_41), .Y(n_105) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_42), .A2(n_264), .B(n_506), .C(n_507), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_43), .B(n_131), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_44), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_45), .B(n_176), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_46), .B(n_132), .Y(n_205) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_47), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_48), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_49), .A2(n_180), .B(n_189), .C(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g262 ( .A(n_50), .Y(n_262) );
OAI22xp5_ASAP7_75t_L g120 ( .A1(n_51), .A2(n_121), .B1(n_122), .B2(n_447), .Y(n_120) );
CKINVDCx16_ASAP7_75t_R g121 ( .A(n_51), .Y(n_121) );
INVx1_ASAP7_75t_L g234 ( .A(n_52), .Y(n_234) );
INVx1_ASAP7_75t_L g514 ( .A(n_53), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_54), .B(n_132), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_55), .Y(n_160) );
CKINVDCx14_ASAP7_75t_R g504 ( .A(n_56), .Y(n_504) );
INVx1_ASAP7_75t_L g138 ( .A(n_57), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_58), .B(n_132), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_59), .B(n_248), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_60), .A2(n_150), .B(n_173), .C(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g157 ( .A(n_61), .Y(n_157) );
OAI22xp5_ASAP7_75t_L g461 ( .A1(n_62), .A2(n_100), .B1(n_462), .B2(n_463), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_62), .Y(n_463) );
INVx1_ASAP7_75t_SL g568 ( .A(n_63), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_64), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_65), .B(n_176), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_66), .B(n_248), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_67), .B(n_177), .Y(n_222) );
INVx1_ASAP7_75t_L g558 ( .A(n_68), .Y(n_558) );
CKINVDCx16_ASAP7_75t_R g258 ( .A(n_69), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_70), .B(n_145), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g170 ( .A1(n_71), .A2(n_140), .B(n_171), .C(n_180), .Y(n_170) );
CKINVDCx16_ASAP7_75t_R g243 ( .A(n_72), .Y(n_243) );
INVx1_ASAP7_75t_L g110 ( .A(n_73), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_74), .A2(n_132), .B(n_503), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_75), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_76), .A2(n_132), .B(n_523), .Y(n_522) );
AOI222xp33_ASAP7_75t_SL g460 ( .A1(n_77), .A2(n_461), .B1(n_464), .B2(n_743), .C1(n_744), .C2(n_748), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_78), .A2(n_131), .B(n_492), .Y(n_491) );
CKINVDCx16_ASAP7_75t_R g477 ( .A(n_79), .Y(n_477) );
INVx1_ASAP7_75t_L g524 ( .A(n_80), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_81), .B(n_148), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_82), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_83), .A2(n_132), .B(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g527 ( .A(n_84), .Y(n_527) );
INVx2_ASAP7_75t_L g155 ( .A(n_85), .Y(n_155) );
INVx1_ASAP7_75t_L g541 ( .A(n_86), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_87), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_88), .B(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g107 ( .A(n_89), .Y(n_107) );
OR2x2_ASAP7_75t_L g452 ( .A(n_89), .B(n_453), .Y(n_452) );
OR2x2_ASAP7_75t_L g467 ( .A(n_89), .B(n_454), .Y(n_467) );
A2O1A1Ixp33_ASAP7_75t_L g556 ( .A1(n_90), .A2(n_140), .B(n_180), .C(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_91), .B(n_132), .Y(n_187) );
INVx1_ASAP7_75t_L g192 ( .A(n_92), .Y(n_192) );
INVxp67_ASAP7_75t_L g246 ( .A(n_93), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_94), .B(n_167), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_95), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g172 ( .A(n_96), .Y(n_172) );
INVx1_ASAP7_75t_L g218 ( .A(n_97), .Y(n_218) );
INVx2_ASAP7_75t_L g517 ( .A(n_98), .Y(n_517) );
AND2x2_ASAP7_75t_L g236 ( .A(n_99), .B(n_154), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_100), .Y(n_462) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_SL g753 ( .A(n_103), .Y(n_753) );
OR2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
OR2x2_ASAP7_75t_L g468 ( .A(n_107), .B(n_454), .Y(n_468) );
NOR2x2_ASAP7_75t_L g750 ( .A(n_107), .B(n_453), .Y(n_750) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
OA21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_117), .B(n_459), .Y(n_111) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g751 ( .A(n_116), .Y(n_751) );
OAI21xp5_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_449), .B(n_457), .Y(n_117) );
INVxp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI22xp5_ASAP7_75t_SL g744 ( .A1(n_122), .A2(n_470), .B1(n_745), .B2(n_746), .Y(n_744) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
BUFx2_ASAP7_75t_L g447 ( .A(n_123), .Y(n_447) );
AND3x1_ASAP7_75t_L g123 ( .A(n_124), .B(n_351), .C(n_408), .Y(n_123) );
NOR3xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_296), .C(n_332), .Y(n_124) );
OAI211xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_198), .B(n_250), .C(n_283), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_162), .Y(n_126) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g253 ( .A(n_128), .B(n_254), .Y(n_253) );
INVx5_ASAP7_75t_L g282 ( .A(n_128), .Y(n_282) );
AND2x2_ASAP7_75t_L g355 ( .A(n_128), .B(n_271), .Y(n_355) );
AND2x2_ASAP7_75t_L g393 ( .A(n_128), .B(n_299), .Y(n_393) );
AND2x2_ASAP7_75t_L g413 ( .A(n_128), .B(n_255), .Y(n_413) );
OR2x6_ASAP7_75t_L g128 ( .A(n_129), .B(n_159), .Y(n_128) );
AOI21xp5_ASAP7_75t_SL g129 ( .A1(n_130), .A2(n_139), .B(n_152), .Y(n_129) );
BUFx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_137), .Y(n_132) );
NAND2x1p5_ASAP7_75t_L g219 ( .A(n_133), .B(n_137), .Y(n_219) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
INVx1_ASAP7_75t_L g150 ( .A(n_134), .Y(n_150) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g141 ( .A(n_135), .Y(n_141) );
INVx1_ASAP7_75t_L g213 ( .A(n_135), .Y(n_213) );
INVx1_ASAP7_75t_L g142 ( .A(n_136), .Y(n_142) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_136), .Y(n_146) );
INVx3_ASAP7_75t_L g177 ( .A(n_136), .Y(n_177) );
INVx1_ASAP7_75t_L g209 ( .A(n_136), .Y(n_209) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_136), .Y(n_224) );
BUFx3_ASAP7_75t_L g151 ( .A(n_137), .Y(n_151) );
INVx4_ASAP7_75t_SL g181 ( .A(n_137), .Y(n_181) );
INVx5_ASAP7_75t_L g190 ( .A(n_140), .Y(n_190) );
AND2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_141), .Y(n_179) );
BUFx3_ASAP7_75t_L g195 ( .A(n_141), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_147), .B(n_149), .Y(n_143) );
INVx2_ASAP7_75t_L g148 ( .A(n_145), .Y(n_148) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx4_ASAP7_75t_L g174 ( .A(n_146), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_L g191 ( .A1(n_148), .A2(n_192), .B(n_193), .C(n_194), .Y(n_191) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_148), .A2(n_194), .B(n_234), .C(n_235), .Y(n_233) );
O2A1O1Ixp5_ASAP7_75t_L g540 ( .A1(n_148), .A2(n_541), .B(n_542), .C(n_543), .Y(n_540) );
O2A1O1Ixp33_ASAP7_75t_L g557 ( .A1(n_148), .A2(n_543), .B(n_558), .C(n_559), .Y(n_557) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_149), .A2(n_176), .B(n_480), .C(n_481), .Y(n_479) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_150), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_153), .B(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g161 ( .A(n_154), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_154), .A2(n_187), .B(n_188), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_154), .A2(n_231), .B(n_232), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_154), .A2(n_219), .B(n_477), .C(n_478), .Y(n_476) );
OA21x2_ASAP7_75t_L g501 ( .A1(n_154), .A2(n_502), .B(n_509), .Y(n_501) );
AND2x2_ASAP7_75t_SL g154 ( .A(n_155), .B(n_156), .Y(n_154) );
AND2x2_ASAP7_75t_L g168 ( .A(n_155), .B(n_156), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
AO21x2_ASAP7_75t_L g536 ( .A1(n_161), .A2(n_537), .B(n_544), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_162), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g162 ( .A(n_163), .B(n_185), .Y(n_162) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_163), .Y(n_294) );
AND2x2_ASAP7_75t_L g308 ( .A(n_163), .B(n_254), .Y(n_308) );
INVx1_ASAP7_75t_L g331 ( .A(n_163), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_163), .B(n_282), .Y(n_370) );
OR2x2_ASAP7_75t_L g407 ( .A(n_163), .B(n_252), .Y(n_407) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_164), .Y(n_343) );
AND2x2_ASAP7_75t_L g350 ( .A(n_164), .B(n_255), .Y(n_350) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g271 ( .A(n_165), .B(n_255), .Y(n_271) );
BUFx2_ASAP7_75t_L g299 ( .A(n_165), .Y(n_299) );
AO21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_169), .B(n_183), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_166), .B(n_184), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_166), .B(n_197), .Y(n_196) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_166), .A2(n_217), .B(n_225), .Y(n_216) );
INVx3_ASAP7_75t_L g248 ( .A(n_166), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_166), .B(n_483), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_166), .B(n_545), .Y(n_544) );
AO21x2_ASAP7_75t_L g553 ( .A1(n_166), .A2(n_554), .B(n_560), .Y(n_553) );
INVx4_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_167), .A2(n_205), .B(n_206), .Y(n_204) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_167), .Y(n_240) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g227 ( .A(n_168), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_170), .B(n_182), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_175), .C(n_178), .Y(n_171) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
OAI22xp33_ASAP7_75t_L g495 ( .A1(n_174), .A2(n_176), .B1(n_496), .B2(n_497), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_174), .B(n_517), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_174), .B(n_527), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_176), .B(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g260 ( .A(n_176), .Y(n_260) );
INVx5_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_177), .B(n_508), .Y(n_507) );
HB1xp67_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx3_ASAP7_75t_L g569 ( .A(n_179), .Y(n_569) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_181), .A2(n_190), .B(n_243), .C(n_244), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_SL g257 ( .A1(n_181), .A2(n_190), .B(n_258), .C(n_259), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_SL g492 ( .A1(n_181), .A2(n_190), .B(n_493), .C(n_494), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_SL g503 ( .A1(n_181), .A2(n_190), .B(n_504), .C(n_505), .Y(n_503) );
O2A1O1Ixp33_ASAP7_75t_SL g513 ( .A1(n_181), .A2(n_190), .B(n_514), .C(n_515), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_SL g523 ( .A1(n_181), .A2(n_190), .B(n_524), .C(n_525), .Y(n_523) );
O2A1O1Ixp33_ASAP7_75t_L g564 ( .A1(n_181), .A2(n_190), .B(n_565), .C(n_566), .Y(n_564) );
INVx5_ASAP7_75t_L g252 ( .A(n_185), .Y(n_252) );
BUFx2_ASAP7_75t_L g275 ( .A(n_185), .Y(n_275) );
AND2x2_ASAP7_75t_L g432 ( .A(n_185), .B(n_286), .Y(n_432) );
OR2x6_ASAP7_75t_L g185 ( .A(n_186), .B(n_196), .Y(n_185) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
HB1xp67_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g264 ( .A(n_195), .Y(n_264) );
INVx1_ASAP7_75t_L g528 ( .A(n_195), .Y(n_528) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NAND2xp33_ASAP7_75t_L g199 ( .A(n_200), .B(n_237), .Y(n_199) );
OAI221xp5_ASAP7_75t_L g332 ( .A1(n_200), .A2(n_333), .B1(n_340), .B2(n_341), .C(n_344), .Y(n_332) );
OR2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_214), .Y(n_200) );
AND2x2_ASAP7_75t_L g238 ( .A(n_201), .B(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_201), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_SL g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g267 ( .A(n_202), .B(n_215), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_202), .B(n_216), .Y(n_277) );
OR2x2_ASAP7_75t_L g288 ( .A(n_202), .B(n_239), .Y(n_288) );
AND2x2_ASAP7_75t_L g291 ( .A(n_202), .B(n_279), .Y(n_291) );
AND2x2_ASAP7_75t_L g307 ( .A(n_202), .B(n_228), .Y(n_307) );
OR2x2_ASAP7_75t_L g323 ( .A(n_202), .B(n_216), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_202), .B(n_239), .Y(n_385) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_203), .B(n_228), .Y(n_377) );
AND2x2_ASAP7_75t_L g380 ( .A(n_203), .B(n_216), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_210), .B(n_211), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_211), .A2(n_222), .B(n_223), .Y(n_221) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
OR2x2_ASAP7_75t_L g301 ( .A(n_214), .B(n_288), .Y(n_301) );
INVx2_ASAP7_75t_L g327 ( .A(n_214), .Y(n_327) );
OR2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_228), .Y(n_214) );
AND2x2_ASAP7_75t_L g249 ( .A(n_215), .B(n_229), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_215), .B(n_239), .Y(n_306) );
OR2x2_ASAP7_75t_L g317 ( .A(n_215), .B(n_229), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_215), .B(n_279), .Y(n_376) );
OAI221xp5_ASAP7_75t_L g409 ( .A1(n_215), .A2(n_410), .B1(n_412), .B2(n_414), .C(n_417), .Y(n_409) );
INVx5_ASAP7_75t_SL g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_216), .B(n_239), .Y(n_348) );
OAI21xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_220), .Y(n_217) );
OAI21xp5_ASAP7_75t_L g537 ( .A1(n_219), .A2(n_538), .B(n_539), .Y(n_537) );
OAI21xp5_ASAP7_75t_L g554 ( .A1(n_219), .A2(n_555), .B(n_556), .Y(n_554) );
INVx4_ASAP7_75t_L g263 ( .A(n_224), .Y(n_263) );
INVx2_ASAP7_75t_L g506 ( .A(n_224), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
INVx2_ASAP7_75t_L g489 ( .A(n_227), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_228), .B(n_279), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_228), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g295 ( .A(n_228), .B(n_267), .Y(n_295) );
OR2x2_ASAP7_75t_L g339 ( .A(n_228), .B(n_239), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_228), .B(n_291), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_228), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g404 ( .A(n_228), .B(n_405), .Y(n_404) );
INVx5_ASAP7_75t_SL g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_SL g268 ( .A(n_229), .B(n_238), .Y(n_268) );
O2A1O1Ixp33_ASAP7_75t_SL g272 ( .A1(n_229), .A2(n_273), .B(n_276), .C(n_280), .Y(n_272) );
OR2x2_ASAP7_75t_L g310 ( .A(n_229), .B(n_306), .Y(n_310) );
OR2x2_ASAP7_75t_L g346 ( .A(n_229), .B(n_288), .Y(n_346) );
OAI311xp33_ASAP7_75t_L g352 ( .A1(n_229), .A2(n_291), .A3(n_353), .B1(n_356), .C1(n_363), .Y(n_352) );
AND2x2_ASAP7_75t_L g403 ( .A(n_229), .B(n_239), .Y(n_403) );
AND2x2_ASAP7_75t_L g411 ( .A(n_229), .B(n_266), .Y(n_411) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_229), .Y(n_429) );
AND2x2_ASAP7_75t_L g446 ( .A(n_229), .B(n_267), .Y(n_446) );
OR2x6_ASAP7_75t_L g229 ( .A(n_230), .B(n_236), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_249), .Y(n_237) );
AND2x2_ASAP7_75t_L g274 ( .A(n_238), .B(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g430 ( .A(n_238), .Y(n_430) );
AND2x2_ASAP7_75t_L g266 ( .A(n_239), .B(n_267), .Y(n_266) );
INVx3_ASAP7_75t_L g279 ( .A(n_239), .Y(n_279) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_239), .Y(n_322) );
INVxp67_ASAP7_75t_L g361 ( .A(n_239), .Y(n_361) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_247), .Y(n_239) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_240), .A2(n_512), .B(n_518), .Y(n_511) );
OA21x2_ASAP7_75t_L g521 ( .A1(n_240), .A2(n_522), .B(n_529), .Y(n_521) );
OA21x2_ASAP7_75t_L g562 ( .A1(n_240), .A2(n_563), .B(n_570), .Y(n_562) );
OA21x2_ASAP7_75t_L g255 ( .A1(n_248), .A2(n_256), .B(n_265), .Y(n_255) );
AND2x2_ASAP7_75t_L g439 ( .A(n_249), .B(n_287), .Y(n_439) );
AOI221xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_266), .B1(n_268), .B2(n_269), .C(n_272), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_252), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g292 ( .A(n_252), .B(n_282), .Y(n_292) );
AND2x2_ASAP7_75t_L g300 ( .A(n_252), .B(n_254), .Y(n_300) );
OR2x2_ASAP7_75t_L g312 ( .A(n_252), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g330 ( .A(n_252), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g354 ( .A(n_252), .B(n_355), .Y(n_354) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_252), .Y(n_374) );
AND2x2_ASAP7_75t_L g426 ( .A(n_252), .B(n_350), .Y(n_426) );
OAI31xp33_ASAP7_75t_L g434 ( .A1(n_252), .A2(n_303), .A3(n_402), .B(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_253), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_SL g398 ( .A(n_253), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_253), .B(n_407), .Y(n_406) );
AND2x4_ASAP7_75t_L g286 ( .A(n_254), .B(n_282), .Y(n_286) );
INVx1_ASAP7_75t_L g373 ( .A(n_254), .Y(n_373) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g423 ( .A(n_255), .B(n_282), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_263), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g543 ( .A(n_264), .Y(n_543) );
INVx1_ASAP7_75t_SL g433 ( .A(n_266), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_267), .B(n_338), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_268), .A2(n_380), .B1(n_418), .B2(n_421), .Y(n_417) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g281 ( .A(n_271), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g340 ( .A(n_271), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_271), .B(n_292), .Y(n_445) );
INVx1_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g415 ( .A(n_274), .B(n_416), .Y(n_415) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_275), .A2(n_334), .B(n_336), .Y(n_333) );
OR2x2_ASAP7_75t_L g341 ( .A(n_275), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g362 ( .A(n_275), .B(n_350), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_275), .B(n_373), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_275), .B(n_413), .Y(n_412) );
OAI221xp5_ASAP7_75t_SL g389 ( .A1(n_276), .A2(n_390), .B1(n_395), .B2(n_398), .C(n_399), .Y(n_389) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
OR2x2_ASAP7_75t_L g366 ( .A(n_277), .B(n_339), .Y(n_366) );
INVx1_ASAP7_75t_L g405 ( .A(n_277), .Y(n_405) );
INVx2_ASAP7_75t_L g381 ( .A(n_278), .Y(n_381) );
INVx1_ASAP7_75t_L g315 ( .A(n_279), .Y(n_315) );
INVx1_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g320 ( .A(n_282), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_282), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g349 ( .A(n_282), .B(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g437 ( .A(n_282), .B(n_407), .Y(n_437) );
AOI222xp33_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_287), .B1(n_289), .B2(n_292), .C1(n_293), .C2(n_295), .Y(n_283) );
INVxp67_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g293 ( .A(n_286), .B(n_294), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_286), .A2(n_336), .B1(n_364), .B2(n_365), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_286), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
OAI21xp33_ASAP7_75t_SL g324 ( .A1(n_295), .A2(n_325), .B(n_328), .Y(n_324) );
OAI211xp5_ASAP7_75t_SL g296 ( .A1(n_297), .A2(n_301), .B(n_302), .C(n_324), .Y(n_296) );
INVxp67_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
AOI221xp5_ASAP7_75t_L g302 ( .A1(n_300), .A2(n_303), .B1(n_308), .B2(n_309), .C(n_311), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_300), .B(n_388), .Y(n_387) );
INVxp67_ASAP7_75t_L g394 ( .A(n_300), .Y(n_394) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
AND2x2_ASAP7_75t_L g396 ( .A(n_305), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g313 ( .A(n_308), .Y(n_313) );
AND2x2_ASAP7_75t_L g319 ( .A(n_308), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_314), .B1(n_318), .B2(n_321), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_315), .B(n_327), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_316), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g416 ( .A(n_320), .Y(n_416) );
AND2x2_ASAP7_75t_L g435 ( .A(n_320), .B(n_350), .Y(n_435) );
OR2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_327), .B(n_384), .Y(n_443) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_330), .B(n_398), .Y(n_441) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g364 ( .A(n_342), .Y(n_364) );
BUFx2_ASAP7_75t_L g388 ( .A(n_343), .Y(n_388) );
OAI21xp5_ASAP7_75t_SL g344 ( .A1(n_345), .A2(n_347), .B(n_349), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NOR3xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_367), .C(n_389), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OAI21xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_359), .B(n_362), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
A2O1A1Ixp33_ASAP7_75t_SL g367 ( .A1(n_368), .A2(n_371), .B(n_375), .C(n_378), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_368), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NOR2xp67_ASAP7_75t_SL g372 ( .A(n_373), .B(n_374), .Y(n_372) );
OR2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
INVx1_ASAP7_75t_SL g397 ( .A(n_377), .Y(n_397) );
OAI21xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_382), .B(n_386), .Y(n_378) );
AND2x4_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
AND2x2_ASAP7_75t_L g402 ( .A(n_380), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_392), .B(n_394), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_402), .B1(n_404), .B2(n_406), .Y(n_399) );
INVx2_ASAP7_75t_SL g420 ( .A(n_407), .Y(n_420) );
NOR3xp33_ASAP7_75t_L g408 ( .A(n_409), .B(n_424), .C(n_436), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVxp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVxp67_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_420), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OAI221xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_427), .B1(n_431), .B2(n_433), .C(n_434), .Y(n_424) );
A2O1A1Ixp33_ASAP7_75t_L g436 ( .A1(n_425), .A2(n_437), .B(n_438), .C(n_440), .Y(n_436) );
INVx1_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
INVxp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_442), .B1(n_444), .B2(n_446), .Y(n_440) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_447), .A2(n_465), .B1(n_468), .B2(n_469), .Y(n_464) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g458 ( .A(n_452), .Y(n_458) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_457), .B(n_460), .C(n_751), .Y(n_459) );
INVx1_ASAP7_75t_L g743 ( .A(n_461), .Y(n_743) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g745 ( .A(n_466), .Y(n_745) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g747 ( .A(n_468), .Y(n_747) );
INVx1_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
OR5x1_ASAP7_75t_L g470 ( .A(n_471), .B(n_637), .C(n_701), .D(n_717), .E(n_732), .Y(n_470) );
NAND4xp25_ASAP7_75t_L g471 ( .A(n_472), .B(n_571), .C(n_598), .D(n_621), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_519), .B(n_530), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_484), .Y(n_473) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx3_ASAP7_75t_SL g550 ( .A(n_475), .Y(n_550) );
AND2x4_ASAP7_75t_L g584 ( .A(n_475), .B(n_573), .Y(n_584) );
OR2x2_ASAP7_75t_L g594 ( .A(n_475), .B(n_552), .Y(n_594) );
OR2x2_ASAP7_75t_L g640 ( .A(n_475), .B(n_487), .Y(n_640) );
AND2x2_ASAP7_75t_L g654 ( .A(n_475), .B(n_551), .Y(n_654) );
AND2x2_ASAP7_75t_L g697 ( .A(n_475), .B(n_587), .Y(n_697) );
AND2x2_ASAP7_75t_L g704 ( .A(n_475), .B(n_562), .Y(n_704) );
AND2x2_ASAP7_75t_L g723 ( .A(n_475), .B(n_613), .Y(n_723) );
AND2x2_ASAP7_75t_L g741 ( .A(n_475), .B(n_583), .Y(n_741) );
OR2x6_ASAP7_75t_L g475 ( .A(n_476), .B(n_482), .Y(n_475) );
INVx1_ASAP7_75t_L g706 ( .A(n_484), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_500), .Y(n_484) );
AND2x2_ASAP7_75t_L g616 ( .A(n_485), .B(n_551), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_485), .B(n_636), .Y(n_635) );
AOI32xp33_ASAP7_75t_L g649 ( .A1(n_485), .A2(n_650), .A3(n_653), .B1(n_655), .B2(n_659), .Y(n_649) );
AND2x2_ASAP7_75t_L g719 ( .A(n_485), .B(n_613), .Y(n_719) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g583 ( .A(n_487), .B(n_552), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_487), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g625 ( .A(n_487), .B(n_572), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_487), .B(n_704), .Y(n_703) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_490), .B(n_498), .Y(n_487) );
INVx1_ASAP7_75t_L g588 ( .A(n_488), .Y(n_588) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OA21x2_ASAP7_75t_L g587 ( .A1(n_491), .A2(n_499), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g590 ( .A(n_500), .B(n_534), .Y(n_590) );
AND2x2_ASAP7_75t_L g666 ( .A(n_500), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_SL g738 ( .A(n_500), .Y(n_738) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_510), .Y(n_500) );
OR2x2_ASAP7_75t_L g533 ( .A(n_501), .B(n_511), .Y(n_533) );
AND2x2_ASAP7_75t_L g547 ( .A(n_501), .B(n_548), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_501), .B(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g597 ( .A(n_501), .Y(n_597) );
AND2x2_ASAP7_75t_L g624 ( .A(n_501), .B(n_511), .Y(n_624) );
BUFx3_ASAP7_75t_L g627 ( .A(n_501), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_501), .B(n_602), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_501), .B(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g578 ( .A(n_510), .Y(n_578) );
AND2x2_ASAP7_75t_L g596 ( .A(n_510), .B(n_576), .Y(n_596) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g607 ( .A(n_511), .B(n_521), .Y(n_607) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_511), .Y(n_620) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_520), .B(n_627), .Y(n_677) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_SL g548 ( .A(n_521), .Y(n_548) );
NAND3xp33_ASAP7_75t_L g595 ( .A(n_521), .B(n_596), .C(n_597), .Y(n_595) );
OR2x2_ASAP7_75t_L g603 ( .A(n_521), .B(n_576), .Y(n_603) );
AND2x2_ASAP7_75t_L g623 ( .A(n_521), .B(n_576), .Y(n_623) );
AND2x2_ASAP7_75t_L g667 ( .A(n_521), .B(n_536), .Y(n_667) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_546), .B(n_549), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_532), .B(n_534), .Y(n_531) );
AND2x2_ASAP7_75t_L g742 ( .A(n_532), .B(n_667), .Y(n_742) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_533), .A2(n_640), .B1(n_682), .B2(n_684), .Y(n_681) );
OR2x2_ASAP7_75t_L g688 ( .A(n_533), .B(n_603), .Y(n_688) );
OR2x2_ASAP7_75t_L g712 ( .A(n_533), .B(n_713), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_533), .B(n_632), .Y(n_725) );
AND2x2_ASAP7_75t_L g618 ( .A(n_534), .B(n_619), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g705 ( .A1(n_534), .A2(n_691), .B(n_706), .Y(n_705) );
AOI32xp33_ASAP7_75t_L g726 ( .A1(n_534), .A2(n_616), .A3(n_727), .B1(n_729), .B2(n_730), .Y(n_726) );
OR2x2_ASAP7_75t_L g737 ( .A(n_534), .B(n_738), .Y(n_737) );
CKINVDCx16_ASAP7_75t_R g534 ( .A(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g605 ( .A(n_535), .B(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_535), .B(n_619), .Y(n_684) );
BUFx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx4_ASAP7_75t_L g576 ( .A(n_536), .Y(n_576) );
AND2x2_ASAP7_75t_L g642 ( .A(n_536), .B(n_607), .Y(n_642) );
AND3x2_ASAP7_75t_L g651 ( .A(n_536), .B(n_547), .C(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g577 ( .A(n_548), .B(n_578), .Y(n_577) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_548), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_548), .B(n_576), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
AND2x2_ASAP7_75t_L g572 ( .A(n_550), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g612 ( .A(n_550), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g630 ( .A(n_550), .B(n_562), .Y(n_630) );
AND2x2_ASAP7_75t_L g648 ( .A(n_550), .B(n_552), .Y(n_648) );
OR2x2_ASAP7_75t_L g662 ( .A(n_550), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g708 ( .A(n_550), .B(n_636), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_551), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_562), .Y(n_551) );
AND2x2_ASAP7_75t_L g609 ( .A(n_552), .B(n_587), .Y(n_609) );
OR2x2_ASAP7_75t_L g663 ( .A(n_552), .B(n_587), .Y(n_663) );
AND2x2_ASAP7_75t_L g716 ( .A(n_552), .B(n_573), .Y(n_716) );
INVx2_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
BUFx2_ASAP7_75t_L g614 ( .A(n_553), .Y(n_614) );
AND2x2_ASAP7_75t_L g636 ( .A(n_553), .B(n_562), .Y(n_636) );
INVx2_ASAP7_75t_L g573 ( .A(n_562), .Y(n_573) );
INVx1_ASAP7_75t_L g593 ( .A(n_562), .Y(n_593) );
AOI211xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_574), .B(n_579), .C(n_591), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_572), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g735 ( .A(n_572), .Y(n_735) );
AND2x2_ASAP7_75t_L g613 ( .A(n_573), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_576), .B(n_577), .Y(n_585) );
INVx1_ASAP7_75t_L g670 ( .A(n_576), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_576), .B(n_597), .Y(n_694) );
AND2x2_ASAP7_75t_L g710 ( .A(n_576), .B(n_624), .Y(n_710) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_577), .B(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g601 ( .A(n_578), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_585), .B1(n_586), .B2(n_589), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_582), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_583), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g608 ( .A(n_584), .B(n_609), .Y(n_608) );
AOI221xp5_ASAP7_75t_SL g673 ( .A1(n_584), .A2(n_626), .B1(n_674), .B2(n_679), .C(n_681), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_584), .B(n_647), .Y(n_680) );
INVx1_ASAP7_75t_L g740 ( .A(n_586), .Y(n_740) );
BUFx3_ASAP7_75t_L g647 ( .A(n_587), .Y(n_647) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AOI21xp33_ASAP7_75t_SL g591 ( .A1(n_592), .A2(n_594), .B(n_595), .Y(n_591) );
INVx1_ASAP7_75t_L g656 ( .A(n_593), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_593), .B(n_647), .Y(n_700) );
INVx1_ASAP7_75t_L g657 ( .A(n_594), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g658 ( .A(n_594), .B(n_647), .Y(n_658) );
INVxp67_ASAP7_75t_L g678 ( .A(n_596), .Y(n_678) );
AND2x2_ASAP7_75t_L g619 ( .A(n_597), .B(n_620), .Y(n_619) );
O2A1O1Ixp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_604), .B(n_608), .C(n_610), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx1_ASAP7_75t_SL g633 ( .A(n_601), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_602), .B(n_633), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_602), .B(n_624), .Y(n_675) );
INVx2_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_605), .A2(n_611), .B1(n_615), .B2(n_617), .Y(n_610) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g626 ( .A(n_607), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g671 ( .A(n_607), .B(n_672), .Y(n_671) );
OAI21xp33_ASAP7_75t_L g674 ( .A1(n_609), .A2(n_675), .B(n_676), .Y(n_674) );
INVx1_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_613), .A2(n_622), .B1(n_625), .B2(n_626), .C(n_628), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_613), .B(n_647), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_613), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g729 ( .A(n_619), .Y(n_729) );
INVxp67_ASAP7_75t_L g652 ( .A(n_620), .Y(n_652) );
INVx1_ASAP7_75t_L g659 ( .A(n_622), .Y(n_659) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
AND2x2_ASAP7_75t_L g698 ( .A(n_623), .B(n_627), .Y(n_698) );
INVx1_ASAP7_75t_L g672 ( .A(n_627), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g702 ( .A(n_627), .B(n_642), .Y(n_702) );
OAI32xp33_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_631), .A3(n_633), .B1(n_634), .B2(n_635), .Y(n_628) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx2_ASAP7_75t_SL g641 ( .A(n_636), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_636), .B(n_668), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_636), .B(n_697), .Y(n_728) );
NAND2x1p5_ASAP7_75t_L g736 ( .A(n_636), .B(n_647), .Y(n_736) );
NAND5xp2_ASAP7_75t_L g637 ( .A(n_638), .B(n_660), .C(n_673), .D(n_685), .E(n_686), .Y(n_637) );
AOI221xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_642), .B1(n_643), .B2(n_645), .C(n_649), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp33_ASAP7_75t_SL g664 ( .A(n_644), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_647), .B(n_716), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_648), .A2(n_661), .B1(n_664), .B2(n_668), .Y(n_660) );
INVx2_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
OAI211xp5_ASAP7_75t_SL g655 ( .A1(n_651), .A2(n_656), .B(n_657), .C(n_658), .Y(n_655) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_SL g683 ( .A(n_663), .Y(n_683) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_672), .B(n_721), .Y(n_731) );
OR2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AOI222xp33_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_689), .B1(n_691), .B2(n_695), .C1(n_698), .C2(n_699), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
OAI221xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B1(n_705), .B2(n_707), .C(n_709), .Y(n_701) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
OAI21xp33_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_711), .B(n_714), .Y(n_709) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g721 ( .A(n_713), .Y(n_721) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
OAI221xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_720), .B1(n_722), .B2(n_724), .C(n_726), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
INVxp67_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
A2O1A1Ixp33_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_736), .B(n_737), .C(n_739), .Y(n_732) );
INVxp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OAI21xp33_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_741), .B(n_742), .Y(n_739) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx3_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
endmodule