module fake_ariane_661_n_8292 (n_83, n_8, n_56, n_60, n_64, n_90, n_38, n_47, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_33, n_19, n_40, n_106, n_12, n_53, n_21, n_66, n_71, n_24, n_7, n_96, n_49, n_20, n_100, n_17, n_50, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_72, n_105, n_44, n_30, n_82, n_31, n_42, n_57, n_70, n_10, n_85, n_6, n_48, n_94, n_101, n_4, n_2, n_32, n_37, n_58, n_65, n_9, n_45, n_11, n_52, n_73, n_77, n_15, n_93, n_23, n_61, n_102, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_35, n_54, n_25, n_8292);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_90;
input n_38;
input n_47;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_33;
input n_19;
input n_40;
input n_106;
input n_12;
input n_53;
input n_21;
input n_66;
input n_71;
input n_24;
input n_7;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_72;
input n_105;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_70;
input n_10;
input n_85;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_9;
input n_45;
input n_11;
input n_52;
input n_73;
input n_77;
input n_15;
input n_93;
input n_23;
input n_61;
input n_102;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_35;
input n_54;
input n_25;

output n_8292;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_7329;
wire n_4030;
wire n_7029;
wire n_6790;
wire n_4770;
wire n_8165;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_6603;
wire n_2679;
wire n_6557;
wire n_5402;
wire n_6581;
wire n_2182;
wire n_5553;
wire n_6002;
wire n_7277;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_5717;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_8139;
wire n_416;
wire n_4962;
wire n_1430;
wire n_7832;
wire n_2002;
wire n_1238;
wire n_2729;
wire n_4302;
wire n_5791;
wire n_7127;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_864;
wire n_5302;
wire n_1096;
wire n_1379;
wire n_2376;
wire n_7922;
wire n_7805;
wire n_2790;
wire n_7542;
wire n_2207;
wire n_7053;
wire n_5712;
wire n_3954;
wire n_6297;
wire n_4982;
wire n_2042;
wire n_462;
wire n_1131;
wire n_8037;
wire n_5479;
wire n_2646;
wire n_8257;
wire n_737;
wire n_2653;
wire n_4610;
wire n_6058;
wire n_232;
wire n_3115;
wire n_4028;
wire n_5263;
wire n_5565;
wire n_6358;
wire n_6293;
wire n_2482;
wire n_1682;
wire n_7001;
wire n_958;
wire n_6129;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_5590;
wire n_2621;
wire n_6524;
wire n_146;
wire n_4853;
wire n_338;
wire n_1909;
wire n_5229;
wire n_6313;
wire n_7464;
wire n_4260;
wire n_903;
wire n_7626;
wire n_3348;
wire n_239;
wire n_3261;
wire n_1761;
wire n_7965;
wire n_7368;
wire n_1690;
wire n_2807;
wire n_6664;
wire n_7562;
wire n_7534;
wire n_1018;
wire n_7428;
wire n_4512;
wire n_6190;
wire n_4132;
wire n_1364;
wire n_7373;
wire n_2390;
wire n_8068;
wire n_6891;
wire n_4500;
wire n_625;
wire n_2322;
wire n_1107;
wire n_331;
wire n_559;
wire n_2663;
wire n_8097;
wire n_5481;
wire n_6539;
wire n_495;
wire n_8114;
wire n_4824;
wire n_7467;
wire n_350;
wire n_8126;
wire n_381;
wire n_5340;
wire n_3545;
wire n_6797;
wire n_7392;
wire n_1428;
wire n_1284;
wire n_4741;
wire n_1241;
wire n_7526;
wire n_561;
wire n_4143;
wire n_4273;
wire n_507;
wire n_901;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_1519;
wire n_7338;
wire n_5896;
wire n_4567;
wire n_786;
wire n_5833;
wire n_6249;
wire n_6887;
wire n_6253;
wire n_6128;
wire n_3552;
wire n_2950;
wire n_6197;
wire n_7200;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_5589;
wire n_3015;
wire n_5744;
wire n_3870;
wire n_6808;
wire n_3749;
wire n_1676;
wire n_1085;
wire n_277;
wire n_5691;
wire n_7937;
wire n_3482;
wire n_7490;
wire n_6295;
wire n_5403;
wire n_823;
wire n_1900;
wire n_620;
wire n_6096;
wire n_4268;
wire n_6338;
wire n_587;
wire n_863;
wire n_6992;
wire n_303;
wire n_3960;
wire n_2433;
wire n_352;
wire n_899;
wire n_3975;
wire n_8035;
wire n_5830;
wire n_365;
wire n_2004;
wire n_4018;
wire n_1495;
wire n_334;
wire n_192;
wire n_3325;
wire n_6681;
wire n_661;
wire n_4227;
wire n_5158;
wire n_5152;
wire n_533;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_1924;
wire n_6542;
wire n_1811;
wire n_6161;
wire n_3612;
wire n_273;
wire n_4505;
wire n_6452;
wire n_1840;
wire n_5247;
wire n_5464;
wire n_7306;
wire n_4476;
wire n_6740;
wire n_6978;
wire n_579;
wire n_7507;
wire n_844;
wire n_1267;
wire n_8176;
wire n_2956;
wire n_5210;
wire n_7215;
wire n_149;
wire n_1213;
wire n_2382;
wire n_7379;
wire n_7441;
wire n_237;
wire n_780;
wire n_5292;
wire n_1918;
wire n_7438;
wire n_4119;
wire n_4443;
wire n_4000;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_6136;
wire n_1140;
wire n_3458;
wire n_570;
wire n_5843;
wire n_7874;
wire n_7108;
wire n_3511;
wire n_2077;
wire n_1121;
wire n_490;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_575;
wire n_7695;
wire n_6156;
wire n_1216;
wire n_4908;
wire n_8098;
wire n_3754;
wire n_8204;
wire n_5060;
wire n_7162;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_7331;
wire n_5913;
wire n_4530;
wire n_1432;
wire n_2245;
wire n_5614;
wire n_5391;
wire n_5452;
wire n_3359;
wire n_7944;
wire n_3841;
wire n_5249;
wire n_249;
wire n_851;
wire n_123;
wire n_444;
wire n_3900;
wire n_3413;
wire n_7850;
wire n_5076;
wire n_3539;
wire n_5757;
wire n_6872;
wire n_6644;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_930;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_5046;
wire n_7607;
wire n_7642;
wire n_1386;
wire n_6236;
wire n_7104;
wire n_8147;
wire n_3506;
wire n_4827;
wire n_6801;
wire n_1842;
wire n_4993;
wire n_7397;
wire n_3678;
wire n_7205;
wire n_366;
wire n_2791;
wire n_1661;
wire n_555;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_6563;
wire n_5968;
wire n_992;
wire n_966;
wire n_3549;
wire n_3914;
wire n_6398;
wire n_5586;
wire n_7461;
wire n_1692;
wire n_2611;
wire n_8075;
wire n_5468;
wire n_3029;
wire n_4745;
wire n_7638;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_5971;
wire n_6319;
wire n_7224;
wire n_6966;
wire n_5056;
wire n_1178;
wire n_2015;
wire n_7259;
wire n_7838;
wire n_5984;
wire n_5204;
wire n_6724;
wire n_6705;
wire n_2877;
wire n_7307;
wire n_6776;
wire n_203;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_150;
wire n_2930;
wire n_7840;
wire n_2745;
wire n_2087;
wire n_619;
wire n_2161;
wire n_746;
wire n_6624;
wire n_1357;
wire n_7888;
wire n_292;
wire n_6710;
wire n_1787;
wire n_6883;
wire n_8108;
wire n_1389;
wire n_8158;
wire n_3172;
wire n_2659;
wire n_4033;
wire n_3747;
wire n_6553;
wire n_4905;
wire n_4508;
wire n_5897;
wire n_4045;
wire n_6261;
wire n_3651;
wire n_1812;
wire n_6659;
wire n_4894;
wire n_428;
wire n_7351;
wire n_3614;
wire n_7256;
wire n_959;
wire n_2257;
wire n_1101;
wire n_1343;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_6893;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_5778;
wire n_7021;
wire n_5179;
wire n_2435;
wire n_6337;
wire n_5680;
wire n_1932;
wire n_6210;
wire n_7583;
wire n_1780;
wire n_2825;
wire n_5685;
wire n_5974;
wire n_5723;
wire n_542;
wire n_5922;
wire n_6378;
wire n_5549;
wire n_1087;
wire n_632;
wire n_2388;
wire n_2273;
wire n_8130;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_7488;
wire n_3700;
wire n_7690;
wire n_4307;
wire n_2795;
wire n_6044;
wire n_1841;
wire n_1680;
wire n_6206;
wire n_7893;
wire n_2954;
wire n_382;
wire n_489;
wire n_4438;
wire n_6538;
wire n_7966;
wire n_251;
wire n_974;
wire n_506;
wire n_3814;
wire n_6996;
wire n_5831;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_7599;
wire n_7231;
wire n_4195;
wire n_7007;
wire n_7717;
wire n_6579;
wire n_5091;
wire n_4866;
wire n_7230;
wire n_1447;
wire n_1220;
wire n_7900;
wire n_2019;
wire n_5708;
wire n_8123;
wire n_698;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_124;
wire n_5454;
wire n_307;
wire n_1209;
wire n_4254;
wire n_646;
wire n_3438;
wire n_8220;
wire n_404;
wire n_2625;
wire n_5373;
wire n_7403;
wire n_1578;
wire n_6665;
wire n_3147;
wire n_299;
wire n_3661;
wire n_7168;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_133;
wire n_1029;
wire n_2649;
wire n_6033;
wire n_6461;
wire n_1247;
wire n_6860;
wire n_522;
wire n_1568;
wire n_2919;
wire n_7322;
wire n_6060;
wire n_3108;
wire n_5983;
wire n_5788;
wire n_367;
wire n_6709;
wire n_2632;
wire n_5557;
wire n_6914;
wire n_4314;
wire n_2980;
wire n_5951;
wire n_1728;
wire n_5647;
wire n_4315;
wire n_6117;
wire n_7287;
wire n_7789;
wire n_3239;
wire n_2631;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_424;
wire n_4857;
wire n_1651;
wire n_3087;
wire n_6009;
wire n_7221;
wire n_5523;
wire n_4637;
wire n_2697;
wire n_1263;
wire n_1817;
wire n_8243;
wire n_3704;
wire n_7963;
wire n_6382;
wire n_670;
wire n_2677;
wire n_4296;
wire n_379;
wire n_138;
wire n_162;
wire n_2483;
wire n_7938;
wire n_5088;
wire n_6615;
wire n_441;
wire n_7294;
wire n_6192;
wire n_5773;
wire n_7414;
wire n_1032;
wire n_1592;
wire n_5392;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_3589;
wire n_6418;
wire n_1743;
wire n_207;
wire n_720;
wire n_6263;
wire n_1943;
wire n_6731;
wire n_8156;
wire n_5138;
wire n_4588;
wire n_6048;
wire n_7185;
wire n_194;
wire n_5149;
wire n_1163;
wire n_3054;
wire n_5280;
wire n_4970;
wire n_6234;
wire n_4153;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_7141;
wire n_2373;
wire n_3881;
wire n_6224;
wire n_5089;
wire n_5775;
wire n_2099;
wire n_3759;
wire n_3323;
wire n_4643;
wire n_6142;
wire n_2617;
wire n_6119;
wire n_6619;
wire n_808;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_1439;
wire n_6759;
wire n_6903;
wire n_3466;
wire n_7416;
wire n_2074;
wire n_5031;
wire n_6768;
wire n_1665;
wire n_7092;
wire n_7233;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_5082;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_5230;
wire n_4555;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_7191;
wire n_2117;
wire n_6189;
wire n_1053;
wire n_5796;
wire n_5296;
wire n_5398;
wire n_1906;
wire n_6761;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_1828;
wire n_1304;
wire n_7202;
wire n_3335;
wire n_5960;
wire n_3007;
wire n_2267;
wire n_7445;
wire n_5858;
wire n_5985;
wire n_604;
wire n_478;
wire n_1349;
wire n_1061;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_7868;
wire n_3370;
wire n_874;
wire n_7654;
wire n_3949;
wire n_2286;
wire n_5192;
wire n_4247;
wire n_707;
wire n_5051;
wire n_5336;
wire n_129;
wire n_126;
wire n_3036;
wire n_2783;
wire n_4583;
wire n_6366;
wire n_1015;
wire n_1162;
wire n_6304;
wire n_4292;
wire n_2118;
wire n_688;
wire n_7176;
wire n_636;
wire n_1490;
wire n_6074;
wire n_7547;
wire n_5552;
wire n_442;
wire n_3764;
wire n_1553;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_1086;
wire n_3025;
wire n_3051;
wire n_986;
wire n_1104;
wire n_2802;
wire n_8030;
wire n_887;
wire n_2125;
wire n_1156;
wire n_4974;
wire n_5123;
wire n_6689;
wire n_2861;
wire n_8245;
wire n_7942;
wire n_4344;
wire n_5242;
wire n_3130;
wire n_1188;
wire n_1498;
wire n_7527;
wire n_4856;
wire n_2618;
wire n_7948;
wire n_7096;
wire n_4216;
wire n_957;
wire n_1242;
wire n_2707;
wire n_5596;
wire n_6482;
wire n_8106;
wire n_2849;
wire n_1489;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_6335;
wire n_5742;
wire n_5127;
wire n_4313;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_1119;
wire n_3713;
wire n_6229;
wire n_1863;
wire n_5933;
wire n_5536;
wire n_4798;
wire n_1500;
wire n_616;
wire n_7293;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_1189;
wire n_5810;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_7144;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_4991;
wire n_7316;
wire n_7508;
wire n_3070;
wire n_1005;
wire n_5818;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_2452;
wire n_4182;
wire n_2827;
wire n_7869;
wire n_3214;
wire n_8166;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5539;
wire n_5009;
wire n_3710;
wire n_1844;
wire n_6943;
wire n_1957;
wire n_1953;
wire n_1219;
wire n_710;
wire n_6631;
wire n_5889;
wire n_7151;
wire n_3944;
wire n_7762;
wire n_5632;
wire n_4729;
wire n_8002;
wire n_6728;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_5613;
wire n_7472;
wire n_4800;
wire n_1373;
wire n_7075;
wire n_1540;
wire n_5427;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_6770;
wire n_5450;
wire n_7611;
wire n_7796;
wire n_6508;
wire n_832;
wire n_7989;
wire n_8047;
wire n_744;
wire n_2821;
wire n_3696;
wire n_7936;
wire n_215;
wire n_1331;
wire n_4781;
wire n_6031;
wire n_1529;
wire n_3531;
wire n_5124;
wire n_655;
wire n_4237;
wire n_5297;
wire n_4828;
wire n_3333;
wire n_4652;
wire n_4114;
wire n_7105;
wire n_7013;
wire n_7655;
wire n_1007;
wire n_1580;
wire n_3135;
wire n_4925;
wire n_5719;
wire n_7254;
wire n_2448;
wire n_2211;
wire n_951;
wire n_8039;
wire n_8193;
wire n_7546;
wire n_5904;
wire n_6628;
wire n_5318;
wire n_5374;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_6456;
wire n_722;
wire n_7407;
wire n_3277;
wire n_4863;
wire n_1766;
wire n_5463;
wire n_1338;
wire n_2978;
wire n_6328;
wire n_6929;
wire n_4859;
wire n_4568;
wire n_3617;
wire n_6012;
wire n_704;
wire n_2958;
wire n_7481;
wire n_1044;
wire n_1714;
wire n_4429;
wire n_6484;
wire n_5435;
wire n_3340;
wire n_5053;
wire n_7182;
wire n_5476;
wire n_5483;
wire n_7605;
wire n_8090;
wire n_1243;
wire n_5511;
wire n_3486;
wire n_6639;
wire n_358;
wire n_608;
wire n_2457;
wire n_2992;
wire n_6124;
wire n_317;
wire n_3197;
wire n_7423;
wire n_3256;
wire n_1878;
wire n_7375;
wire n_7076;
wire n_7689;
wire n_6344;
wire n_8189;
wire n_266;
wire n_7736;
wire n_6435;
wire n_3646;
wire n_5829;
wire n_2520;
wire n_7419;
wire n_811;
wire n_6600;
wire n_7010;
wire n_791;
wire n_5881;
wire n_3864;
wire n_4694;
wire n_8192;
wire n_1025;
wire n_4664;
wire n_6201;
wire n_3450;
wire n_687;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_480;
wire n_7918;
wire n_642;
wire n_1406;
wire n_6555;
wire n_5073;
wire n_4306;
wire n_6360;
wire n_6735;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_6803;
wire n_4288;
wire n_3452;
wire n_474;
wire n_4098;
wire n_2691;
wire n_5894;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_695;
wire n_2991;
wire n_5419;
wire n_386;
wire n_1596;
wire n_4289;
wire n_4972;
wire n_197;
wire n_2723;
wire n_1476;
wire n_6036;
wire n_7346;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_678;
wire n_651;
wire n_2850;
wire n_1874;
wire n_5077;
wire n_6102;
wire n_3780;
wire n_1657;
wire n_6650;
wire n_6573;
wire n_6904;
wire n_3753;
wire n_6329;
wire n_7385;
wire n_1488;
wire n_6244;
wire n_4846;
wire n_1330;
wire n_906;
wire n_6204;
wire n_2295;
wire n_5225;
wire n_283;
wire n_7295;
wire n_4076;
wire n_7824;
wire n_7148;
wire n_3142;
wire n_7169;
wire n_3129;
wire n_374;
wire n_3843;
wire n_3495;
wire n_6756;
wire n_4805;
wire n_2606;
wire n_7600;
wire n_2386;
wire n_5826;
wire n_4822;
wire n_6946;
wire n_7947;
wire n_5931;
wire n_8146;
wire n_1829;
wire n_4635;
wire n_7847;
wire n_8154;
wire n_1450;
wire n_5532;
wire n_7311;
wire n_3740;
wire n_6804;
wire n_5441;
wire n_6179;
wire n_2417;
wire n_6059;
wire n_1815;
wire n_7039;
wire n_8027;
wire n_7807;
wire n_1493;
wire n_2911;
wire n_515;
wire n_8063;
wire n_3313;
wire n_2354;
wire n_6427;
wire n_4281;
wire n_3945;
wire n_5994;
wire n_3726;
wire n_4419;
wire n_5405;
wire n_7660;
wire n_1256;
wire n_5365;
wire n_3560;
wire n_3345;
wire n_5772;
wire n_6442;
wire n_8241;
wire n_140;
wire n_6188;
wire n_3421;
wire n_1448;
wire n_1009;
wire n_230;
wire n_3548;
wire n_4906;
wire n_6846;
wire n_4630;
wire n_8261;
wire n_6840;
wire n_142;
wire n_6645;
wire n_4829;
wire n_6749;
wire n_6915;
wire n_7831;
wire n_8138;
wire n_2612;
wire n_5259;
wire n_3236;
wire n_1995;
wire n_7455;
wire n_8273;
wire n_1397;
wire n_5921;
wire n_6247;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_4966;
wire n_2250;
wire n_8235;
wire n_1117;
wire n_6104;
wire n_3321;
wire n_1303;
wire n_4188;
wire n_2001;
wire n_7509;
wire n_6205;
wire n_2506;
wire n_2413;
wire n_4825;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_2626;
wire n_7497;
wire n_7315;
wire n_2892;
wire n_6939;
wire n_2605;
wire n_7887;
wire n_2804;
wire n_5884;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_5728;
wire n_1035;
wire n_3475;
wire n_4878;
wire n_2070;
wire n_426;
wire n_6706;
wire n_7431;
wire n_8140;
wire n_398;
wire n_3842;
wire n_1367;
wire n_4202;
wire n_6909;
wire n_2044;
wire n_5679;
wire n_6487;
wire n_166;
wire n_8117;
wire n_3886;
wire n_825;
wire n_732;
wire n_2619;
wire n_7521;
wire n_1192;
wire n_5141;
wire n_3098;
wire n_6627;
wire n_4503;
wire n_8129;
wire n_1291;
wire n_7253;
wire n_5208;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_7569;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_7452;
wire n_6551;
wire n_3386;
wire n_400;
wire n_7972;
wire n_7505;
wire n_3921;
wire n_282;
wire n_467;
wire n_2177;
wire n_6516;
wire n_2766;
wire n_7524;
wire n_4196;
wire n_1197;
wire n_7318;
wire n_2613;
wire n_7411;
wire n_7326;
wire n_5667;
wire n_168;
wire n_1517;
wire n_2647;
wire n_8005;
wire n_5508;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_5879;
wire n_1671;
wire n_6500;
wire n_5027;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_3380;
wire n_5688;
wire n_2826;
wire n_5825;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_8221;
wire n_7573;
wire n_6630;
wire n_5629;
wire n_5759;
wire n_2411;
wire n_4631;
wire n_8191;
wire n_6798;
wire n_5999;
wire n_1504;
wire n_2110;
wire n_7498;
wire n_7895;
wire n_6421;
wire n_5377;
wire n_6180;
wire n_8225;
wire n_3822;
wire n_889;
wire n_7453;
wire n_4355;
wire n_3818;
wire n_7932;
wire n_7890;
wire n_5599;
wire n_3587;
wire n_2608;
wire n_6004;
wire n_1948;
wire n_6652;
wire n_7183;
wire n_4155;
wire n_810;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_6275;
wire n_6395;
wire n_3497;
wire n_6403;
wire n_4542;
wire n_5451;
wire n_6578;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_6350;
wire n_5460;
wire n_4685;
wire n_565;
wire n_3927;
wire n_6141;
wire n_2068;
wire n_3595;
wire n_6875;
wire n_7189;
wire n_1194;
wire n_4060;
wire n_1647;
wire n_6194;
wire n_1454;
wire n_2459;
wire n_941;
wire n_3396;
wire n_5517;
wire n_5807;
wire n_5426;
wire n_6475;
wire n_4093;
wire n_452;
wire n_5693;
wire n_5695;
wire n_4123;
wire n_4294;
wire n_1521;
wire n_1940;
wire n_3683;
wire n_6502;
wire n_6944;
wire n_4452;
wire n_284;
wire n_3887;
wire n_3195;
wire n_5587;
wire n_4722;
wire n_6318;
wire n_8163;
wire n_6805;
wire n_3048;
wire n_3339;
wire n_4126;
wire n_4164;
wire n_7240;
wire n_5030;
wire n_409;
wire n_2963;
wire n_5674;
wire n_2561;
wire n_7499;
wire n_1056;
wire n_526;
wire n_5584;
wire n_674;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_6075;
wire n_6559;
wire n_4088;
wire n_2669;
wire n_3911;
wire n_6068;
wire n_3802;
wire n_4366;
wire n_1584;
wire n_6541;
wire n_6248;
wire n_848;
wire n_5125;
wire n_4922;
wire n_6066;
wire n_6080;
wire n_629;
wire n_4733;
wire n_7927;
wire n_161;
wire n_1814;
wire n_7219;
wire n_2441;
wire n_8081;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_216;
wire n_6150;
wire n_6638;
wire n_7063;
wire n_7402;
wire n_6351;
wire n_4509;
wire n_4935;
wire n_2073;
wire n_7382;
wire n_4004;
wire n_5238;
wire n_750;
wire n_834;
wire n_3630;
wire n_1612;
wire n_800;
wire n_1910;
wire n_5906;
wire n_7767;
wire n_2189;
wire n_5732;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_2602;
wire n_5780;
wire n_724;
wire n_2931;
wire n_3433;
wire n_8284;
wire n_5556;
wire n_6006;
wire n_3597;
wire n_6474;
wire n_5743;
wire n_6481;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_5633;
wire n_7510;
wire n_3786;
wire n_875;
wire n_6022;
wire n_6991;
wire n_2828;
wire n_7434;
wire n_1626;
wire n_5950;
wire n_1335;
wire n_1715;
wire n_4204;
wire n_7691;
wire n_296;
wire n_3553;
wire n_5323;
wire n_7745;
wire n_6744;
wire n_3645;
wire n_793;
wire n_5705;
wire n_6927;
wire n_7335;
wire n_132;
wire n_4996;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_7735;
wire n_6116;
wire n_8074;
wire n_494;
wire n_3550;
wire n_7956;
wire n_5510;
wire n_7495;
wire n_7651;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1805;
wire n_4068;
wire n_5440;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_2443;
wire n_3610;
wire n_185;
wire n_5011;
wire n_6757;
wire n_7536;
wire n_1554;
wire n_3279;
wire n_5513;
wire n_5875;
wire n_972;
wire n_7734;
wire n_4262;
wire n_2923;
wire n_164;
wire n_2843;
wire n_3714;
wire n_184;
wire n_7671;
wire n_4832;
wire n_8033;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_6485;
wire n_5848;
wire n_118;
wire n_1679;
wire n_5834;
wire n_7926;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_5784;
wire n_3125;
wire n_5128;
wire n_2356;
wire n_5618;
wire n_6495;
wire n_7528;
wire n_6209;
wire n_4672;
wire n_8094;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_783;
wire n_4053;
wire n_1127;
wire n_7413;
wire n_7993;
wire n_7821;
wire n_160;
wire n_7620;
wire n_119;
wire n_1008;
wire n_3963;
wire n_581;
wire n_3091;
wire n_6274;
wire n_1024;
wire n_176;
wire n_5157;
wire n_4496;
wire n_2518;
wire n_936;
wire n_4596;
wire n_5178;
wire n_3105;
wire n_6237;
wire n_1525;
wire n_4628;
wire n_6802;
wire n_7343;
wire n_5982;
wire n_1775;
wire n_908;
wire n_1036;
wire n_7109;
wire n_8028;
wire n_341;
wire n_4083;
wire n_1270;
wire n_109;
wire n_1272;
wire n_549;
wire n_2794;
wire n_6155;
wire n_2901;
wire n_7506;
wire n_3940;
wire n_6809;
wire n_6099;
wire n_3225;
wire n_3621;
wire n_5529;
wire n_244;
wire n_7561;
wire n_3473;
wire n_6349;
wire n_3680;
wire n_6716;
wire n_3565;
wire n_7885;
wire n_6905;
wire n_7722;
wire n_5388;
wire n_7470;
wire n_5824;
wire n_8025;
wire n_5354;
wire n_2453;
wire n_7898;
wire n_3331;
wire n_1788;
wire n_6203;
wire n_2138;
wire n_6407;
wire n_3040;
wire n_4230;
wire n_6899;
wire n_7980;
wire n_7817;
wire n_6413;
wire n_445;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_7070;
wire n_2000;
wire n_5276;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_3211;
wire n_7299;
wire n_917;
wire n_5196;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_8029;
wire n_2215;
wire n_3847;
wire n_6960;
wire n_4073;
wire n_1261;
wire n_7249;
wire n_5763;
wire n_3633;
wire n_857;
wire n_363;
wire n_6061;
wire n_1235;
wire n_2584;
wire n_4001;
wire n_1462;
wire n_5701;
wire n_7002;
wire n_1064;
wire n_633;
wire n_1446;
wire n_1701;
wire n_6273;
wire n_7094;
wire n_7396;
wire n_3111;
wire n_731;
wire n_1813;
wire n_315;
wire n_2997;
wire n_7018;
wire n_1573;
wire n_6746;
wire n_3258;
wire n_758;
wire n_3691;
wire n_2252;
wire n_6174;
wire n_6545;
wire n_7773;
wire n_6763;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_7297;
wire n_784;
wire n_4339;
wire n_5907;
wire n_7730;
wire n_8134;
wire n_6013;
wire n_6182;
wire n_6754;
wire n_4690;
wire n_2987;
wire n_6279;
wire n_1473;
wire n_1076;
wire n_1348;
wire n_5895;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_2103;
wire n_4169;
wire n_4024;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_7637;
wire n_2522;
wire n_3632;
wire n_309;
wire n_1344;
wire n_115;
wire n_485;
wire n_4064;
wire n_6131;
wire n_3351;
wire n_5478;
wire n_435;
wire n_6113;
wire n_1141;
wire n_3457;
wire n_6477;
wire n_5384;
wire n_7486;
wire n_840;
wire n_2324;
wire n_6575;
wire n_5283;
wire n_3454;
wire n_5961;
wire n_7544;
wire n_2139;
wire n_7613;
wire n_7995;
wire n_8113;
wire n_2521;
wire n_5686;
wire n_6391;
wire n_2740;
wire n_1991;
wire n_7140;
wire n_614;
wire n_4066;
wire n_6252;
wire n_6426;
wire n_4681;
wire n_8253;
wire n_3303;
wire n_7910;
wire n_6592;
wire n_4414;
wire n_2541;
wire n_5094;
wire n_3232;
wire n_1113;
wire n_248;
wire n_7741;
wire n_3768;
wire n_4295;
wire n_1615;
wire n_4100;
wire n_228;
wire n_6668;
wire n_1265;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_4087;
wire n_8232;
wire n_1409;
wire n_1684;
wire n_1148;
wire n_1588;
wire n_1673;
wire n_4473;
wire n_4619;
wire n_6670;
wire n_5371;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_7679;
wire n_3018;
wire n_7698;
wire n_1875;
wire n_6962;
wire n_2429;
wire n_6779;
wire n_5286;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_1039;
wire n_5676;
wire n_5949;
wire n_5040;
wire n_6901;
wire n_1150;
wire n_7800;
wire n_4266;
wire n_6336;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_6503;
wire n_7835;
wire n_1136;
wire n_458;
wire n_1190;
wire n_6049;
wire n_5885;
wire n_3628;
wire n_7100;
wire n_4777;
wire n_7243;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_7415;
wire n_5399;
wire n_658;
wire n_362;
wire n_2846;
wire n_3371;
wire n_4918;
wire n_5856;
wire n_8016;
wire n_3872;
wire n_5760;
wire n_7747;
wire n_4415;
wire n_5110;
wire n_1964;
wire n_3659;
wire n_7552;
wire n_3928;
wire n_1777;
wire n_3366;
wire n_6998;
wire n_7395;
wire n_5844;
wire n_6298;
wire n_8132;
wire n_7650;
wire n_3441;
wire n_199;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_7535;
wire n_708;
wire n_6609;
wire n_2545;
wire n_2513;
wire n_7635;
wire n_4408;
wire n_2115;
wire n_8259;
wire n_2017;
wire n_1810;
wire n_1347;
wire n_4976;
wire n_860;
wire n_6525;
wire n_3555;
wire n_5938;
wire n_7274;
wire n_3534;
wire n_450;
wire n_4548;
wire n_7819;
wire n_2670;
wire n_6494;
wire n_3556;
wire n_896;
wire n_4574;
wire n_8160;
wire n_2644;
wire n_6132;
wire n_4557;
wire n_3071;
wire n_1698;
wire n_1337;
wire n_774;
wire n_2148;
wire n_5548;
wire n_7788;
wire n_6974;
wire n_1168;
wire n_4663;
wire n_219;
wire n_5840;
wire n_6882;
wire n_3296;
wire n_3794;
wire n_3762;
wire n_4624;
wire n_656;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_6498;
wire n_6562;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_8229;
wire n_415;
wire n_4686;
wire n_2384;
wire n_7794;
wire n_1705;
wire n_768;
wire n_3707;
wire n_1091;
wire n_3895;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_5917;
wire n_6965;
wire n_2058;
wire n_3231;
wire n_1846;
wire n_7630;
wire n_4161;
wire n_110;
wire n_304;
wire n_6168;
wire n_5304;
wire n_5437;
wire n_6963;
wire n_6951;
wire n_1581;
wire n_946;
wire n_757;
wire n_5355;
wire n_2047;
wire n_3058;
wire n_375;
wire n_113;
wire n_1655;
wire n_3398;
wire n_1146;
wire n_3709;
wire n_6284;
wire n_998;
wire n_3592;
wire n_5321;
wire n_7454;
wire n_2536;
wire n_1604;
wire n_3399;
wire n_4772;
wire n_6931;
wire n_6521;
wire n_5915;
wire n_7276;
wire n_174;
wire n_6379;
wire n_1368;
wire n_963;
wire n_7085;
wire n_6306;
wire n_4120;
wire n_925;
wire n_7753;
wire n_6834;
wire n_2880;
wire n_1313;
wire n_1001;
wire n_3722;
wire n_4716;
wire n_1115;
wire n_4654;
wire n_1339;
wire n_1051;
wire n_5116;
wire n_3771;
wire n_7225;
wire n_719;
wire n_7541;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_7913;
wire n_8020;
wire n_7946;
wire n_1010;
wire n_2830;
wire n_5500;
wire n_4622;
wire n_4757;
wire n_803;
wire n_1871;
wire n_6471;
wire n_6949;
wire n_5669;
wire n_5672;
wire n_4016;
wire n_3334;
wire n_5621;
wire n_6760;
wire n_2940;
wire n_548;
wire n_3427;
wire n_3162;
wire n_5966;
wire n_5569;
wire n_4591;
wire n_5515;
wire n_6589;
wire n_3083;
wire n_4570;
wire n_7014;
wire n_2491;
wire n_7920;
wire n_1931;
wire n_5559;
wire n_2259;
wire n_5337;
wire n_849;
wire n_5059;
wire n_4655;
wire n_7459;
wire n_1820;
wire n_7841;
wire n_7160;
wire n_7324;
wire n_8205;
wire n_6046;
wire n_7054;
wire n_1233;
wire n_4493;
wire n_6055;
wire n_7161;
wire n_1808;
wire n_6364;
wire n_6091;
wire n_6348;
wire n_1635;
wire n_1704;
wire n_4896;
wire n_8041;
wire n_4851;
wire n_6848;
wire n_2479;
wire n_886;
wire n_7837;
wire n_359;
wire n_6788;
wire n_1308;
wire n_6144;
wire n_1451;
wire n_1487;
wire n_675;
wire n_5528;
wire n_7806;
wire n_5605;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_6896;
wire n_2484;
wire n_5753;
wire n_8076;
wire n_5358;
wire n_1469;
wire n_4901;
wire n_3480;
wire n_1355;
wire n_7201;
wire n_4213;
wire n_4127;
wire n_6221;
wire n_2500;
wire n_7676;
wire n_8177;
wire n_2334;
wire n_5467;
wire n_7241;
wire n_1169;
wire n_789;
wire n_3181;
wire n_5493;
wire n_1916;
wire n_6285;
wire n_610;
wire n_7644;
wire n_4602;
wire n_1713;
wire n_7816;
wire n_1436;
wire n_2818;
wire n_4900;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_3745;
wire n_6748;
wire n_7430;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_1515;
wire n_817;
wire n_5901;
wire n_1566;
wire n_2837;
wire n_717;
wire n_952;
wire n_2446;
wire n_6582;
wire n_4116;
wire n_7724;
wire n_5360;
wire n_7269;
wire n_7047;
wire n_2671;
wire n_2702;
wire n_6937;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_1138;
wire n_214;
wire n_4103;
wire n_2529;
wire n_8101;
wire n_2374;
wire n_5439;
wire n_6115;
wire n_1225;
wire n_3154;
wire n_137;
wire n_1366;
wire n_3938;
wire n_2278;
wire n_6272;
wire n_7067;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_4416;
wire n_7879;
wire n_6607;
wire n_4439;
wire n_520;
wire n_870;
wire n_4985;
wire n_3382;
wire n_7117;
wire n_3930;
wire n_3808;
wire n_5471;
wire n_2248;
wire n_813;
wire n_4660;
wire n_3081;
wire n_6446;
wire n_5497;
wire n_5519;
wire n_6071;
wire n_995;
wire n_2579;
wire n_1961;
wire n_1535;
wire n_6849;
wire n_2960;
wire n_3270;
wire n_871;
wire n_6807;
wire n_2844;
wire n_8197;
wire n_402;
wire n_1979;
wire n_6616;
wire n_6719;
wire n_829;
wire n_4814;
wire n_8019;
wire n_339;
wire n_6178;
wire n_6677;
wire n_2221;
wire n_7875;
wire n_5502;
wire n_8248;
wire n_1283;
wire n_7550;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_7302;
wire n_2781;
wire n_6191;
wire n_2442;
wire n_7238;
wire n_6862;
wire n_3657;
wire n_5706;
wire n_2634;
wire n_2746;
wire n_7292;
wire n_242;
wire n_645;
wire n_7804;
wire n_5098;
wire n_721;
wire n_1084;
wire n_6000;
wire n_6774;
wire n_6443;
wire n_1276;
wire n_8263;
wire n_5145;
wire n_6072;
wire n_2878;
wire n_7248;
wire n_3830;
wire n_3252;
wire n_6647;
wire n_8040;
wire n_5466;
wire n_1528;
wire n_6941;
wire n_7239;
wire n_6552;
wire n_7826;
wire n_3315;
wire n_6094;
wire n_3523;
wire n_8102;
wire n_3999;
wire n_518;
wire n_8196;
wire n_7112;
wire n_3420;
wire n_3859;
wire n_868;
wire n_5213;
wire n_3474;
wire n_5738;
wire n_2458;
wire n_7971;
wire n_5592;
wire n_5620;
wire n_3150;
wire n_5491;
wire n_1542;
wire n_4831;
wire n_4782;
wire n_1539;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_5953;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_5703;
wire n_6886;
wire n_7078;
wire n_1636;
wire n_4597;
wire n_8152;
wire n_8269;
wire n_4546;
wire n_5187;
wire n_7006;
wire n_4031;
wire n_5119;
wire n_1254;
wire n_4147;
wire n_1703;
wire n_3073;
wire n_6531;
wire n_3571;
wire n_238;
wire n_4576;
wire n_7577;
wire n_7354;
wire n_6098;
wire n_5995;
wire n_3297;
wire n_8144;
wire n_5148;
wire n_3003;
wire n_6726;
wire n_6983;
wire n_7513;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_7812;
wire n_5330;
wire n_6935;
wire n_1560;
wire n_2899;
wire n_6984;
wire n_6778;
wire n_8058;
wire n_6897;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5526;
wire n_5202;
wire n_3817;
wire n_6345;
wire n_6386;
wire n_2722;
wire n_3728;
wire n_6596;
wire n_612;
wire n_333;
wire n_5107;
wire n_7165;
wire n_512;
wire n_4680;
wire n_5067;
wire n_6830;
wire n_1012;
wire n_2061;
wire n_2685;
wire n_5987;
wire n_2512;
wire n_1790;
wire n_2788;
wire n_6642;
wire n_6291;
wire n_6510;
wire n_1443;
wire n_5264;
wire n_2595;
wire n_1465;
wire n_3084;
wire n_705;
wire n_6781;
wire n_7667;
wire n_4593;
wire n_8024;
wire n_7123;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_461;
wire n_3554;
wire n_6509;
wire n_2717;
wire n_6376;
wire n_1391;
wire n_8107;
wire n_2981;
wire n_225;
wire n_1006;
wire n_546;
wire n_4995;
wire n_1159;
wire n_6514;
wire n_5873;
wire n_4498;
wire n_772;
wire n_6741;
wire n_1245;
wire n_6434;
wire n_5741;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_6593;
wire n_676;
wire n_7827;
wire n_3758;
wire n_7631;
wire n_6690;
wire n_5423;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_3777;
wire n_1872;
wire n_1585;
wire n_3767;
wire n_6056;
wire n_5926;
wire n_5866;
wire n_212;
wire n_3692;
wire n_1351;
wire n_3234;
wire n_2216;
wire n_8122;
wire n_2426;
wire n_652;
wire n_6947;
wire n_4850;
wire n_1260;
wire n_3716;
wire n_7157;
wire n_2926;
wire n_4937;
wire n_798;
wire n_5574;
wire n_3391;
wire n_5877;
wire n_912;
wire n_6375;
wire n_460;
wire n_7781;
wire n_4786;
wire n_6042;
wire n_8238;
wire n_5203;
wire n_7908;
wire n_7091;
wire n_4354;
wire n_6429;
wire n_4235;
wire n_3159;
wire n_6315;
wire n_7855;
wire n_2855;
wire n_794;
wire n_2848;
wire n_7886;
wire n_7675;
wire n_6775;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_288;
wire n_1292;
wire n_7774;
wire n_6970;
wire n_1026;
wire n_6948;
wire n_3460;
wire n_1610;
wire n_5155;
wire n_2202;
wire n_306;
wire n_2952;
wire n_3530;
wire n_6133;
wire n_6920;
wire n_2693;
wire n_7409;
wire n_5408;
wire n_5812;
wire n_5540;
wire n_7381;
wire n_5804;
wire n_3240;
wire n_7999;
wire n_5066;
wire n_931;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_7087;
wire n_967;
wire n_5130;
wire n_4175;
wire n_6241;
wire n_1079;
wire n_5200;
wire n_3393;
wire n_2836;
wire n_7873;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_5992;
wire n_2172;
wire n_2601;
wire n_1880;
wire n_2365;
wire n_5684;
wire n_1399;
wire n_7228;
wire n_5981;
wire n_7784;
wire n_1855;
wire n_6632;
wire n_2333;
wire n_3629;
wire n_4948;
wire n_5413;
wire n_1903;
wire n_2147;
wire n_7713;
wire n_6623;
wire n_4020;
wire n_5150;
wire n_5111;
wire n_1226;
wire n_2224;
wire n_6933;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_3046;
wire n_2921;
wire n_1240;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_5444;
wire n_8031;
wire n_3257;
wire n_5737;
wire n_8015;
wire n_425;
wire n_3730;
wire n_5615;
wire n_3979;
wire n_6908;
wire n_5097;
wire n_2695;
wire n_7084;
wire n_2598;
wire n_3727;
wire n_6083;
wire n_6537;
wire n_976;
wire n_4003;
wire n_1832;
wire n_767;
wire n_6390;
wire n_7640;
wire n_2302;
wire n_6799;
wire n_3014;
wire n_7912;
wire n_2294;
wire n_6278;
wire n_2274;
wire n_7195;
wire n_5640;
wire n_3342;
wire n_2895;
wire n_6101;
wire n_7298;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_5550;
wire n_397;
wire n_3375;
wire n_2768;
wire n_351;
wire n_155;
wire n_3760;
wire n_5661;
wire n_7641;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_5306;
wire n_5905;
wire n_7949;
wire n_6112;
wire n_2728;
wire n_2025;
wire n_3744;
wire n_5457;
wire n_5159;
wire n_4022;
wire n_7115;
wire n_1020;
wire n_7764;
wire n_172;
wire n_2495;
wire n_1058;
wire n_4336;
wire n_8128;
wire n_7520;
wire n_5314;
wire n_7616;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_6412;
wire n_1279;
wire n_6271;
wire n_7235;
wire n_2511;
wire n_564;
wire n_6572;
wire n_3981;
wire n_7271;
wire n_2681;
wire n_7222;
wire n_1689;
wire n_2535;
wire n_1255;
wire n_3031;
wire n_345;
wire n_6930;
wire n_2335;
wire n_5482;
wire n_3215;
wire n_1401;
wire n_3138;
wire n_776;
wire n_2860;
wire n_2041;
wire n_1933;
wire n_6584;
wire n_4494;
wire n_130;
wire n_6387;
wire n_466;
wire n_4201;
wire n_346;
wire n_6470;
wire n_7206;
wire n_552;
wire n_5287;
wire n_8272;
wire n_4719;
wire n_5651;
wire n_264;
wire n_3577;
wire n_6625;
wire n_4074;
wire n_7383;
wire n_3994;
wire n_4636;
wire n_6826;
wire n_3185;
wire n_4983;
wire n_1217;
wire n_327;
wire n_2662;
wire n_4386;
wire n_6341;
wire n_6374;
wire n_3917;
wire n_1231;
wire n_5623;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_8178;
wire n_5524;
wire n_7854;
wire n_926;
wire n_2296;
wire n_5735;
wire n_7959;
wire n_8234;
wire n_6363;
wire n_6588;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_7897;
wire n_186;
wire n_4225;
wire n_6811;
wire n_6687;
wire n_4658;
wire n_7135;
wire n_6037;
wire n_4186;
wire n_1501;
wire n_2241;
wire n_6865;
wire n_7211;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_2531;
wire n_7132;
wire n_1570;
wire n_7533;
wire n_3377;
wire n_6722;
wire n_1518;
wire n_6420;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_7766;
wire n_855;
wire n_2059;
wire n_8184;
wire n_4713;
wire n_5787;
wire n_6911;
wire n_1287;
wire n_1611;
wire n_120;
wire n_7129;
wire n_7080;
wire n_3374;
wire n_4870;
wire n_6981;
wire n_7776;
wire n_4818;
wire n_8001;
wire n_7436;
wire n_7020;
wire n_5935;
wire n_8064;
wire n_6696;
wire n_4916;
wire n_5967;
wire n_6095;
wire n_4323;
wire n_6045;
wire n_529;
wire n_1899;
wire n_5934;
wire n_5376;
wire n_3508;
wire n_6300;
wire n_6653;
wire n_6372;
wire n_4129;
wire n_7120;
wire n_7978;
wire n_5488;
wire n_1105;
wire n_6900;
wire n_5727;
wire n_3599;
wire n_6660;
wire n_8131;
wire n_5988;
wire n_6424;
wire n_5646;
wire n_7448;
wire n_4480;
wire n_5711;
wire n_3734;
wire n_6787;
wire n_7694;
wire n_5832;
wire n_6254;
wire n_7460;
wire n_3401;
wire n_983;
wire n_7142;
wire n_6423;
wire n_6526;
wire n_699;
wire n_3542;
wire n_301;
wire n_3263;
wire n_5891;
wire n_8150;
wire n_2523;
wire n_1945;
wire n_2418;
wire n_1377;
wire n_1614;
wire n_5328;
wire n_3819;
wire n_3222;
wire n_325;
wire n_1740;
wire n_4616;
wire n_5016;
wire n_6011;
wire n_7465;
wire n_5470;
wire n_1092;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_6176;
wire n_1963;
wire n_3868;
wire n_729;
wire n_8230;
wire n_6222;
wire n_2218;
wire n_1122;
wire n_7760;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_6969;
wire n_390;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_6587;
wire n_6688;
wire n_6505;
wire n_5362;
wire n_8209;
wire n_388;
wire n_2754;
wire n_4580;
wire n_6762;
wire n_1218;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_7629;
wire n_6987;
wire n_877;
wire n_3995;
wire n_7567;
wire n_3908;
wire n_6453;
wire n_6308;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_1089;
wire n_7449;
wire n_8151;
wire n_1502;
wire n_3501;
wire n_1478;
wire n_2555;
wire n_3216;
wire n_3568;
wire n_2708;
wire n_6187;
wire n_735;
wire n_6597;
wire n_4844;
wire n_6220;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_845;
wire n_7479;
wire n_7882;
wire n_1649;
wire n_2470;
wire n_7517;
wire n_1297;
wire n_3551;
wire n_417;
wire n_1708;
wire n_5037;
wire n_7305;
wire n_5650;
wire n_5729;
wire n_5581;
wire n_4677;
wire n_5189;
wire n_8070;
wire n_4525;
wire n_6149;
wire n_3364;
wire n_2643;
wire n_755;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_7878;
wire n_4369;
wire n_3826;
wire n_5648;
wire n_278;
wire n_2266;
wire n_6439;
wire n_4324;
wire n_842;
wire n_148;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_6547;
wire n_7177;
wire n_7902;
wire n_742;
wire n_5160;
wire n_1719;
wire n_2742;
wire n_769;
wire n_3671;
wire n_2366;
wire n_5762;
wire n_1753;
wire n_5484;
wire n_1372;
wire n_476;
wire n_1895;
wire n_7353;
wire n_4104;
wire n_8054;
wire n_982;
wire n_3791;
wire n_915;
wire n_6478;
wire n_2008;
wire n_454;
wire n_298;
wire n_4989;
wire n_5874;
wire n_3064;
wire n_3199;
wire n_2127;
wire n_7050;
wire n_3151;
wire n_7590;
wire n_6906;
wire n_403;
wire n_3016;
wire n_2460;
wire n_6739;
wire n_1319;
wire n_3669;
wire n_3367;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_606;
wire n_4528;
wire n_2772;
wire n_1700;
wire n_659;
wire n_1332;
wire n_7818;
wire n_509;
wire n_7645;
wire n_5385;
wire n_7482;
wire n_1747;
wire n_3990;
wire n_5622;
wire n_1171;
wire n_5635;
wire n_4069;
wire n_3582;
wire n_7907;
wire n_4280;
wire n_1867;
wire n_6034;
wire n_5609;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_4811;
wire n_2696;
wire n_5595;
wire n_5256;
wire n_4779;
wire n_521;
wire n_5910;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_5380;
wire n_1400;
wire n_7862;
wire n_3735;
wire n_7565;
wire n_7410;
wire n_6422;
wire n_1527;
wire n_1513;
wire n_3656;
wire n_7721;
wire n_4524;
wire n_8061;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_5568;
wire n_5941;
wire n_4891;
wire n_2629;
wire n_3369;
wire n_1257;
wire n_1954;
wire n_6604;
wire n_3964;
wire n_6611;
wire n_5364;
wire n_3302;
wire n_5597;
wire n_2486;
wire n_1897;
wire n_6999;
wire n_8072;
wire n_8086;
wire n_5469;
wire n_2137;
wire n_3685;
wire n_6019;
wire n_7539;
wire n_6440;
wire n_4977;
wire n_2492;
wire n_6976;
wire n_7608;
wire n_7234;
wire n_2939;
wire n_3425;
wire n_4876;
wire n_241;
wire n_5021;
wire n_1449;
wire n_2900;
wire n_797;
wire n_2912;
wire n_5936;
wire n_595;
wire n_1405;
wire n_3813;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_6784;
wire n_1757;
wire n_1950;
wire n_2264;
wire n_805;
wire n_5928;
wire n_2032;
wire n_2090;
wire n_7830;
wire n_8050;
wire n_3124;
wire n_3811;
wire n_295;
wire n_4200;
wire n_190;
wire n_2249;
wire n_5785;
wire n_3411;
wire n_5222;
wire n_6165;
wire n_3463;
wire n_2785;
wire n_730;
wire n_4938;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_6114;
wire n_1856;
wire n_463;
wire n_1524;
wire n_2928;
wire n_5505;
wire n_1118;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_1293;
wire n_961;
wire n_469;
wire n_726;
wire n_5504;
wire n_878;
wire n_7348;
wire n_4118;
wire n_6829;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_8010;
wire n_3157;
wire n_1180;
wire n_1697;
wire n_2730;
wire n_6464;
wire n_5129;
wire n_806;
wire n_1350;
wire n_7320;
wire n_4704;
wire n_2720;
wire n_649;
wire n_1561;
wire n_5494;
wire n_5970;
wire n_2405;
wire n_6838;
wire n_2700;
wire n_6368;
wire n_1616;
wire n_7935;
wire n_2416;
wire n_8143;
wire n_2064;
wire n_3640;
wire n_5663;
wire n_5161;
wire n_7933;
wire n_1557;
wire n_6640;
wire n_7155;
wire n_6166;
wire n_4744;
wire n_5378;
wire n_5626;
wire n_349;
wire n_4706;
wire n_3879;
wire n_2022;
wire n_4343;
wire n_6850;
wire n_1505;
wire n_2408;
wire n_4764;
wire n_5389;
wire n_7743;
wire n_4990;
wire n_2986;
wire n_949;
wire n_2454;
wire n_6550;
wire n_6656;
wire n_8153;
wire n_6972;
wire n_3591;
wire n_198;
wire n_2760;
wire n_4919;
wire n_1208;
wire n_7043;
wire n_7986;
wire n_3317;
wire n_8049;
wire n_7266;
wire n_5653;
wire n_4835;
wire n_1151;
wire n_554;
wire n_4420;
wire n_7996;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_354;
wire n_5266;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_5800;
wire n_1133;
wire n_883;
wire n_4372;
wire n_5396;
wire n_4097;
wire n_4162;
wire n_5766;
wire n_5293;
wire n_779;
wire n_4790;
wire n_594;
wire n_7035;
wire n_4173;
wire n_5309;
wire n_6047;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_422;
wire n_1269;
wire n_8277;
wire n_7442;
wire n_4727;
wire n_1547;
wire n_1438;
wire n_6568;
wire n_3654;
wire n_5627;
wire n_1047;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_7153;
wire n_6258;
wire n_1288;
wire n_7939;
wire n_7715;
wire n_2173;
wire n_3982;
wire n_7350;
wire n_3647;
wire n_7314;
wire n_6026;
wire n_1143;
wire n_3973;
wire n_8052;
wire n_4799;
wire n_8082;
wire n_5882;
wire n_6700;
wire n_7136;
wire n_4534;
wire n_5636;
wire n_4960;
wire n_7699;
wire n_1153;
wire n_271;
wire n_465;
wire n_1103;
wire n_5707;
wire n_5594;
wire n_3738;
wire n_894;
wire n_5697;
wire n_1380;
wire n_562;
wire n_2020;
wire n_7580;
wire n_5606;
wire n_6727;
wire n_2310;
wire n_510;
wire n_5911;
wire n_7340;
wire n_8080;
wire n_256;
wire n_3600;
wire n_7303;
wire n_1023;
wire n_914;
wire n_7870;
wire n_689;
wire n_6139;
wire n_7568;
wire n_7399;
wire n_5382;
wire n_4327;
wire n_7387;
wire n_3190;
wire n_3027;
wire n_6454;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_497;
wire n_3733;
wire n_1165;
wire n_3967;
wire n_6333;
wire n_7004;
wire n_455;
wire n_588;
wire n_638;
wire n_4370;
wire n_5638;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_1417;
wire n_3096;
wire n_7207;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_7167;
wire n_2234;
wire n_1341;
wire n_5849;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_1603;
wire n_5841;
wire n_7146;
wire n_7030;
wire n_4478;
wire n_8203;
wire n_413;
wire n_2935;
wire n_4246;
wire n_715;
wire n_7618;
wire n_1066;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_685;
wire n_4061;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_4754;
wire n_1534;
wire n_8268;
wire n_8171;
wire n_1290;
wire n_4375;
wire n_617;
wire n_2396;
wire n_3368;
wire n_1559;
wire n_8008;
wire n_7633;
wire n_3117;
wire n_4684;
wire n_743;
wire n_1546;
wire n_3384;
wire n_5279;
wire n_7159;
wire n_2592;
wire n_3490;
wire n_7280;
wire n_962;
wire n_5043;
wire n_7339;
wire n_7597;
wire n_4241;
wire n_1622;
wire n_3113;
wire n_2751;
wire n_4183;
wire n_7768;
wire n_918;
wire n_1968;
wire n_5645;
wire n_639;
wire n_5020;
wire n_673;
wire n_6455;
wire n_2842;
wire n_7615;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_8271;
wire n_3720;
wire n_6183;
wire n_6107;
wire n_6476;
wire n_5232;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_8228;
wire n_1193;
wire n_1345;
wire n_5035;
wire n_3037;
wire n_1336;
wire n_1033;
wire n_5453;
wire n_4333;
wire n_5339;
wire n_6003;
wire n_5443;
wire n_8133;
wire n_7612;
wire n_1166;
wire n_2007;
wire n_3363;
wire n_6636;
wire n_1158;
wire n_1803;
wire n_872;
wire n_3522;
wire n_8172;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_6554;
wire n_5631;
wire n_3481;
wire n_280;
wire n_6994;
wire n_7401;
wire n_5101;
wire n_6020;
wire n_2236;
wire n_6185;
wire n_692;
wire n_7594;
wire n_7711;
wire n_7321;
wire n_4457;
wire n_223;
wire n_2150;
wire n_6785;
wire n_1816;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_6870;
wire n_3305;
wire n_6643;
wire n_7574;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_8226;
wire n_6695;
wire n_7529;
wire n_3354;
wire n_5608;
wire n_6501;
wire n_2204;
wire n_1481;
wire n_2040;
wire n_6466;
wire n_2151;
wire n_2455;
wire n_827;
wire n_3437;
wire n_6467;
wire n_2231;
wire n_4212;
wire n_622;
wire n_4584;
wire n_7522;
wire n_7188;
wire n_8088;
wire n_5702;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_4477;
wire n_5806;
wire n_4110;
wire n_5182;
wire n_1221;
wire n_4217;
wire n_5277;
wire n_792;
wire n_1262;
wire n_6507;
wire n_1942;
wire n_6618;
wire n_2951;
wire n_4048;
wire n_3807;
wire n_6213;
wire n_1579;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_229;
wire n_923;
wire n_1124;
wire n_7872;
wire n_1326;
wire n_3969;
wire n_6873;
wire n_7958;
wire n_2282;
wire n_4605;
wire n_8118;
wire n_981;
wire n_3873;
wire n_4649;
wire n_5747;
wire n_7101;
wire n_1204;
wire n_7843;
wire n_994;
wire n_2428;
wire n_1360;
wire n_6063;
wire n_2858;
wire n_3076;
wire n_7578;
wire n_3410;
wire n_5415;
wire n_856;
wire n_7261;
wire n_4999;
wire n_4592;
wire n_1564;
wire n_6993;
wire n_508;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_8100;
wire n_1858;
wire n_353;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_1361;
wire n_6767;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_5687;
wire n_1411;
wire n_1359;
wire n_6558;
wire n_6755;
wire n_6153;
wire n_3536;
wire n_1721;
wire n_7263;
wire n_3782;
wire n_1317;
wire n_6608;
wire n_6202;
wire n_6780;
wire n_7688;
wire n_3594;
wire n_5383;
wire n_2385;
wire n_6635;
wire n_7245;
wire n_7925;
wire n_7310;
wire n_294;
wire n_6359;
wire n_5690;
wire n_1980;
wire n_5740;
wire n_7093;
wire n_4177;
wire n_2501;
wire n_7585;
wire n_1385;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_7418;
wire n_6353;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_6577;
wire n_7772;
wire n_2028;
wire n_919;
wire n_3114;
wire n_2092;
wire n_6082;
wire n_3622;
wire n_2817;
wire n_2773;
wire n_2402;
wire n_1458;
wire n_679;
wire n_220;
wire n_3047;
wire n_3163;
wire n_5361;
wire n_7312;
wire n_7514;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_6105;
wire n_387;
wire n_826;
wire n_5512;
wire n_7738;
wire n_2808;
wire n_2344;
wire n_3520;
wire n_2392;
wire n_7609;
wire n_3272;
wire n_3122;
wire n_5898;
wire n_7113;
wire n_6548;
wire n_607;
wire n_8213;
wire n_5923;
wire n_3687;
wire n_2787;
wire n_6657;
wire n_5617;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_5946;
wire n_1268;
wire n_2676;
wire n_7282;
wire n_372;
wire n_2770;
wire n_4550;
wire n_4347;
wire n_7921;
wire n_702;
wire n_5193;
wire n_4933;
wire n_968;
wire n_4144;
wire n_5514;
wire n_5611;
wire n_2375;
wire n_3278;
wire n_5579;
wire n_4167;
wire n_6380;
wire n_3608;
wire n_4895;
wire n_1282;
wire n_6163;
wire n_7170;
wire n_4726;
wire n_5573;
wire n_5143;
wire n_5836;
wire n_1755;
wire n_5188;
wire n_6674;
wire n_5049;
wire n_2212;
wire n_7489;
wire n_6331;
wire n_5308;
wire n_311;
wire n_4434;
wire n_5068;
wire n_7863;
wire n_6493;
wire n_7363;
wire n_7281;
wire n_5739;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_7968;
wire n_6023;
wire n_7820;
wire n_269;
wire n_816;
wire n_7833;
wire n_1322;
wire n_3829;
wire n_4510;
wire n_7750;
wire n_5057;
wire n_446;
wire n_6196;
wire n_5425;
wire n_5273;
wire n_5839;
wire n_2469;
wire n_7588;
wire n_1125;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_7697;
wire n_5887;
wire n_7808;
wire n_3068;
wire n_1629;
wire n_7603;
wire n_1094;
wire n_6321;
wire n_5683;
wire n_1510;
wire n_3002;
wire n_7192;
wire n_1099;
wire n_5248;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_759;
wire n_567;
wire n_4156;
wire n_1727;
wire n_3693;
wire n_5880;
wire n_8012;
wire n_3132;
wire n_5002;
wire n_5487;
wire n_5649;
wire n_5531;
wire n_831;
wire n_3681;
wire n_5666;
wire n_3970;
wire n_778;
wire n_2351;
wire n_1619;
wire n_7988;
wire n_550;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_6824;
wire n_6954;
wire n_6450;
wire n_1152;
wire n_6995;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_1236;
wire n_4579;
wire n_6347;
wire n_6496;
wire n_4776;
wire n_671;
wire n_8105;
wire n_2704;
wire n_1334;
wire n_6745;
wire n_7943;
wire n_3729;
wire n_6698;
wire n_4471;
wire n_6968;
wire n_7377;
wire n_4392;
wire n_3103;
wire n_488;
wire n_6064;
wire n_505;
wire n_2048;
wire n_7723;
wire n_498;
wire n_3028;
wire n_4691;
wire n_7904;
wire n_3148;
wire n_3775;
wire n_5682;
wire n_684;
wire n_5461;
wire n_7296;
wire n_3966;
wire n_4397;
wire n_6164;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_5730;
wire n_6292;
wire n_7759;
wire n_6743;
wire n_4165;
wire n_2056;
wire n_5754;
wire n_2852;
wire n_2515;
wire n_6330;
wire n_1600;
wire n_1144;
wire n_7178;
wire n_838;
wire n_1941;
wire n_7045;
wire n_175;
wire n_3637;
wire n_1017;
wire n_734;
wire n_4893;
wire n_2240;
wire n_7777;
wire n_4258;
wire n_5756;
wire n_310;
wire n_7693;
wire n_709;
wire n_2917;
wire n_3194;
wire n_2085;
wire n_2432;
wire n_5033;
wire n_6015;
wire n_1686;
wire n_6408;
wire n_4232;
wire n_5075;
wire n_8078;
wire n_2097;
wire n_662;
wire n_3461;
wire n_7682;
wire n_7300;
wire n_939;
wire n_1410;
wire n_2297;
wire n_6861;
wire n_4203;
wire n_5789;
wire n_5400;
wire n_1325;
wire n_7558;
wire n_1223;
wire n_5347;
wire n_2957;
wire n_572;
wire n_8103;
wire n_1983;
wire n_7798;
wire n_4767;
wire n_4569;
wire n_948;
wire n_448;
wire n_6528;
wire n_3820;
wire n_5144;
wire n_6895;
wire n_3072;
wire n_2961;
wire n_5509;
wire n_4468;
wire n_1923;
wire n_3848;
wire n_7400;
wire n_3631;
wire n_7393;
wire n_6590;
wire n_8116;
wire n_6523;
wire n_5169;
wire n_4885;
wire n_7475;
wire n_1479;
wire n_4698;
wire n_1031;
wire n_3674;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_5349;
wire n_6472;
wire n_3763;
wire n_933;
wire n_6389;
wire n_3499;
wire n_5534;
wire n_1821;
wire n_3947;
wire n_3910;
wire n_492;
wire n_252;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_2995;
wire n_6073;
wire n_4533;
wire n_4287;
wire n_3228;
wire n_8286;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_1186;
wire n_6869;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_7672;
wire n_4556;
wire n_6137;
wire n_2205;
wire n_2183;
wire n_389;
wire n_1724;
wire n_3088;
wire n_1707;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_1126;
wire n_5079;
wire n_8247;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_895;
wire n_1639;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_5751;
wire n_626;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_7712;
wire n_6885;
wire n_7681;
wire n_5039;
wire n_1818;
wire n_6613;
wire n_6580;
wire n_4265;
wire n_6404;
wire n_6120;
wire n_3557;
wire n_1598;
wire n_2269;
wire n_7491;
wire n_265;
wire n_1583;
wire n_4612;
wire n_5997;
wire n_5375;
wire n_5438;
wire n_7150;
wire n_7954;
wire n_7974;
wire n_1264;
wire n_6602;
wire n_6530;
wire n_7915;
wire n_4958;
wire n_1827;
wire n_4149;
wire n_6135;
wire n_246;
wire n_1752;
wire n_2361;
wire n_4538;
wire n_3030;
wire n_3505;
wire n_5563;
wire n_3075;
wire n_1102;
wire n_2239;
wire n_6942;
wire n_7860;
wire n_6892;
wire n_1296;
wire n_4730;
wire n_7357;
wire n_8112;
wire n_8060;
wire n_6782;
wire n_4421;
wire n_6230;
wire n_2464;
wire n_3697;
wire n_882;
wire n_8244;
wire n_2304;
wire n_2514;
wire n_6977;
wire n_7229;
wire n_8096;
wire n_7336;
wire n_5932;
wire n_289;
wire n_112;
wire n_6598;
wire n_6795;
wire n_6121;
wire n_457;
wire n_1299;
wire n_3430;
wire n_5919;
wire n_2063;
wire n_3489;
wire n_5012;
wire n_6614;
wire n_6506;
wire n_2079;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_3484;
wire n_6001;
wire n_411;
wire n_4971;
wire n_2095;
wire n_7493;
wire n_5664;
wire n_2738;
wire n_6406;
wire n_5890;
wire n_2590;
wire n_4661;
wire n_2797;
wire n_357;
wire n_3041;
wire n_412;
wire n_5823;
wire n_1421;
wire n_2423;
wire n_2208;
wire n_5944;
wire n_5422;
wire n_6989;
wire n_8145;
wire n_8237;
wire n_6299;
wire n_7424;
wire n_5246;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_1069;
wire n_4305;
wire n_2037;
wire n_2953;
wire n_573;
wire n_2823;
wire n_7273;
wire n_7901;
wire n_3684;
wire n_5725;
wire n_5404;
wire n_913;
wire n_1681;
wire n_4834;
wire n_1507;
wire n_5332;
wire n_7149;
wire n_589;
wire n_2866;
wire n_7116;
wire n_3153;
wire n_1174;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_8211;
wire n_3268;
wire n_2559;
wire n_5616;
wire n_1383;
wire n_603;
wire n_8055;
wire n_373;
wire n_4259;
wire n_5870;
wire n_7909;
wire n_2030;
wire n_6053;
wire n_850;
wire n_6233;
wire n_4299;
wire n_5625;
wire n_245;
wire n_319;
wire n_6758;
wire n_2407;
wire n_690;
wire n_5367;
wire n_525;
wire n_2243;
wire n_6629;
wire n_5288;
wire n_2694;
wire n_6356;
wire n_5601;
wire n_3742;
wire n_4965;
wire n_7601;
wire n_1837;
wire n_7033;
wire n_4178;
wire n_6010;
wire n_189;
wire n_8157;
wire n_2006;
wire n_4953;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_7147;
wire n_7596;
wire n_5294;
wire n_8161;
wire n_5570;
wire n_6411;
wire n_2731;
wire n_3703;
wire n_5670;
wire n_5411;
wire n_1246;
wire n_5265;
wire n_5955;
wire n_7549;
wire n_2123;
wire n_2238;
wire n_4802;
wire n_4793;
wire n_6032;
wire n_1196;
wire n_5733;
wire n_3435;
wire n_410;
wire n_2380;
wire n_1187;
wire n_4897;
wire n_6918;
wire n_1298;
wire n_1745;
wire n_4674;
wire n_568;
wire n_4796;
wire n_8290;
wire n_1088;
wire n_7138;
wire n_766;
wire n_6401;
wire n_7279;
wire n_5184;
wire n_7976;
wire n_377;
wire n_2750;
wire n_2547;
wire n_7617;
wire n_279;
wire n_945;
wire n_4575;
wire n_3665;
wire n_3063;
wire n_8062;
wire n_3281;
wire n_7137;
wire n_3535;
wire n_5061;
wire n_2288;
wire n_3858;
wire n_7700;
wire n_4653;
wire n_8275;
wire n_7474;
wire n_4589;
wire n_7124;
wire n_5978;
wire n_6853;
wire n_3220;
wire n_4581;
wire n_6008;
wire n_500;
wire n_665;
wire n_4625;
wire n_7098;
wire n_6181;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_3679;
wire n_738;
wire n_5575;
wire n_6654;
wire n_7661;
wire n_672;
wire n_4968;
wire n_7801;
wire n_6907;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_4038;
wire n_3856;
wire n_5316;
wire n_7876;
wire n_2735;
wire n_953;
wire n_4214;
wire n_143;
wire n_1888;
wire n_5290;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_557;
wire n_3419;
wire n_7323;
wire n_989;
wire n_5048;
wire n_2233;
wire n_5363;
wire n_5665;
wire n_6517;
wire n_795;
wire n_4892;
wire n_6339;
wire n_1936;
wire n_3890;
wire n_6170;
wire n_7247;
wire n_6394;
wire n_8048;
wire n_821;
wire n_770;
wire n_5607;
wire n_1514;
wire n_7929;
wire n_486;
wire n_2782;
wire n_569;
wire n_3929;
wire n_971;
wire n_4353;
wire n_2201;
wire n_8212;
wire n_4950;
wire n_1650;
wire n_7755;
wire n_6504;
wire n_4176;
wire n_7556;
wire n_222;
wire n_4124;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_5462;
wire n_6814;
wire n_7216;
wire n_4488;
wire n_5278;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_3756;
wire n_8043;
wire n_8223;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_8159;
wire n_5845;
wire n_4608;
wire n_6691;
wire n_432;
wire n_293;
wire n_3948;
wire n_4839;
wire n_1074;
wire n_5969;
wire n_1765;
wire n_108;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_206;
wire n_2332;
wire n_2391;
wire n_6343;
wire n_6005;
wire n_611;
wire n_1295;
wire n_2060;
wire n_3883;
wire n_1013;
wire n_6686;
wire n_4032;
wire n_2571;
wire n_136;
wire n_6437;
wire n_5736;
wire n_4929;
wire n_2874;
wire n_6029;
wire n_6536;
wire n_6684;
wire n_4117;
wire n_300;
wire n_6025;
wire n_3049;
wire n_3634;
wire n_5436;
wire n_7962;
wire n_2341;
wire n_1654;
wire n_6697;
wire n_3066;
wire n_2045;
wire n_6085;
wire n_3913;
wire n_5341;
wire n_2575;
wire n_3739;
wire n_1230;
wire n_5140;
wire n_376;
wire n_1597;
wire n_2942;
wire n_6062;
wire n_1771;
wire n_4541;
wire n_6715;
wire n_3271;
wire n_3164;
wire n_3861;
wire n_5096;
wire n_2043;
wire n_6771;
wire n_7905;
wire n_4171;
wire n_5847;
wire n_7204;
wire n_7022;
wire n_6383;
wire n_4815;
wire n_4665;
wire n_5639;
wire n_6877;
wire n_7308;
wire n_7476;
wire n_4884;
wire n_3580;
wire n_1437;
wire n_8249;
wire n_4276;
wire n_1378;
wire n_5268;
wire n_5050;
wire n_209;
wire n_5240;
wire n_5503;
wire n_1461;
wire n_5718;
wire n_7208;
wire n_7718;
wire n_1876;
wire n_1830;
wire n_5001;
wire n_6567;
wire n_503;
wire n_5658;
wire n_1112;
wire n_700;
wire n_4174;
wire n_6868;
wire n_7290;
wire n_5131;
wire n_6813;
wire n_7756;
wire n_5546;
wire n_6294;
wire n_7795;
wire n_7822;
wire n_5174;
wire n_2145;
wire n_4801;
wire n_6079;
wire n_6260;
wire n_680;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_6520;
wire n_7623;
wire n_380;
wire n_3119;
wire n_6671;
wire n_4740;
wire n_1108;
wire n_1274;
wire n_7632;
wire n_4394;
wire n_257;
wire n_5544;
wire n_6637;
wire n_6444;
wire n_475;
wire n_6729;
wire n_5660;
wire n_6958;
wire n_8073;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_5541;
wire n_6314;
wire n_577;
wire n_5610;
wire n_407;
wire n_916;
wire n_2810;
wire n_6703;
wire n_1884;
wire n_1555;
wire n_762;
wire n_1253;
wire n_1468;
wire n_4378;
wire n_5166;
wire n_2683;
wire n_6065;
wire n_7265;
wire n_4180;
wire n_4459;
wire n_6878;
wire n_3624;
wire n_6725;
wire n_8181;
wire n_5808;
wire n_1182;
wire n_6527;
wire n_4594;
wire n_8045;
wire n_7289;
wire n_7538;
wire n_2748;
wire n_4642;
wire n_6913;
wire n_1376;
wire n_7473;
wire n_7242;
wire n_6533;
wire n_513;
wire n_179;
wire n_7164;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_8022;
wire n_3544;
wire n_6845;
wire n_5300;
wire n_8227;
wire n_7853;
wire n_2072;
wire n_3852;
wire n_5233;
wire n_5381;
wire n_436;
wire n_5770;
wire n_7483;
wire n_5710;
wire n_324;
wire n_1491;
wire n_2628;
wire n_7389;
wire n_3219;
wire n_111;
wire n_274;
wire n_1083;
wire n_5333;
wire n_5799;
wire n_6265;
wire n_4914;
wire n_3510;
wire n_7046;
wire n_7834;
wire n_4587;
wire n_1139;
wire n_3688;
wire n_5008;
wire n_1312;
wire n_3871;
wire n_892;
wire n_3757;
wire n_1567;
wire n_563;
wire n_2219;
wire n_6148;
wire n_2100;
wire n_8255;
wire n_3666;
wire n_5538;
wire n_990;
wire n_6357;
wire n_867;
wire n_8216;
wire n_3479;
wire n_944;
wire n_5499;
wire n_749;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_6522;
wire n_7811;
wire n_4285;
wire n_7097;
wire n_7000;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_650;
wire n_3741;
wire n_5582;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_5675;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_5109;
wire n_7880;
wire n_712;
wire n_909;
wire n_6713;
wire n_8149;
wire n_1392;
wire n_2066;
wire n_5281;
wire n_2762;
wire n_6087;
wire n_964;
wire n_7851;
wire n_2220;
wire n_7342;
wire n_7044;
wire n_7810;
wire n_6108;
wire n_7664;
wire n_6100;
wire n_6800;
wire n_7364;
wire n_6866;
wire n_7114;
wire n_6373;
wire n_4433;
wire n_2829;
wire n_7332;
wire n_5862;
wire n_471;
wire n_7477;
wire n_1914;
wire n_8208;
wire n_2253;
wire n_7468;
wire n_5886;
wire n_7714;
wire n_7899;
wire n_6415;
wire n_6783;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_1633;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_2328;
wire n_7845;
wire n_347;
wire n_2434;
wire n_183;
wire n_1234;
wire n_3936;
wire n_479;
wire n_5564;
wire n_2261;
wire n_3082;
wire n_5162;
wire n_5442;
wire n_2473;
wire n_5802;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_6340;
wire n_7858;
wire n_3867;
wire n_3397;
wire n_6103;
wire n_1646;
wire n_6513;
wire n_6392;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_1237;
wire n_6720;
wire n_5883;
wire n_1095;
wire n_3078;
wire n_6078;
wire n_3971;
wire n_370;
wire n_7680;
wire n_5630;
wire n_6666;
wire n_286;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_1531;
wire n_2113;
wire n_6815;
wire n_1387;
wire n_6207;
wire n_6381;
wire n_3711;
wire n_5054;
wire n_6571;
wire n_3171;
wire n_5929;
wire n_7710;
wire n_5394;
wire n_4751;
wire n_4242;
wire n_5975;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_1496;
wire n_2812;
wire n_3300;
wire n_7061;
wire n_8104;
wire n_7066;
wire n_5496;
wire n_7485;
wire n_3104;
wire n_7174;
wire n_8014;
wire n_6661;
wire n_4122;
wire n_2132;
wire n_4522;
wire n_5991;
wire n_4952;
wire n_6967;
wire n_4426;
wire n_5956;
wire n_5699;
wire n_4362;
wire n_3267;
wire n_6017;
wire n_3946;
wire n_5920;
wire n_2112;
wire n_2640;
wire n_6125;
wire n_5000;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_4089;
wire n_3513;
wire n_1173;
wire n_3498;
wire n_5132;
wire n_2350;
wire n_6414;
wire n_5535;
wire n_1068;
wire n_1198;
wire n_4506;
wire n_6097;
wire n_7783;
wire n_7662;
wire n_6057;
wire n_6936;
wire n_487;
wire n_4728;
wire n_7171;
wire n_7990;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_7003;
wire n_8137;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_3863;
wire n_6302;
wire n_2327;
wire n_158;
wire n_3882;
wire n_3916;
wire n_6922;
wire n_1365;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_405;
wire n_3332;
wire n_8069;
wire n_7501;
wire n_320;
wire n_6432;
wire n_7984;
wire n_2055;
wire n_2998;
wire n_7366;
wire n_1423;
wire n_8173;
wire n_4359;
wire n_481;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_7589;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_218;
wire n_6880;
wire n_6223;
wire n_5176;
wire n_4039;
wire n_5793;
wire n_6926;
wire n_1798;
wire n_8091;
wire n_3057;
wire n_1608;
wire n_5761;
wire n_6699;
wire n_547;
wire n_439;
wire n_677;
wire n_3983;
wire n_8254;
wire n_703;
wire n_3318;
wire n_7232;
wire n_3385;
wire n_7511;
wire n_326;
wire n_227;
wire n_3773;
wire n_3494;
wire n_1278;
wire n_6957;
wire n_5074;
wire n_7917;
wire n_3788;
wire n_3939;
wire n_590;
wire n_727;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_6694;
wire n_545;
wire n_2496;
wire n_3260;
wire n_536;
wire n_3349;
wire n_6449;
wire n_4348;
wire n_1602;
wire n_7422;
wire n_3139;
wire n_427;
wire n_3801;
wire n_5681;
wire n_2338;
wire n_5261;
wire n_1080;
wire n_3636;
wire n_6591;
wire n_7466;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_7621;
wire n_8274;
wire n_2057;
wire n_6594;
wire n_6342;
wire n_1205;
wire n_6195;
wire n_163;
wire n_2716;
wire n_6441;
wire n_7158;
wire n_7572;
wire n_314;
wire n_2944;
wire n_2780;
wire n_3439;
wire n_1120;
wire n_7500;
wire n_1202;
wire n_4084;
wire n_627;
wire n_7985;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_233;
wire n_2774;
wire n_6354;
wire n_2799;
wire n_5748;
wire n_4393;
wire n_321;
wire n_6662;
wire n_7494;
wire n_3984;
wire n_1586;
wire n_1431;
wire n_4389;
wire n_6433;
wire n_1763;
wire n_6200;
wire n_5641;
wire n_8071;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_6902;
wire n_4615;
wire n_3044;
wire n_3492;
wire n_7197;
wire n_3737;
wire n_6369;
wire n_5657;
wire n_297;
wire n_2379;
wire n_3579;
wire n_1667;
wire n_888;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_1677;
wire n_5244;
wire n_5765;
wire n_5114;
wire n_4551;
wire n_178;
wire n_551;
wire n_4521;
wire n_6956;
wire n_7587;
wire n_2284;
wire n_6451;
wire n_3005;
wire n_7704;
wire n_5420;
wire n_6497;
wire n_7865;
wire n_2283;
wire n_5206;
wire n_582;
wire n_2526;
wire n_1097;
wire n_1711;
wire n_4387;
wire n_534;
wire n_2508;
wire n_3186;
wire n_6701;
wire n_2594;
wire n_1239;
wire n_5298;
wire n_3417;
wire n_8246;
wire n_560;
wire n_890;
wire n_3626;
wire n_451;
wire n_4598;
wire n_4464;
wire n_5106;
wire n_7881;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_1081;
wire n_2119;
wire n_2493;
wire n_5080;
wire n_535;
wire n_7032;
wire n_4565;
wire n_3392;
wire n_1800;
wire n_7198;
wire n_6884;
wire n_7752;
wire n_5081;
wire n_8201;
wire n_6921;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_7953;
wire n_6106;
wire n_6876;
wire n_3512;
wire n_1860;
wire n_1734;
wire n_8046;
wire n_4552;
wire n_7193;
wire n_6287;
wire n_2840;
wire n_6172;
wire n_4482;
wire n_837;
wire n_812;
wire n_4172;
wire n_5957;
wire n_4040;
wire n_3024;
wire n_5567;
wire n_5406;
wire n_6362;
wire n_4328;
wire n_1854;
wire n_666;
wire n_5191;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_6067;
wire n_2893;
wire n_6833;
wire n_4940;
wire n_785;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_7126;
wire n_5867;
wire n_456;
wire n_1394;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_7496;
wire n_6430;
wire n_873;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_6296;
wire n_4112;
wire n_342;
wire n_5602;
wire n_2035;
wire n_4928;
wire n_7196;
wire n_2614;
wire n_7360;
wire n_5428;
wire n_6325;
wire n_2494;
wire n_1538;
wire n_4865;
wire n_6678;
wire n_7982;
wire n_2128;
wire n_4071;
wire n_6564;
wire n_7268;
wire n_8174;
wire n_8187;
wire n_4436;
wire n_5786;
wire n_5822;
wire n_3586;
wire n_5817;
wire n_4160;
wire n_6109;
wire n_6385;
wire n_1668;
wire n_5798;
wire n_4137;
wire n_1078;
wire n_8032;
wire n_5417;
wire n_4545;
wire n_8200;
wire n_4758;
wire n_1161;
wire n_8036;
wire n_5713;
wire n_4840;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_618;
wire n_1191;
wire n_4535;
wire n_7518;
wire n_4385;
wire n_7779;
wire n_1215;
wire n_3748;
wire n_4731;
wire n_7575;
wire n_2337;
wire n_7073;
wire n_8092;
wire n_1786;
wire n_6309;
wire n_3732;
wire n_211;
wire n_1804;
wire n_408;
wire n_8135;
wire n_6519;
wire n_4671;
wire n_2272;
wire n_5989;
wire n_4766;
wire n_5571;
wire n_592;
wire n_4558;
wire n_1318;
wire n_1632;
wire n_1769;
wire n_7349;
wire n_1929;
wire n_4319;
wire n_6585;
wire n_7786;
wire n_2929;
wire n_4358;
wire n_1526;
wire n_7579;
wire n_7122;
wire n_4874;
wire n_180;
wire n_2656;
wire n_4904;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1258;
wire n_640;
wire n_1733;
wire n_6490;
wire n_7867;
wire n_4651;
wire n_943;
wire n_3167;
wire n_4748;
wire n_7624;
wire n_1807;
wire n_1123;
wire n_2857;
wire n_7828;
wire n_1784;
wire n_4618;
wire n_6721;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_752;
wire n_985;
wire n_5506;
wire n_7543;
wire n_5475;
wire n_8042;
wire n_7727;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_5908;
wire n_1352;
wire n_5431;
wire n_643;
wire n_8034;
wire n_226;
wire n_7778;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_7019;
wire n_682;
wire n_5315;
wire n_2633;
wire n_3708;
wire n_5752;
wire n_2907;
wire n_1429;
wire n_2353;
wire n_7702;
wire n_2528;
wire n_1778;
wire n_5746;
wire n_686;
wire n_1154;
wire n_584;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_1130;
wire n_3718;
wire n_6685;
wire n_756;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_4666;
wire n_4082;
wire n_3140;
wire n_2320;
wire n_979;
wire n_3976;
wire n_3381;
wire n_897;
wire n_2546;
wire n_2813;
wire n_7952;
wire n_7347;
wire n_3736;
wire n_6016;
wire n_4466;
wire n_891;
wire n_885;
wire n_1659;
wire n_3955;
wire n_5366;
wire n_5322;
wire n_1864;
wire n_5414;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_7791;
wire n_6971;
wire n_3336;
wire n_7739;
wire n_396;
wire n_7945;
wire n_7656;
wire n_5903;
wire n_7199;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_714;
wire n_3605;
wire n_5307;
wire n_2170;
wire n_4721;
wire n_6549;
wire n_725;
wire n_1577;
wire n_5003;
wire n_3840;
wire n_6540;
wire n_7166;
wire n_2198;
wire n_6658;
wire n_5369;
wire n_6683;
wire n_3067;
wire n_154;
wire n_3809;
wire n_4921;
wire n_473;
wire n_1852;
wire n_801;
wire n_5912;
wire n_5745;
wire n_7923;
wire n_6086;
wire n_4377;
wire n_818;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_5803;
wire n_6327;
wire n_5593;
wire n_5270;
wire n_5853;
wire n_6171;
wire n_3468;
wire n_5779;
wire n_1877;
wire n_272;
wire n_7213;
wire n_4301;
wire n_5313;
wire n_2133;
wire n_6820;
wire n_2497;
wire n_879;
wire n_5446;
wire n_7610;
wire n_7107;
wire n_4561;
wire n_1541;
wire n_597;
wire n_3291;
wire n_7456;
wire n_8095;
wire n_7369;
wire n_1472;
wire n_1050;
wire n_7548;
wire n_2578;
wire n_152;
wire n_1201;
wire n_7598;
wire n_1185;
wire n_2475;
wire n_7250;
wire n_7823;
wire n_4715;
wire n_6157;
wire n_2715;
wire n_335;
wire n_2665;
wire n_4879;
wire n_344;
wire n_5044;
wire n_210;
wire n_1090;
wire n_3755;
wire n_4536;
wire n_6676;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_5459;
wire n_224;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_7525;
wire n_4418;
wire n_7924;
wire n_3341;
wire n_4125;
wire n_5390;
wire n_5351;
wire n_5267;
wire n_1116;
wire n_5024;
wire n_7012;
wire n_3043;
wire n_2747;
wire n_1511;
wire n_276;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_538;
wire n_2845;
wire n_4151;
wire n_6923;
wire n_2036;
wire n_7649;
wire n_4412;
wire n_843;
wire n_8009;
wire n_8195;
wire n_3358;
wire n_6704;
wire n_7634;
wire n_2003;
wire n_2533;
wire n_1307;
wire n_7406;
wire n_4682;
wire n_1128;
wire n_6673;
wire n_2419;
wire n_2330;
wire n_6534;
wire n_5078;
wire n_4810;
wire n_7659;
wire n_6162;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_1955;
wire n_3289;
wire n_6127;
wire n_1440;
wire n_6246;
wire n_1370;
wire n_305;
wire n_5005;
wire n_6126;
wire n_7372;
wire n_1549;
wire n_7427;
wire n_6151;
wire n_6828;
wire n_6841;
wire n_7844;
wire n_5207;
wire n_7934;
wire n_361;
wire n_2658;
wire n_5624;
wire n_3620;
wire n_4601;
wire n_1065;
wire n_4518;
wire n_2767;
wire n_7009;
wire n_5474;
wire n_3376;
wire n_181;
wire n_7371;
wire n_1362;
wire n_3123;
wire n_5447;
wire n_2692;
wire n_683;
wire n_7463;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_5700;
wire n_5755;
wire n_2862;
wire n_4325;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_4711;
wire n_6889;
wire n_2749;
wire n_5962;
wire n_660;
wire n_464;
wire n_4413;
wire n_1210;
wire n_3307;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_6723;
wire n_7398;
wire n_1038;
wire n_3723;
wire n_7941;
wire n_4135;
wire n_6154;
wire n_5223;
wire n_5662;
wire n_414;
wire n_571;
wire n_3880;
wire n_5801;
wire n_3904;
wire n_6054;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_7011;
wire n_3405;
wire n_2313;
wire n_6393;
wire n_7074;
wire n_613;
wire n_1022;
wire n_5465;
wire n_171;
wire n_3532;
wire n_5154;
wire n_5721;
wire n_2609;
wire n_8169;
wire n_6184;
wire n_8018;
wire n_1767;
wire n_4138;
wire n_1040;
wire n_3131;
wire n_7083;
wire n_316;
wire n_125;
wire n_1973;
wire n_1444;
wire n_820;
wire n_8260;
wire n_254;
wire n_2882;
wire n_7143;
wire n_2303;
wire n_7701;
wire n_7969;
wire n_8279;
wire n_4384;
wire n_4639;
wire n_1664;
wire n_6312;
wire n_4577;
wire n_7683;
wire n_532;
wire n_2154;
wire n_7669;
wire n_1986;
wire n_6711;
wire n_2624;
wire n_6818;
wire n_6438;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_984;
wire n_5087;
wire n_1552;
wire n_2938;
wire n_7209;
wire n_2498;
wire n_6193;
wire n_3992;
wire n_8023;
wire n_7330;
wire n_6007;
wire n_621;
wire n_6734;
wire n_6535;
wire n_8053;
wire n_8059;
wire n_1772;
wire n_6879;
wire n_493;
wire n_1311;
wire n_3106;
wire n_7190;
wire n_6208;
wire n_2881;
wire n_6303;
wire n_3092;
wire n_6014;
wire n_4270;
wire n_7692;
wire n_697;
wire n_4620;
wire n_5397;
wire n_6255;
wire n_6457;
wire n_4924;
wire n_4044;
wire n_6270;
wire n_2305;
wire n_5996;
wire n_880;
wire n_5566;
wire n_3304;
wire n_7288;
wire n_4388;
wire n_7362;
wire n_7082;
wire n_7237;
wire n_3247;
wire n_7131;
wire n_6276;
wire n_739;
wire n_1028;
wire n_530;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_7042;
wire n_2809;
wire n_5652;
wire n_975;
wire n_1645;
wire n_5805;
wire n_7304;
wire n_932;
wire n_6266;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_5492;
wire n_8077;
wire n_2465;
wire n_5501;
wire n_6934;
wire n_7386;
wire n_2972;
wire n_7391;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_7754;
wire n_3178;
wire n_268;
wire n_7023;
wire n_2251;
wire n_5758;
wire n_5842;
wire n_3100;
wire n_3721;
wire n_7404;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_6147;
wire n_5692;
wire n_6765;
wire n_4973;
wire n_7981;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_191;
wire n_2487;
wire n_5473;
wire n_1834;
wire n_1011;
wire n_2534;
wire n_6352;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_6211;
wire n_8109;
wire n_116;
wire n_3576;
wire n_5562;
wire n_4858;
wire n_1445;
wire n_6093;
wire n_5370;
wire n_7378;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_5458;
wire n_7877;
wire n_7787;
wire n_7836;
wire n_8007;
wire n_2387;
wire n_4318;
wire n_332;
wire n_5227;
wire n_830;
wire n_5902;
wire n_987;
wire n_2510;
wire n_6402;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_2793;
wire n_5282;
wire n_6764;
wire n_7871;
wire n_541;
wire n_499;
wire n_2639;
wire n_7016;
wire n_4738;
wire n_2603;
wire n_5386;
wire n_1167;
wire n_6215;
wire n_4554;
wire n_7571;
wire n_8252;
wire n_4526;
wire n_4105;
wire n_969;
wire n_3663;
wire n_1663;
wire n_6955;
wire n_7563;
wire n_5952;
wire n_7180;
wire n_2086;
wire n_1926;
wire n_6569;
wire n_1630;
wire n_7919;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_8278;
wire n_443;
wire n_3431;
wire n_8180;
wire n_3355;
wire n_7031;
wire n_1738;
wire n_5716;
wire n_406;
wire n_3897;
wire n_7103;
wire n_139;
wire n_6605;
wire n_1735;
wire n_391;
wire n_5888;
wire n_4005;
wire n_8270;
wire n_8231;
wire n_4181;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_6832;
wire n_5980;
wire n_956;
wire n_765;
wire n_4092;
wire n_122;
wire n_4875;
wire n_7771;
wire n_4255;
wire n_2758;
wire n_385;
wire n_6544;
wire n_6469;
wire n_5036;
wire n_1271;
wire n_6332;
wire n_2186;
wire n_5790;
wire n_399;
wire n_7130;
wire n_6680;
wire n_4647;
wire n_3575;
wire n_6310;
wire n_8264;
wire n_2471;
wire n_7134;
wire n_3042;
wire n_8288;
wire n_1067;
wire n_1323;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_900;
wire n_5485;
wire n_5525;
wire n_7102;
wire n_6259;
wire n_3004;
wire n_1551;
wire n_5271;
wire n_4849;
wire n_2039;
wire n_7133;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_3838;
wire n_6289;
wire n_6651;
wire n_4059;
wire n_6565;
wire n_5194;
wire n_5445;
wire n_2734;
wire n_8067;
wire n_5948;
wire n_7227;
wire n_4499;
wire n_4504;
wire n_3598;
wire n_4917;
wire n_7706;
wire n_7813;
wire n_8142;
wire n_2420;
wire n_7992;
wire n_7643;
wire n_153;
wire n_648;
wire n_6836;
wire n_3273;
wire n_2918;
wire n_6595;
wire n_835;
wire n_6186;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_401;
wire n_7628;
wire n_1792;
wire n_5628;
wire n_504;
wire n_5245;
wire n_2062;
wire n_483;
wire n_4489;
wire n_822;
wire n_1459;
wire n_2153;
wire n_5329;
wire n_8224;
wire n_5472;
wire n_6035;
wire n_839;
wire n_1754;
wire n_7236;
wire n_4833;
wire n_3394;
wire n_6405;
wire n_2235;
wire n_5850;
wire n_1575;
wire n_8242;
wire n_6786;
wire n_4564;
wire n_1848;
wire n_1172;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_3581;
wire n_8110;
wire n_5072;
wire n_3778;
wire n_6769;
wire n_6844;
wire n_4322;
wire n_6361;
wire n_2260;
wire n_323;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_2206;
wire n_997;
wire n_635;
wire n_6766;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_5940;
wire n_3001;
wire n_5260;
wire n_6751;
wire n_4981;
wire n_6232;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_7519;
wire n_7802;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_7457;
wire n_5372;
wire n_6736;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_5860;
wire n_2422;
wire n_6416;
wire n_654;
wire n_2933;
wire n_7515;
wire n_3387;
wire n_7639;
wire n_6214;
wire n_3952;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_1059;
wire n_7049;
wire n_7884;
wire n_6945;
wire n_6143;
wire n_2736;
wire n_6491;
wire n_7749;
wire n_7592;
wire n_3825;
wire n_4198;
wire n_7172;
wire n_539;
wire n_8283;
wire n_977;
wire n_449;
wire n_2339;
wire n_392;
wire n_6225;
wire n_2532;
wire n_4373;
wire n_7914;
wire n_1866;
wire n_2664;
wire n_4154;
wire n_7344;
wire n_5859;
wire n_6447;
wire n_4390;
wire n_459;
wire n_1782;
wire n_7892;
wire n_1558;
wire n_4107;
wire n_2519;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_7325;
wire n_2360;
wire n_4453;
wire n_6219;
wire n_723;
wire n_1393;
wire n_7674;
wire n_6175;
wire n_6445;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3032;
wire n_5612;
wire n_4886;
wire n_6198;
wire n_5172;
wire n_881;
wire n_1019;
wire n_1477;
wire n_6499;
wire n_1982;
wire n_7983;
wire n_641;
wire n_5311;
wire n_910;
wire n_290;
wire n_5164;
wire n_4964;
wire n_6842;
wire n_4700;
wire n_4002;
wire n_217;
wire n_7361;
wire n_1114;
wire n_1742;
wire n_4679;
wire n_6397;
wire n_3815;
wire n_6827;
wire n_201;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_1273;
wire n_2982;
wire n_5495;
wire n_6281;
wire n_4483;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_5547;
wire n_4693;
wire n_1043;
wire n_6822;
wire n_5121;
wire n_4956;
wire n_255;
wire n_2869;
wire n_5379;
wire n_7079;
wire n_4487;
wire n_5878;
wire n_2674;
wire n_5820;
wire n_1737;
wire n_7309;
wire n_7119;
wire n_1613;
wire n_3026;
wire n_7184;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_7696;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_196;
wire n_3244;
wire n_1779;
wire n_2562;
wire n_954;
wire n_3112;
wire n_2051;
wire n_3196;
wire n_231;
wire n_5964;
wire n_2673;
wire n_6076;
wire n_4678;
wire n_664;
wire n_1591;
wire n_5301;
wire n_5126;
wire n_6732;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_6817;
wire n_1967;
wire n_5776;
wire n_2179;
wire n_1280;
wire n_544;
wire n_7646;
wire n_3779;
wire n_599;
wire n_6982;
wire n_537;
wire n_1063;
wire n_7291;
wire n_991;
wire n_2275;
wire n_7668;
wire n_7435;
wire n_4606;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_5603;
wire n_938;
wire n_1891;
wire n_6560;
wire n_6634;
wire n_5348;
wire n_583;
wire n_1000;
wire n_313;
wire n_4868;
wire n_7017;
wire n_378;
wire n_4072;
wire n_7848;
wire n_2792;
wire n_4465;
wire n_8127;
wire n_2596;
wire n_5217;
wire n_3986;
wire n_5558;
wire n_3725;
wire n_7861;
wire n_472;
wire n_4026;
wire n_4245;
wire n_5520;
wire n_2524;
wire n_7889;
wire n_208;
wire n_3894;
wire n_1702;
wire n_5909;
wire n_4852;
wire n_275;
wire n_7554;
wire n_3202;
wire n_4290;
wire n_4945;
wire n_5750;
wire n_7648;
wire n_147;
wire n_1232;
wire n_1211;
wire n_996;
wire n_1082;
wire n_1725;
wire n_5654;
wire n_2318;
wire n_866;
wire n_2819;
wire n_1722;
wire n_2229;
wire n_7653;
wire n_6400;
wire n_1644;
wire n_7846;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_131;
wire n_2255;
wire n_5554;
wire n_1252;
wire n_3045;
wire n_250;
wire n_773;
wire n_5135;
wire n_7551;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_6655;
wire n_718;
wire n_1434;
wire n_8093;
wire n_1905;
wire n_1569;
wire n_5448;
wire n_2573;
wire n_6480;
wire n_7737;
wire n_5837;
wire n_2336;
wire n_5412;
wire n_523;
wire n_1662;
wire n_3249;
wire n_3483;
wire n_6621;
wire n_6851;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_782;
wire n_2915;
wire n_7606;
wire n_7420;
wire n_8115;
wire n_4869;
wire n_3213;
wire n_5533;
wire n_4047;
wire n_1244;
wire n_1796;
wire n_484;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_6226;
wire n_1574;
wire n_3033;
wire n_893;
wire n_1582;
wire n_8182;
wire n_1981;
wire n_2824;
wire n_7973;
wire n_7545;
wire n_5327;
wire n_4417;
wire n_796;
wire n_127;
wire n_531;
wire n_1374;
wire n_2089;
wire n_7896;
wire n_6283;
wire n_4688;
wire n_7156;
wire n_4939;
wire n_5900;
wire n_8186;
wire n_7319;
wire n_1486;
wire n_3619;
wire n_6158;
wire n_4013;
wire n_3434;
wire n_4342;
wire n_691;
wire n_6819;
wire n_4903;
wire n_6122;
wire n_2131;
wire n_3853;
wire n_8233;
wire n_4382;
wire n_2509;
wire n_423;
wire n_4085;
wire n_6898;
wire n_6570;
wire n_5486;
wire n_2135;
wire n_8282;
wire n_7260;
wire n_6894;
wire n_4475;
wire n_6843;
wire n_5851;
wire n_7516;
wire n_5432;
wire n_6928;
wire n_6317;
wire n_6707;
wire n_7244;
wire n_187;
wire n_1463;
wire n_4626;
wire n_7625;
wire n_4997;
wire n_8183;
wire n_5065;
wire n_6806;
wire n_924;
wire n_7991;
wire n_781;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_6835;
wire n_7286;
wire n_2436;
wire n_3517;
wire n_6269;
wire n_7857;
wire n_7970;
wire n_1706;
wire n_2461;
wire n_8258;
wire n_3719;
wire n_117;
wire n_7154;
wire n_524;
wire n_634;
wire n_1214;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_5295;
wire n_6088;
wire n_1181;
wire n_1999;
wire n_7194;
wire n_4841;
wire n_4683;
wire n_5173;
wire n_2873;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_5655;
wire n_3383;
wire n_1835;
wire n_7175;
wire n_5855;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_7163;
wire n_3797;
wire n_1836;
wire n_7027;
wire n_3416;
wire n_5861;
wire n_4600;
wire n_1453;
wire n_6964;
wire n_3943;
wire n_3145;
wire n_7964;
wire n_5749;
wire n_6320;
wire n_6316;
wire n_419;
wire n_7068;
wire n_2908;
wire n_270;
wire n_4106;
wire n_285;
wire n_2156;
wire n_1184;
wire n_202;
wire n_8162;
wire n_754;
wire n_2323;
wire n_1073;
wire n_4549;
wire n_7327;
wire n_1277;
wire n_1746;
wire n_6610;
wire n_1062;
wire n_5998;
wire n_4702;
wire n_5102;
wire n_4954;
wire n_740;
wire n_167;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_6752;
wire n_6959;
wire n_6250;
wire n_3283;
wire n_259;
wire n_4331;
wire n_7317;
wire n_4159;
wire n_7864;
wire n_3451;
wire n_8051;
wire n_4734;
wire n_6675;
wire n_7955;
wire n_2832;
wire n_1688;
wire n_5827;
wire n_2370;
wire n_1944;
wire n_7384;
wire n_267;
wire n_2914;
wire n_5656;
wire n_7218;
wire n_1988;
wire n_5678;
wire n_6561;
wire n_6858;
wire n_5865;
wire n_6050;
wire n_7512;
wire n_1718;
wire n_7814;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_200;
wire n_2539;
wire n_5555;
wire n_2078;
wire n_1145;
wire n_4809;
wire n_7152;
wire n_787;
wire n_4012;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_5212;
wire n_4760;
wire n_1207;
wire n_6823;
wire n_3606;
wire n_7062;
wire n_7090;
wire n_8202;
wire n_2232;
wire n_1847;
wire n_5815;
wire n_4320;
wire n_5084;
wire n_7223;
wire n_5251;
wire n_1314;
wire n_1512;
wire n_5965;
wire n_884;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_6796;
wire n_5407;
wire n_2988;
wire n_4560;
wire n_7761;
wire n_8141;
wire n_3230;
wire n_3793;
wire n_859;
wire n_5042;
wire n_8199;
wire n_7055;
wire n_6024;
wire n_4768;
wire n_1889;
wire n_6090;
wire n_693;
wire n_5368;
wire n_929;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_8004;
wire n_3607;
wire n_1637;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_7388;
wire n_1751;
wire n_7056;
wire n_7437;
wire n_6489;
wire n_5310;
wire n_2769;
wire n_438;
wire n_1548;
wire n_4987;
wire n_6714;
wire n_440;
wire n_7849;
wire n_7726;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_7417;
wire n_2739;
wire n_3962;
wire n_4988;
wire n_7446;
wire n_6038;
wire n_2902;
wire n_6030;
wire n_6245;
wire n_4360;
wire n_1544;
wire n_6791;
wire n_6620;
wire n_4540;
wire n_6821;
wire n_2094;
wire n_5588;
wire n_3854;
wire n_8198;
wire n_1354;
wire n_6583;
wire n_2349;
wire n_3652;
wire n_7859;
wire n_3449;
wire n_1021;
wire n_3089;
wire n_4854;
wire n_491;
wire n_1595;
wire n_8017;
wire n_1142;
wire n_5477;
wire n_260;
wire n_2727;
wire n_942;
wire n_7523;
wire n_5234;
wire n_1416;
wire n_6890;
wire n_7559;
wire n_7576;
wire n_6988;
wire n_1599;
wire n_5871;
wire n_4747;
wire n_8000;
wire n_3472;
wire n_2527;
wire n_6052;
wire n_7769;
wire n_7257;
wire n_3126;
wire n_2759;
wire n_6973;
wire n_5007;
wire n_4881;
wire n_2038;
wire n_6488;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_4357;
wire n_7729;
wire n_2806;
wire n_4502;
wire n_287;
wire n_3191;
wire n_1716;
wire n_302;
wire n_7005;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_7081;
wire n_7742;
wire n_5253;
wire n_3588;
wire n_355;
wire n_6280;
wire n_1590;
wire n_3280;
wire n_4115;
wire n_5274;
wire n_6399;
wire n_5418;
wire n_5019;
wire n_5939;
wire n_1819;
wire n_135;
wire n_3095;
wire n_947;
wire n_7341;
wire n_5792;
wire n_3698;
wire n_4513;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_4775;
wire n_6256;
wire n_482;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_8250;
wire n_7264;
wire n_7842;
wire n_2499;
wire n_2549;
wire n_6648;
wire n_7492;
wire n_804;
wire n_6649;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_6910;
wire n_3885;
wire n_955;
wire n_4264;
wire n_5954;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_514;
wire n_6431;
wire n_418;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_8266;
wire n_3839;
wire n_7285;
wire n_5490;
wire n_5694;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_6324;
wire n_5489;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_3120;
wire n_6512;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_4794;
wire n_4843;
wire n_669;
wire n_5580;
wire n_5215;
wire n_337;
wire n_437;
wire n_3937;
wire n_4763;
wire n_1418;
wire n_6243;
wire n_5795;
wire n_5715;
wire n_4170;
wire n_5561;
wire n_8267;
wire n_2462;
wire n_7051;
wire n_6773;
wire n_2155;
wire n_6231;
wire n_615;
wire n_7503;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_517;
wire n_8124;
wire n_3604;
wire n_5430;
wire n_6041;
wire n_824;
wire n_159;
wire n_7997;
wire n_5659;
wire n_6859;
wire n_7716;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_144;
wire n_3792;
wire n_7950;
wire n_6323;
wire n_5720;
wire n_4267;
wire n_8214;
wire n_7793;
wire n_2083;
wire n_815;
wire n_5598;
wire n_2753;
wire n_1340;
wire n_470;
wire n_3021;
wire n_7746;
wire n_477;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_7570;
wire n_2898;
wire n_1825;
wire n_6912;
wire n_3567;
wire n_7425;
wire n_2682;
wire n_5854;
wire n_5958;
wire n_5585;
wire n_5112;
wire n_5326;
wire n_1627;
wire n_5783;
wire n_7829;
wire n_6837;
wire n_6747;
wire n_2903;
wire n_5303;
wire n_3812;
wire n_3127;
wire n_6916;
wire n_1731;
wire n_799;
wire n_7894;
wire n_1147;
wire n_7957;
wire n_8262;
wire n_2378;
wire n_5530;
wire n_6718;
wire n_8289;
wire n_965;
wire n_5809;
wire n_934;
wire n_2213;
wire n_7121;
wire n_7531;
wire n_6410;
wire n_356;
wire n_6473;
wire n_8087;
wire n_4056;
wire n_4806;
wire n_7961;
wire n_1674;
wire n_5993;
wire n_4015;
wire n_6574;
wire n_2924;
wire n_6492;
wire n_4445;
wire n_7687;
wire n_4462;
wire n_5299;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_1042;
wire n_3170;
wire n_2311;
wire n_6857;
wire n_1455;
wire n_2287;
wire n_836;
wire n_3415;
wire n_6975;
wire n_7763;
wire n_3464;
wire n_6290;
wire n_3414;
wire n_6646;
wire n_205;
wire n_7703;
wire n_7928;
wire n_4234;
wire n_760;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_3467;
wire n_5821;
wire n_713;
wire n_3179;
wire n_598;
wire n_6622;
wire n_5522;
wire n_4836;
wire n_3889;
wire n_7665;
wire n_5262;
wire n_7677;
wire n_3262;
wire n_5319;
wire n_927;
wire n_7469;
wire n_261;
wire n_3699;
wire n_6118;
wire n_706;
wire n_2120;
wire n_7125;
wire n_7856;
wire n_6028;
wire n_6663;
wire n_6532;
wire n_1419;
wire n_3816;
wire n_8099;
wire n_3528;
wire n_6267;
wire n_6682;
wire n_4207;
wire n_8085;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_4725;
wire n_348;
wire n_2312;
wire n_7203;
wire n_7797;
wire n_1826;
wire n_5943;
wire n_6556;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_6216;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_637;
wire n_7128;
wire n_5335;
wire n_1259;
wire n_6365;
wire n_7111;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_5284;
wire n_4978;
wire n_5771;
wire n_3246;
wire n_3299;
wire n_980;
wire n_1618;
wire n_1869;
wire n_3623;
wire n_905;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_6950;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_5516;
wire n_7284;
wire n_3615;
wire n_8276;
wire n_7057;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_3200;
wire n_6167;
wire n_3642;
wire n_145;
wire n_2146;
wire n_5583;
wire n_4274;
wire n_3276;
wire n_7064;
wire n_5433;
wire n_3682;
wire n_7278;
wire n_5429;
wire n_6772;
wire n_7088;
wire n_7799;
wire n_5698;
wire n_5731;
wire n_4007;
wire n_1456;
wire n_1879;
wire n_6159;
wire n_2129;
wire n_5857;
wire n_7048;
wire n_7979;
wire n_6617;
wire n_553;
wire n_7725;
wire n_814;
wire n_578;
wire n_5120;
wire n_3572;
wire n_2975;
wire n_2399;
wire n_1134;
wire n_4075;
wire n_3471;
wire n_1484;
wire n_647;
wire n_2027;
wire n_2932;
wire n_6217;
wire n_600;
wire n_3118;
wire n_5560;
wire n_4441;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_5455;
wire n_502;
wire n_6777;
wire n_6742;
wire n_1467;
wire n_7447;
wire n_5209;
wire n_247;
wire n_6307;
wire n_5704;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_5916;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_6479;
wire n_5099;
wire n_681;
wire n_3286;
wire n_5781;
wire n_5619;
wire n_2023;
wire n_3974;
wire n_7365;
wire n_3443;
wire n_2599;
wire n_3988;
wire n_7792;
wire n_5022;
wire n_8089;
wire n_6370;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_7275;
wire n_5353;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_6856;
wire n_1098;
wire n_3009;
wire n_777;
wire n_7095;
wire n_7390;
wire n_6140;
wire n_6111;
wire n_5219;
wire n_920;
wire n_3951;
wire n_5518;
wire n_3035;
wire n_4261;
wire n_7037;
wire n_1132;
wire n_8125;
wire n_501;
wire n_1823;
wire n_6240;
wire n_5236;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_6693;
wire n_6712;
wire n_7530;
wire n_1402;
wire n_3957;
wire n_3418;
wire n_1607;
wire n_7471;
wire n_6465;
wire n_221;
wire n_8188;
wire n_5673;
wire n_861;
wire n_5814;
wire n_1666;
wire n_6586;
wire n_7058;
wire n_5103;
wire n_4648;
wire n_8011;
wire n_2214;
wire n_6730;
wire n_6367;
wire n_2256;
wire n_281;
wire n_3326;
wire n_262;
wire n_8222;
wire n_6069;
wire n_2732;
wire n_1883;
wire n_6515;
wire n_8206;
wire n_4094;
wire n_2776;
wire n_6077;
wire n_3224;
wire n_1969;
wire n_5671;
wire n_7429;
wire n_6940;
wire n_8065;
wire n_527;
wire n_2949;
wire n_7008;
wire n_6468;
wire n_7709;
wire n_4269;
wire n_1927;
wire n_7540;
wire n_7581;
wire n_343;
wire n_1222;
wire n_7139;
wire n_3803;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_7782;
wire n_7432;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_8155;
wire n_2449;
wire n_4428;
wire n_745;
wire n_6483;
wire n_1572;
wire n_7770;
wire n_4463;
wire n_5357;
wire n_8175;
wire n_7173;
wire n_3648;
wire n_6576;
wire n_6810;
wire n_1975;
wire n_5421;
wire n_1388;
wire n_1266;
wire n_4396;
wire n_1990;
wire n_6708;
wire n_8026;
wire n_6667;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1075;
wire n_6040;
wire n_1890;
wire n_6847;
wire n_6305;
wire n_4034;
wire n_4228;
wire n_1227;
wire n_7251;
wire n_3166;
wire n_7356;
wire n_3649;
wire n_7412;
wire n_3065;
wire n_8168;
wire n_7212;
wire n_5045;
wire n_5237;
wire n_7751;
wire n_7951;
wire n_657;
wire n_7060;
wire n_3924;
wire n_3997;
wire n_7591;
wire n_3564;
wire n_862;
wire n_6750;
wire n_2637;
wire n_5769;
wire n_7444;
wire n_7911;
wire n_3795;
wire n_7595;
wire n_4931;
wire n_2306;
wire n_7790;
wire n_2071;
wire n_7426;
wire n_430;
wire n_3953;
wire n_7502;
wire n_4400;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_5434;
wire n_1532;
wire n_6855;
wire n_8170;
wire n_1030;
wire n_5181;
wire n_6239;
wire n_3208;
wire n_5768;
wire n_1342;
wire n_6199;
wire n_2737;
wire n_3282;
wire n_8120;
wire n_852;
wire n_2916;
wire n_7252;
wire n_1060;
wire n_5963;
wire n_4424;
wire n_4351;
wire n_6543;
wire n_7532;
wire n_4192;
wire n_8003;
wire n_1748;
wire n_1301;
wire n_6789;
wire n_5972;
wire n_3400;
wire n_7065;
wire n_1466;
wire n_8083;
wire n_6177;
wire n_8057;
wire n_2581;
wire n_5937;
wire n_1783;
wire n_5146;
wire n_7367;
wire n_8164;
wire n_7267;
wire n_7405;
wire n_4646;
wire n_4221;
wire n_1037;
wire n_3650;
wire n_1329;
wire n_6825;
wire n_7614;
wire n_1993;
wire n_1545;
wire n_6460;
wire n_134;
wire n_4035;
wire n_6952;
wire n_1480;
wire n_3670;
wire n_6173;
wire n_2540;
wire n_4190;
wire n_1605;
wire n_3060;
wire n_6218;
wire n_7685;
wire n_6486;
wire n_2984;
wire n_4009;
wire n_157;
wire n_7619;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_6852;
wire n_624;
wire n_5577;
wire n_876;
wire n_5872;
wire n_7883;
wire n_6692;
wire n_5017;
wire n_736;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_7220;
wire n_7560;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_5976;
wire n_4717;
wire n_6888;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_602;
wire n_854;
wire n_8256;
wire n_2091;
wire n_393;
wire n_4312;
wire n_5424;
wire n_3789;
wire n_7270;
wire n_1658;
wire n_1072;
wire n_1305;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_2725;
wire n_2667;
wire n_3746;
wire n_7731;
wire n_6626;
wire n_4537;
wire n_1046;
wire n_5838;
wire n_7034;
wire n_3694;
wire n_6854;
wire n_7940;
wire n_771;
wire n_6793;
wire n_5456;
wire n_3893;
wire n_4847;
wire n_5846;
wire n_2307;
wire n_421;
wire n_3702;
wire n_5930;
wire n_1984;
wire n_3453;
wire n_1556;
wire n_7537;
wire n_6980;
wire n_7040;
wire n_5345;
wire n_2815;
wire n_4427;
wire n_7458;
wire n_1824;
wire n_7740;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_6794;
wire n_819;
wire n_1971;
wire n_2945;
wire n_586;
wire n_1324;
wire n_3543;
wire n_7179;
wire n_1776;
wire n_3448;
wire n_7433;
wire n_4279;
wire n_605;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_6334;
wire n_6257;
wire n_4152;
wire n_6874;
wire n_5537;
wire n_2698;
wire n_5572;
wire n_4783;
wire n_7658;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_5409;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_807;
wire n_5142;
wire n_6355;
wire n_7015;
wire n_6039;
wire n_6286;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_7226;
wire n_7987;
wire n_1987;
wire n_7217;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_6377;
wire n_802;
wire n_5401;
wire n_4595;
wire n_960;
wire n_7272;
wire n_8215;
wire n_2352;
wire n_5201;
wire n_5816;
wire n_790;
wire n_5551;
wire n_5416;
wire n_4404;
wire n_2377;
wire n_151;
wire n_7906;
wire n_2652;
wire n_5498;
wire n_5543;
wire n_4054;
wire n_6018;
wire n_7765;
wire n_1286;
wire n_6021;
wire n_4617;
wire n_1685;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_5797;
wire n_6511;
wire n_7815;
wire n_1052;
wire n_4732;
wire n_2076;
wire n_2203;
wire n_5942;
wire n_5764;
wire n_1426;
wire n_4969;
wire n_8121;
wire n_5252;
wire n_5777;
wire n_7785;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_6867;
wire n_4140;
wire n_5171;
wire n_566;
wire n_7728;
wire n_8280;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_7255;
wire n_3309;
wire n_169;
wire n_7181;
wire n_173;
wire n_2796;
wire n_858;
wire n_5393;
wire n_4817;
wire n_6863;
wire n_7352;
wire n_7355;
wire n_2136;
wire n_433;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_7328;
wire n_2771;
wire n_6322;
wire n_7359;
wire n_2403;
wire n_2947;
wire n_5643;
wire n_253;
wire n_928;
wire n_3769;
wire n_7825;
wire n_1565;
wire n_4437;
wire n_6419;
wire n_128;
wire n_7916;
wire n_3055;
wire n_8194;
wire n_420;
wire n_4070;
wire n_5346;
wire n_7283;
wire n_748;
wire n_7903;
wire n_7089;
wire n_1045;
wire n_8217;
wire n_1881;
wire n_2635;
wire n_7604;
wire n_7647;
wire n_2999;
wire n_988;
wire n_4139;
wire n_4769;
wire n_6130;
wire n_330;
wire n_5868;
wire n_6417;
wire n_328;
wire n_368;
wire n_8285;
wire n_7145;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_7803;
wire n_2713;
wire n_1422;
wire n_1965;
wire n_644;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_6979;
wire n_5986;
wire n_6932;
wire n_2934;
wire n_7258;
wire n_5104;
wire n_6961;
wire n_576;
wire n_511;
wire n_7622;
wire n_429;
wire n_7839;
wire n_6792;
wire n_7720;
wire n_2210;
wire n_4368;
wire n_5794;
wire n_8136;
wire n_3141;
wire n_2053;
wire n_5272;
wire n_3476;
wire n_6919;
wire n_1049;
wire n_141;
wire n_4430;
wire n_6123;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_7440;
wire n_1356;
wire n_6831;
wire n_1773;
wire n_3175;
wire n_4544;
wire n_2666;
wire n_5578;
wire n_312;
wire n_728;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_7809;
wire n_3255;
wire n_2588;
wire n_5722;
wire n_5811;
wire n_935;
wire n_7072;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_911;
wire n_623;
wire n_3509;
wire n_1403;
wire n_5395;
wire n_453;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_6458;
wire n_543;
wire n_6986;
wire n_3456;
wire n_4532;
wire n_236;
wire n_601;
wire n_7564;
wire n_628;
wire n_5863;
wire n_8185;
wire n_6633;
wire n_3790;
wire n_7775;
wire n_907;
wire n_7118;
wire n_7960;
wire n_6152;
wire n_5734;
wire n_8281;
wire n_847;
wire n_747;
wire n_1135;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_107;
wire n_6169;
wire n_5774;
wire n_7069;
wire n_5199;
wire n_6546;
wire n_4257;
wire n_4282;
wire n_7636;
wire n_4341;
wire n_1694;
wire n_6925;
wire n_7186;
wire n_593;
wire n_1695;
wire n_4027;
wire n_4309;
wire n_5480;
wire n_4650;
wire n_6428;
wire n_609;
wire n_6924;
wire n_3077;
wire n_4944;
wire n_8066;
wire n_7666;
wire n_6425;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_4994;
wire n_7967;
wire n_5977;
wire n_519;
wire n_384;
wire n_3533;
wire n_5175;
wire n_7246;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_3409;
wire n_4381;
wire n_8239;
wire n_3583;
wire n_4316;
wire n_7301;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_1157;
wire n_7262;
wire n_234;
wire n_5959;
wire n_8056;
wire n_8210;
wire n_3563;
wire n_5945;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_3689;
wire n_7584;
wire n_7748;
wire n_1789;
wire n_763;
wire n_6301;
wire n_2174;
wire n_540;
wire n_5668;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_1687;
wire n_6282;
wire n_7686;
wire n_4934;
wire n_4703;
wire n_2638;
wire n_2046;
wire n_7059;
wire n_6985;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_5600;
wire n_395;
wire n_6737;
wire n_1587;
wire n_213;
wire n_2340;
wire n_4804;
wire n_2444;
wire n_4888;
wire n_1014;
wire n_5767;
wire n_6459;
wire n_1427;
wire n_7670;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_2199;
wire n_6384;
wire n_4669;
wire n_114;
wire n_5228;
wire n_1100;
wire n_585;
wire n_1617;
wire n_2600;
wire n_7443;
wire n_3436;
wire n_5973;
wire n_7484;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_5869;
wire n_5914;
wire n_2114;
wire n_6753;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_1175;
wire n_4887;
wire n_3751;
wire n_3402;
wire n_1621;
wire n_6448;
wire n_5186;
wire n_7930;
wire n_7487;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_580;
wire n_3664;
wire n_4218;
wire n_434;
wire n_4687;
wire n_7077;
wire n_394;
wire n_1381;
wire n_3686;
wire n_1183;
wire n_4720;
wire n_2889;
wire n_6043;
wire n_6268;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_5604;
wire n_3470;
wire n_243;
wire n_7663;
wire n_5221;
wire n_7024;
wire n_1407;
wire n_8148;
wire n_6145;
wire n_2865;
wire n_5925;
wire n_6529;
wire n_973;
wire n_5591;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_8236;
wire n_7214;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_1176;
wire n_3677;
wire n_1054;
wire n_7977;
wire n_121;
wire n_5387;
wire n_3292;
wire n_6311;
wire n_8167;
wire n_3989;
wire n_7652;
wire n_4644;
wire n_4752;
wire n_4746;
wire n_7566;
wire n_1057;
wire n_4131;
wire n_5449;
wire n_4215;
wire n_978;
wire n_2488;
wire n_1509;
wire n_828;
wire n_6134;
wire n_322;
wire n_4158;
wire n_6812;
wire n_3079;
wire n_5190;
wire n_6733;
wire n_3269;
wire n_558;
wire n_5325;
wire n_4231;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_653;
wire n_6262;
wire n_4926;
wire n_2050;
wire n_8207;
wire n_6938;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_5876;
wire n_5344;
wire n_2550;
wire n_556;
wire n_170;
wire n_1536;
wire n_3177;
wire n_6160;
wire n_4667;
wire n_5813;
wire n_6235;
wire n_1471;
wire n_6212;
wire n_3440;
wire n_6816;
wire n_3658;
wire n_7374;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1620;
wire n_2542;
wire n_5892;
wire n_7678;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_788;
wire n_7110;
wire n_5714;
wire n_2169;
wire n_6953;
wire n_7975;
wire n_6089;
wire n_591;
wire n_5634;
wire n_5133;
wire n_7553;
wire n_5305;
wire n_7086;
wire n_2175;
wire n_1625;
wire n_5990;
wire n_5689;
wire n_7732;
wire n_7891;
wire n_4578;
wire n_318;
wire n_5644;
wire n_3644;
wire n_8038;
wire n_8190;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_6138;
wire n_528;
wire n_1922;
wire n_940;
wire n_1537;
wire n_4877;
wire n_2065;
wire n_8179;
wire n_7038;
wire n_7994;
wire n_4470;
wire n_4187;
wire n_8287;
wire n_1904;
wire n_8111;
wire n_4998;
wire n_5576;
wire n_2395;
wire n_2868;
wire n_7345;
wire n_1530;
wire n_4057;
wire n_6070;
wire n_5852;
wire n_5918;
wire n_631;
wire n_8021;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_7041;
wire n_6717;
wire n_7593;
wire n_8265;
wire n_898;
wire n_6881;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_6871;
wire n_2967;
wire n_5343;
wire n_6672;
wire n_7757;
wire n_1093;
wire n_8251;
wire n_7866;
wire n_6518;
wire n_7334;
wire n_4021;
wire n_6396;
wire n_7028;
wire n_3379;
wire n_4379;
wire n_5947;
wire n_6242;
wire n_336;
wire n_6601;
wire n_2268;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_5835;
wire n_668;
wire n_2111;
wire n_3743;
wire n_8079;
wire n_5542;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_5527;
wire n_2897;
wire n_4812;
wire n_4497;
wire n_6606;
wire n_2583;
wire n_8291;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_701;
wire n_1003;
wire n_7758;
wire n_4472;
wire n_2699;
wire n_5819;
wire n_3901;
wire n_291;
wire n_5180;
wire n_1640;
wire n_2973;
wire n_5893;
wire n_2710;
wire n_7705;
wire n_6092;
wire n_6462;
wire n_2505;
wire n_4519;
wire n_5025;
wire n_2397;
wire n_240;
wire n_369;
wire n_7333;
wire n_3878;
wire n_4197;
wire n_6669;
wire n_8006;
wire n_2721;
wire n_1892;
wire n_6251;
wire n_2615;
wire n_4787;
wire n_8218;
wire n_1212;
wire n_7337;
wire n_4310;
wire n_5726;
wire n_3933;
wire n_7439;
wire n_4566;
wire n_4371;
wire n_188;
wire n_1902;
wire n_5828;
wire n_2784;
wire n_7210;
wire n_7744;
wire n_3898;
wire n_694;
wire n_6228;
wire n_6702;
wire n_7358;
wire n_8240;
wire n_4749;
wire n_7707;
wire n_5924;
wire n_1845;
wire n_7733;
wire n_921;
wire n_5545;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_5083;
wire n_7684;
wire n_3253;
wire n_2088;
wire n_1275;
wire n_6997;
wire n_4238;
wire n_6371;
wire n_904;
wire n_7673;
wire n_2005;
wire n_1696;
wire n_7187;
wire n_8013;
wire n_2108;
wire n_3824;
wire n_2246;
wire n_7313;
wire n_5899;
wire n_3846;
wire n_5122;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_6641;
wire n_3845;
wire n_6463;
wire n_3203;
wire n_383;
wire n_4986;
wire n_1316;
wire n_4668;
wire n_950;
wire n_711;
wire n_6264;
wire n_5782;
wire n_8119;
wire n_630;
wire n_4168;
wire n_1369;
wire n_7036;
wire n_4298;
wire n_7370;
wire n_7931;
wire n_4743;
wire n_1781;
wire n_4250;
wire n_3143;
wire n_8044;
wire n_3690;
wire n_3229;
wire n_5864;
wire n_235;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_5637;
wire n_4211;
wire n_6084;
wire n_3094;
wire n_741;
wire n_7480;
wire n_371;
wire n_5185;
wire n_2964;
wire n_308;
wire n_5032;
wire n_6990;
wire n_865;
wire n_7071;
wire n_3312;
wire n_5034;
wire n_1041;
wire n_2451;
wire n_2913;
wire n_6288;
wire n_993;
wire n_1862;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_7380;
wire n_2839;
wire n_3237;
wire n_7708;
wire n_4128;
wire n_4036;
wire n_5269;
wire n_3655;
wire n_2955;
wire n_5709;
wire n_1764;
wire n_4807;
wire n_6277;
wire n_5115;
wire n_7376;
wire n_902;
wire n_1723;
wire n_3918;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_596;
wire n_6409;
wire n_4095;
wire n_1310;
wire n_5927;
wire n_4485;
wire n_7657;
wire n_6388;
wire n_574;
wire n_3593;
wire n_6839;
wire n_5163;
wire n_1229;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_1896;
wire n_6864;
wire n_1516;
wire n_4890;
wire n_8084;
wire n_2485;
wire n_6679;
wire n_6051;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_8219;
wire n_5507;
wire n_195;
wire n_4573;
wire n_1328;
wire n_4943;
wire n_2875;
wire n_6599;
wire n_3519;
wire n_2209;
wire n_7504;
wire n_4042;
wire n_7099;
wire n_7586;
wire n_4244;
wire n_1928;
wire n_5642;
wire n_4708;
wire n_4883;
wire n_6227;
wire n_4553;
wire n_7052;
wire n_1634;
wire n_1203;
wire n_1699;
wire n_6738;
wire n_5226;
wire n_2081;
wire n_937;
wire n_1474;
wire n_1631;
wire n_7602;
wire n_156;
wire n_6566;
wire n_1794;
wire n_5696;
wire n_7998;
wire n_1375;
wire n_3053;
wire n_5014;
wire n_7106;
wire n_6346;
wire n_204;
wire n_7557;
wire n_3772;
wire n_7408;
wire n_2891;
wire n_496;
wire n_4335;
wire n_7026;
wire n_3128;
wire n_6146;
wire n_5677;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_1002;
wire n_7394;
wire n_263;
wire n_4516;
wire n_5235;
wire n_360;
wire n_1129;
wire n_7627;
wire n_6436;
wire n_1464;
wire n_7719;
wire n_2798;
wire n_7450;
wire n_165;
wire n_3217;
wire n_6081;
wire n_1249;
wire n_329;
wire n_7852;
wire n_5724;
wire n_3821;
wire n_340;
wire n_3201;
wire n_7462;
wire n_7780;
wire n_3503;
wire n_5979;
wire n_6027;
wire n_1870;
wire n_4467;
wire n_177;
wire n_364;
wire n_258;
wire n_7582;
wire n_5521;
wire n_431;
wire n_2654;
wire n_7421;
wire n_3935;
wire n_1861;
wire n_1228;
wire n_2319;
wire n_2965;
wire n_4955;
wire n_7555;
wire n_5410;
wire n_1251;
wire n_1989;
wire n_447;
wire n_2689;
wire n_6110;
wire n_1762;
wire n_6238;
wire n_7025;
wire n_3798;
wire n_3080;
wire n_5241;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_5331;
wire n_7478;
wire n_3308;
wire n_6326;
wire n_841;
wire n_3204;
wire n_7451;
wire n_4134;
wire n_5018;
wire n_6917;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;
wire n_6612;
wire n_5258;

BUFx3_ASAP7_75t_L g107 ( 
.A(n_37),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_78),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_35),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_61),
.Y(n_112)
);

INVxp67_ASAP7_75t_SL g113 ( 
.A(n_52),
.Y(n_113)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_73),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_30),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_43),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_92),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_37),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_93),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_83),
.Y(n_122)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_73),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_65),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_40),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_24),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_96),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_57),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_29),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_106),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_103),
.Y(n_131)
);

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_24),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_70),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_14),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_23),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_8),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_33),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_71),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_18),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_42),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_94),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_11),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_59),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_34),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_6),
.Y(n_146)
);

BUFx10_ASAP7_75t_L g147 ( 
.A(n_29),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_19),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_43),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_98),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_7),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_20),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_86),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_47),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_19),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_53),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_95),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_52),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_39),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_51),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_51),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_32),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_34),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_42),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_5),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_22),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_41),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_70),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_62),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_72),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_33),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_15),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_36),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_62),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_20),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_71),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_2),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_13),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_8),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_4),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_91),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_18),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_60),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_13),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_47),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_23),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_3),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_41),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_6),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_66),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_1),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_15),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_22),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_101),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_30),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_10),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_84),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_1),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_3),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_61),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_11),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_68),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_27),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_64),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_100),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_104),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_69),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_4),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_27),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_36),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_46),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_192),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_148),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_160),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_148),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_111),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_152),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

INVxp67_ASAP7_75t_SL g222 ( 
.A(n_142),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_111),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_192),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_142),
.Y(n_225)
);

INVxp33_ASAP7_75t_SL g226 ( 
.A(n_160),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_152),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_142),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_143),
.Y(n_229)
);

INVxp67_ASAP7_75t_SL g230 ( 
.A(n_143),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_167),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_153),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_143),
.Y(n_233)
);

INVxp33_ASAP7_75t_L g234 ( 
.A(n_160),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_167),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_153),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_107),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_179),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_109),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_179),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_179),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_118),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_109),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_107),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_223),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_216),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_107),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g249 ( 
.A(n_214),
.Y(n_249)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_223),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_214),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_223),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_118),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_121),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_223),
.Y(n_257)
);

AND2x4_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_218),
.Y(n_258)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_223),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_215),
.Y(n_260)
);

AND2x4_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_163),
.Y(n_261)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_223),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_215),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_223),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_218),
.Y(n_265)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_218),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_218),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_213),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_215),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_121),
.Y(n_270)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_237),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_213),
.B(n_144),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_213),
.Y(n_273)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_237),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_217),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_237),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_217),
.B(n_144),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_217),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_219),
.B(n_150),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_219),
.B(n_150),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_219),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g282 ( 
.A(n_258),
.B(n_243),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_247),
.B(n_237),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_278),
.Y(n_285)
);

INVx6_ASAP7_75t_L g286 ( 
.A(n_261),
.Y(n_286)
);

AND2x4_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_274),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_278),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_278),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_265),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_265),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_265),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_268),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_244),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_268),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_247),
.B(n_243),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_265),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_268),
.Y(n_300)
);

AND2x4_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_222),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_258),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_276),
.B(n_243),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_247),
.B(n_234),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_249),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_260),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_271),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_247),
.B(n_234),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_244),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_268),
.B(n_221),
.Y(n_310)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_244),
.Y(n_311)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_244),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_268),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_244),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_268),
.B(n_221),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_268),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_265),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_263),
.A2(n_226),
.B1(n_269),
.B2(n_260),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_271),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_268),
.Y(n_320)
);

BUFx8_ASAP7_75t_L g321 ( 
.A(n_249),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_244),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_268),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_258),
.Y(n_324)
);

AND2x4_ASAP7_75t_L g325 ( 
.A(n_271),
.B(n_222),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_247),
.B(n_222),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_258),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_281),
.B(n_221),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_276),
.B(n_220),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_258),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_244),
.Y(n_331)
);

INVx6_ASAP7_75t_L g332 ( 
.A(n_261),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_281),
.B(n_252),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_265),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_244),
.Y(n_335)
);

OA21x2_ASAP7_75t_L g336 ( 
.A1(n_272),
.A2(n_158),
.B(n_151),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_258),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_258),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_258),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_258),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_265),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_265),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_258),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_260),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_245),
.B(n_230),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_281),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_281),
.Y(n_347)
);

AND2x6_ASAP7_75t_L g348 ( 
.A(n_261),
.B(n_111),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_263),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_281),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_265),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_263),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_265),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_265),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_281),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_281),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_252),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_276),
.B(n_220),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_252),
.B(n_224),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_252),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_265),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_273),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_276),
.B(n_224),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_273),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_261),
.B(n_254),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_263),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_265),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_273),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_244),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_265),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_271),
.B(n_239),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_261),
.B(n_224),
.Y(n_372)
);

AND2x4_ASAP7_75t_L g373 ( 
.A(n_271),
.B(n_230),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_267),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_267),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_273),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_261),
.B(n_230),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_245),
.B(n_220),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_273),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_269),
.A2(n_232),
.B1(n_236),
.B2(n_175),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_273),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_261),
.B(n_227),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_261),
.Y(n_383)
);

AND2x2_ASAP7_75t_SL g384 ( 
.A(n_269),
.B(n_111),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_244),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_269),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_245),
.B(n_248),
.Y(n_387)
);

NAND2x1_ASAP7_75t_L g388 ( 
.A(n_261),
.B(n_111),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_273),
.Y(n_389)
);

NAND2xp33_ASAP7_75t_SL g390 ( 
.A(n_253),
.B(n_141),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_245),
.B(n_227),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_245),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_273),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_285),
.Y(n_394)
);

NAND3xp33_ASAP7_75t_L g395 ( 
.A(n_324),
.B(n_279),
.C(n_277),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_384),
.B(n_253),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_285),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_288),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_384),
.B(n_253),
.Y(n_399)
);

NAND2xp33_ASAP7_75t_SL g400 ( 
.A(n_386),
.B(n_253),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_346),
.B(n_255),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_288),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_289),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_346),
.B(n_255),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_289),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_293),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_293),
.Y(n_407)
);

INVxp33_ASAP7_75t_SL g408 ( 
.A(n_349),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_357),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_357),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_384),
.B(n_245),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_287),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_360),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_384),
.B(n_253),
.Y(n_414)
);

CKINVDCx11_ASAP7_75t_R g415 ( 
.A(n_366),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_303),
.B(n_249),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_360),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_306),
.B(n_239),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_347),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_L g420 ( 
.A1(n_336),
.A2(n_226),
.B1(n_271),
.B2(n_274),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_347),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_350),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_350),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_355),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_355),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_356),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_282),
.B(n_273),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_356),
.Y(n_428)
);

AO21x2_ASAP7_75t_L g429 ( 
.A1(n_303),
.A2(n_256),
.B(n_255),
.Y(n_429)
);

BUFx6f_ASAP7_75t_SL g430 ( 
.A(n_282),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_294),
.Y(n_431)
);

NAND2xp33_ASAP7_75t_L g432 ( 
.A(n_365),
.B(n_273),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_333),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_333),
.B(n_255),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_294),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_296),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_329),
.B(n_358),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_287),
.Y(n_438)
);

NOR2x1p5_ASAP7_75t_L g439 ( 
.A(n_298),
.B(n_249),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_296),
.Y(n_440)
);

NOR2x1p5_ASAP7_75t_L g441 ( 
.A(n_298),
.B(n_249),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_324),
.B(n_256),
.Y(n_442)
);

INVx2_ASAP7_75t_SL g443 ( 
.A(n_348),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_282),
.B(n_273),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_297),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_328),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_327),
.B(n_256),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_282),
.B(n_273),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_329),
.B(n_358),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_297),
.B(n_273),
.Y(n_450)
);

AOI21x1_ASAP7_75t_L g451 ( 
.A1(n_365),
.A2(n_257),
.B(n_254),
.Y(n_451)
);

OAI22xp33_ASAP7_75t_L g452 ( 
.A1(n_318),
.A2(n_256),
.B1(n_270),
.B2(n_185),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_306),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_328),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_359),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_359),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_300),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_327),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_378),
.B(n_249),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_330),
.B(n_270),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_300),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_302),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_330),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_287),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_313),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_337),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_287),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_306),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_337),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_338),
.Y(n_470)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_305),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_392),
.B(n_249),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_338),
.B(n_270),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_387),
.B(n_248),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_339),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_339),
.Y(n_476)
);

BUFx6f_ASAP7_75t_SL g477 ( 
.A(n_287),
.Y(n_477)
);

BUFx6f_ASAP7_75t_SL g478 ( 
.A(n_348),
.Y(n_478)
);

AND2x6_ASAP7_75t_L g479 ( 
.A(n_321),
.B(n_261),
.Y(n_479)
);

AOI21x1_ASAP7_75t_L g480 ( 
.A1(n_310),
.A2(n_315),
.B(n_364),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_340),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_386),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_313),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_302),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_378),
.B(n_271),
.Y(n_485)
);

INVxp33_ASAP7_75t_L g486 ( 
.A(n_380),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_340),
.B(n_270),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_343),
.Y(n_488)
);

OR2x6_ASAP7_75t_L g489 ( 
.A(n_302),
.B(n_272),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_391),
.B(n_386),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_316),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_302),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_343),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_316),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_391),
.B(n_271),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_310),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_305),
.B(n_271),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_363),
.B(n_277),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_315),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_320),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_320),
.B(n_273),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_323),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_383),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_383),
.Y(n_504)
);

NOR2x1p5_ASAP7_75t_L g505 ( 
.A(n_298),
.B(n_113),
.Y(n_505)
);

AND3x2_ASAP7_75t_L g506 ( 
.A(n_344),
.B(n_113),
.C(n_248),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_323),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_283),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_383),
.Y(n_509)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_348),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_363),
.B(n_277),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_345),
.B(n_279),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_283),
.Y(n_513)
);

INVx2_ASAP7_75t_SL g514 ( 
.A(n_348),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_283),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_372),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_372),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_345),
.B(n_279),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_383),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_345),
.B(n_271),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_387),
.B(n_273),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_341),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_387),
.B(n_275),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_286),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_366),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_286),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_301),
.B(n_275),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_341),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_341),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_348),
.Y(n_530)
);

INVx5_ASAP7_75t_L g531 ( 
.A(n_295),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_392),
.B(n_286),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_286),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_286),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_326),
.B(n_271),
.Y(n_535)
);

OR2x6_ASAP7_75t_L g536 ( 
.A(n_286),
.B(n_332),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_336),
.A2(n_301),
.B1(n_373),
.B2(n_325),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_332),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_332),
.Y(n_539)
);

NAND3xp33_ASAP7_75t_L g540 ( 
.A(n_377),
.B(n_280),
.C(n_272),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_332),
.B(n_248),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_332),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_332),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_388),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_342),
.Y(n_545)
);

NAND3xp33_ASAP7_75t_L g546 ( 
.A(n_377),
.B(n_280),
.C(n_272),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_301),
.B(n_275),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_326),
.B(n_271),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_388),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_307),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_342),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_307),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_321),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_307),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_301),
.B(n_325),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_388),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_301),
.B(n_271),
.Y(n_557)
);

INVx5_ASAP7_75t_L g558 ( 
.A(n_295),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_342),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_351),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_348),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_295),
.Y(n_562)
);

INVx8_ASAP7_75t_L g563 ( 
.A(n_348),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_295),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_325),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_326),
.B(n_271),
.Y(n_566)
);

INVx5_ASAP7_75t_L g567 ( 
.A(n_295),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_325),
.B(n_275),
.Y(n_568)
);

BUFx6f_ASAP7_75t_SL g569 ( 
.A(n_348),
.Y(n_569)
);

NOR2x1p5_ASAP7_75t_L g570 ( 
.A(n_304),
.B(n_235),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_351),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_325),
.B(n_275),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_373),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_373),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_348),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_351),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_375),
.Y(n_577)
);

BUFx10_ASAP7_75t_L g578 ( 
.A(n_373),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_375),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_373),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_336),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_375),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_319),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_304),
.B(n_308),
.Y(n_584)
);

CKINVDCx6p67_ASAP7_75t_R g585 ( 
.A(n_344),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_295),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_290),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_321),
.B(n_275),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_336),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_284),
.B(n_274),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_336),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_318),
.A2(n_168),
.B1(n_175),
.B2(n_185),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g593 ( 
.A(n_352),
.B(n_248),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_336),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_319),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_290),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_319),
.Y(n_597)
);

INVx8_ASAP7_75t_L g598 ( 
.A(n_348),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_352),
.B(n_248),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_290),
.Y(n_600)
);

AND2x6_ASAP7_75t_L g601 ( 
.A(n_321),
.B(n_244),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_284),
.B(n_304),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_290),
.Y(n_603)
);

BUFx10_ASAP7_75t_L g604 ( 
.A(n_321),
.Y(n_604)
);

BUFx10_ASAP7_75t_L g605 ( 
.A(n_364),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_284),
.B(n_274),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_291),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_291),
.Y(n_608)
);

INVxp33_ASAP7_75t_L g609 ( 
.A(n_380),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_308),
.B(n_274),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_382),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_291),
.Y(n_612)
);

AND2x2_ASAP7_75t_SL g613 ( 
.A(n_308),
.B(n_151),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_291),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_292),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_292),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_390),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_382),
.B(n_274),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_292),
.Y(n_619)
);

INVxp33_ASAP7_75t_L g620 ( 
.A(n_390),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_371),
.Y(n_621)
);

BUFx4f_ASAP7_75t_L g622 ( 
.A(n_295),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_295),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_311),
.B(n_275),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_292),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_299),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_299),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_299),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_299),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_317),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_371),
.B(n_274),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_317),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_317),
.Y(n_633)
);

NOR2x1p5_ASAP7_75t_L g634 ( 
.A(n_362),
.B(n_235),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_317),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_311),
.B(n_227),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_334),
.A2(n_274),
.B1(n_205),
.B2(n_168),
.Y(n_637)
);

INVx5_ASAP7_75t_L g638 ( 
.A(n_309),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_334),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_311),
.B(n_275),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_334),
.B(n_274),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_L g642 ( 
.A(n_334),
.B(n_275),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_353),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_353),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_353),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_353),
.B(n_274),
.Y(n_646)
);

INVx5_ASAP7_75t_L g647 ( 
.A(n_309),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_411),
.B(n_274),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_411),
.B(n_274),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_415),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_431),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_411),
.B(n_274),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_397),
.Y(n_653)
);

XNOR2x1_ASAP7_75t_L g654 ( 
.A(n_592),
.B(n_232),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_397),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_437),
.B(n_274),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_585),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_398),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_431),
.Y(n_659)
);

AND2x2_ASAP7_75t_SL g660 ( 
.A(n_613),
.B(n_158),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_398),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_536),
.B(n_274),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_403),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_403),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_405),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_408),
.B(n_236),
.Y(n_666)
);

INVxp33_ASAP7_75t_L g667 ( 
.A(n_525),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_458),
.Y(n_668)
);

AND2x2_ASAP7_75t_SL g669 ( 
.A(n_613),
.B(n_195),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_458),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_463),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_578),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_463),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_466),
.Y(n_674)
);

XNOR2xp5_ASAP7_75t_L g675 ( 
.A(n_592),
.B(n_452),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_431),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_466),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_469),
.Y(n_678)
);

XOR2xp5_ASAP7_75t_L g679 ( 
.A(n_452),
.B(n_205),
.Y(n_679)
);

AND2x2_ASAP7_75t_SL g680 ( 
.A(n_613),
.B(n_195),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_536),
.B(n_274),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_469),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_SL g683 ( 
.A(n_471),
.B(n_141),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_474),
.B(n_280),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_474),
.B(n_280),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_578),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_470),
.Y(n_687)
);

CKINVDCx20_ASAP7_75t_R g688 ( 
.A(n_585),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_L g689 ( 
.A1(n_540),
.A2(n_361),
.B(n_354),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_405),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_406),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_536),
.B(n_225),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_406),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_394),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_620),
.B(n_231),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_437),
.B(n_231),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_510),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_512),
.B(n_231),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_435),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_394),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_474),
.B(n_225),
.Y(n_701)
);

NAND2x1p5_ASAP7_75t_L g702 ( 
.A(n_510),
.B(n_266),
.Y(n_702)
);

INVxp67_ASAP7_75t_SL g703 ( 
.A(n_462),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_394),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_536),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_585),
.B(n_206),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_402),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_402),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_584),
.B(n_512),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_402),
.Y(n_710)
);

INVxp67_ASAP7_75t_SL g711 ( 
.A(n_462),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_525),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_453),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_407),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_578),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_518),
.B(n_311),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_407),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_536),
.B(n_225),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_407),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g720 ( 
.A(n_453),
.B(n_156),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_617),
.B(n_418),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_410),
.Y(n_722)
);

INVxp33_ASAP7_75t_SL g723 ( 
.A(n_468),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_SL g724 ( 
.A(n_471),
.B(n_206),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_410),
.Y(n_725)
);

AND2x6_ASAP7_75t_L g726 ( 
.A(n_553),
.B(n_354),
.Y(n_726)
);

INVxp33_ASAP7_75t_L g727 ( 
.A(n_418),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_584),
.B(n_228),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_435),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_435),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_536),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_462),
.B(n_228),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_413),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_413),
.Y(n_734)
);

BUFx8_ASAP7_75t_L g735 ( 
.A(n_430),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_409),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_409),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_622),
.A2(n_311),
.B(n_354),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_409),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_417),
.Y(n_740)
);

OAI21xp5_ASAP7_75t_L g741 ( 
.A1(n_540),
.A2(n_361),
.B(n_354),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_518),
.B(n_207),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_417),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_417),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_419),
.Y(n_745)
);

NOR2xp67_ASAP7_75t_L g746 ( 
.A(n_418),
.B(n_266),
.Y(n_746)
);

AOI21x1_ASAP7_75t_L g747 ( 
.A1(n_449),
.A2(n_367),
.B(n_361),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_419),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_436),
.Y(n_749)
);

XOR2x2_ASAP7_75t_L g750 ( 
.A(n_637),
.B(n_156),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_423),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_484),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_423),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_436),
.Y(n_754)
);

INVxp33_ASAP7_75t_L g755 ( 
.A(n_468),
.Y(n_755)
);

XNOR2xp5_ASAP7_75t_L g756 ( 
.A(n_486),
.B(n_207),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_424),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_541),
.B(n_188),
.Y(n_758)
);

XOR2xp5_ASAP7_75t_L g759 ( 
.A(n_609),
.B(n_114),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_436),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_424),
.Y(n_761)
);

NOR2xp67_ASAP7_75t_L g762 ( 
.A(n_546),
.B(n_266),
.Y(n_762)
);

XNOR2xp5_ASAP7_75t_L g763 ( 
.A(n_505),
.B(n_114),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_428),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_617),
.B(n_188),
.Y(n_765)
);

INVxp67_ASAP7_75t_SL g766 ( 
.A(n_484),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_428),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_421),
.Y(n_768)
);

OAI21xp5_ASAP7_75t_L g769 ( 
.A1(n_546),
.A2(n_367),
.B(n_361),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_421),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_421),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_422),
.Y(n_772)
);

INVx1_ASAP7_75t_SL g773 ( 
.A(n_482),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_422),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_422),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_425),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_541),
.B(n_203),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_440),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_425),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_425),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_584),
.B(n_228),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_482),
.B(n_203),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_426),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_440),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_426),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_426),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_500),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_498),
.B(n_367),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_500),
.Y(n_789)
);

CKINVDCx20_ASAP7_75t_R g790 ( 
.A(n_400),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_470),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_498),
.B(n_367),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_602),
.B(n_229),
.Y(n_793)
);

AND2x4_ASAP7_75t_L g794 ( 
.A(n_484),
.B(n_229),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_475),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_578),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_475),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_578),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_476),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_476),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_505),
.B(n_229),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_622),
.A2(n_434),
.B(n_404),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_481),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_553),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_481),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_488),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_488),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_440),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_493),
.Y(n_809)
);

NAND2xp33_ASAP7_75t_SL g810 ( 
.A(n_439),
.B(n_112),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_445),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_493),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_445),
.Y(n_813)
);

XOR2xp5_ASAP7_75t_L g814 ( 
.A(n_637),
.B(n_115),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_445),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_599),
.B(n_233),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_565),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_565),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_573),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_573),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_599),
.B(n_489),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_489),
.B(n_233),
.Y(n_822)
);

INVxp33_ASAP7_75t_L g823 ( 
.A(n_570),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_574),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_511),
.B(n_370),
.Y(n_825)
);

XNOR2xp5_ASAP7_75t_L g826 ( 
.A(n_439),
.B(n_115),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_574),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_SL g828 ( 
.A(n_471),
.B(n_147),
.Y(n_828)
);

INVxp67_ASAP7_75t_SL g829 ( 
.A(n_562),
.Y(n_829)
);

INVxp33_ASAP7_75t_L g830 ( 
.A(n_570),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_489),
.B(n_233),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_489),
.B(n_238),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_580),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_580),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_457),
.Y(n_835)
);

CKINVDCx16_ASAP7_75t_R g836 ( 
.A(n_430),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_510),
.B(n_131),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_563),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_489),
.B(n_238),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_489),
.B(n_238),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_516),
.B(n_240),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_457),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_516),
.B(n_240),
.Y(n_843)
);

XOR2xp5_ASAP7_75t_L g844 ( 
.A(n_396),
.B(n_132),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_457),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_461),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_414),
.B(n_132),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_461),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_461),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_618),
.A2(n_374),
.B(n_370),
.Y(n_850)
);

XNOR2xp5_ASAP7_75t_L g851 ( 
.A(n_441),
.B(n_133),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_555),
.B(n_240),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_517),
.B(n_241),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_465),
.Y(n_854)
);

XOR2xp5_ASAP7_75t_L g855 ( 
.A(n_396),
.B(n_133),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_465),
.Y(n_856)
);

XNOR2x2_ASAP7_75t_L g857 ( 
.A(n_399),
.B(n_108),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_465),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_399),
.B(n_136),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_483),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_483),
.Y(n_861)
);

INVxp67_ASAP7_75t_SL g862 ( 
.A(n_562),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_412),
.Y(n_863)
);

INVxp67_ASAP7_75t_L g864 ( 
.A(n_593),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_517),
.B(n_241),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_593),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_483),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_491),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_491),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_491),
.Y(n_870)
);

CKINVDCx16_ASAP7_75t_R g871 ( 
.A(n_430),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_555),
.B(n_241),
.Y(n_872)
);

AND2x2_ASAP7_75t_SL g873 ( 
.A(n_416),
.B(n_108),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_449),
.B(n_136),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_593),
.B(n_275),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_494),
.Y(n_876)
);

XNOR2x2_ASAP7_75t_L g877 ( 
.A(n_416),
.B(n_110),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_494),
.Y(n_878)
);

CKINVDCx16_ASAP7_75t_R g879 ( 
.A(n_430),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_494),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_502),
.Y(n_881)
);

INVx2_ASAP7_75t_SL g882 ( 
.A(n_563),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_511),
.B(n_370),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_502),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_502),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_507),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_507),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_507),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_401),
.Y(n_889)
);

XOR2xp5_ASAP7_75t_L g890 ( 
.A(n_621),
.B(n_537),
.Y(n_890)
);

AND2x6_ASAP7_75t_SL g891 ( 
.A(n_532),
.B(n_110),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_563),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_477),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_490),
.B(n_138),
.Y(n_894)
);

CKINVDCx20_ASAP7_75t_R g895 ( 
.A(n_553),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_401),
.Y(n_896)
);

INVxp33_ASAP7_75t_L g897 ( 
.A(n_532),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_404),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_433),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_433),
.Y(n_900)
);

INVxp33_ASAP7_75t_L g901 ( 
.A(n_610),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_622),
.A2(n_374),
.B(n_370),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_446),
.Y(n_903)
);

XOR2x2_ASAP7_75t_L g904 ( 
.A(n_506),
.B(n_112),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_446),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_454),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_492),
.B(n_138),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_557),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_454),
.Y(n_909)
);

XOR2xp5_ASAP7_75t_L g910 ( 
.A(n_537),
.B(n_395),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_455),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_492),
.B(n_204),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_471),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_477),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_492),
.B(n_204),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_455),
.Y(n_916)
);

XOR2xp5_ASAP7_75t_L g917 ( 
.A(n_395),
.B(n_211),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_456),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_456),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_412),
.B(n_438),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_520),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_520),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_557),
.B(n_374),
.Y(n_923)
);

OR2x2_ASAP7_75t_L g924 ( 
.A(n_610),
.B(n_162),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_521),
.Y(n_925)
);

OR2x2_ASAP7_75t_L g926 ( 
.A(n_590),
.B(n_162),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_492),
.B(n_211),
.Y(n_927)
);

NOR2xp67_ASAP7_75t_L g928 ( 
.A(n_471),
.B(n_266),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_524),
.B(n_526),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_521),
.Y(n_930)
);

XNOR2xp5_ASAP7_75t_L g931 ( 
.A(n_441),
.B(n_116),
.Y(n_931)
);

CKINVDCx20_ASAP7_75t_R g932 ( 
.A(n_604),
.Y(n_932)
);

NAND2x1p5_ASAP7_75t_L g933 ( 
.A(n_510),
.B(n_266),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_523),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_523),
.Y(n_935)
);

XOR2xp5_ASAP7_75t_L g936 ( 
.A(n_420),
.B(n_119),
.Y(n_936)
);

XNOR2xp5_ASAP7_75t_SL g937 ( 
.A(n_506),
.B(n_420),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_477),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_544),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_544),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_549),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_549),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_556),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_524),
.B(n_526),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_556),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_533),
.B(n_123),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_496),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_508),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_496),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_499),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_499),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_434),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_477),
.Y(n_953)
);

XNOR2xp5_ASAP7_75t_L g954 ( 
.A(n_634),
.B(n_124),
.Y(n_954)
);

INVxp33_ASAP7_75t_SL g955 ( 
.A(n_472),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_557),
.B(n_374),
.Y(n_956)
);

CKINVDCx20_ASAP7_75t_R g957 ( 
.A(n_604),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_557),
.B(n_266),
.Y(n_958)
);

XOR2xp5_ASAP7_75t_L g959 ( 
.A(n_557),
.B(n_125),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_412),
.B(n_266),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_533),
.B(n_128),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_503),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_519),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_709),
.B(n_412),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_696),
.A2(n_472),
.B(n_447),
.C(n_460),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_752),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_952),
.B(n_442),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_660),
.B(n_510),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_709),
.B(n_660),
.Y(n_969)
);

O2A1O1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_874),
.A2(n_447),
.B(n_460),
.C(n_442),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_669),
.B(n_438),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_669),
.B(n_530),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_680),
.B(n_530),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_752),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_723),
.B(n_534),
.Y(n_975)
);

AOI22xp33_ASAP7_75t_L g976 ( 
.A1(n_680),
.A2(n_606),
.B1(n_590),
.B2(n_548),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_952),
.B(n_473),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_955),
.B(n_530),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_653),
.Y(n_979)
);

AO221x1_ASAP7_75t_L g980 ( 
.A1(n_877),
.A2(n_212),
.B1(n_209),
.B2(n_134),
.C(n_137),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_684),
.B(n_438),
.Y(n_981)
);

NAND3xp33_ASAP7_75t_L g982 ( 
.A(n_721),
.B(n_495),
.C(n_485),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_653),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_889),
.B(n_473),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_955),
.B(n_530),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_889),
.B(n_487),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_910),
.A2(n_487),
.B1(n_589),
.B2(n_581),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_948),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_896),
.B(n_429),
.Y(n_989)
);

NAND2x1p5_ASAP7_75t_L g990 ( 
.A(n_705),
.B(n_530),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_723),
.B(n_897),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_896),
.B(n_429),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_683),
.B(n_561),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_698),
.A2(n_606),
.B(n_611),
.C(n_459),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_724),
.B(n_561),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_655),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_802),
.A2(n_589),
.B(n_581),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_706),
.B(n_534),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_948),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_684),
.B(n_438),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_773),
.B(n_561),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_672),
.B(n_561),
.Y(n_1002)
);

OR2x2_ASAP7_75t_L g1003 ( 
.A(n_866),
.B(n_429),
.Y(n_1003)
);

BUFx8_ASAP7_75t_L g1004 ( 
.A(n_705),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_898),
.B(n_429),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_672),
.B(n_561),
.Y(n_1006)
);

AND2x6_ASAP7_75t_SL g1007 ( 
.A(n_666),
.B(n_126),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_651),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_898),
.B(n_921),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_921),
.B(n_611),
.Y(n_1010)
);

INVx2_ASAP7_75t_SL g1011 ( 
.A(n_731),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_788),
.A2(n_622),
.B(n_792),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_727),
.B(n_538),
.Y(n_1013)
);

AOI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_873),
.A2(n_444),
.B1(n_448),
.B2(n_427),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_655),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_922),
.B(n_685),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_658),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_742),
.B(n_538),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_750),
.A2(n_675),
.B1(n_679),
.B2(n_814),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_922),
.B(n_611),
.Y(n_1020)
);

OAI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_790),
.A2(n_598),
.B1(n_563),
.B2(n_504),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_685),
.B(n_503),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_658),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_697),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_686),
.B(n_503),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_899),
.B(n_503),
.Y(n_1026)
);

AOI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_873),
.A2(n_444),
.B1(n_448),
.B2(n_427),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_686),
.B(n_504),
.Y(n_1028)
);

INVx2_ASAP7_75t_SL g1029 ( 
.A(n_731),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_697),
.Y(n_1030)
);

AOI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_750),
.A2(n_548),
.B1(n_566),
.B2(n_535),
.Y(n_1031)
);

INVx2_ASAP7_75t_SL g1032 ( 
.A(n_893),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_675),
.B(n_539),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_899),
.B(n_504),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_765),
.B(n_539),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_651),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_864),
.B(n_542),
.Y(n_1037)
);

AOI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_679),
.A2(n_566),
.B1(n_535),
.B2(n_464),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_661),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_958),
.B(n_464),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_661),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_910),
.A2(n_509),
.B1(n_504),
.B2(n_519),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_890),
.B(n_542),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_890),
.B(n_758),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_755),
.B(n_543),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_814),
.A2(n_464),
.B1(n_467),
.B2(n_631),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_659),
.Y(n_1047)
);

NAND2xp33_ASAP7_75t_SL g1048 ( 
.A(n_715),
.B(n_478),
.Y(n_1048)
);

NAND2xp33_ASAP7_75t_L g1049 ( 
.A(n_715),
.B(n_563),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_697),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_777),
.B(n_543),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_659),
.Y(n_1052)
);

INVxp67_ASAP7_75t_L g1053 ( 
.A(n_713),
.Y(n_1053)
);

NAND3xp33_ASAP7_75t_L g1054 ( 
.A(n_859),
.B(n_782),
.C(n_894),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_663),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_667),
.B(n_464),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_911),
.A2(n_636),
.B(n_443),
.C(n_575),
.Y(n_1057)
);

OAI22xp33_ASAP7_75t_SL g1058 ( 
.A1(n_828),
.A2(n_588),
.B1(n_594),
.B2(n_591),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_663),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_911),
.B(n_509),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_796),
.B(n_509),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_958),
.B(n_467),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_916),
.B(n_509),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_664),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_821),
.A2(n_588),
.B1(n_467),
.B2(n_634),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_676),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_916),
.B(n_467),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_664),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_918),
.B(n_527),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_918),
.B(n_527),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_919),
.B(n_547),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_919),
.B(n_547),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_665),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_801),
.B(n_900),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_900),
.B(n_443),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_796),
.B(n_443),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_903),
.B(n_514),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_903),
.B(n_514),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_676),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_905),
.B(n_514),
.Y(n_1080)
);

AO22x1_ASAP7_75t_L g1081 ( 
.A1(n_735),
.A2(n_479),
.B1(n_601),
.B2(n_594),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_665),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_901),
.B(n_568),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_825),
.A2(n_623),
.B(n_564),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_905),
.B(n_906),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_906),
.B(n_575),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_844),
.B(n_568),
.Y(n_1087)
);

INVx2_ASAP7_75t_SL g1088 ( 
.A(n_893),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_798),
.B(n_575),
.Y(n_1089)
);

BUFx8_ASAP7_75t_L g1090 ( 
.A(n_662),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_844),
.B(n_572),
.Y(n_1091)
);

AOI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_821),
.A2(n_478),
.B1(n_569),
.B2(n_572),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_923),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_798),
.B(n_562),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_699),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_847),
.A2(n_212),
.B(n_209),
.C(n_166),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_909),
.B(n_563),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_699),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_863),
.B(n_562),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_923),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_863),
.B(n_712),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_729),
.Y(n_1102)
);

INVx2_ASAP7_75t_SL g1103 ( 
.A(n_914),
.Y(n_1103)
);

INVxp67_ASAP7_75t_SL g1104 ( 
.A(n_703),
.Y(n_1104)
);

O2A1O1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_926),
.A2(n_166),
.B(n_112),
.C(n_618),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_958),
.B(n_631),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_909),
.B(n_598),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_947),
.B(n_598),
.Y(n_1108)
);

NOR3xp33_ASAP7_75t_L g1109 ( 
.A(n_810),
.B(n_134),
.C(n_126),
.Y(n_1109)
);

INVx5_ASAP7_75t_L g1110 ( 
.A(n_726),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_729),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_947),
.B(n_598),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_855),
.B(n_550),
.Y(n_1113)
);

AOI221xp5_ASAP7_75t_L g1114 ( 
.A1(n_917),
.A2(n_145),
.B1(n_201),
.B2(n_199),
.C(n_186),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_914),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_949),
.B(n_598),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_712),
.B(n_920),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_730),
.Y(n_1118)
);

OR2x2_ASAP7_75t_L g1119 ( 
.A(n_720),
.B(n_591),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_949),
.B(n_598),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_950),
.B(n_550),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_950),
.B(n_550),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_648),
.B(n_631),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_951),
.B(n_550),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_855),
.B(n_552),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_951),
.B(n_552),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_690),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_920),
.B(n_562),
.Y(n_1128)
);

OR2x6_ASAP7_75t_L g1129 ( 
.A(n_939),
.B(n_497),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_791),
.B(n_552),
.Y(n_1130)
);

INVx2_ASAP7_75t_SL g1131 ( 
.A(n_938),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_826),
.B(n_562),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_791),
.B(n_552),
.Y(n_1133)
);

NAND2x1p5_ASAP7_75t_L g1134 ( 
.A(n_923),
.B(n_623),
.Y(n_1134)
);

NOR2xp67_ASAP7_75t_L g1135 ( 
.A(n_787),
.B(n_554),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_795),
.B(n_554),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_735),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_795),
.B(n_554),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_826),
.B(n_562),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_851),
.B(n_564),
.Y(n_1140)
);

OR2x2_ASAP7_75t_L g1141 ( 
.A(n_720),
.B(n_926),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_648),
.B(n_641),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_797),
.B(n_554),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_797),
.B(n_583),
.Y(n_1144)
);

INVx1_ASAP7_75t_SL g1145 ( 
.A(n_956),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_851),
.B(n_564),
.Y(n_1146)
);

BUFx8_ASAP7_75t_L g1147 ( 
.A(n_662),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_799),
.B(n_583),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_730),
.Y(n_1149)
);

AOI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_917),
.A2(n_478),
.B1(n_569),
.B2(n_479),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_735),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_799),
.B(n_583),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_800),
.B(n_583),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_690),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_956),
.Y(n_1155)
);

NAND2xp33_ASAP7_75t_L g1156 ( 
.A(n_838),
.B(n_564),
.Y(n_1156)
);

NOR3xp33_ASAP7_75t_L g1157 ( 
.A(n_946),
.B(n_137),
.C(n_135),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_800),
.B(n_595),
.Y(n_1158)
);

AND2x4_ASAP7_75t_SL g1159 ( 
.A(n_662),
.B(n_604),
.Y(n_1159)
);

OR2x2_ASAP7_75t_L g1160 ( 
.A(n_924),
.B(n_597),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_806),
.B(n_691),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_956),
.Y(n_1162)
);

OR2x2_ASAP7_75t_L g1163 ( 
.A(n_924),
.B(n_597),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_691),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_806),
.B(n_595),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_749),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_650),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_693),
.B(n_595),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_693),
.B(n_595),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_654),
.A2(n_478),
.B1(n_569),
.B2(n_641),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_681),
.B(n_931),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_722),
.A2(n_569),
.B1(n_586),
.B2(n_564),
.Y(n_1172)
);

AND2x4_ASAP7_75t_SL g1173 ( 
.A(n_681),
.B(n_604),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_681),
.B(n_931),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_722),
.B(n_632),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_959),
.B(n_480),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_725),
.B(n_632),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_725),
.B(n_632),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_649),
.B(n_641),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_733),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_649),
.B(n_480),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_733),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_652),
.B(n_607),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_749),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_734),
.B(n_607),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_657),
.B(n_564),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_688),
.B(n_564),
.Y(n_1187)
);

INVx2_ASAP7_75t_SL g1188 ( 
.A(n_938),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_654),
.A2(n_479),
.B1(n_646),
.B2(n_147),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_652),
.B(n_614),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_692),
.B(n_586),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_801),
.B(n_614),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_953),
.Y(n_1193)
);

INVx2_ASAP7_75t_SL g1194 ( 
.A(n_953),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_960),
.Y(n_1195)
);

NAND3xp33_ASAP7_75t_L g1196 ( 
.A(n_907),
.B(n_432),
.C(n_636),
.Y(n_1196)
);

OAI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_823),
.A2(n_171),
.B1(n_169),
.B2(n_184),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_883),
.A2(n_623),
.B(n_586),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_701),
.B(n_627),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_701),
.B(n_627),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_754),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_754),
.Y(n_1202)
);

INVxp33_ASAP7_75t_SL g1203 ( 
.A(n_954),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_728),
.B(n_628),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_760),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_734),
.A2(n_645),
.B(n_630),
.C(n_646),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_728),
.B(n_628),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_781),
.B(n_635),
.Y(n_1208)
);

INVx2_ASAP7_75t_SL g1209 ( 
.A(n_908),
.Y(n_1209)
);

BUFx5_ASAP7_75t_L g1210 ( 
.A(n_726),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_959),
.B(n_450),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_692),
.B(n_586),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_936),
.A2(n_479),
.B1(n_181),
.B2(n_157),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_745),
.A2(n_586),
.B1(n_623),
.B2(n_645),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_891),
.B(n_450),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_936),
.A2(n_479),
.B1(n_147),
.B2(n_601),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_759),
.A2(n_479),
.B1(n_147),
.B2(n_601),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_760),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_SL g1219 ( 
.A(n_692),
.B(n_586),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_960),
.B(n_838),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_880),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_787),
.B(n_635),
.Y(n_1222)
);

INVxp67_ASAP7_75t_L g1223 ( 
.A(n_759),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_726),
.Y(n_1224)
);

INVx2_ASAP7_75t_SL g1225 ( 
.A(n_960),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_778),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_778),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_880),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_882),
.B(n_479),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_781),
.B(n_644),
.Y(n_1230)
);

OR2x2_ASAP7_75t_L g1231 ( 
.A(n_718),
.B(n_644),
.Y(n_1231)
);

NOR2x1p5_ASAP7_75t_L g1232 ( 
.A(n_817),
.B(n_630),
.Y(n_1232)
);

BUFx4_ASAP7_75t_L g1233 ( 
.A(n_937),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_718),
.B(n_479),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_718),
.B(n_479),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_784),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_763),
.B(n_501),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_852),
.B(n_587),
.Y(n_1238)
);

NAND2xp33_ASAP7_75t_L g1239 ( 
.A(n_882),
.B(n_586),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_763),
.B(n_501),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_852),
.B(n_587),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_746),
.B(n_531),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_954),
.B(n_531),
.Y(n_1243)
);

OR2x6_ASAP7_75t_L g1244 ( 
.A(n_939),
.B(n_587),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_881),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_852),
.B(n_872),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_738),
.A2(n_623),
.B(n_558),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_830),
.B(n_451),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_695),
.B(n_451),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_784),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_872),
.B(n_596),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_756),
.B(n_630),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_808),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_745),
.A2(n_645),
.B1(n_166),
.B2(n_172),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_804),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_808),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_811),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_789),
.B(n_596),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_756),
.B(n_630),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_818),
.B(n_596),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_877),
.A2(n_147),
.B1(n_601),
.B2(n_515),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_789),
.B(n_600),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_819),
.B(n_600),
.Y(n_1263)
);

OR2x2_ASAP7_75t_L g1264 ( 
.A(n_822),
.B(n_600),
.Y(n_1264)
);

INVx2_ASAP7_75t_SL g1265 ( 
.A(n_895),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_913),
.B(n_531),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_904),
.A2(n_857),
.B1(n_872),
.B2(n_824),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_820),
.B(n_603),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_811),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_827),
.B(n_603),
.Y(n_1270)
);

NOR2xp67_ASAP7_75t_L g1271 ( 
.A(n_881),
.B(n_624),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_813),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_884),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_726),
.Y(n_1274)
);

A2O1A1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_912),
.A2(n_545),
.B(n_528),
.C(n_551),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_892),
.B(n_531),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_892),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_822),
.A2(n_155),
.B1(n_146),
.B2(n_140),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_813),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_748),
.B(n_603),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_711),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_748),
.B(n_608),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_751),
.B(n_608),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_815),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_766),
.B(n_531),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_884),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_885),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_751),
.B(n_608),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_962),
.B(n_531),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_962),
.B(n_531),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_885),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_886),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_753),
.B(n_612),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_886),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_833),
.B(n_612),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_753),
.B(n_612),
.Y(n_1296)
);

NAND3xp33_ASAP7_75t_L g1297 ( 
.A(n_915),
.B(n_640),
.C(n_624),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_757),
.B(n_615),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_834),
.B(n_601),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_887),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_732),
.B(n_531),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_757),
.B(n_615),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_815),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_835),
.Y(n_1304)
);

AOI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_831),
.A2(n_839),
.B1(n_840),
.B2(n_832),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_761),
.B(n_615),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_835),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_961),
.B(n_616),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_846),
.Y(n_1309)
);

AND2x4_ASAP7_75t_SL g1310 ( 
.A(n_875),
.B(n_604),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_887),
.Y(n_1311)
);

INVx8_ASAP7_75t_L g1312 ( 
.A(n_726),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_888),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_846),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_761),
.B(n_616),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_SL g1316 ( 
.A(n_732),
.B(n_558),
.Y(n_1316)
);

OR2x2_ASAP7_75t_L g1317 ( 
.A(n_831),
.B(n_616),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_732),
.B(n_558),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_888),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_925),
.B(n_619),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_764),
.B(n_619),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_764),
.B(n_619),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_849),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_849),
.Y(n_1324)
);

AOI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_832),
.A2(n_177),
.B1(n_176),
.B2(n_174),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_694),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_794),
.B(n_558),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_794),
.B(n_558),
.Y(n_1328)
);

AOI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_839),
.A2(n_164),
.B1(n_129),
.B2(n_183),
.Y(n_1329)
);

AND2x4_ASAP7_75t_SL g1330 ( 
.A(n_875),
.B(n_605),
.Y(n_1330)
);

INVxp33_ASAP7_75t_L g1331 ( 
.A(n_840),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_816),
.B(n_625),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_SL g1333 ( 
.A(n_794),
.B(n_558),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_867),
.Y(n_1334)
);

O2A1O1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_656),
.A2(n_180),
.B(n_139),
.C(n_149),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_767),
.B(n_625),
.Y(n_1336)
);

NAND2xp33_ASAP7_75t_L g1337 ( 
.A(n_726),
.B(n_601),
.Y(n_1337)
);

AND2x6_ASAP7_75t_SL g1338 ( 
.A(n_927),
.B(n_135),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_816),
.B(n_625),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_L g1340 ( 
.A(n_925),
.B(n_626),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_930),
.B(n_626),
.Y(n_1341)
);

NOR2x1p5_ASAP7_75t_L g1342 ( 
.A(n_668),
.B(n_163),
.Y(n_1342)
);

NOR2xp67_ASAP7_75t_L g1343 ( 
.A(n_767),
.B(n_640),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_670),
.B(n_558),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_793),
.Y(n_1345)
);

INVxp67_ASAP7_75t_L g1346 ( 
.A(n_793),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_902),
.A2(n_567),
.B(n_558),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_930),
.B(n_626),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_SL g1349 ( 
.A(n_671),
.B(n_567),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_694),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_700),
.Y(n_1351)
);

AOI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_934),
.A2(n_601),
.B1(n_193),
.B2(n_161),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_673),
.B(n_629),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_841),
.B(n_629),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_934),
.B(n_629),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_700),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_SL g1357 ( 
.A(n_674),
.B(n_567),
.Y(n_1357)
);

NAND2xp33_ASAP7_75t_SL g1358 ( 
.A(n_677),
.B(n_633),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_678),
.B(n_633),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_682),
.B(n_633),
.Y(n_1360)
);

AND2x6_ASAP7_75t_L g1361 ( 
.A(n_940),
.B(n_941),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_704),
.Y(n_1362)
);

INVx4_ASAP7_75t_L g1363 ( 
.A(n_726),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_841),
.B(n_843),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_904),
.A2(n_601),
.B1(n_515),
.B2(n_508),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_867),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_704),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_707),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_707),
.Y(n_1369)
);

OR2x2_ASAP7_75t_SL g1370 ( 
.A(n_836),
.B(n_139),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_687),
.B(n_639),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_803),
.B(n_805),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_708),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_702),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_807),
.B(n_639),
.Y(n_1375)
);

NOR3xp33_ASAP7_75t_L g1376 ( 
.A(n_837),
.B(n_159),
.C(n_149),
.Y(n_1376)
);

NAND2x1_ASAP7_75t_L g1377 ( 
.A(n_708),
.B(n_508),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_768),
.Y(n_1378)
);

INVx2_ASAP7_75t_SL g1379 ( 
.A(n_871),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_702),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_768),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_809),
.B(n_639),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_812),
.B(n_643),
.Y(n_1383)
);

INVx2_ASAP7_75t_SL g1384 ( 
.A(n_879),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_857),
.A2(n_601),
.B1(n_522),
.B2(n_513),
.Y(n_1385)
);

INVx4_ASAP7_75t_L g1386 ( 
.A(n_702),
.Y(n_1386)
);

AOI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_935),
.A2(n_944),
.B1(n_929),
.B2(n_762),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_843),
.A2(n_172),
.B1(n_159),
.B2(n_161),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_853),
.B(n_643),
.Y(n_1389)
);

INVx8_ASAP7_75t_L g1390 ( 
.A(n_932),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_710),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_853),
.B(n_643),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_SL g1393 ( 
.A(n_935),
.B(n_842),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_865),
.B(n_513),
.Y(n_1394)
);

NOR3xp33_ASAP7_75t_L g1395 ( 
.A(n_865),
.B(n_170),
.C(n_165),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_963),
.B(n_513),
.Y(n_1396)
);

BUFx6f_ASAP7_75t_L g1397 ( 
.A(n_933),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_937),
.A2(n_571),
.B1(n_515),
.B2(n_522),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_710),
.B(n_522),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_770),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_957),
.Y(n_1401)
);

NOR3xp33_ASAP7_75t_L g1402 ( 
.A(n_714),
.B(n_165),
.C(n_170),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_829),
.A2(n_647),
.B(n_567),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1378),
.Y(n_1404)
);

INVx2_ASAP7_75t_SL g1405 ( 
.A(n_1110),
.Y(n_1405)
);

AOI21xp33_ASAP7_75t_L g1406 ( 
.A1(n_1054),
.A2(n_717),
.B(n_714),
.Y(n_1406)
);

AO22x2_ASAP7_75t_L g1407 ( 
.A1(n_987),
.A2(n_945),
.B1(n_943),
.B2(n_942),
.Y(n_1407)
);

AOI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1172),
.A2(n_747),
.B(n_719),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1221),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1214),
.A2(n_862),
.B(n_850),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1054),
.A2(n_737),
.B1(n_717),
.B2(n_719),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1214),
.A2(n_638),
.B(n_567),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1221),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1156),
.A2(n_638),
.B(n_567),
.Y(n_1414)
);

BUFx4f_ASAP7_75t_L g1415 ( 
.A(n_1361),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1363),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1239),
.A2(n_638),
.B(n_567),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_SL g1418 ( 
.A(n_998),
.B(n_845),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_SL g1419 ( 
.A(n_1213),
.B(n_1016),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1113),
.B(n_940),
.Y(n_1420)
);

AND2x6_ASAP7_75t_L g1421 ( 
.A(n_1224),
.B(n_941),
.Y(n_1421)
);

INVx11_ASAP7_75t_L g1422 ( 
.A(n_1090),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1012),
.A2(n_638),
.B(n_567),
.Y(n_1423)
);

NOR2x1_ASAP7_75t_L g1424 ( 
.A(n_982),
.B(n_736),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_965),
.A2(n_716),
.B(n_689),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_1110),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1084),
.A2(n_1198),
.B(n_1358),
.Y(n_1427)
);

AOI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_984),
.A2(n_647),
.B(n_638),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1016),
.B(n_736),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_984),
.B(n_737),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_986),
.B(n_1364),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_986),
.A2(n_647),
.B(n_638),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1364),
.B(n_739),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1297),
.A2(n_769),
.B(n_741),
.Y(n_1434)
);

BUFx4f_ASAP7_75t_L g1435 ( 
.A(n_1361),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_969),
.B(n_1123),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1125),
.B(n_942),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_991),
.B(n_943),
.Y(n_1438)
);

O2A1O1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1157),
.A2(n_739),
.B(n_743),
.C(n_740),
.Y(n_1439)
);

BUFx4f_ASAP7_75t_L g1440 ( 
.A(n_1361),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1009),
.B(n_740),
.Y(n_1441)
);

O2A1O1Ixp5_ASAP7_75t_L g1442 ( 
.A1(n_1249),
.A2(n_1308),
.B(n_1187),
.C(n_1186),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1009),
.B(n_743),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1228),
.Y(n_1444)
);

OAI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1297),
.A2(n_1196),
.B(n_970),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_967),
.B(n_744),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1337),
.A2(n_647),
.B(n_638),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1247),
.A2(n_647),
.B(n_638),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_977),
.B(n_744),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_969),
.B(n_945),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1312),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1123),
.B(n_848),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1213),
.A2(n_775),
.B1(n_770),
.B2(n_774),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1087),
.B(n_854),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1049),
.A2(n_647),
.B(n_771),
.Y(n_1455)
);

INVx2_ASAP7_75t_SL g1456 ( 
.A(n_1110),
.Y(n_1456)
);

INVx4_ASAP7_75t_L g1457 ( 
.A(n_1312),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1172),
.A2(n_647),
.B(n_771),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1010),
.B(n_772),
.Y(n_1459)
);

AOI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_997),
.A2(n_647),
.B(n_772),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1010),
.B(n_774),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1020),
.B(n_775),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1020),
.B(n_776),
.Y(n_1463)
);

OAI21xp33_ASAP7_75t_L g1464 ( 
.A1(n_1278),
.A2(n_163),
.B(n_173),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_997),
.A2(n_779),
.B(n_776),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1022),
.B(n_779),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1347),
.A2(n_783),
.B(n_780),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1022),
.B(n_780),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1378),
.Y(n_1469)
);

INVxp67_ASAP7_75t_L g1470 ( 
.A(n_1252),
.Y(n_1470)
);

INVx1_ASAP7_75t_SL g1471 ( 
.A(n_1145),
.Y(n_1471)
);

AOI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1081),
.A2(n_747),
.B(n_783),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1196),
.A2(n_1339),
.B(n_1332),
.Y(n_1473)
);

BUFx8_ASAP7_75t_L g1474 ( 
.A(n_971),
.Y(n_1474)
);

OAI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_994),
.A2(n_786),
.B(n_785),
.Y(n_1475)
);

AOI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1121),
.A2(n_786),
.B(n_785),
.Y(n_1476)
);

A2O1A1Ixp33_ASAP7_75t_L g1477 ( 
.A1(n_1018),
.A2(n_928),
.B(n_856),
.C(n_878),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_981),
.B(n_858),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1121),
.A2(n_1124),
.B(n_1122),
.Y(n_1479)
);

AOI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1122),
.A2(n_551),
.B(n_545),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1378),
.Y(n_1481)
);

INVx4_ASAP7_75t_L g1482 ( 
.A(n_1312),
.Y(n_1482)
);

OR2x6_ASAP7_75t_L g1483 ( 
.A(n_1312),
.B(n_860),
.Y(n_1483)
);

AOI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1124),
.A2(n_551),
.B(n_545),
.Y(n_1484)
);

O2A1O1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_1096),
.A2(n_861),
.B(n_876),
.C(n_870),
.Y(n_1485)
);

O2A1O1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_987),
.A2(n_1035),
.B(n_1053),
.C(n_1160),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_981),
.B(n_868),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1228),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1142),
.B(n_869),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1000),
.B(n_528),
.Y(n_1490)
);

AOI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1126),
.A2(n_528),
.B(n_559),
.Y(n_1491)
);

AOI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1126),
.A2(n_560),
.B(n_559),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1091),
.B(n_131),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1185),
.A2(n_560),
.B(n_559),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1142),
.B(n_267),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1275),
.A2(n_529),
.B(n_571),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1179),
.B(n_267),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1000),
.B(n_529),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_L g1499 ( 
.A(n_1312),
.Y(n_1499)
);

AOI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1185),
.A2(n_571),
.B(n_560),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1245),
.Y(n_1501)
);

OAI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1206),
.A2(n_529),
.B(n_582),
.Y(n_1502)
);

AOI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1222),
.A2(n_576),
.B(n_577),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1222),
.A2(n_576),
.B(n_577),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1381),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1097),
.A2(n_1108),
.B(n_1107),
.Y(n_1506)
);

AOI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1097),
.A2(n_576),
.B(n_577),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1183),
.B(n_579),
.Y(n_1508)
);

AOI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1107),
.A2(n_579),
.B(n_582),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1183),
.B(n_579),
.Y(n_1510)
);

A2O1A1Ixp33_ASAP7_75t_L g1511 ( 
.A1(n_1176),
.A2(n_582),
.B(n_191),
.C(n_173),
.Y(n_1511)
);

AOI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1108),
.A2(n_1116),
.B(n_1112),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1141),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1042),
.A2(n_178),
.B1(n_180),
.B2(n_187),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1237),
.B(n_117),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1190),
.B(n_933),
.Y(n_1516)
);

AO21x1_ASAP7_75t_L g1517 ( 
.A1(n_1058),
.A2(n_933),
.B(n_642),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1179),
.B(n_267),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_1167),
.Y(n_1519)
);

BUFx6f_ASAP7_75t_L g1520 ( 
.A(n_1110),
.Y(n_1520)
);

NAND2x1p5_ASAP7_75t_L g1521 ( 
.A(n_1110),
.B(n_267),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1141),
.Y(n_1522)
);

OAI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_989),
.A2(n_381),
.B(n_393),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_964),
.B(n_267),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1019),
.A2(n_1044),
.B1(n_980),
.B2(n_1267),
.Y(n_1525)
);

AOI21xp33_ASAP7_75t_L g1526 ( 
.A1(n_1058),
.A2(n_189),
.B(n_191),
.Y(n_1526)
);

AOI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1033),
.A2(n_193),
.B1(n_208),
.B2(n_202),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_SL g1528 ( 
.A(n_1021),
.B(n_605),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1190),
.B(n_605),
.Y(n_1529)
);

AOI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1112),
.A2(n_369),
.B(n_322),
.Y(n_1530)
);

OAI21x1_ASAP7_75t_L g1531 ( 
.A1(n_989),
.A2(n_381),
.B(n_393),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1245),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1085),
.B(n_605),
.Y(n_1533)
);

OAI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_992),
.A2(n_389),
.B(n_379),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1273),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1116),
.A2(n_314),
.B(n_322),
.Y(n_1536)
);

AOI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1120),
.A2(n_314),
.B(n_322),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1381),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_L g1539 ( 
.A(n_1240),
.B(n_120),
.Y(n_1539)
);

OAI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_992),
.A2(n_368),
.B(n_389),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1273),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1085),
.B(n_605),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1354),
.B(n_267),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1120),
.A2(n_385),
.B(n_309),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_964),
.B(n_267),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1354),
.B(n_267),
.Y(n_1546)
);

OAI321xp33_ASAP7_75t_L g1547 ( 
.A1(n_1217),
.A2(n_196),
.A3(n_194),
.B1(n_190),
.B2(n_189),
.C(n_187),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1161),
.B(n_267),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1338),
.B(n_122),
.Y(n_1549)
);

OAI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1005),
.A2(n_1057),
.B(n_1181),
.Y(n_1550)
);

BUFx6f_ASAP7_75t_L g1551 ( 
.A(n_1110),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1361),
.Y(n_1552)
);

INVxp67_ASAP7_75t_L g1553 ( 
.A(n_1259),
.Y(n_1553)
);

O2A1O1Ixp33_ASAP7_75t_SL g1554 ( 
.A1(n_978),
.A2(n_379),
.B(n_376),
.C(n_368),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1381),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1161),
.B(n_267),
.Y(n_1556)
);

NAND2x1p5_ASAP7_75t_L g1557 ( 
.A(n_1363),
.B(n_267),
.Y(n_1557)
);

O2A1O1Ixp33_ASAP7_75t_L g1558 ( 
.A1(n_1160),
.A2(n_210),
.B(n_208),
.C(n_202),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1286),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1211),
.B(n_267),
.Y(n_1560)
);

BUFx12f_ASAP7_75t_L g1561 ( 
.A(n_1370),
.Y(n_1561)
);

AOI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1258),
.A2(n_385),
.B(n_314),
.Y(n_1562)
);

OAI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1005),
.A2(n_1181),
.B(n_1042),
.Y(n_1563)
);

A2O1A1Ixp33_ASAP7_75t_L g1564 ( 
.A1(n_1215),
.A2(n_190),
.B(n_200),
.C(n_197),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1199),
.B(n_267),
.Y(n_1565)
);

O2A1O1Ixp33_ASAP7_75t_L g1566 ( 
.A1(n_1163),
.A2(n_200),
.B(n_197),
.C(n_196),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_SL g1567 ( 
.A(n_1163),
.B(n_975),
.Y(n_1567)
);

BUFx24_ASAP7_75t_L g1568 ( 
.A(n_1370),
.Y(n_1568)
);

AOI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1081),
.A2(n_376),
.B(n_254),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1286),
.Y(n_1570)
);

AOI21xp5_ASAP7_75t_L g1571 ( 
.A1(n_1258),
.A2(n_385),
.B(n_369),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1106),
.B(n_266),
.Y(n_1572)
);

A2O1A1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1335),
.A2(n_1352),
.B(n_1387),
.C(n_1083),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1287),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_SL g1575 ( 
.A(n_1387),
.B(n_309),
.Y(n_1575)
);

BUFx3_ASAP7_75t_L g1576 ( 
.A(n_1090),
.Y(n_1576)
);

BUFx3_ASAP7_75t_L g1577 ( 
.A(n_1090),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_SL g1578 ( 
.A(n_1074),
.B(n_1220),
.Y(n_1578)
);

NAND2xp33_ASAP7_75t_L g1579 ( 
.A(n_1361),
.B(n_309),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1200),
.B(n_275),
.Y(n_1580)
);

OAI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1014),
.A2(n_257),
.B(n_254),
.Y(n_1581)
);

AOI21x1_ASAP7_75t_L g1582 ( 
.A1(n_1377),
.A2(n_254),
.B(n_257),
.Y(n_1582)
);

AOI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1262),
.A2(n_385),
.B(n_369),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1287),
.Y(n_1584)
);

AOI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_980),
.A2(n_210),
.B1(n_194),
.B2(n_178),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_1220),
.B(n_309),
.Y(n_1586)
);

OAI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1014),
.A2(n_257),
.B(n_254),
.Y(n_1587)
);

AOI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1262),
.A2(n_385),
.B(n_369),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1204),
.B(n_275),
.Y(n_1589)
);

NOR2xp67_ASAP7_75t_L g1590 ( 
.A(n_1400),
.B(n_254),
.Y(n_1590)
);

OAI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1027),
.A2(n_1343),
.B(n_982),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1207),
.B(n_275),
.Y(n_1592)
);

INVxp67_ASAP7_75t_L g1593 ( 
.A(n_1255),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1280),
.A2(n_385),
.B(n_369),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_1203),
.Y(n_1595)
);

NOR2x2_ASAP7_75t_L g1596 ( 
.A(n_1390),
.B(n_257),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1013),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1280),
.A2(n_385),
.B(n_369),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1338),
.B(n_1043),
.Y(n_1599)
);

AOI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1282),
.A2(n_1288),
.B(n_1283),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1331),
.B(n_127),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1363),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1208),
.B(n_1230),
.Y(n_1603)
);

AOI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1282),
.A2(n_385),
.B(n_369),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1093),
.B(n_275),
.Y(n_1605)
);

A2O1A1Ixp33_ASAP7_75t_L g1606 ( 
.A1(n_1352),
.A2(n_130),
.B(n_154),
.C(n_182),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1305),
.A2(n_275),
.B1(n_257),
.B2(n_266),
.Y(n_1607)
);

AOI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1283),
.A2(n_369),
.B(n_309),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1093),
.B(n_1162),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1291),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1093),
.B(n_257),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1093),
.B(n_266),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1162),
.B(n_266),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1162),
.B(n_266),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1223),
.B(n_198),
.Y(n_1615)
);

AOI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1288),
.A2(n_335),
.B(n_331),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1400),
.Y(n_1617)
);

BUFx4f_ASAP7_75t_L g1618 ( 
.A(n_1361),
.Y(n_1618)
);

AOI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1293),
.A2(n_335),
.B(n_331),
.Y(n_1619)
);

BUFx3_ASAP7_75t_L g1620 ( 
.A(n_1090),
.Y(n_1620)
);

AOI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1293),
.A2(n_335),
.B(n_331),
.Y(n_1621)
);

OAI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1027),
.A2(n_362),
.B(n_266),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1220),
.B(n_309),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1291),
.Y(n_1624)
);

BUFx6f_ASAP7_75t_L g1625 ( 
.A(n_1224),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1045),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_SL g1627 ( 
.A1(n_1233),
.A2(n_266),
.B1(n_2),
.B2(n_5),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_1255),
.B(n_0),
.Y(n_1628)
);

AOI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_971),
.A2(n_266),
.B1(n_335),
.B2(n_331),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1162),
.B(n_266),
.Y(n_1630)
);

AO21x1_ASAP7_75t_L g1631 ( 
.A1(n_1320),
.A2(n_1341),
.B(n_1340),
.Y(n_1631)
);

AOI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1296),
.A2(n_335),
.B(n_331),
.Y(n_1632)
);

AOI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1296),
.A2(n_335),
.B(n_331),
.Y(n_1633)
);

OAI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1343),
.A2(n_362),
.B(n_312),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_976),
.B(n_362),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1192),
.B(n_362),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_979),
.B(n_335),
.Y(n_1637)
);

AOI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1377),
.A2(n_335),
.B(n_331),
.Y(n_1638)
);

AOI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1298),
.A2(n_331),
.B(n_322),
.Y(n_1639)
);

AOI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1298),
.A2(n_322),
.B(n_314),
.Y(n_1640)
);

OAI321xp33_ASAP7_75t_L g1641 ( 
.A1(n_1261),
.A2(n_0),
.A3(n_7),
.B1(n_9),
.B2(n_10),
.C(n_12),
.Y(n_1641)
);

INVx11_ASAP7_75t_L g1642 ( 
.A(n_1147),
.Y(n_1642)
);

AOI21x1_ASAP7_75t_L g1643 ( 
.A1(n_1244),
.A2(n_322),
.B(n_314),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1056),
.Y(n_1644)
);

AOI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1395),
.A2(n_322),
.B1(n_314),
.B2(n_244),
.Y(n_1645)
);

AOI21xp33_ASAP7_75t_L g1646 ( 
.A1(n_1105),
.A2(n_1119),
.B(n_1398),
.Y(n_1646)
);

BUFx2_ASAP7_75t_L g1647 ( 
.A(n_1361),
.Y(n_1647)
);

AOI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1302),
.A2(n_322),
.B(n_314),
.Y(n_1648)
);

CKINVDCx8_ASAP7_75t_R g1649 ( 
.A(n_1390),
.Y(n_1649)
);

AOI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1302),
.A2(n_314),
.B(n_244),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1265),
.B(n_9),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1305),
.A2(n_264),
.B1(n_251),
.B2(n_246),
.Y(n_1652)
);

AOI21x1_ASAP7_75t_L g1653 ( 
.A1(n_1244),
.A2(n_312),
.B(n_264),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1265),
.B(n_1007),
.Y(n_1654)
);

INVx4_ASAP7_75t_L g1655 ( 
.A(n_1361),
.Y(n_1655)
);

O2A1O1Ixp33_ASAP7_75t_L g1656 ( 
.A1(n_1388),
.A2(n_12),
.B(n_14),
.C(n_16),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1400),
.Y(n_1657)
);

AOI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1306),
.A2(n_251),
.B(n_264),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1306),
.A2(n_251),
.B(n_264),
.Y(n_1659)
);

AND2x6_ASAP7_75t_L g1660 ( 
.A(n_1224),
.B(n_264),
.Y(n_1660)
);

BUFx3_ASAP7_75t_L g1661 ( 
.A(n_1147),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_979),
.B(n_264),
.Y(n_1662)
);

AND2x4_ASAP7_75t_L g1663 ( 
.A(n_1220),
.B(n_88),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_988),
.Y(n_1664)
);

BUFx4f_ASAP7_75t_L g1665 ( 
.A(n_990),
.Y(n_1665)
);

OAI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1271),
.A2(n_312),
.B(n_250),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_SL g1667 ( 
.A(n_1065),
.B(n_251),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1315),
.A2(n_251),
.B(n_264),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_983),
.B(n_264),
.Y(n_1669)
);

OAI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1271),
.A2(n_312),
.B(n_250),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_983),
.B(n_264),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_996),
.B(n_264),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1315),
.A2(n_251),
.B(n_264),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1345),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1321),
.A2(n_251),
.B(n_264),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1321),
.A2(n_1336),
.B(n_1322),
.Y(n_1676)
);

AOI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1322),
.A2(n_251),
.B(n_264),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1292),
.Y(n_1678)
);

NOR2xp33_ASAP7_75t_L g1679 ( 
.A(n_1007),
.B(n_1117),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_996),
.B(n_264),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_SL g1681 ( 
.A(n_1363),
.B(n_312),
.Y(n_1681)
);

AOI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1336),
.A2(n_1133),
.B(n_1130),
.Y(n_1682)
);

AOI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1130),
.A2(n_251),
.B(n_264),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1015),
.B(n_251),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_SL g1685 ( 
.A(n_1274),
.B(n_312),
.Y(n_1685)
);

BUFx2_ASAP7_75t_L g1686 ( 
.A(n_1244),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1133),
.A2(n_251),
.B(n_246),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1015),
.B(n_1017),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1209),
.Y(n_1689)
);

AOI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1136),
.A2(n_251),
.B(n_246),
.Y(n_1690)
);

BUFx3_ASAP7_75t_L g1691 ( 
.A(n_1147),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1106),
.B(n_16),
.Y(n_1692)
);

AOI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1136),
.A2(n_251),
.B(n_246),
.Y(n_1693)
);

AOI21x1_ASAP7_75t_L g1694 ( 
.A1(n_1244),
.A2(n_312),
.B(n_251),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_988),
.Y(n_1695)
);

AOI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1138),
.A2(n_251),
.B(n_246),
.Y(n_1696)
);

AOI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1138),
.A2(n_246),
.B(n_244),
.Y(n_1697)
);

OAI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1389),
.A2(n_312),
.B(n_262),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1017),
.B(n_246),
.Y(n_1699)
);

INVxp67_ASAP7_75t_L g1700 ( 
.A(n_1401),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1023),
.B(n_1039),
.Y(n_1701)
);

O2A1O1Ixp33_ASAP7_75t_SL g1702 ( 
.A1(n_985),
.A2(n_17),
.B(n_21),
.C(n_25),
.Y(n_1702)
);

AOI21x1_ASAP7_75t_L g1703 ( 
.A1(n_1244),
.A2(n_246),
.B(n_244),
.Y(n_1703)
);

INVx11_ASAP7_75t_L g1704 ( 
.A(n_1147),
.Y(n_1704)
);

O2A1O1Ixp33_ASAP7_75t_L g1705 ( 
.A1(n_1388),
.A2(n_17),
.B(n_21),
.C(n_25),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1401),
.B(n_26),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1143),
.A2(n_246),
.B(n_259),
.Y(n_1707)
);

OR2x6_ASAP7_75t_L g1708 ( 
.A(n_1274),
.B(n_246),
.Y(n_1708)
);

BUFx6f_ASAP7_75t_L g1709 ( 
.A(n_1274),
.Y(n_1709)
);

AOI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1143),
.A2(n_246),
.B(n_259),
.Y(n_1710)
);

AOI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1144),
.A2(n_246),
.B(n_259),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1195),
.B(n_26),
.Y(n_1712)
);

NOR3xp33_ASAP7_75t_L g1713 ( 
.A(n_1114),
.B(n_28),
.C(n_31),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1023),
.B(n_246),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1195),
.B(n_28),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1039),
.B(n_1041),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_SL g1717 ( 
.A(n_1065),
.B(n_246),
.Y(n_1717)
);

AOI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1144),
.A2(n_246),
.B(n_259),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1041),
.B(n_1055),
.Y(n_1719)
);

AOI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1148),
.A2(n_262),
.B(n_259),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1292),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1055),
.B(n_31),
.Y(n_1722)
);

AOI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1031),
.A2(n_262),
.B1(n_259),
.B2(n_250),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1059),
.B(n_32),
.Y(n_1724)
);

BUFx12f_ASAP7_75t_L g1725 ( 
.A(n_1032),
.Y(n_1725)
);

INVx3_ASAP7_75t_L g1726 ( 
.A(n_1229),
.Y(n_1726)
);

OAI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1392),
.A2(n_262),
.B(n_259),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_988),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1401),
.B(n_35),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1059),
.B(n_38),
.Y(n_1730)
);

AOI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1148),
.A2(n_262),
.B(n_259),
.Y(n_1731)
);

INVx3_ASAP7_75t_L g1732 ( 
.A(n_1229),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_SL g1733 ( 
.A(n_966),
.B(n_262),
.Y(n_1733)
);

O2A1O1Ixp5_ASAP7_75t_L g1734 ( 
.A1(n_1344),
.A2(n_38),
.B(n_39),
.C(n_40),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1195),
.B(n_44),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1064),
.B(n_44),
.Y(n_1736)
);

AOI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1152),
.A2(n_262),
.B(n_259),
.Y(n_1737)
);

AOI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1152),
.A2(n_262),
.B(n_259),
.Y(n_1738)
);

INVx3_ASAP7_75t_L g1739 ( 
.A(n_1229),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_SL g1740 ( 
.A(n_966),
.B(n_262),
.Y(n_1740)
);

AOI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1153),
.A2(n_262),
.B(n_259),
.Y(n_1741)
);

AOI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1153),
.A2(n_262),
.B(n_259),
.Y(n_1742)
);

AOI21xp5_ASAP7_75t_L g1743 ( 
.A1(n_1158),
.A2(n_262),
.B(n_259),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1294),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_999),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_SL g1746 ( 
.A(n_1137),
.B(n_1151),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_1209),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_999),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1100),
.B(n_105),
.Y(n_1749)
);

CKINVDCx10_ASAP7_75t_R g1750 ( 
.A(n_1129),
.Y(n_1750)
);

AOI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1158),
.A2(n_262),
.B(n_259),
.Y(n_1751)
);

NOR3xp33_ASAP7_75t_L g1752 ( 
.A(n_1197),
.B(n_45),
.C(n_46),
.Y(n_1752)
);

AOI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1165),
.A2(n_262),
.B(n_259),
.Y(n_1753)
);

AOI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1038),
.A2(n_262),
.B1(n_259),
.B2(n_250),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1294),
.Y(n_1755)
);

CKINVDCx8_ASAP7_75t_R g1756 ( 
.A(n_1390),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1064),
.B(n_45),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1300),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1300),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_SL g1760 ( 
.A(n_974),
.B(n_262),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1068),
.B(n_48),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1068),
.B(n_48),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1073),
.B(n_49),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1073),
.B(n_49),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_999),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1231),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1189),
.A2(n_250),
.B1(n_53),
.B2(n_54),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1008),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_SL g1769 ( 
.A(n_1137),
.B(n_250),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1311),
.Y(n_1770)
);

BUFx2_ASAP7_75t_L g1771 ( 
.A(n_1281),
.Y(n_1771)
);

BUFx4f_ASAP7_75t_L g1772 ( 
.A(n_990),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1082),
.B(n_1127),
.Y(n_1773)
);

INVx4_ASAP7_75t_L g1774 ( 
.A(n_1100),
.Y(n_1774)
);

BUFx2_ASAP7_75t_L g1775 ( 
.A(n_1281),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1008),
.Y(n_1776)
);

BUFx12f_ASAP7_75t_L g1777 ( 
.A(n_1032),
.Y(n_1777)
);

BUFx3_ASAP7_75t_L g1778 ( 
.A(n_1100),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1082),
.B(n_50),
.Y(n_1779)
);

OAI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1394),
.A2(n_250),
.B(n_54),
.Y(n_1780)
);

O2A1O1Ixp5_ASAP7_75t_L g1781 ( 
.A1(n_1349),
.A2(n_50),
.B(n_55),
.C(n_56),
.Y(n_1781)
);

AOI21xp5_ASAP7_75t_L g1782 ( 
.A1(n_1165),
.A2(n_250),
.B(n_56),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1003),
.B(n_1119),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1008),
.Y(n_1784)
);

BUFx6f_ASAP7_75t_L g1785 ( 
.A(n_1397),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1127),
.B(n_55),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1311),
.Y(n_1787)
);

OAI21xp33_ASAP7_75t_L g1788 ( 
.A1(n_1278),
.A2(n_1329),
.B(n_1325),
.Y(n_1788)
);

AOI33xp33_ASAP7_75t_L g1789 ( 
.A1(n_1325),
.A2(n_57),
.A3(n_58),
.B1(n_59),
.B2(n_63),
.B3(n_64),
.Y(n_1789)
);

NOR3xp33_ASAP7_75t_L g1790 ( 
.A(n_1109),
.B(n_58),
.C(n_63),
.Y(n_1790)
);

BUFx3_ASAP7_75t_L g1791 ( 
.A(n_1100),
.Y(n_1791)
);

AOI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1168),
.A2(n_250),
.B(n_66),
.Y(n_1792)
);

AOI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1346),
.A2(n_250),
.B1(n_67),
.B2(n_68),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1154),
.B(n_65),
.Y(n_1794)
);

NOR3xp33_ASAP7_75t_L g1795 ( 
.A(n_1101),
.B(n_67),
.C(n_69),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1313),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_SL g1797 ( 
.A(n_974),
.B(n_1100),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1154),
.B(n_1164),
.Y(n_1798)
);

AND2x4_ASAP7_75t_L g1799 ( 
.A(n_1100),
.B(n_87),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1164),
.B(n_72),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1003),
.B(n_74),
.Y(n_1801)
);

CKINVDCx16_ASAP7_75t_R g1802 ( 
.A(n_1137),
.Y(n_1802)
);

OAI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1372),
.A2(n_74),
.B1(n_250),
.B2(n_76),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1180),
.B(n_250),
.Y(n_1804)
);

NAND2x1p5_ASAP7_75t_L g1805 ( 
.A(n_1386),
.B(n_250),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1168),
.A2(n_250),
.B(n_77),
.Y(n_1806)
);

HB1xp67_ASAP7_75t_L g1807 ( 
.A(n_1231),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1169),
.A2(n_250),
.B(n_85),
.Y(n_1808)
);

AOI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1246),
.A2(n_250),
.B1(n_89),
.B2(n_90),
.Y(n_1809)
);

A2O1A1Ixp33_ASAP7_75t_L g1810 ( 
.A1(n_1248),
.A2(n_75),
.B(n_97),
.C(n_102),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1180),
.B(n_1182),
.Y(n_1811)
);

O2A1O1Ixp5_ASAP7_75t_L g1812 ( 
.A1(n_1357),
.A2(n_1242),
.B(n_972),
.C(n_973),
.Y(n_1812)
);

AOI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1169),
.A2(n_1177),
.B(n_1175),
.Y(n_1813)
);

AOI21xp5_ASAP7_75t_L g1814 ( 
.A1(n_1175),
.A2(n_1178),
.B(n_1177),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_SL g1815 ( 
.A(n_1155),
.B(n_1135),
.Y(n_1815)
);

AOI21x1_ASAP7_75t_L g1816 ( 
.A1(n_1094),
.A2(n_1393),
.B(n_1099),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_SL g1817 ( 
.A(n_1155),
.B(n_1135),
.Y(n_1817)
);

BUFx8_ASAP7_75t_L g1818 ( 
.A(n_1195),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1036),
.Y(n_1819)
);

AOI21xp5_ASAP7_75t_L g1820 ( 
.A1(n_1178),
.A2(n_1077),
.B(n_1075),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1036),
.Y(n_1821)
);

INVx4_ASAP7_75t_L g1822 ( 
.A(n_1155),
.Y(n_1822)
);

AND2x6_ASAP7_75t_SL g1823 ( 
.A(n_1129),
.B(n_1234),
.Y(n_1823)
);

BUFx2_ASAP7_75t_L g1824 ( 
.A(n_1129),
.Y(n_1824)
);

AOI21xp33_ASAP7_75t_L g1825 ( 
.A1(n_1216),
.A2(n_1365),
.B(n_1254),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1182),
.B(n_1264),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1372),
.A2(n_1072),
.B1(n_1071),
.B2(n_1070),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_SL g1828 ( 
.A(n_1155),
.B(n_1088),
.Y(n_1828)
);

HB1xp67_ASAP7_75t_L g1829 ( 
.A(n_1264),
.Y(n_1829)
);

AOI22xp33_ASAP7_75t_L g1830 ( 
.A1(n_1170),
.A2(n_1171),
.B1(n_1174),
.B2(n_1146),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1317),
.B(n_1145),
.Y(n_1831)
);

BUFx6f_ASAP7_75t_L g1832 ( 
.A(n_1397),
.Y(n_1832)
);

AOI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1075),
.A2(n_1078),
.B(n_1077),
.Y(n_1833)
);

BUFx4f_ASAP7_75t_L g1834 ( 
.A(n_990),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1036),
.Y(n_1835)
);

AOI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1078),
.A2(n_1086),
.B(n_1080),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1313),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1047),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_L g1839 ( 
.A(n_1088),
.B(n_1103),
.Y(n_1839)
);

OAI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1069),
.A2(n_1329),
.B1(n_1150),
.B2(n_1317),
.Y(n_1840)
);

AOI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1080),
.A2(n_1086),
.B(n_1353),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1047),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1319),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1047),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1067),
.B(n_1026),
.Y(n_1845)
);

AO21x1_ASAP7_75t_L g1846 ( 
.A1(n_1348),
.A2(n_1355),
.B(n_1048),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1155),
.B(n_1103),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1011),
.B(n_1029),
.Y(n_1848)
);

OAI21xp5_ASAP7_75t_L g1849 ( 
.A1(n_1051),
.A2(n_1396),
.B(n_1263),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1319),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1026),
.B(n_1034),
.Y(n_1851)
);

AOI21xp5_ASAP7_75t_L g1852 ( 
.A1(n_1353),
.A2(n_1360),
.B(n_1359),
.Y(n_1852)
);

AO21x1_ASAP7_75t_L g1853 ( 
.A1(n_1260),
.A2(n_1270),
.B(n_1268),
.Y(n_1853)
);

AOI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1359),
.A2(n_1371),
.B(n_1360),
.Y(n_1854)
);

AOI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1046),
.A2(n_1402),
.B1(n_968),
.B2(n_1129),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1052),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1034),
.B(n_1326),
.Y(n_1857)
);

AOI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1371),
.A2(n_1382),
.B(n_1375),
.Y(n_1858)
);

AOI21xp5_ASAP7_75t_L g1859 ( 
.A1(n_1375),
.A2(n_1383),
.B(n_1382),
.Y(n_1859)
);

AOI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1383),
.A2(n_1403),
.B(n_1295),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1326),
.Y(n_1861)
);

BUFx4f_ASAP7_75t_L g1862 ( 
.A(n_1134),
.Y(n_1862)
);

AOI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1060),
.A2(n_1063),
.B(n_1399),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1350),
.Y(n_1864)
);

NOR2xp67_ASAP7_75t_L g1865 ( 
.A(n_1150),
.B(n_1350),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1052),
.Y(n_1866)
);

INVx3_ASAP7_75t_L g1867 ( 
.A(n_1229),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1351),
.B(n_1356),
.Y(n_1868)
);

BUFx12f_ASAP7_75t_L g1869 ( 
.A(n_1115),
.Y(n_1869)
);

BUFx6f_ASAP7_75t_L g1870 ( 
.A(n_1397),
.Y(n_1870)
);

AOI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1330),
.A2(n_1104),
.B(n_1285),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1351),
.B(n_1356),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1362),
.B(n_1367),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_SL g1874 ( 
.A(n_1155),
.B(n_1115),
.Y(n_1874)
);

INVx11_ASAP7_75t_L g1875 ( 
.A(n_1004),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1362),
.B(n_1367),
.Y(n_1876)
);

AND2x4_ASAP7_75t_L g1877 ( 
.A(n_1159),
.B(n_1173),
.Y(n_1877)
);

AOI21xp5_ASAP7_75t_L g1878 ( 
.A1(n_1330),
.A2(n_1050),
.B(n_1030),
.Y(n_1878)
);

NOR2x1_ASAP7_75t_L g1879 ( 
.A(n_1151),
.B(n_1232),
.Y(n_1879)
);

INVx3_ASAP7_75t_L g1880 ( 
.A(n_1299),
.Y(n_1880)
);

AOI21xp5_ASAP7_75t_L g1881 ( 
.A1(n_1330),
.A2(n_1050),
.B(n_1030),
.Y(n_1881)
);

INVx3_ASAP7_75t_L g1882 ( 
.A(n_1299),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_SL g1883 ( 
.A(n_1131),
.B(n_1188),
.Y(n_1883)
);

O2A1O1Ixp33_ASAP7_75t_L g1884 ( 
.A1(n_1254),
.A2(n_1037),
.B(n_1219),
.C(n_1212),
.Y(n_1884)
);

AOI21xp5_ASAP7_75t_L g1885 ( 
.A1(n_1024),
.A2(n_1050),
.B(n_1030),
.Y(n_1885)
);

INVx3_ASAP7_75t_L g1886 ( 
.A(n_1299),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1368),
.B(n_1369),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_SL g1888 ( 
.A(n_1131),
.B(n_1188),
.Y(n_1888)
);

INVx4_ASAP7_75t_L g1889 ( 
.A(n_1134),
.Y(n_1889)
);

HB1xp67_ASAP7_75t_L g1890 ( 
.A(n_1195),
.Y(n_1890)
);

BUFx2_ASAP7_75t_L g1891 ( 
.A(n_1129),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1368),
.B(n_1369),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1024),
.A2(n_1050),
.B(n_1030),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1373),
.Y(n_1894)
);

OAI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1238),
.A2(n_1241),
.B(n_1251),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1373),
.B(n_1391),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1391),
.Y(n_1897)
);

O2A1O1Ixp33_ASAP7_75t_L g1898 ( 
.A1(n_1191),
.A2(n_1376),
.B(n_1301),
.C(n_1327),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1193),
.B(n_1194),
.Y(n_1899)
);

NAND2x1p5_ASAP7_75t_L g1900 ( 
.A(n_1386),
.B(n_1397),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1195),
.B(n_1040),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1011),
.B(n_1029),
.Y(n_1902)
);

OAI21xp5_ASAP7_75t_L g1903 ( 
.A1(n_1385),
.A2(n_1128),
.B(n_1299),
.Y(n_1903)
);

AOI21xp5_ASAP7_75t_L g1904 ( 
.A1(n_1024),
.A2(n_1276),
.B(n_1290),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1225),
.B(n_1040),
.Y(n_1905)
);

AOI21xp5_ASAP7_75t_L g1906 ( 
.A1(n_1024),
.A2(n_1289),
.B(n_1333),
.Y(n_1906)
);

AOI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1316),
.A2(n_1318),
.B(n_1328),
.Y(n_1907)
);

NOR2xp33_ASAP7_75t_L g1908 ( 
.A(n_1193),
.B(n_1194),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1225),
.B(n_1040),
.Y(n_1909)
);

AOI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1002),
.A2(n_1006),
.B(n_1134),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1040),
.B(n_1062),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1052),
.Y(n_1912)
);

AOI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1025),
.A2(n_1028),
.B(n_1061),
.Y(n_1913)
);

OAI21xp5_ASAP7_75t_L g1914 ( 
.A1(n_1092),
.A2(n_1089),
.B(n_1076),
.Y(n_1914)
);

INVx3_ASAP7_75t_L g1915 ( 
.A(n_1210),
.Y(n_1915)
);

INVx3_ASAP7_75t_L g1916 ( 
.A(n_1210),
.Y(n_1916)
);

AOI21xp5_ASAP7_75t_L g1917 ( 
.A1(n_1310),
.A2(n_1266),
.B(n_1092),
.Y(n_1917)
);

INVx4_ASAP7_75t_L g1918 ( 
.A(n_1210),
.Y(n_1918)
);

OAI21xp5_ASAP7_75t_L g1919 ( 
.A1(n_1235),
.A2(n_1001),
.B(n_1366),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1062),
.B(n_1232),
.Y(n_1920)
);

AOI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1310),
.A2(n_993),
.B(n_995),
.Y(n_1921)
);

INVx1_ASAP7_75t_SL g1922 ( 
.A(n_1062),
.Y(n_1922)
);

AOI21xp5_ASAP7_75t_L g1923 ( 
.A1(n_1310),
.A2(n_1277),
.B(n_1314),
.Y(n_1923)
);

OAI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1066),
.A2(n_1227),
.B(n_1279),
.Y(n_1924)
);

OAI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1066),
.A2(n_1227),
.B(n_1279),
.Y(n_1925)
);

OAI21xp5_ASAP7_75t_L g1926 ( 
.A1(n_1066),
.A2(n_1227),
.B(n_1279),
.Y(n_1926)
);

AOI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1277),
.A2(n_1205),
.B(n_1314),
.Y(n_1927)
);

AOI21xp5_ASAP7_75t_L g1928 ( 
.A1(n_1277),
.A2(n_1205),
.B(n_1314),
.Y(n_1928)
);

AOI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1277),
.A2(n_1236),
.B(n_1323),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_SL g1930 ( 
.A(n_1277),
.B(n_1397),
.Y(n_1930)
);

OAI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1079),
.A2(n_1226),
.B(n_1269),
.Y(n_1931)
);

AOI21xp5_ASAP7_75t_L g1932 ( 
.A1(n_1277),
.A2(n_1236),
.B(n_1323),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1159),
.B(n_1173),
.Y(n_1933)
);

INVx5_ASAP7_75t_L g1934 ( 
.A(n_1397),
.Y(n_1934)
);

AND2x2_ASAP7_75t_SL g1935 ( 
.A(n_1233),
.B(n_1159),
.Y(n_1935)
);

AOI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1079),
.A2(n_1218),
.B(n_1334),
.Y(n_1936)
);

AOI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1079),
.A2(n_1218),
.B(n_1334),
.Y(n_1937)
);

AOI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1095),
.A2(n_1250),
.B(n_1366),
.Y(n_1938)
);

NOR3xp33_ASAP7_75t_L g1939 ( 
.A(n_1243),
.B(n_1140),
.C(n_1139),
.Y(n_1939)
);

AOI33xp33_ASAP7_75t_L g1940 ( 
.A1(n_1379),
.A2(n_1384),
.A3(n_1062),
.B1(n_1342),
.B2(n_1098),
.B3(n_1102),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1095),
.B(n_1256),
.Y(n_1941)
);

AOI21xp5_ASAP7_75t_L g1942 ( 
.A1(n_1095),
.A2(n_1256),
.B(n_1098),
.Y(n_1942)
);

A2O1A1Ixp33_ASAP7_75t_L g1943 ( 
.A1(n_1342),
.A2(n_1374),
.B(n_1380),
.C(n_1132),
.Y(n_1943)
);

A2O1A1Ixp33_ASAP7_75t_L g1944 ( 
.A1(n_1374),
.A2(n_1380),
.B(n_1173),
.C(n_1102),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_SL g1945 ( 
.A(n_1374),
.B(n_1380),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1374),
.B(n_1380),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1098),
.B(n_1256),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1102),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1111),
.A2(n_1257),
.B(n_1118),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1111),
.B(n_1257),
.Y(n_1950)
);

AOI21xp5_ASAP7_75t_L g1951 ( 
.A1(n_1111),
.A2(n_1257),
.B(n_1118),
.Y(n_1951)
);

INVx4_ASAP7_75t_L g1952 ( 
.A(n_1210),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1118),
.B(n_1269),
.Y(n_1953)
);

INVx3_ASAP7_75t_L g1954 ( 
.A(n_1210),
.Y(n_1954)
);

AOI21xp5_ASAP7_75t_L g1955 ( 
.A1(n_1149),
.A2(n_1272),
.B(n_1334),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1149),
.B(n_1269),
.Y(n_1956)
);

BUFx6f_ASAP7_75t_L g1957 ( 
.A(n_1386),
.Y(n_1957)
);

NOR2xp67_ASAP7_75t_L g1958 ( 
.A(n_1149),
.B(n_1272),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1166),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1166),
.B(n_1272),
.Y(n_1960)
);

INVx1_ASAP7_75t_SL g1961 ( 
.A(n_1390),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1166),
.B(n_1284),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1184),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1184),
.Y(n_1964)
);

AOI21xp5_ASAP7_75t_L g1965 ( 
.A1(n_1184),
.A2(n_1284),
.B(n_1324),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1201),
.B(n_1303),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1201),
.Y(n_1967)
);

OAI21xp5_ASAP7_75t_L g1968 ( 
.A1(n_1201),
.A2(n_1303),
.B(n_1366),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_SL g1969 ( 
.A(n_1386),
.B(n_1210),
.Y(n_1969)
);

OAI22xp5_ASAP7_75t_L g1970 ( 
.A1(n_1390),
.A2(n_1151),
.B1(n_1384),
.B2(n_1379),
.Y(n_1970)
);

AOI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1202),
.A2(n_1253),
.B(n_1205),
.Y(n_1971)
);

OAI22xp5_ASAP7_75t_L g1972 ( 
.A1(n_1202),
.A2(n_1284),
.B1(n_1323),
.B2(n_1218),
.Y(n_1972)
);

AOI21xp5_ASAP7_75t_L g1973 ( 
.A1(n_1202),
.A2(n_1253),
.B(n_1309),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1324),
.B(n_1253),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1226),
.B(n_1324),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1309),
.B(n_1250),
.Y(n_1976)
);

OAI21xp5_ASAP7_75t_L g1977 ( 
.A1(n_1226),
.A2(n_1303),
.B(n_1307),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1309),
.B(n_1236),
.Y(n_1978)
);

OAI21xp33_ASAP7_75t_L g1979 ( 
.A1(n_1250),
.A2(n_1304),
.B(n_1307),
.Y(n_1979)
);

INVx3_ASAP7_75t_L g1980 ( 
.A(n_1210),
.Y(n_1980)
);

AOI21xp5_ASAP7_75t_L g1981 ( 
.A1(n_1304),
.A2(n_1307),
.B(n_1210),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1304),
.B(n_1004),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1004),
.B(n_1210),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1004),
.B(n_1016),
.Y(n_1984)
);

NOR2xp33_ASAP7_75t_L g1985 ( 
.A(n_1054),
.B(n_408),
.Y(n_1985)
);

OAI21xp5_ASAP7_75t_L g1986 ( 
.A1(n_1012),
.A2(n_437),
.B(n_802),
.Y(n_1986)
);

AOI22xp33_ASAP7_75t_L g1987 ( 
.A1(n_1019),
.A2(n_679),
.B1(n_750),
.B2(n_669),
.Y(n_1987)
);

AOI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1214),
.A2(n_622),
.B(n_802),
.Y(n_1988)
);

A2O1A1Ixp33_ASAP7_75t_L g1989 ( 
.A1(n_1054),
.A2(n_669),
.B(n_680),
.C(n_660),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1016),
.B(n_984),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1221),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1221),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_SL g1993 ( 
.A(n_998),
.B(n_660),
.Y(n_1993)
);

OAI21xp33_ASAP7_75t_L g1994 ( 
.A1(n_1054),
.A2(n_955),
.B(n_669),
.Y(n_1994)
);

A2O1A1Ixp33_ASAP7_75t_L g1995 ( 
.A1(n_1054),
.A2(n_669),
.B(n_680),
.C(n_660),
.Y(n_1995)
);

INVx1_ASAP7_75t_SL g1996 ( 
.A(n_1145),
.Y(n_1996)
);

AOI21x1_ASAP7_75t_L g1997 ( 
.A1(n_1569),
.A2(n_1427),
.B(n_1458),
.Y(n_1997)
);

AOI21xp5_ASAP7_75t_L g1998 ( 
.A1(n_1579),
.A2(n_1455),
.B(n_1412),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1450),
.B(n_1436),
.Y(n_1999)
);

AOI21xp5_ASAP7_75t_L g2000 ( 
.A1(n_1455),
.A2(n_1412),
.B(n_1415),
.Y(n_2000)
);

AOI22xp5_ASAP7_75t_L g2001 ( 
.A1(n_1788),
.A2(n_1995),
.B1(n_1989),
.B2(n_1993),
.Y(n_2001)
);

NOR3xp33_ASAP7_75t_L g2002 ( 
.A(n_1788),
.B(n_1705),
.C(n_1656),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_SL g2003 ( 
.A(n_1420),
.B(n_1437),
.Y(n_2003)
);

AOI21xp5_ASAP7_75t_L g2004 ( 
.A1(n_1415),
.A2(n_1440),
.B(n_1435),
.Y(n_2004)
);

AOI21xp5_ASAP7_75t_L g2005 ( 
.A1(n_1415),
.A2(n_1440),
.B(n_1435),
.Y(n_2005)
);

NOR2xp33_ASAP7_75t_L g2006 ( 
.A(n_1985),
.B(n_1595),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1404),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1407),
.Y(n_2008)
);

OR2x6_ASAP7_75t_L g2009 ( 
.A(n_1655),
.B(n_1407),
.Y(n_2009)
);

NOR2xp67_ASAP7_75t_L g2010 ( 
.A(n_1655),
.B(n_1923),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_SL g2011 ( 
.A(n_1454),
.B(n_1994),
.Y(n_2011)
);

AND2x4_ASAP7_75t_L g2012 ( 
.A(n_1726),
.B(n_1732),
.Y(n_2012)
);

A2O1A1Ixp33_ASAP7_75t_L g2013 ( 
.A1(n_1994),
.A2(n_1515),
.B(n_1539),
.C(n_1464),
.Y(n_2013)
);

O2A1O1Ixp33_ASAP7_75t_L g2014 ( 
.A1(n_1493),
.A2(n_1573),
.B(n_1713),
.C(n_1705),
.Y(n_2014)
);

AOI22xp5_ASAP7_75t_L g2015 ( 
.A1(n_1987),
.A2(n_1527),
.B1(n_1599),
.B2(n_1514),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1990),
.B(n_1783),
.Y(n_2016)
);

NAND2xp33_ASAP7_75t_L g2017 ( 
.A(n_1533),
.B(n_1542),
.Y(n_2017)
);

NOR2xp33_ASAP7_75t_L g2018 ( 
.A(n_1679),
.B(n_1654),
.Y(n_2018)
);

NOR2xp33_ASAP7_75t_L g2019 ( 
.A(n_1615),
.B(n_1470),
.Y(n_2019)
);

NOR2xp33_ASAP7_75t_L g2020 ( 
.A(n_1553),
.B(n_1700),
.Y(n_2020)
);

NOR2xp33_ASAP7_75t_L g2021 ( 
.A(n_1519),
.B(n_1644),
.Y(n_2021)
);

AOI22xp5_ASAP7_75t_L g2022 ( 
.A1(n_1527),
.A2(n_1514),
.B1(n_1525),
.B2(n_1464),
.Y(n_2022)
);

OAI22xp5_ASAP7_75t_L g2023 ( 
.A1(n_1415),
.A2(n_1440),
.B1(n_1618),
.B2(n_1435),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1407),
.Y(n_2024)
);

INVx4_ASAP7_75t_L g2025 ( 
.A(n_1435),
.Y(n_2025)
);

AO21x1_ASAP7_75t_L g2026 ( 
.A1(n_1803),
.A2(n_1419),
.B(n_1453),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_SL g2027 ( 
.A(n_1440),
.B(n_1618),
.Y(n_2027)
);

OAI22xp5_ASAP7_75t_L g2028 ( 
.A1(n_1618),
.A2(n_1585),
.B1(n_1407),
.B2(n_1990),
.Y(n_2028)
);

BUFx3_ASAP7_75t_L g2029 ( 
.A(n_1576),
.Y(n_2029)
);

AOI21xp5_ASAP7_75t_L g2030 ( 
.A1(n_1618),
.A2(n_1417),
.B(n_1414),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1783),
.B(n_1431),
.Y(n_2031)
);

OAI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_1442),
.A2(n_1473),
.B(n_1849),
.Y(n_2032)
);

AOI22xp5_ASAP7_75t_L g2033 ( 
.A1(n_1585),
.A2(n_1855),
.B1(n_1752),
.B2(n_1840),
.Y(n_2033)
);

OAI21xp5_ASAP7_75t_L g2034 ( 
.A1(n_1473),
.A2(n_1849),
.B(n_1780),
.Y(n_2034)
);

AOI21x1_ASAP7_75t_L g2035 ( 
.A1(n_1569),
.A2(n_1427),
.B(n_1458),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_SL g2036 ( 
.A(n_1940),
.B(n_1486),
.Y(n_2036)
);

AND2x4_ASAP7_75t_L g2037 ( 
.A(n_1726),
.B(n_1732),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1404),
.Y(n_2038)
);

OAI22xp5_ASAP7_75t_L g2039 ( 
.A1(n_1407),
.A2(n_1431),
.B1(n_1793),
.B2(n_1603),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1826),
.B(n_1827),
.Y(n_2040)
);

NOR2xp33_ASAP7_75t_SL g2041 ( 
.A(n_1655),
.B(n_1552),
.Y(n_2041)
);

OAI22xp5_ASAP7_75t_L g2042 ( 
.A1(n_1793),
.A2(n_1603),
.B1(n_1647),
.B2(n_1552),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1826),
.B(n_1827),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1991),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1857),
.B(n_1441),
.Y(n_2045)
);

INVx3_ASAP7_75t_L g2046 ( 
.A(n_1655),
.Y(n_2046)
);

OAI22xp5_ASAP7_75t_L g2047 ( 
.A1(n_1647),
.A2(n_1855),
.B1(n_1656),
.B2(n_1566),
.Y(n_2047)
);

AOI21xp5_ASAP7_75t_L g2048 ( 
.A1(n_1414),
.A2(n_1417),
.B(n_1447),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1857),
.B(n_1441),
.Y(n_2049)
);

AO22x1_ASAP7_75t_L g2050 ( 
.A1(n_1474),
.A2(n_1421),
.B1(n_1591),
.B2(n_1577),
.Y(n_2050)
);

OAI22xp5_ASAP7_75t_L g2051 ( 
.A1(n_1558),
.A2(n_1566),
.B1(n_1652),
.B2(n_1542),
.Y(n_2051)
);

NOR2xp33_ASAP7_75t_L g2052 ( 
.A(n_1513),
.B(n_1522),
.Y(n_2052)
);

O2A1O1Ixp33_ASAP7_75t_L g2053 ( 
.A1(n_1564),
.A2(n_1558),
.B(n_1790),
.C(n_1606),
.Y(n_2053)
);

AOI21xp5_ASAP7_75t_L g2054 ( 
.A1(n_1447),
.A2(n_1528),
.B(n_1460),
.Y(n_2054)
);

OA21x2_ASAP7_75t_L g2055 ( 
.A1(n_1986),
.A2(n_1445),
.B(n_1531),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1443),
.B(n_1430),
.Y(n_2056)
);

BUFx2_ASAP7_75t_L g2057 ( 
.A(n_1771),
.Y(n_2057)
);

AOI21x1_ASAP7_75t_L g2058 ( 
.A1(n_1408),
.A2(n_1472),
.B(n_1638),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_SL g2059 ( 
.A(n_1486),
.B(n_1862),
.Y(n_2059)
);

AOI21xp5_ASAP7_75t_L g2060 ( 
.A1(n_1460),
.A2(n_1860),
.B(n_1676),
.Y(n_2060)
);

BUFx12f_ASAP7_75t_L g2061 ( 
.A(n_1561),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1443),
.B(n_1430),
.Y(n_2062)
);

NOR2xp33_ASAP7_75t_L g2063 ( 
.A(n_1593),
.B(n_1970),
.Y(n_2063)
);

OAI22xp5_ASAP7_75t_L g2064 ( 
.A1(n_1652),
.A2(n_1533),
.B1(n_1433),
.B2(n_1567),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1851),
.B(n_1429),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1851),
.B(n_1429),
.Y(n_2066)
);

NAND2x1p5_ASAP7_75t_L g2067 ( 
.A(n_1934),
.B(n_1665),
.Y(n_2067)
);

AOI21xp5_ASAP7_75t_L g2068 ( 
.A1(n_1860),
.A2(n_1676),
.B(n_1600),
.Y(n_2068)
);

AOI21xp5_ASAP7_75t_L g2069 ( 
.A1(n_1600),
.A2(n_1410),
.B(n_1841),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1459),
.B(n_1461),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1409),
.Y(n_2071)
);

OAI21xp33_ASAP7_75t_L g2072 ( 
.A1(n_1789),
.A2(n_1445),
.B(n_1780),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1404),
.Y(n_2073)
);

AOI21xp5_ASAP7_75t_L g2074 ( 
.A1(n_1410),
.A2(n_1841),
.B(n_1852),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1459),
.B(n_1461),
.Y(n_2075)
);

OAI21xp5_ASAP7_75t_L g2076 ( 
.A1(n_1411),
.A2(n_1425),
.B(n_1424),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1462),
.B(n_1463),
.Y(n_2077)
);

BUFx6f_ASAP7_75t_L g2078 ( 
.A(n_1426),
.Y(n_2078)
);

BUFx2_ASAP7_75t_L g2079 ( 
.A(n_1771),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1462),
.B(n_1463),
.Y(n_2080)
);

NOR2xp33_ASAP7_75t_L g2081 ( 
.A(n_1970),
.B(n_1839),
.Y(n_2081)
);

NOR3xp33_ASAP7_75t_L g2082 ( 
.A(n_1641),
.B(n_1795),
.C(n_1729),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_1450),
.B(n_1436),
.Y(n_2083)
);

AOI21xp5_ASAP7_75t_L g2084 ( 
.A1(n_1852),
.A2(n_1858),
.B(n_1854),
.Y(n_2084)
);

INVx3_ASAP7_75t_L g2085 ( 
.A(n_1421),
.Y(n_2085)
);

A2O1A1Ixp33_ASAP7_75t_L g2086 ( 
.A1(n_1825),
.A2(n_1511),
.B(n_1591),
.C(n_1549),
.Y(n_2086)
);

NOR2xp33_ASAP7_75t_L g2087 ( 
.A(n_1899),
.B(n_1908),
.Y(n_2087)
);

NOR2xp33_ASAP7_75t_L g2088 ( 
.A(n_1961),
.B(n_1802),
.Y(n_2088)
);

AOI21xp5_ASAP7_75t_L g2089 ( 
.A1(n_1854),
.A2(n_1859),
.B(n_1858),
.Y(n_2089)
);

AOI21xp5_ASAP7_75t_L g2090 ( 
.A1(n_1859),
.A2(n_1836),
.B(n_1833),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1409),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1688),
.B(n_1701),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_1452),
.B(n_1413),
.Y(n_2093)
);

BUFx3_ASAP7_75t_L g2094 ( 
.A(n_1576),
.Y(n_2094)
);

AOI33xp33_ASAP7_75t_L g2095 ( 
.A1(n_1627),
.A2(n_1767),
.A3(n_1692),
.B1(n_1702),
.B2(n_1488),
.B3(n_1413),
.Y(n_2095)
);

INVx1_ASAP7_75t_SL g2096 ( 
.A(n_1775),
.Y(n_2096)
);

AOI33xp33_ASAP7_75t_L g2097 ( 
.A1(n_1692),
.A2(n_1488),
.A3(n_1444),
.B1(n_1535),
.B2(n_1532),
.B3(n_1501),
.Y(n_2097)
);

AOI21xp5_ASAP7_75t_L g2098 ( 
.A1(n_1833),
.A2(n_1836),
.B(n_1988),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1688),
.B(n_1701),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_SL g2100 ( 
.A(n_1862),
.B(n_1984),
.Y(n_2100)
);

AND2x4_ASAP7_75t_L g2101 ( 
.A(n_1726),
.B(n_1732),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1716),
.B(n_1719),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_SL g2103 ( 
.A(n_1862),
.B(n_1984),
.Y(n_2103)
);

INVx1_ASAP7_75t_SL g2104 ( 
.A(n_1775),
.Y(n_2104)
);

BUFx10_ASAP7_75t_L g2105 ( 
.A(n_1438),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1716),
.B(n_1719),
.Y(n_2106)
);

BUFx3_ASAP7_75t_L g2107 ( 
.A(n_1576),
.Y(n_2107)
);

AO32x1_ASAP7_75t_L g2108 ( 
.A1(n_1411),
.A2(n_1803),
.A3(n_1972),
.B1(n_1453),
.B2(n_1840),
.Y(n_2108)
);

NOR2xp33_ASAP7_75t_L g2109 ( 
.A(n_1961),
.B(n_1802),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1469),
.Y(n_2110)
);

NOR2xp33_ASAP7_75t_L g2111 ( 
.A(n_1706),
.B(n_1626),
.Y(n_2111)
);

HB1xp67_ASAP7_75t_L g2112 ( 
.A(n_1674),
.Y(n_2112)
);

A2O1A1Ixp33_ASAP7_75t_L g2113 ( 
.A1(n_1825),
.A2(n_1547),
.B(n_1526),
.C(n_1646),
.Y(n_2113)
);

AOI21xp5_ASAP7_75t_L g2114 ( 
.A1(n_1988),
.A2(n_1986),
.B(n_1448),
.Y(n_2114)
);

AOI21xp5_ASAP7_75t_L g2115 ( 
.A1(n_1448),
.A2(n_1682),
.B(n_1479),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1469),
.Y(n_2116)
);

AOI21xp5_ASAP7_75t_L g2117 ( 
.A1(n_1682),
.A2(n_1479),
.B(n_1423),
.Y(n_2117)
);

BUFx3_ASAP7_75t_L g2118 ( 
.A(n_1577),
.Y(n_2118)
);

NOR2xp33_ASAP7_75t_L g2119 ( 
.A(n_1766),
.B(n_1807),
.Y(n_2119)
);

NOR2xp33_ASAP7_75t_L g2120 ( 
.A(n_1597),
.B(n_1561),
.Y(n_2120)
);

INVx5_ASAP7_75t_L g2121 ( 
.A(n_1421),
.Y(n_2121)
);

BUFx2_ASAP7_75t_L g2122 ( 
.A(n_1686),
.Y(n_2122)
);

NAND2x1p5_ASAP7_75t_L g2123 ( 
.A(n_1934),
.B(n_1665),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_SL g2124 ( 
.A(n_1862),
.B(n_1665),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1444),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_1452),
.B(n_1501),
.Y(n_2126)
);

AOI21xp5_ASAP7_75t_L g2127 ( 
.A1(n_1423),
.A2(n_1820),
.B(n_1432),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1773),
.B(n_1798),
.Y(n_2128)
);

OAI21xp5_ASAP7_75t_L g2129 ( 
.A1(n_1425),
.A2(n_1424),
.B(n_1720),
.Y(n_2129)
);

O2A1O1Ixp33_ASAP7_75t_L g2130 ( 
.A1(n_1641),
.A2(n_1651),
.B(n_1628),
.C(n_1898),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1773),
.B(n_1798),
.Y(n_2131)
);

NOR2xp33_ASAP7_75t_L g2132 ( 
.A(n_1561),
.B(n_1725),
.Y(n_2132)
);

A2O1A1Ixp33_ASAP7_75t_L g2133 ( 
.A1(n_1547),
.A2(n_1526),
.B(n_1646),
.C(n_1809),
.Y(n_2133)
);

AO22x1_ASAP7_75t_L g2134 ( 
.A1(n_1474),
.A2(n_1421),
.B1(n_1620),
.B2(n_1577),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1811),
.B(n_1868),
.Y(n_2135)
);

AOI21xp5_ASAP7_75t_L g2136 ( 
.A1(n_1820),
.A2(n_1432),
.B(n_1428),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_SL g2137 ( 
.A(n_1665),
.B(n_1772),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_1811),
.B(n_1868),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1469),
.Y(n_2139)
);

NOR2xp33_ASAP7_75t_L g2140 ( 
.A(n_1725),
.B(n_1777),
.Y(n_2140)
);

AOI21xp5_ASAP7_75t_L g2141 ( 
.A1(n_1428),
.A2(n_1813),
.B(n_1814),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_SL g2142 ( 
.A(n_1772),
.B(n_1834),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_1532),
.B(n_1535),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_1541),
.B(n_1559),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_1481),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1481),
.Y(n_2146)
);

OAI22xp5_ASAP7_75t_SL g2147 ( 
.A1(n_1568),
.A2(n_1935),
.B1(n_1649),
.B2(n_1756),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1541),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_SL g2149 ( 
.A(n_1772),
.B(n_1834),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1559),
.Y(n_2150)
);

INVx3_ASAP7_75t_L g2151 ( 
.A(n_1421),
.Y(n_2151)
);

A2O1A1Ixp33_ASAP7_75t_SL g2152 ( 
.A1(n_1782),
.A2(n_1792),
.B(n_1434),
.C(n_1806),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_1570),
.B(n_1574),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1481),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1872),
.B(n_1873),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_1505),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_SL g2157 ( 
.A(n_1772),
.B(n_1834),
.Y(n_2157)
);

NAND3xp33_ASAP7_75t_SL g2158 ( 
.A(n_1853),
.B(n_1746),
.C(n_1601),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_1872),
.B(n_1873),
.Y(n_2159)
);

NOR2xp33_ASAP7_75t_L g2160 ( 
.A(n_1725),
.B(n_1777),
.Y(n_2160)
);

INVx4_ASAP7_75t_L g2161 ( 
.A(n_1421),
.Y(n_2161)
);

O2A1O1Ixp33_ASAP7_75t_L g2162 ( 
.A1(n_1898),
.A2(n_1884),
.B(n_1888),
.C(n_1883),
.Y(n_2162)
);

NOR2xp33_ASAP7_75t_SL g2163 ( 
.A(n_1935),
.B(n_1746),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_SL g2164 ( 
.A(n_1834),
.B(n_1853),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_1876),
.B(n_1887),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_1876),
.B(n_1887),
.Y(n_2166)
);

OAI22xp5_ASAP7_75t_L g2167 ( 
.A1(n_1433),
.A2(n_1645),
.B1(n_1724),
.B2(n_1722),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_1892),
.B(n_1896),
.Y(n_2168)
);

INVx2_ASAP7_75t_SL g2169 ( 
.A(n_1875),
.Y(n_2169)
);

AOI21xp5_ASAP7_75t_L g2170 ( 
.A1(n_1813),
.A2(n_1814),
.B(n_1863),
.Y(n_2170)
);

OAI22xp5_ASAP7_75t_L g2171 ( 
.A1(n_1645),
.A2(n_1722),
.B1(n_1730),
.B2(n_1724),
.Y(n_2171)
);

AOI21xp5_ASAP7_75t_L g2172 ( 
.A1(n_1863),
.A2(n_1681),
.B(n_1571),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_1892),
.B(n_1896),
.Y(n_2173)
);

AND2x4_ASAP7_75t_L g2174 ( 
.A(n_1726),
.B(n_1732),
.Y(n_2174)
);

NOR2xp33_ASAP7_75t_L g2175 ( 
.A(n_1777),
.B(n_1869),
.Y(n_2175)
);

AOI22xp5_ASAP7_75t_L g2176 ( 
.A1(n_1578),
.A2(n_1489),
.B1(n_1418),
.B2(n_1607),
.Y(n_2176)
);

NOR2xp33_ASAP7_75t_L g2177 ( 
.A(n_1869),
.B(n_1689),
.Y(n_2177)
);

HB1xp67_ASAP7_75t_L g2178 ( 
.A(n_1747),
.Y(n_2178)
);

NOR2xp33_ASAP7_75t_SL g2179 ( 
.A(n_1935),
.B(n_1457),
.Y(n_2179)
);

AOI21xp5_ASAP7_75t_L g2180 ( 
.A1(n_1681),
.A2(n_1571),
.B(n_1562),
.Y(n_2180)
);

AOI21xp5_ASAP7_75t_L g2181 ( 
.A1(n_1562),
.A2(n_1588),
.B(n_1583),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_1446),
.B(n_1449),
.Y(n_2182)
);

HB1xp67_ASAP7_75t_L g2183 ( 
.A(n_1829),
.Y(n_2183)
);

A2O1A1Ixp33_ASAP7_75t_L g2184 ( 
.A1(n_1809),
.A2(n_1917),
.B(n_1865),
.C(n_1884),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_1570),
.B(n_1574),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_1446),
.B(n_1449),
.Y(n_2186)
);

OAI22xp5_ASAP7_75t_L g2187 ( 
.A1(n_1730),
.A2(n_1736),
.B1(n_1761),
.B2(n_1757),
.Y(n_2187)
);

OAI22xp5_ASAP7_75t_L g2188 ( 
.A1(n_1736),
.A2(n_1757),
.B1(n_1762),
.B2(n_1761),
.Y(n_2188)
);

O2A1O1Ixp33_ASAP7_75t_L g2189 ( 
.A1(n_1810),
.A2(n_1762),
.B(n_1764),
.C(n_1763),
.Y(n_2189)
);

AOI21xp5_ASAP7_75t_L g2190 ( 
.A1(n_1583),
.A2(n_1594),
.B(n_1588),
.Y(n_2190)
);

OAI22xp5_ASAP7_75t_L g2191 ( 
.A1(n_1763),
.A2(n_1764),
.B1(n_1786),
.B2(n_1779),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1845),
.B(n_1466),
.Y(n_2192)
);

AOI21xp5_ASAP7_75t_L g2193 ( 
.A1(n_1594),
.A2(n_1604),
.B(n_1598),
.Y(n_2193)
);

AOI21xp5_ASAP7_75t_L g2194 ( 
.A1(n_1598),
.A2(n_1608),
.B(n_1604),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_SL g2195 ( 
.A(n_1846),
.B(n_1663),
.Y(n_2195)
);

O2A1O1Ixp33_ASAP7_75t_SL g2196 ( 
.A1(n_1779),
.A2(n_1786),
.B(n_1800),
.C(n_1794),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_1845),
.B(n_1466),
.Y(n_2197)
);

NOR2xp33_ASAP7_75t_L g2198 ( 
.A(n_1869),
.B(n_1920),
.Y(n_2198)
);

OAI22xp5_ASAP7_75t_L g2199 ( 
.A1(n_1794),
.A2(n_1800),
.B1(n_1529),
.B2(n_1801),
.Y(n_2199)
);

NAND2x1p5_ASAP7_75t_L g2200 ( 
.A(n_1934),
.B(n_1889),
.Y(n_2200)
);

AOI21xp5_ASAP7_75t_L g2201 ( 
.A1(n_1608),
.A2(n_1619),
.B(n_1616),
.Y(n_2201)
);

OAI22xp5_ASAP7_75t_L g2202 ( 
.A1(n_1529),
.A2(n_1801),
.B1(n_1478),
.B2(n_1487),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_1468),
.B(n_1831),
.Y(n_2203)
);

AO21x1_ASAP7_75t_L g2204 ( 
.A1(n_1575),
.A2(n_1792),
.B(n_1782),
.Y(n_2204)
);

AND2x4_ASAP7_75t_L g2205 ( 
.A(n_1739),
.B(n_1867),
.Y(n_2205)
);

OR2x6_ASAP7_75t_SL g2206 ( 
.A(n_1983),
.B(n_1982),
.Y(n_2206)
);

AOI21xp5_ASAP7_75t_L g2207 ( 
.A1(n_1616),
.A2(n_1621),
.B(n_1619),
.Y(n_2207)
);

NOR3xp33_ASAP7_75t_L g2208 ( 
.A(n_1734),
.B(n_1781),
.C(n_1879),
.Y(n_2208)
);

AOI21xp5_ASAP7_75t_L g2209 ( 
.A1(n_1621),
.A2(n_1633),
.B(n_1632),
.Y(n_2209)
);

AOI21x1_ASAP7_75t_L g2210 ( 
.A1(n_1408),
.A2(n_1472),
.B(n_1638),
.Y(n_2210)
);

CKINVDCx5p33_ASAP7_75t_R g2211 ( 
.A(n_1422),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_1468),
.B(n_1831),
.Y(n_2212)
);

BUFx6f_ASAP7_75t_L g2213 ( 
.A(n_1426),
.Y(n_2213)
);

OAI22xp5_ASAP7_75t_L g2214 ( 
.A1(n_1478),
.A2(n_1487),
.B1(n_1756),
.B2(n_1649),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_1505),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_1505),
.Y(n_2216)
);

OAI21xp33_ASAP7_75t_L g2217 ( 
.A1(n_1434),
.A2(n_1406),
.B(n_1635),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_1538),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_1489),
.B(n_1584),
.Y(n_2219)
);

O2A1O1Ixp5_ASAP7_75t_L g2220 ( 
.A1(n_1846),
.A2(n_1631),
.B(n_1517),
.C(n_1720),
.Y(n_2220)
);

AOI21xp5_ASAP7_75t_L g2221 ( 
.A1(n_1632),
.A2(n_1639),
.B(n_1633),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_1584),
.B(n_1610),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1610),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_1624),
.B(n_1678),
.Y(n_2224)
);

AOI21xp5_ASAP7_75t_L g2225 ( 
.A1(n_1639),
.A2(n_1648),
.B(n_1640),
.Y(n_2225)
);

A2O1A1Ixp33_ASAP7_75t_L g2226 ( 
.A1(n_1917),
.A2(n_1865),
.B(n_1808),
.C(n_1806),
.Y(n_2226)
);

AOI21xp5_ASAP7_75t_L g2227 ( 
.A1(n_1640),
.A2(n_1648),
.B(n_1878),
.Y(n_2227)
);

NAND2xp33_ASAP7_75t_L g2228 ( 
.A(n_1421),
.B(n_1879),
.Y(n_2228)
);

NOR2x1_ASAP7_75t_L g2229 ( 
.A(n_1889),
.B(n_1983),
.Y(n_2229)
);

AOI21xp5_ASAP7_75t_L g2230 ( 
.A1(n_1878),
.A2(n_1881),
.B(n_1465),
.Y(n_2230)
);

NOR2xp33_ASAP7_75t_L g2231 ( 
.A(n_1920),
.B(n_1911),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_1538),
.Y(n_2232)
);

BUFx12f_ASAP7_75t_L g2233 ( 
.A(n_1818),
.Y(n_2233)
);

AOI21xp5_ASAP7_75t_L g2234 ( 
.A1(n_1881),
.A2(n_1465),
.B(n_1467),
.Y(n_2234)
);

OAI22xp5_ASAP7_75t_L g2235 ( 
.A1(n_1649),
.A2(n_1756),
.B1(n_1607),
.B2(n_1686),
.Y(n_2235)
);

NAND3xp33_ASAP7_75t_L g2236 ( 
.A(n_1406),
.B(n_1439),
.C(n_1485),
.Y(n_2236)
);

AOI21xp5_ASAP7_75t_L g2237 ( 
.A1(n_1467),
.A2(n_1685),
.B(n_1500),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_1624),
.B(n_1678),
.Y(n_2238)
);

AOI21xp5_ASAP7_75t_L g2239 ( 
.A1(n_1685),
.A2(n_1500),
.B(n_1494),
.Y(n_2239)
);

AND2x2_ASAP7_75t_L g2240 ( 
.A(n_1721),
.B(n_1744),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_1721),
.B(n_1744),
.Y(n_2241)
);

AOI22x1_ASAP7_75t_L g2242 ( 
.A1(n_1885),
.A2(n_1893),
.B1(n_1808),
.B2(n_1913),
.Y(n_2242)
);

BUFx6f_ASAP7_75t_L g2243 ( 
.A(n_1426),
.Y(n_2243)
);

OAI22xp5_ASAP7_75t_L g2244 ( 
.A1(n_1755),
.A2(n_1759),
.B1(n_1770),
.B2(n_1758),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_1538),
.Y(n_2245)
);

BUFx6f_ASAP7_75t_L g2246 ( 
.A(n_1426),
.Y(n_2246)
);

INVx2_ASAP7_75t_SL g2247 ( 
.A(n_1875),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_1555),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_1755),
.B(n_1758),
.Y(n_2249)
);

O2A1O1Ixp33_ASAP7_75t_L g2250 ( 
.A1(n_1485),
.A2(n_1477),
.B(n_1847),
.C(n_1828),
.Y(n_2250)
);

OAI22xp5_ASAP7_75t_L g2251 ( 
.A1(n_1759),
.A2(n_1787),
.B1(n_1796),
.B2(n_1770),
.Y(n_2251)
);

AOI21xp5_ASAP7_75t_L g2252 ( 
.A1(n_1494),
.A2(n_1504),
.B(n_1503),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_SL g2253 ( 
.A(n_1663),
.B(n_1631),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1787),
.Y(n_2254)
);

O2A1O1Ixp33_ASAP7_75t_L g2255 ( 
.A1(n_1874),
.A2(n_1439),
.B(n_1740),
.C(n_1733),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1796),
.Y(n_2256)
);

AND2x4_ASAP7_75t_L g2257 ( 
.A(n_1739),
.B(n_1867),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1555),
.Y(n_2258)
);

INVxp33_ASAP7_75t_SL g2259 ( 
.A(n_1712),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_SL g2260 ( 
.A(n_1663),
.B(n_1957),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_1837),
.B(n_1843),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_1837),
.B(n_1843),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_1850),
.B(n_1861),
.Y(n_2263)
);

NAND2x1p5_ASAP7_75t_L g2264 ( 
.A(n_1934),
.B(n_1889),
.Y(n_2264)
);

HB1xp67_ASAP7_75t_L g2265 ( 
.A(n_1848),
.Y(n_2265)
);

O2A1O1Ixp33_ASAP7_75t_L g2266 ( 
.A1(n_1760),
.A2(n_1560),
.B(n_1812),
.C(n_1635),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_SL g2267 ( 
.A(n_1663),
.B(n_1957),
.Y(n_2267)
);

OR2x6_ASAP7_75t_SL g2268 ( 
.A(n_1982),
.B(n_1848),
.Y(n_2268)
);

AOI21xp5_ASAP7_75t_L g2269 ( 
.A1(n_1503),
.A2(n_1504),
.B(n_1523),
.Y(n_2269)
);

HB1xp67_ASAP7_75t_L g2270 ( 
.A(n_1902),
.Y(n_2270)
);

AOI21xp5_ASAP7_75t_L g2271 ( 
.A1(n_1650),
.A2(n_1484),
.B(n_1480),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_1850),
.B(n_1861),
.Y(n_2272)
);

OAI21xp5_ASAP7_75t_L g2273 ( 
.A1(n_1731),
.A2(n_1738),
.B(n_1737),
.Y(n_2273)
);

AOI22x1_ASAP7_75t_L g2274 ( 
.A1(n_1885),
.A2(n_1893),
.B1(n_1913),
.B2(n_1506),
.Y(n_2274)
);

AOI21xp5_ASAP7_75t_L g2275 ( 
.A1(n_1650),
.A2(n_1484),
.B(n_1480),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_SL g2276 ( 
.A(n_1957),
.B(n_1871),
.Y(n_2276)
);

AOI21xp5_ASAP7_75t_L g2277 ( 
.A1(n_1491),
.A2(n_1492),
.B(n_1530),
.Y(n_2277)
);

A2O1A1Ixp33_ASAP7_75t_L g2278 ( 
.A1(n_1914),
.A2(n_1871),
.B(n_1921),
.C(n_1923),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_1864),
.B(n_1894),
.Y(n_2279)
);

NOR2xp67_ASAP7_75t_SL g2280 ( 
.A(n_1620),
.B(n_1661),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_1864),
.B(n_1894),
.Y(n_2281)
);

BUFx12f_ASAP7_75t_L g2282 ( 
.A(n_1818),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_SL g2283 ( 
.A(n_1957),
.B(n_1889),
.Y(n_2283)
);

OAI21xp5_ASAP7_75t_L g2284 ( 
.A1(n_1731),
.A2(n_1738),
.B(n_1737),
.Y(n_2284)
);

OAI22xp5_ASAP7_75t_L g2285 ( 
.A1(n_1897),
.A2(n_1992),
.B1(n_1991),
.B2(n_1498),
.Y(n_2285)
);

NOR2xp33_ASAP7_75t_L g2286 ( 
.A(n_1911),
.B(n_1750),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_SL g2287 ( 
.A(n_1957),
.B(n_1749),
.Y(n_2287)
);

CKINVDCx5p33_ASAP7_75t_R g2288 ( 
.A(n_1422),
.Y(n_2288)
);

OAI21xp33_ASAP7_75t_L g2289 ( 
.A1(n_1490),
.A2(n_1498),
.B(n_1581),
.Y(n_2289)
);

INVxp67_ASAP7_75t_L g2290 ( 
.A(n_1890),
.Y(n_2290)
);

AOI21xp5_ASAP7_75t_L g2291 ( 
.A1(n_1491),
.A2(n_1492),
.B(n_1530),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_1897),
.B(n_1992),
.Y(n_2292)
);

NAND3xp33_ASAP7_75t_L g2293 ( 
.A(n_1919),
.B(n_1907),
.C(n_1742),
.Y(n_2293)
);

CKINVDCx20_ASAP7_75t_R g2294 ( 
.A(n_1818),
.Y(n_2294)
);

AOI21xp5_ASAP7_75t_L g2295 ( 
.A1(n_1536),
.A2(n_1544),
.B(n_1537),
.Y(n_2295)
);

O2A1O1Ixp33_ASAP7_75t_L g2296 ( 
.A1(n_1475),
.A2(n_1623),
.B(n_1586),
.C(n_1907),
.Y(n_2296)
);

AOI22x1_ASAP7_75t_L g2297 ( 
.A1(n_1506),
.A2(n_1512),
.B1(n_1904),
.B2(n_1537),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_1555),
.B(n_1617),
.Y(n_2298)
);

OAI22x1_ASAP7_75t_L g2299 ( 
.A1(n_1824),
.A2(n_1891),
.B1(n_1922),
.B2(n_1717),
.Y(n_2299)
);

AO21x1_ASAP7_75t_L g2300 ( 
.A1(n_1512),
.A2(n_1475),
.B(n_1667),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_1617),
.B(n_1657),
.Y(n_2301)
);

CKINVDCx5p33_ASAP7_75t_R g2302 ( 
.A(n_1642),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_1617),
.Y(n_2303)
);

A2O1A1Ixp33_ASAP7_75t_L g2304 ( 
.A1(n_1914),
.A2(n_1921),
.B(n_1563),
.C(n_1943),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_L g2305 ( 
.A(n_1657),
.B(n_1960),
.Y(n_2305)
);

AOI21xp5_ASAP7_75t_L g2306 ( 
.A1(n_1536),
.A2(n_1544),
.B(n_1476),
.Y(n_2306)
);

AOI21xp5_ASAP7_75t_L g2307 ( 
.A1(n_1523),
.A2(n_1540),
.B(n_1534),
.Y(n_2307)
);

O2A1O1Ixp33_ASAP7_75t_L g2308 ( 
.A1(n_1815),
.A2(n_1817),
.B(n_1490),
.C(n_1510),
.Y(n_2308)
);

OR2x2_ASAP7_75t_L g2309 ( 
.A(n_1563),
.B(n_1824),
.Y(n_2309)
);

INVx4_ASAP7_75t_SL g2310 ( 
.A(n_1421),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_1657),
.B(n_1960),
.Y(n_2311)
);

BUFx6f_ASAP7_75t_SL g2312 ( 
.A(n_1620),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_1664),
.Y(n_2313)
);

AOI21x1_ASAP7_75t_L g2314 ( 
.A1(n_1643),
.A2(n_1582),
.B(n_1707),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_1664),
.Y(n_2315)
);

AOI21xp5_ASAP7_75t_L g2316 ( 
.A1(n_1534),
.A2(n_1540),
.B(n_1476),
.Y(n_2316)
);

AOI22xp5_ASAP7_75t_L g2317 ( 
.A1(n_1516),
.A2(n_1922),
.B1(n_1891),
.B2(n_1712),
.Y(n_2317)
);

AOI21xp5_ASAP7_75t_L g2318 ( 
.A1(n_1483),
.A2(n_1708),
.B(n_1634),
.Y(n_2318)
);

BUFx4f_ASAP7_75t_L g2319 ( 
.A(n_1421),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_SL g2320 ( 
.A(n_1957),
.B(n_1749),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_1912),
.Y(n_2321)
);

OAI21x1_ASAP7_75t_L g2322 ( 
.A1(n_1981),
.A2(n_1582),
.B(n_1707),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_1664),
.Y(n_2323)
);

A2O1A1Ixp33_ASAP7_75t_L g2324 ( 
.A1(n_1903),
.A2(n_1622),
.B(n_1723),
.C(n_1550),
.Y(n_2324)
);

AOI21xp5_ASAP7_75t_L g2325 ( 
.A1(n_1483),
.A2(n_1708),
.B(n_1634),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_1695),
.Y(n_2326)
);

OAI21xp33_ASAP7_75t_L g2327 ( 
.A1(n_1581),
.A2(n_1587),
.B(n_1497),
.Y(n_2327)
);

OAI22xp5_ASAP7_75t_L g2328 ( 
.A1(n_1508),
.A2(n_1510),
.B1(n_1516),
.B2(n_1483),
.Y(n_2328)
);

NAND3xp33_ASAP7_75t_SL g2329 ( 
.A(n_1715),
.B(n_1735),
.C(n_1769),
.Y(n_2329)
);

AOI21xp5_ASAP7_75t_L g2330 ( 
.A1(n_1483),
.A2(n_1708),
.B(n_1637),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_1508),
.B(n_1471),
.Y(n_2331)
);

OAI22xp5_ASAP7_75t_SL g2332 ( 
.A1(n_1830),
.A2(n_1750),
.B1(n_1691),
.B2(n_1661),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_1695),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_SL g2334 ( 
.A(n_1749),
.B(n_1799),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_1471),
.B(n_1996),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_1695),
.Y(n_2336)
);

O2A1O1Ixp33_ASAP7_75t_L g2337 ( 
.A1(n_1741),
.A2(n_1743),
.B(n_1751),
.C(n_1742),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_1996),
.B(n_1902),
.Y(n_2338)
);

AOI22xp5_ASAP7_75t_L g2339 ( 
.A1(n_1715),
.A2(n_1735),
.B1(n_1769),
.B2(n_1622),
.Y(n_2339)
);

AOI21xp5_ASAP7_75t_L g2340 ( 
.A1(n_1483),
.A2(n_1708),
.B(n_1637),
.Y(n_2340)
);

AOI21xp5_ASAP7_75t_L g2341 ( 
.A1(n_1483),
.A2(n_1708),
.B(n_1587),
.Y(n_2341)
);

AOI21xp5_ASAP7_75t_L g2342 ( 
.A1(n_1708),
.A2(n_1502),
.B(n_1507),
.Y(n_2342)
);

AOI21xp5_ASAP7_75t_L g2343 ( 
.A1(n_1502),
.A2(n_1509),
.B(n_1507),
.Y(n_2343)
);

AOI21xp5_ASAP7_75t_L g2344 ( 
.A1(n_1509),
.A2(n_1981),
.B(n_1556),
.Y(n_2344)
);

AO22x1_ASAP7_75t_L g2345 ( 
.A1(n_1474),
.A2(n_1691),
.B1(n_1661),
.B2(n_1939),
.Y(n_2345)
);

OAI22xp5_ASAP7_75t_L g2346 ( 
.A1(n_1548),
.A2(n_1556),
.B1(n_1609),
.B2(n_1565),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_1895),
.B(n_1609),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_1895),
.B(n_1941),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_1728),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_1941),
.B(n_1947),
.Y(n_2350)
);

INVx4_ASAP7_75t_L g2351 ( 
.A(n_1625),
.Y(n_2351)
);

AOI21xp5_ASAP7_75t_L g2352 ( 
.A1(n_1548),
.A2(n_1659),
.B(n_1658),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_1728),
.Y(n_2353)
);

AOI21xp5_ASAP7_75t_L g2354 ( 
.A1(n_1658),
.A2(n_1668),
.B(n_1659),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_1947),
.B(n_1950),
.Y(n_2355)
);

OAI21xp5_ASAP7_75t_L g2356 ( 
.A1(n_1741),
.A2(n_1751),
.B(n_1743),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_SL g2357 ( 
.A(n_1749),
.B(n_1799),
.Y(n_2357)
);

OAI22xp5_ASAP7_75t_L g2358 ( 
.A1(n_1565),
.A2(n_1543),
.B1(n_1546),
.B2(n_1629),
.Y(n_2358)
);

OR2x6_ASAP7_75t_L g2359 ( 
.A(n_1625),
.B(n_1709),
.Y(n_2359)
);

O2A1O1Ixp33_ASAP7_75t_L g2360 ( 
.A1(n_1753),
.A2(n_1711),
.B(n_1710),
.C(n_1718),
.Y(n_2360)
);

NOR2x1_ASAP7_75t_R g2361 ( 
.A(n_1691),
.B(n_1457),
.Y(n_2361)
);

AOI21x1_ASAP7_75t_L g2362 ( 
.A1(n_1643),
.A2(n_1711),
.B(n_1710),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_1950),
.B(n_1953),
.Y(n_2363)
);

O2A1O1Ixp33_ASAP7_75t_L g2364 ( 
.A1(n_1753),
.A2(n_1718),
.B(n_1554),
.C(n_1612),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_1953),
.B(n_1956),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_1728),
.Y(n_2366)
);

BUFx12f_ASAP7_75t_L g2367 ( 
.A(n_1818),
.Y(n_2367)
);

A2O1A1Ixp33_ASAP7_75t_SL g2368 ( 
.A1(n_1904),
.A2(n_1906),
.B(n_1683),
.C(n_1687),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_SL g2369 ( 
.A(n_1799),
.B(n_1877),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_SL g2370 ( 
.A(n_1799),
.B(n_1877),
.Y(n_2370)
);

CKINVDCx5p33_ASAP7_75t_R g2371 ( 
.A(n_1642),
.Y(n_2371)
);

NOR3xp33_ASAP7_75t_L g2372 ( 
.A(n_1797),
.B(n_1822),
.C(n_1774),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_1956),
.B(n_1962),
.Y(n_2373)
);

NOR2xp33_ASAP7_75t_L g2374 ( 
.A(n_1774),
.B(n_1822),
.Y(n_2374)
);

NOR2xp33_ASAP7_75t_L g2375 ( 
.A(n_1774),
.B(n_1822),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_1962),
.B(n_1966),
.Y(n_2376)
);

BUFx6f_ASAP7_75t_L g2377 ( 
.A(n_1426),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_1745),
.Y(n_2378)
);

NOR2xp33_ASAP7_75t_L g2379 ( 
.A(n_1774),
.B(n_1822),
.Y(n_2379)
);

CKINVDCx14_ASAP7_75t_R g2380 ( 
.A(n_1901),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_SL g2381 ( 
.A(n_1877),
.B(n_1933),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_1966),
.B(n_1974),
.Y(n_2382)
);

INVx2_ASAP7_75t_SL g2383 ( 
.A(n_1934),
.Y(n_2383)
);

OR2x6_ASAP7_75t_L g2384 ( 
.A(n_1625),
.B(n_1709),
.Y(n_2384)
);

AOI21xp5_ASAP7_75t_L g2385 ( 
.A1(n_1668),
.A2(n_1675),
.B(n_1673),
.Y(n_2385)
);

OAI22xp5_ASAP7_75t_L g2386 ( 
.A1(n_1543),
.A2(n_1546),
.B1(n_1629),
.B2(n_1592),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_1974),
.B(n_1975),
.Y(n_2387)
);

AOI21xp5_ASAP7_75t_L g2388 ( 
.A1(n_1673),
.A2(n_1677),
.B(n_1675),
.Y(n_2388)
);

BUFx2_ASAP7_75t_L g2389 ( 
.A(n_1870),
.Y(n_2389)
);

BUFx3_ASAP7_75t_L g2390 ( 
.A(n_1474),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_1975),
.B(n_1976),
.Y(n_2391)
);

A2O1A1Ixp33_ASAP7_75t_L g2392 ( 
.A1(n_1903),
.A2(n_1723),
.B(n_1550),
.C(n_1754),
.Y(n_2392)
);

NOR2xp33_ASAP7_75t_R g2393 ( 
.A(n_1778),
.B(n_1791),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_1976),
.B(n_1978),
.Y(n_2394)
);

AOI21x1_ASAP7_75t_L g2395 ( 
.A1(n_1703),
.A2(n_1694),
.B(n_1653),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_1978),
.B(n_1963),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_1963),
.B(n_1964),
.Y(n_2397)
);

NOR3xp33_ASAP7_75t_L g2398 ( 
.A(n_1930),
.B(n_1816),
.C(n_1613),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_1745),
.Y(n_2399)
);

OAI22xp5_ASAP7_75t_L g2400 ( 
.A1(n_1580),
.A2(n_1592),
.B1(n_1589),
.B2(n_1704),
.Y(n_2400)
);

NOR2xp33_ASAP7_75t_L g2401 ( 
.A(n_1704),
.B(n_1901),
.Y(n_2401)
);

OAI22xp5_ASAP7_75t_L g2402 ( 
.A1(n_1580),
.A2(n_1589),
.B1(n_1636),
.B2(n_1518),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_1745),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_1748),
.Y(n_2404)
);

AOI21xp5_ASAP7_75t_L g2405 ( 
.A1(n_1677),
.A2(n_1687),
.B(n_1683),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_SL g2406 ( 
.A(n_1877),
.B(n_1933),
.Y(n_2406)
);

INVx4_ASAP7_75t_L g2407 ( 
.A(n_1625),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_1964),
.B(n_1748),
.Y(n_2408)
);

BUFx4f_ASAP7_75t_L g2409 ( 
.A(n_1451),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_1748),
.B(n_1765),
.Y(n_2410)
);

NOR2xp33_ASAP7_75t_L g2411 ( 
.A(n_1739),
.B(n_1867),
.Y(n_2411)
);

INVx11_ASAP7_75t_L g2412 ( 
.A(n_1660),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_1765),
.Y(n_2413)
);

AND2x4_ASAP7_75t_L g2414 ( 
.A(n_1739),
.B(n_1867),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_1765),
.Y(n_2415)
);

NOR2xp33_ASAP7_75t_L g2416 ( 
.A(n_1572),
.B(n_1905),
.Y(n_2416)
);

OAI22xp5_ASAP7_75t_L g2417 ( 
.A1(n_1636),
.A2(n_1495),
.B1(n_1518),
.B2(n_1497),
.Y(n_2417)
);

AOI22xp5_ASAP7_75t_L g2418 ( 
.A1(n_1572),
.A2(n_1909),
.B1(n_1905),
.B2(n_1754),
.Y(n_2418)
);

INVx5_ASAP7_75t_L g2419 ( 
.A(n_1660),
.Y(n_2419)
);

NOR2xp67_ASAP7_75t_L g2420 ( 
.A(n_1934),
.B(n_1927),
.Y(n_2420)
);

A2O1A1Ixp33_ASAP7_75t_L g2421 ( 
.A1(n_1919),
.A2(n_1944),
.B(n_1666),
.C(n_1670),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_1768),
.B(n_1776),
.Y(n_2422)
);

AOI21xp5_ASAP7_75t_L g2423 ( 
.A1(n_1690),
.A2(n_1693),
.B(n_1696),
.Y(n_2423)
);

AOI21xp5_ASAP7_75t_L g2424 ( 
.A1(n_1690),
.A2(n_1693),
.B(n_1696),
.Y(n_2424)
);

AND2x2_ASAP7_75t_SL g2425 ( 
.A(n_1625),
.B(n_1709),
.Y(n_2425)
);

OA22x2_ASAP7_75t_L g2426 ( 
.A1(n_1909),
.A2(n_1880),
.B1(n_1886),
.B2(n_1882),
.Y(n_2426)
);

INVx4_ASAP7_75t_L g2427 ( 
.A(n_1625),
.Y(n_2427)
);

OR2x6_ASAP7_75t_L g2428 ( 
.A(n_1625),
.B(n_1709),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_SL g2429 ( 
.A(n_1933),
.B(n_1709),
.Y(n_2429)
);

AOI21xp5_ASAP7_75t_L g2430 ( 
.A1(n_1697),
.A2(n_1496),
.B(n_1416),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_1768),
.B(n_1776),
.Y(n_2431)
);

OAI21xp5_ASAP7_75t_L g2432 ( 
.A1(n_1531),
.A2(n_1697),
.B(n_1698),
.Y(n_2432)
);

AOI21xp5_ASAP7_75t_L g2433 ( 
.A1(n_1496),
.A2(n_1602),
.B(n_1416),
.Y(n_2433)
);

OAI22xp5_ASAP7_75t_L g2434 ( 
.A1(n_1495),
.A2(n_1611),
.B1(n_1699),
.B2(n_1669),
.Y(n_2434)
);

INVx4_ASAP7_75t_L g2435 ( 
.A(n_1709),
.Y(n_2435)
);

AOI21xp5_ASAP7_75t_L g2436 ( 
.A1(n_1531),
.A2(n_1602),
.B(n_1416),
.Y(n_2436)
);

AOI21xp5_ASAP7_75t_L g2437 ( 
.A1(n_1416),
.A2(n_1602),
.B(n_1918),
.Y(n_2437)
);

NAND2x1_ASAP7_75t_L g2438 ( 
.A(n_1602),
.B(n_1915),
.Y(n_2438)
);

BUFx4f_ASAP7_75t_L g2439 ( 
.A(n_1451),
.Y(n_2439)
);

BUFx6f_ASAP7_75t_L g2440 ( 
.A(n_1426),
.Y(n_2440)
);

CKINVDCx5p33_ASAP7_75t_R g2441 ( 
.A(n_1778),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_SL g2442 ( 
.A(n_1933),
.B(n_1709),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_1768),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_1776),
.Y(n_2444)
);

NOR2xp33_ASAP7_75t_L g2445 ( 
.A(n_1880),
.B(n_1882),
.Y(n_2445)
);

AOI21xp5_ASAP7_75t_L g2446 ( 
.A1(n_1918),
.A2(n_1952),
.B(n_1969),
.Y(n_2446)
);

OAI22xp5_ASAP7_75t_L g2447 ( 
.A1(n_1611),
.A2(n_1680),
.B1(n_1714),
.B2(n_1662),
.Y(n_2447)
);

AOI21xp5_ASAP7_75t_L g2448 ( 
.A1(n_1918),
.A2(n_1952),
.B(n_1405),
.Y(n_2448)
);

NOR2x1_ASAP7_75t_L g2449 ( 
.A(n_1880),
.B(n_1882),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_1784),
.B(n_1819),
.Y(n_2450)
);

BUFx8_ASAP7_75t_L g2451 ( 
.A(n_1451),
.Y(n_2451)
);

INVx3_ASAP7_75t_L g2452 ( 
.A(n_1426),
.Y(n_2452)
);

AOI21xp5_ASAP7_75t_L g2453 ( 
.A1(n_1918),
.A2(n_1952),
.B(n_1405),
.Y(n_2453)
);

OAI22x1_ASAP7_75t_L g2454 ( 
.A1(n_1945),
.A2(n_1946),
.B1(n_1900),
.B2(n_1816),
.Y(n_2454)
);

INVx4_ASAP7_75t_L g2455 ( 
.A(n_1934),
.Y(n_2455)
);

AO32x2_ASAP7_75t_L g2456 ( 
.A1(n_1972),
.A2(n_1952),
.A3(n_1456),
.B1(n_1405),
.B2(n_1517),
.Y(n_2456)
);

OAI22xp5_ASAP7_75t_L g2457 ( 
.A1(n_1662),
.A2(n_1680),
.B1(n_1669),
.B2(n_1672),
.Y(n_2457)
);

AOI21xp5_ASAP7_75t_L g2458 ( 
.A1(n_1456),
.A2(n_1910),
.B(n_1521),
.Y(n_2458)
);

OAI22xp5_ASAP7_75t_L g2459 ( 
.A1(n_1671),
.A2(n_1672),
.B1(n_1699),
.B2(n_1684),
.Y(n_2459)
);

BUFx2_ASAP7_75t_L g2460 ( 
.A(n_1870),
.Y(n_2460)
);

INVx4_ASAP7_75t_L g2461 ( 
.A(n_1451),
.Y(n_2461)
);

O2A1O1Ixp33_ASAP7_75t_L g2462 ( 
.A1(n_1612),
.A2(n_1614),
.B(n_1630),
.C(n_1613),
.Y(n_2462)
);

AOI21xp5_ASAP7_75t_L g2463 ( 
.A1(n_1456),
.A2(n_1910),
.B(n_1521),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_1784),
.Y(n_2464)
);

AOI21xp5_ASAP7_75t_L g2465 ( 
.A1(n_1521),
.A2(n_1557),
.B(n_1906),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_1784),
.Y(n_2466)
);

AOI21xp5_ASAP7_75t_L g2467 ( 
.A1(n_1557),
.A2(n_1927),
.B(n_1928),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_1819),
.B(n_1821),
.Y(n_2468)
);

AOI21xp5_ASAP7_75t_L g2469 ( 
.A1(n_1557),
.A2(n_1928),
.B(n_1929),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_SL g2470 ( 
.A(n_1870),
.B(n_1785),
.Y(n_2470)
);

AOI21xp5_ASAP7_75t_L g2471 ( 
.A1(n_1929),
.A2(n_1932),
.B(n_1915),
.Y(n_2471)
);

AND2x2_ASAP7_75t_L g2472 ( 
.A(n_1778),
.B(n_1791),
.Y(n_2472)
);

AND2x2_ASAP7_75t_L g2473 ( 
.A(n_1791),
.B(n_1524),
.Y(n_2473)
);

NOR2xp33_ASAP7_75t_L g2474 ( 
.A(n_1880),
.B(n_1882),
.Y(n_2474)
);

BUFx2_ASAP7_75t_L g2475 ( 
.A(n_1870),
.Y(n_2475)
);

BUFx6f_ASAP7_75t_L g2476 ( 
.A(n_1551),
.Y(n_2476)
);

A2O1A1Ixp33_ASAP7_75t_L g2477 ( 
.A1(n_1666),
.A2(n_1670),
.B(n_1727),
.C(n_1590),
.Y(n_2477)
);

NOR2xp33_ASAP7_75t_L g2478 ( 
.A(n_1886),
.B(n_1630),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_1819),
.B(n_1856),
.Y(n_2479)
);

AOI21xp5_ASAP7_75t_L g2480 ( 
.A1(n_1932),
.A2(n_1980),
.B(n_1915),
.Y(n_2480)
);

CKINVDCx10_ASAP7_75t_R g2481 ( 
.A(n_1596),
.Y(n_2481)
);

OR2x6_ASAP7_75t_L g2482 ( 
.A(n_1457),
.B(n_1482),
.Y(n_2482)
);

AOI21xp5_ASAP7_75t_L g2483 ( 
.A1(n_1915),
.A2(n_1980),
.B(n_1954),
.Y(n_2483)
);

OAI22xp5_ASAP7_75t_L g2484 ( 
.A1(n_1671),
.A2(n_1714),
.B1(n_1684),
.B2(n_1886),
.Y(n_2484)
);

AOI21xp5_ASAP7_75t_L g2485 ( 
.A1(n_1916),
.A2(n_1980),
.B(n_1954),
.Y(n_2485)
);

AND2x4_ASAP7_75t_L g2486 ( 
.A(n_1886),
.B(n_1785),
.Y(n_2486)
);

AO221x2_ASAP7_75t_L g2487 ( 
.A1(n_1823),
.A2(n_1605),
.B1(n_1727),
.B2(n_1698),
.C(n_1804),
.Y(n_2487)
);

NOR2xp33_ASAP7_75t_L g2488 ( 
.A(n_1614),
.B(n_1823),
.Y(n_2488)
);

AND2x2_ASAP7_75t_L g2489 ( 
.A(n_1524),
.B(n_1545),
.Y(n_2489)
);

BUFx6f_ASAP7_75t_L g2490 ( 
.A(n_1551),
.Y(n_2490)
);

OAI22xp5_ASAP7_75t_L g2491 ( 
.A1(n_1605),
.A2(n_1457),
.B1(n_1482),
.B2(n_1804),
.Y(n_2491)
);

OAI22xp5_ASAP7_75t_L g2492 ( 
.A1(n_1482),
.A2(n_1545),
.B1(n_1590),
.B2(n_1451),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_SL g2493 ( 
.A(n_1870),
.B(n_1785),
.Y(n_2493)
);

AOI21xp5_ASAP7_75t_L g2494 ( 
.A1(n_1916),
.A2(n_1980),
.B(n_1954),
.Y(n_2494)
);

AOI21xp5_ASAP7_75t_L g2495 ( 
.A1(n_1916),
.A2(n_1954),
.B(n_1551),
.Y(n_2495)
);

AND2x4_ASAP7_75t_L g2496 ( 
.A(n_1785),
.B(n_1832),
.Y(n_2496)
);

AOI21xp5_ASAP7_75t_L g2497 ( 
.A1(n_1916),
.A2(n_1551),
.B(n_1520),
.Y(n_2497)
);

INVx3_ASAP7_75t_SL g2498 ( 
.A(n_1870),
.Y(n_2498)
);

AOI21xp5_ASAP7_75t_L g2499 ( 
.A1(n_1551),
.A2(n_1520),
.B(n_1482),
.Y(n_2499)
);

A2O1A1Ixp33_ASAP7_75t_L g2500 ( 
.A1(n_1958),
.A2(n_1979),
.B(n_1973),
.C(n_1971),
.Y(n_2500)
);

NOR2x1_ASAP7_75t_L g2501 ( 
.A(n_1958),
.B(n_1870),
.Y(n_2501)
);

O2A1O1Ixp33_ASAP7_75t_L g2502 ( 
.A1(n_1805),
.A2(n_1925),
.B(n_1977),
.C(n_1924),
.Y(n_2502)
);

INVx3_ASAP7_75t_L g2503 ( 
.A(n_1551),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_1821),
.B(n_1844),
.Y(n_2504)
);

BUFx2_ASAP7_75t_R g2505 ( 
.A(n_1900),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_1821),
.B(n_1844),
.Y(n_2506)
);

BUFx2_ASAP7_75t_L g2507 ( 
.A(n_1785),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_1835),
.Y(n_2508)
);

AO32x2_ASAP7_75t_L g2509 ( 
.A1(n_1979),
.A2(n_1973),
.A3(n_1971),
.B1(n_1965),
.B2(n_1955),
.Y(n_2509)
);

AND2x2_ASAP7_75t_L g2510 ( 
.A(n_1785),
.B(n_1832),
.Y(n_2510)
);

AOI21xp5_ASAP7_75t_L g2511 ( 
.A1(n_1551),
.A2(n_1520),
.B(n_1936),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_1835),
.Y(n_2512)
);

OAI21x1_ASAP7_75t_L g2513 ( 
.A1(n_1703),
.A2(n_1694),
.B(n_1653),
.Y(n_2513)
);

NOR2xp67_ASAP7_75t_L g2514 ( 
.A(n_1936),
.B(n_1937),
.Y(n_2514)
);

AOI21xp5_ASAP7_75t_L g2515 ( 
.A1(n_1520),
.A2(n_1951),
.B(n_1938),
.Y(n_2515)
);

NOR2xp33_ASAP7_75t_L g2516 ( 
.A(n_1832),
.B(n_1900),
.Y(n_2516)
);

AOI22xp5_ASAP7_75t_L g2517 ( 
.A1(n_1451),
.A2(n_1499),
.B1(n_1832),
.B2(n_1660),
.Y(n_2517)
);

INVx1_ASAP7_75t_SL g2518 ( 
.A(n_1832),
.Y(n_2518)
);

BUFx6f_ASAP7_75t_L g2519 ( 
.A(n_1520),
.Y(n_2519)
);

AND2x2_ASAP7_75t_L g2520 ( 
.A(n_1832),
.B(n_1967),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_1835),
.B(n_1856),
.Y(n_2521)
);

NAND2x1p5_ASAP7_75t_L g2522 ( 
.A(n_1520),
.B(n_1499),
.Y(n_2522)
);

NOR2xp67_ASAP7_75t_L g2523 ( 
.A(n_1937),
.B(n_1942),
.Y(n_2523)
);

INVx2_ASAP7_75t_L g2524 ( 
.A(n_1838),
.Y(n_2524)
);

A2O1A1Ixp33_ASAP7_75t_L g2525 ( 
.A1(n_1938),
.A2(n_1965),
.B(n_1955),
.C(n_1951),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_1838),
.B(n_1967),
.Y(n_2526)
);

INVx4_ASAP7_75t_L g2527 ( 
.A(n_1499),
.Y(n_2527)
);

AOI21xp5_ASAP7_75t_L g2528 ( 
.A1(n_1942),
.A2(n_1949),
.B(n_1499),
.Y(n_2528)
);

INVx3_ASAP7_75t_L g2529 ( 
.A(n_1499),
.Y(n_2529)
);

INVxp67_ASAP7_75t_L g2530 ( 
.A(n_1838),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_1842),
.B(n_1967),
.Y(n_2531)
);

OAI22xp5_ASAP7_75t_L g2532 ( 
.A1(n_1499),
.A2(n_1805),
.B1(n_1959),
.B2(n_1842),
.Y(n_2532)
);

AOI21xp5_ASAP7_75t_L g2533 ( 
.A1(n_1949),
.A2(n_1925),
.B(n_1968),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_1842),
.B(n_1959),
.Y(n_2534)
);

OAI21x1_ASAP7_75t_L g2535 ( 
.A1(n_1924),
.A2(n_1926),
.B(n_1968),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_1844),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_1856),
.B(n_1959),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_L g2538 ( 
.A(n_1866),
.B(n_1948),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_1866),
.B(n_1948),
.Y(n_2539)
);

AOI21xp5_ASAP7_75t_L g2540 ( 
.A1(n_1977),
.A2(n_1926),
.B(n_1931),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_1866),
.Y(n_2541)
);

AOI21xp5_ASAP7_75t_L g2542 ( 
.A1(n_1931),
.A2(n_1948),
.B(n_1660),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_1660),
.B(n_1805),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_SL g2544 ( 
.A(n_1660),
.B(n_1420),
.Y(n_2544)
);

O2A1O1Ixp33_ASAP7_75t_L g2545 ( 
.A1(n_1660),
.A2(n_1788),
.B(n_1995),
.C(n_1989),
.Y(n_2545)
);

OAI21xp5_ASAP7_75t_L g2546 ( 
.A1(n_1660),
.A2(n_1054),
.B(n_1989),
.Y(n_2546)
);

OAI22xp5_ASAP7_75t_L g2547 ( 
.A1(n_1660),
.A2(n_660),
.B1(n_680),
.B2(n_669),
.Y(n_2547)
);

OAI22xp5_ASAP7_75t_L g2548 ( 
.A1(n_1989),
.A2(n_660),
.B1(n_680),
.B2(n_669),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_1404),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_1404),
.Y(n_2550)
);

OR2x2_ASAP7_75t_L g2551 ( 
.A(n_1783),
.B(n_1771),
.Y(n_2551)
);

A2O1A1Ixp33_ASAP7_75t_L g2552 ( 
.A1(n_1788),
.A2(n_660),
.B(n_680),
.C(n_669),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_SL g2553 ( 
.A(n_1420),
.B(n_1437),
.Y(n_2553)
);

AOI22xp33_ASAP7_75t_L g2554 ( 
.A1(n_1987),
.A2(n_679),
.B1(n_1788),
.B2(n_675),
.Y(n_2554)
);

AOI21xp5_ASAP7_75t_L g2555 ( 
.A1(n_1579),
.A2(n_1455),
.B(n_1412),
.Y(n_2555)
);

AOI21xp5_ASAP7_75t_L g2556 ( 
.A1(n_1579),
.A2(n_1455),
.B(n_1412),
.Y(n_2556)
);

O2A1O1Ixp33_ASAP7_75t_L g2557 ( 
.A1(n_1788),
.A2(n_1989),
.B(n_1995),
.C(n_1054),
.Y(n_2557)
);

AOI21xp5_ASAP7_75t_L g2558 ( 
.A1(n_1579),
.A2(n_1455),
.B(n_1412),
.Y(n_2558)
);

AOI22xp5_ASAP7_75t_L g2559 ( 
.A1(n_1788),
.A2(n_660),
.B1(n_680),
.B2(n_669),
.Y(n_2559)
);

O2A1O1Ixp33_ASAP7_75t_L g2560 ( 
.A1(n_1788),
.A2(n_1989),
.B(n_1995),
.C(n_1054),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_1990),
.B(n_1783),
.Y(n_2561)
);

OAI22xp5_ASAP7_75t_L g2562 ( 
.A1(n_1989),
.A2(n_660),
.B1(n_680),
.B2(n_669),
.Y(n_2562)
);

HB1xp67_ASAP7_75t_L g2563 ( 
.A(n_1513),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_1404),
.Y(n_2564)
);

NAND2x1p5_ASAP7_75t_L g2565 ( 
.A(n_1415),
.B(n_1435),
.Y(n_2565)
);

AOI21xp5_ASAP7_75t_L g2566 ( 
.A1(n_1579),
.A2(n_1455),
.B(n_1412),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_1990),
.B(n_1783),
.Y(n_2567)
);

INVx3_ASAP7_75t_L g2568 ( 
.A(n_1655),
.Y(n_2568)
);

AOI22x1_ASAP7_75t_L g2569 ( 
.A1(n_1445),
.A2(n_1782),
.B1(n_1792),
.B2(n_1986),
.Y(n_2569)
);

INVxp67_ASAP7_75t_L g2570 ( 
.A(n_1513),
.Y(n_2570)
);

BUFx12f_ASAP7_75t_L g2571 ( 
.A(n_1519),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_SL g2572 ( 
.A(n_1420),
.B(n_1437),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_L g2573 ( 
.A(n_1990),
.B(n_1783),
.Y(n_2573)
);

OAI22xp5_ASAP7_75t_L g2574 ( 
.A1(n_1989),
.A2(n_660),
.B1(n_680),
.B2(n_669),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_SL g2575 ( 
.A(n_1420),
.B(n_1437),
.Y(n_2575)
);

BUFx2_ASAP7_75t_L g2576 ( 
.A(n_1771),
.Y(n_2576)
);

OAI22xp5_ASAP7_75t_L g2577 ( 
.A1(n_1989),
.A2(n_660),
.B1(n_680),
.B2(n_669),
.Y(n_2577)
);

O2A1O1Ixp33_ASAP7_75t_L g2578 ( 
.A1(n_1788),
.A2(n_1989),
.B(n_1995),
.C(n_1054),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_L g2579 ( 
.A(n_1990),
.B(n_1783),
.Y(n_2579)
);

OAI22xp5_ASAP7_75t_L g2580 ( 
.A1(n_1989),
.A2(n_660),
.B1(n_680),
.B2(n_669),
.Y(n_2580)
);

NAND3xp33_ASAP7_75t_L g2581 ( 
.A(n_1989),
.B(n_1054),
.C(n_1995),
.Y(n_2581)
);

AOI33xp33_ASAP7_75t_L g2582 ( 
.A1(n_1527),
.A2(n_188),
.A3(n_203),
.B1(n_156),
.B2(n_1114),
.B3(n_1525),
.Y(n_2582)
);

OAI21xp5_ASAP7_75t_L g2583 ( 
.A1(n_1989),
.A2(n_1054),
.B(n_1995),
.Y(n_2583)
);

INVx2_ASAP7_75t_SL g2584 ( 
.A(n_1875),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_1407),
.Y(n_2585)
);

AOI21xp5_ASAP7_75t_L g2586 ( 
.A1(n_1579),
.A2(n_1455),
.B(n_1412),
.Y(n_2586)
);

AO22x1_ASAP7_75t_L g2587 ( 
.A1(n_1514),
.A2(n_1474),
.B1(n_1421),
.B2(n_1591),
.Y(n_2587)
);

AOI22xp5_ASAP7_75t_L g2588 ( 
.A1(n_1788),
.A2(n_660),
.B1(n_680),
.B2(n_669),
.Y(n_2588)
);

AND2x4_ASAP7_75t_L g2589 ( 
.A(n_2310),
.B(n_2085),
.Y(n_2589)
);

AOI21x1_ASAP7_75t_L g2590 ( 
.A1(n_2058),
.A2(n_2210),
.B(n_2035),
.Y(n_2590)
);

NAND3xp33_ASAP7_75t_L g2591 ( 
.A(n_2013),
.B(n_2082),
.C(n_2002),
.Y(n_2591)
);

INVx4_ASAP7_75t_L g2592 ( 
.A(n_2319),
.Y(n_2592)
);

AO31x2_ASAP7_75t_L g2593 ( 
.A1(n_2026),
.A2(n_2074),
.A3(n_2300),
.B(n_2069),
.Y(n_2593)
);

INVx2_ASAP7_75t_SL g2594 ( 
.A(n_2121),
.Y(n_2594)
);

OAI21x1_ASAP7_75t_L g2595 ( 
.A1(n_2098),
.A2(n_2115),
.B(n_2117),
.Y(n_2595)
);

OAI21x1_ASAP7_75t_L g2596 ( 
.A1(n_2115),
.A2(n_2117),
.B(n_2127),
.Y(n_2596)
);

OAI21x1_ASAP7_75t_L g2597 ( 
.A1(n_2127),
.A2(n_2060),
.B(n_2136),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_SL g2598 ( 
.A(n_2003),
.B(n_2553),
.Y(n_2598)
);

AOI21xp5_ASAP7_75t_L g2599 ( 
.A1(n_1998),
.A2(n_2556),
.B(n_2555),
.Y(n_2599)
);

OAI21x1_ASAP7_75t_L g2600 ( 
.A1(n_2136),
.A2(n_2114),
.B(n_2141),
.Y(n_2600)
);

NAND3x1_ASAP7_75t_L g2601 ( 
.A(n_2583),
.B(n_2001),
.C(n_2559),
.Y(n_2601)
);

AOI21xp5_ASAP7_75t_L g2602 ( 
.A1(n_2586),
.A2(n_2555),
.B(n_1998),
.Y(n_2602)
);

INVx3_ASAP7_75t_L g2603 ( 
.A(n_2161),
.Y(n_2603)
);

INVx1_ASAP7_75t_SL g2604 ( 
.A(n_2096),
.Y(n_2604)
);

OAI21xp5_ASAP7_75t_L g2605 ( 
.A1(n_2014),
.A2(n_2562),
.B(n_2548),
.Y(n_2605)
);

OAI22xp5_ASAP7_75t_L g2606 ( 
.A1(n_2559),
.A2(n_2588),
.B1(n_2562),
.B2(n_2574),
.Y(n_2606)
);

OAI22x1_ASAP7_75t_L g2607 ( 
.A1(n_2588),
.A2(n_2001),
.B1(n_2033),
.B2(n_2015),
.Y(n_2607)
);

AO21x1_ASAP7_75t_L g2608 ( 
.A1(n_2548),
.A2(n_2577),
.B(n_2574),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2040),
.B(n_2043),
.Y(n_2609)
);

AOI21xp5_ASAP7_75t_L g2610 ( 
.A1(n_2586),
.A2(n_2558),
.B(n_2556),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2321),
.Y(n_2611)
);

OAI21xp5_ASAP7_75t_L g2612 ( 
.A1(n_2577),
.A2(n_2580),
.B(n_2552),
.Y(n_2612)
);

AOI21xp5_ASAP7_75t_L g2613 ( 
.A1(n_2558),
.A2(n_2566),
.B(n_2000),
.Y(n_2613)
);

AO31x2_ASAP7_75t_L g2614 ( 
.A1(n_2026),
.A2(n_2300),
.A3(n_2226),
.B(n_2204),
.Y(n_2614)
);

AO31x2_ASAP7_75t_L g2615 ( 
.A1(n_2204),
.A2(n_2090),
.A3(n_2068),
.B(n_2170),
.Y(n_2615)
);

AO31x2_ASAP7_75t_L g2616 ( 
.A1(n_2084),
.A2(n_2089),
.A3(n_2184),
.B(n_2525),
.Y(n_2616)
);

NAND3x1_ASAP7_75t_L g2617 ( 
.A(n_2583),
.B(n_2033),
.C(n_2015),
.Y(n_2617)
);

INVxp67_ASAP7_75t_L g2618 ( 
.A(n_2021),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2321),
.Y(n_2619)
);

AOI21x1_ASAP7_75t_L g2620 ( 
.A1(n_2058),
.A2(n_2210),
.B(n_2035),
.Y(n_2620)
);

NAND2x1p5_ASAP7_75t_L g2621 ( 
.A(n_2319),
.B(n_2121),
.Y(n_2621)
);

NOR2x1_ASAP7_75t_SL g2622 ( 
.A(n_2009),
.B(n_2121),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2040),
.B(n_2043),
.Y(n_2623)
);

OAI21x1_ASAP7_75t_L g2624 ( 
.A1(n_2114),
.A2(n_1997),
.B(n_2277),
.Y(n_2624)
);

NAND3xp33_ASAP7_75t_L g2625 ( 
.A(n_2581),
.B(n_2130),
.C(n_2557),
.Y(n_2625)
);

AOI21xp5_ASAP7_75t_L g2626 ( 
.A1(n_2566),
.A2(n_2000),
.B(n_2048),
.Y(n_2626)
);

AOI221x1_ASAP7_75t_L g2627 ( 
.A1(n_2580),
.A2(n_2072),
.B1(n_2086),
.B2(n_2158),
.C(n_2133),
.Y(n_2627)
);

AND2x2_ASAP7_75t_L g2628 ( 
.A(n_1999),
.B(n_2083),
.Y(n_2628)
);

AOI21xp5_ASAP7_75t_L g2629 ( 
.A1(n_2547),
.A2(n_2030),
.B(n_2172),
.Y(n_2629)
);

BUFx6f_ASAP7_75t_L g2630 ( 
.A(n_2078),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_L g2631 ( 
.A(n_2016),
.B(n_2561),
.Y(n_2631)
);

INVx3_ASAP7_75t_L g2632 ( 
.A(n_2161),
.Y(n_2632)
);

BUFx6f_ASAP7_75t_L g2633 ( 
.A(n_2078),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2016),
.B(n_2561),
.Y(n_2634)
);

OAI21x1_ASAP7_75t_SL g2635 ( 
.A1(n_2547),
.A2(n_2578),
.B(n_2560),
.Y(n_2635)
);

OAI21x1_ASAP7_75t_L g2636 ( 
.A1(n_1997),
.A2(n_2291),
.B(n_2277),
.Y(n_2636)
);

BUFx2_ASAP7_75t_L g2637 ( 
.A(n_2009),
.Y(n_2637)
);

OAI21x1_ASAP7_75t_L g2638 ( 
.A1(n_2291),
.A2(n_2295),
.B(n_2190),
.Y(n_2638)
);

NAND2xp33_ASAP7_75t_L g2639 ( 
.A(n_2211),
.B(n_2288),
.Y(n_2639)
);

OAI21x1_ASAP7_75t_L g2640 ( 
.A1(n_2295),
.A2(n_2193),
.B(n_2181),
.Y(n_2640)
);

NOR2xp33_ASAP7_75t_L g2641 ( 
.A(n_2087),
.B(n_2572),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_L g2642 ( 
.A(n_2567),
.B(n_2573),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_2007),
.Y(n_2643)
);

OAI21x1_ASAP7_75t_L g2644 ( 
.A1(n_2194),
.A2(n_2207),
.B(n_2201),
.Y(n_2644)
);

AOI21xp5_ASAP7_75t_L g2645 ( 
.A1(n_2237),
.A2(n_2234),
.B(n_2054),
.Y(n_2645)
);

OAI21xp5_ASAP7_75t_L g2646 ( 
.A1(n_2236),
.A2(n_2189),
.B(n_2581),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2044),
.Y(n_2647)
);

INVx1_ASAP7_75t_SL g2648 ( 
.A(n_2096),
.Y(n_2648)
);

AOI21xp5_ASAP7_75t_L g2649 ( 
.A1(n_2180),
.A2(n_2230),
.B(n_2239),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_2567),
.B(n_2573),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_L g2651 ( 
.A(n_2579),
.B(n_2192),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_L g2652 ( 
.A(n_2579),
.B(n_2192),
.Y(n_2652)
);

AND2x2_ASAP7_75t_L g2653 ( 
.A(n_1999),
.B(n_2083),
.Y(n_2653)
);

OAI21xp5_ASAP7_75t_L g2654 ( 
.A1(n_2236),
.A2(n_2575),
.B(n_2113),
.Y(n_2654)
);

AOI21x1_ASAP7_75t_L g2655 ( 
.A1(n_2314),
.A2(n_2362),
.B(n_2395),
.Y(n_2655)
);

A2O1A1Ixp33_ASAP7_75t_L g2656 ( 
.A1(n_2053),
.A2(n_2545),
.B(n_2582),
.C(n_2072),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_L g2657 ( 
.A(n_2197),
.B(n_2065),
.Y(n_2657)
);

OAI21x1_ASAP7_75t_L g2658 ( 
.A1(n_2209),
.A2(n_2225),
.B(n_2221),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2197),
.B(n_2065),
.Y(n_2659)
);

OAI21x1_ASAP7_75t_L g2660 ( 
.A1(n_2306),
.A2(n_2252),
.B(n_2271),
.Y(n_2660)
);

AOI221xp5_ASAP7_75t_L g2661 ( 
.A1(n_2039),
.A2(n_2047),
.B1(n_2554),
.B2(n_2051),
.C(n_2064),
.Y(n_2661)
);

OAI21xp5_ASAP7_75t_L g2662 ( 
.A1(n_2034),
.A2(n_2076),
.B(n_2051),
.Y(n_2662)
);

BUFx6f_ASAP7_75t_L g2663 ( 
.A(n_2078),
.Y(n_2663)
);

AND2x2_ASAP7_75t_L g2664 ( 
.A(n_2093),
.B(n_2126),
.Y(n_2664)
);

NAND2x2_ASAP7_75t_L g2665 ( 
.A(n_2169),
.B(n_2247),
.Y(n_2665)
);

AOI21xp5_ASAP7_75t_L g2666 ( 
.A1(n_2316),
.A2(n_2343),
.B(n_2319),
.Y(n_2666)
);

AOI21xp5_ASAP7_75t_L g2667 ( 
.A1(n_2319),
.A2(n_2076),
.B(n_2108),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_2066),
.B(n_2182),
.Y(n_2668)
);

OAI21x1_ASAP7_75t_L g2669 ( 
.A1(n_2306),
.A2(n_2275),
.B(n_2271),
.Y(n_2669)
);

AO21x1_ASAP7_75t_L g2670 ( 
.A1(n_2039),
.A2(n_2047),
.B(n_2028),
.Y(n_2670)
);

BUFx3_ASAP7_75t_L g2671 ( 
.A(n_2206),
.Y(n_2671)
);

OAI21x1_ASAP7_75t_SL g2672 ( 
.A1(n_2162),
.A2(n_2034),
.B(n_2546),
.Y(n_2672)
);

OAI21x1_ASAP7_75t_L g2673 ( 
.A1(n_2275),
.A2(n_2227),
.B(n_2297),
.Y(n_2673)
);

NOR2xp33_ASAP7_75t_L g2674 ( 
.A(n_2019),
.B(n_2006),
.Y(n_2674)
);

A2O1A1Ixp33_ASAP7_75t_L g2675 ( 
.A1(n_2022),
.A2(n_2304),
.B(n_2028),
.C(n_2253),
.Y(n_2675)
);

AOI21xp5_ASAP7_75t_L g2676 ( 
.A1(n_2108),
.A2(n_2152),
.B(n_2269),
.Y(n_2676)
);

OAI21x1_ASAP7_75t_L g2677 ( 
.A1(n_2297),
.A2(n_2471),
.B(n_2385),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2007),
.Y(n_2678)
);

OAI21x1_ASAP7_75t_L g2679 ( 
.A1(n_2354),
.A2(n_2388),
.B(n_2405),
.Y(n_2679)
);

INVx5_ASAP7_75t_L g2680 ( 
.A(n_2009),
.Y(n_2680)
);

OAI21x1_ASAP7_75t_L g2681 ( 
.A1(n_2423),
.A2(n_2424),
.B(n_2242),
.Y(n_2681)
);

AND2x2_ASAP7_75t_L g2682 ( 
.A(n_2093),
.B(n_2126),
.Y(n_2682)
);

OAI21xp5_ASAP7_75t_L g2683 ( 
.A1(n_2011),
.A2(n_2171),
.B(n_2022),
.Y(n_2683)
);

OR2x2_ASAP7_75t_L g2684 ( 
.A(n_2551),
.B(n_2008),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2066),
.B(n_2182),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2044),
.Y(n_2686)
);

AOI22xp5_ASAP7_75t_L g2687 ( 
.A1(n_2042),
.A2(n_2111),
.B1(n_2036),
.B2(n_2332),
.Y(n_2687)
);

AOI21xp5_ASAP7_75t_L g2688 ( 
.A1(n_2108),
.A2(n_2342),
.B(n_2017),
.Y(n_2688)
);

OAI21xp5_ASAP7_75t_L g2689 ( 
.A1(n_2171),
.A2(n_2032),
.B(n_2187),
.Y(n_2689)
);

INVx3_ASAP7_75t_L g2690 ( 
.A(n_2161),
.Y(n_2690)
);

OAI21x1_ASAP7_75t_SL g2691 ( 
.A1(n_2546),
.A2(n_2004),
.B(n_2005),
.Y(n_2691)
);

AO22x2_ASAP7_75t_L g2692 ( 
.A1(n_2008),
.A2(n_2585),
.B1(n_2024),
.B2(n_2042),
.Y(n_2692)
);

OR2x2_ASAP7_75t_L g2693 ( 
.A(n_2551),
.B(n_2024),
.Y(n_2693)
);

BUFx3_ASAP7_75t_L g2694 ( 
.A(n_2206),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_L g2695 ( 
.A(n_2186),
.B(n_2031),
.Y(n_2695)
);

OAI21x1_ASAP7_75t_L g2696 ( 
.A1(n_2242),
.A2(n_2322),
.B(n_2274),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2186),
.B(n_2031),
.Y(n_2697)
);

OAI21x1_ASAP7_75t_L g2698 ( 
.A1(n_2322),
.A2(n_2274),
.B(n_2273),
.Y(n_2698)
);

INVx4_ASAP7_75t_L g2699 ( 
.A(n_2121),
.Y(n_2699)
);

AOI21xp33_ASAP7_75t_L g2700 ( 
.A1(n_2569),
.A2(n_2167),
.B(n_2187),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_2045),
.B(n_2049),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_SL g2702 ( 
.A(n_2105),
.B(n_2081),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_L g2703 ( 
.A(n_2045),
.B(n_2049),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2203),
.B(n_2212),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2203),
.B(n_2212),
.Y(n_2705)
);

OAI21x1_ASAP7_75t_SL g2706 ( 
.A1(n_2004),
.A2(n_2005),
.B(n_2188),
.Y(n_2706)
);

BUFx10_ASAP7_75t_L g2707 ( 
.A(n_2140),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2092),
.B(n_2099),
.Y(n_2708)
);

INVx2_ASAP7_75t_SL g2709 ( 
.A(n_2121),
.Y(n_2709)
);

O2A1O1Ixp33_ASAP7_75t_L g2710 ( 
.A1(n_2188),
.A2(n_2191),
.B(n_2196),
.C(n_2032),
.Y(n_2710)
);

OAI21x1_ASAP7_75t_L g2711 ( 
.A1(n_2273),
.A2(n_2356),
.B(n_2284),
.Y(n_2711)
);

OAI21x1_ASAP7_75t_L g2712 ( 
.A1(n_2284),
.A2(n_2356),
.B(n_2362),
.Y(n_2712)
);

NAND2xp33_ASAP7_75t_L g2713 ( 
.A(n_2302),
.B(n_2371),
.Y(n_2713)
);

OAI21x1_ASAP7_75t_L g2714 ( 
.A1(n_2528),
.A2(n_2344),
.B(n_2515),
.Y(n_2714)
);

INVxp67_ASAP7_75t_L g2715 ( 
.A(n_2112),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2071),
.Y(n_2716)
);

AO31x2_ASAP7_75t_L g2717 ( 
.A1(n_2500),
.A2(n_2278),
.A3(n_2346),
.B(n_2484),
.Y(n_2717)
);

OAI21x1_ASAP7_75t_L g2718 ( 
.A1(n_2314),
.A2(n_2360),
.B(n_2337),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2071),
.Y(n_2719)
);

BUFx2_ASAP7_75t_L g2720 ( 
.A(n_2009),
.Y(n_2720)
);

NAND2x1_ASAP7_75t_L g2721 ( 
.A(n_2009),
.B(n_2161),
.Y(n_2721)
);

INVx3_ASAP7_75t_L g2722 ( 
.A(n_2085),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_L g2723 ( 
.A(n_2092),
.B(n_2099),
.Y(n_2723)
);

NOR2xp33_ASAP7_75t_L g2724 ( 
.A(n_2020),
.B(n_2018),
.Y(n_2724)
);

A2O1A1Ixp33_ASAP7_75t_L g2725 ( 
.A1(n_2392),
.A2(n_2195),
.B(n_2095),
.C(n_2324),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2102),
.B(n_2106),
.Y(n_2726)
);

OAI21x1_ASAP7_75t_L g2727 ( 
.A1(n_2569),
.A2(n_2469),
.B(n_2467),
.Y(n_2727)
);

NOR2xp33_ASAP7_75t_L g2728 ( 
.A(n_2571),
.B(n_2177),
.Y(n_2728)
);

INVxp67_ASAP7_75t_SL g2729 ( 
.A(n_2335),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_L g2730 ( 
.A(n_2102),
.B(n_2106),
.Y(n_2730)
);

AOI221x1_ASAP7_75t_L g2731 ( 
.A1(n_2191),
.A2(n_2208),
.B1(n_2398),
.B2(n_2217),
.C(n_2167),
.Y(n_2731)
);

BUFx2_ASAP7_75t_L g2732 ( 
.A(n_2389),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2128),
.B(n_2131),
.Y(n_2733)
);

A2O1A1Ixp33_ASAP7_75t_L g2734 ( 
.A1(n_2220),
.A2(n_2064),
.B(n_2199),
.C(n_2250),
.Y(n_2734)
);

OAI21x1_ASAP7_75t_L g2735 ( 
.A1(n_2352),
.A2(n_2480),
.B(n_2430),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2128),
.B(n_2131),
.Y(n_2736)
);

OAI22x1_ASAP7_75t_L g2737 ( 
.A1(n_2585),
.A2(n_2317),
.B1(n_2164),
.B2(n_2339),
.Y(n_2737)
);

OAI21x1_ASAP7_75t_L g2738 ( 
.A1(n_2511),
.A2(n_2436),
.B(n_2542),
.Y(n_2738)
);

OAI21xp5_ASAP7_75t_L g2739 ( 
.A1(n_2307),
.A2(n_2400),
.B(n_2296),
.Y(n_2739)
);

AOI21xp5_ASAP7_75t_L g2740 ( 
.A1(n_2108),
.A2(n_2368),
.B(n_2341),
.Y(n_2740)
);

AND2x2_ASAP7_75t_L g2741 ( 
.A(n_2143),
.B(n_2144),
.Y(n_2741)
);

BUFx2_ASAP7_75t_L g2742 ( 
.A(n_2389),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2135),
.B(n_2138),
.Y(n_2743)
);

BUFx8_ASAP7_75t_L g2744 ( 
.A(n_2312),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2135),
.B(n_2138),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2155),
.B(n_2159),
.Y(n_2746)
);

AO21x1_ASAP7_75t_L g2747 ( 
.A1(n_2199),
.A2(n_2059),
.B(n_2202),
.Y(n_2747)
);

OAI21xp5_ASAP7_75t_L g2748 ( 
.A1(n_2400),
.A2(n_2266),
.B(n_2293),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2155),
.B(n_2159),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2165),
.B(n_2166),
.Y(n_2750)
);

OAI22x1_ASAP7_75t_L g2751 ( 
.A1(n_2317),
.A2(n_2339),
.B1(n_2063),
.B2(n_2108),
.Y(n_2751)
);

AO22x1_ASAP7_75t_L g2752 ( 
.A1(n_2121),
.A2(n_2390),
.B1(n_2488),
.B2(n_2259),
.Y(n_2752)
);

AOI21xp5_ASAP7_75t_L g2753 ( 
.A1(n_2108),
.A2(n_2433),
.B(n_2465),
.Y(n_2753)
);

AO31x2_ASAP7_75t_L g2754 ( 
.A1(n_2346),
.A2(n_2484),
.A3(n_2491),
.B(n_2285),
.Y(n_2754)
);

OAI21x1_ASAP7_75t_L g2755 ( 
.A1(n_2436),
.A2(n_2542),
.B(n_2533),
.Y(n_2755)
);

OR2x2_ASAP7_75t_L g2756 ( 
.A(n_2309),
.B(n_2057),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2165),
.B(n_2166),
.Y(n_2757)
);

OA21x2_ASAP7_75t_L g2758 ( 
.A1(n_2129),
.A2(n_2217),
.B(n_2432),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2091),
.Y(n_2759)
);

AOI21xp5_ASAP7_75t_L g2760 ( 
.A1(n_2458),
.A2(n_2463),
.B(n_2267),
.Y(n_2760)
);

BUFx2_ASAP7_75t_L g2761 ( 
.A(n_2460),
.Y(n_2761)
);

BUFx3_ASAP7_75t_L g2762 ( 
.A(n_2029),
.Y(n_2762)
);

BUFx2_ASAP7_75t_L g2763 ( 
.A(n_2460),
.Y(n_2763)
);

AOI21xp5_ASAP7_75t_L g2764 ( 
.A1(n_2260),
.A2(n_2340),
.B(n_2330),
.Y(n_2764)
);

OAI21x1_ASAP7_75t_L g2765 ( 
.A1(n_2446),
.A2(n_2453),
.B(n_2448),
.Y(n_2765)
);

AOI21xp5_ASAP7_75t_L g2766 ( 
.A1(n_2276),
.A2(n_2023),
.B(n_2587),
.Y(n_2766)
);

OAI21x1_ASAP7_75t_L g2767 ( 
.A1(n_2513),
.A2(n_2395),
.B(n_2432),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_2168),
.B(n_2173),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2168),
.B(n_2173),
.Y(n_2769)
);

OAI21x1_ASAP7_75t_L g2770 ( 
.A1(n_2513),
.A2(n_2437),
.B(n_2499),
.Y(n_2770)
);

OAI21x1_ASAP7_75t_SL g2771 ( 
.A1(n_2214),
.A2(n_2255),
.B(n_2023),
.Y(n_2771)
);

OAI21x1_ASAP7_75t_L g2772 ( 
.A1(n_2129),
.A2(n_2495),
.B(n_2497),
.Y(n_2772)
);

INVx3_ASAP7_75t_L g2773 ( 
.A(n_2085),
.Y(n_2773)
);

OAI21x1_ASAP7_75t_L g2774 ( 
.A1(n_2535),
.A2(n_2485),
.B(n_2483),
.Y(n_2774)
);

INVxp67_ASAP7_75t_SL g2775 ( 
.A(n_2335),
.Y(n_2775)
);

BUFx2_ASAP7_75t_L g2776 ( 
.A(n_2475),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2056),
.B(n_2062),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_L g2778 ( 
.A(n_2056),
.B(n_2062),
.Y(n_2778)
);

OAI21xp33_ASAP7_75t_SL g2779 ( 
.A1(n_2097),
.A2(n_2426),
.B(n_2357),
.Y(n_2779)
);

OAI21x1_ASAP7_75t_L g2780 ( 
.A1(n_2535),
.A2(n_2494),
.B(n_2540),
.Y(n_2780)
);

AOI21x1_ASAP7_75t_L g2781 ( 
.A1(n_2587),
.A2(n_2523),
.B(n_2514),
.Y(n_2781)
);

AOI211x1_ASAP7_75t_L g2782 ( 
.A1(n_2202),
.A2(n_2219),
.B(n_2338),
.C(n_2251),
.Y(n_2782)
);

O2A1O1Ixp5_ASAP7_75t_L g2783 ( 
.A1(n_2544),
.A2(n_2235),
.B(n_2050),
.C(n_2491),
.Y(n_2783)
);

OAI21x1_ASAP7_75t_L g2784 ( 
.A1(n_2540),
.A2(n_2364),
.B(n_2438),
.Y(n_2784)
);

CKINVDCx11_ASAP7_75t_R g2785 ( 
.A(n_2571),
.Y(n_2785)
);

AOI21xp33_ASAP7_75t_L g2786 ( 
.A1(n_2293),
.A2(n_2055),
.B(n_2235),
.Y(n_2786)
);

OAI21xp5_ASAP7_75t_L g2787 ( 
.A1(n_2421),
.A2(n_2402),
.B(n_2477),
.Y(n_2787)
);

OAI21x1_ASAP7_75t_L g2788 ( 
.A1(n_2438),
.A2(n_2325),
.B(n_2318),
.Y(n_2788)
);

BUFx5_ASAP7_75t_L g2789 ( 
.A(n_2425),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2070),
.B(n_2075),
.Y(n_2790)
);

INVx3_ASAP7_75t_L g2791 ( 
.A(n_2085),
.Y(n_2791)
);

BUFx2_ASAP7_75t_L g2792 ( 
.A(n_2475),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2070),
.B(n_2075),
.Y(n_2793)
);

AND2x2_ASAP7_75t_L g2794 ( 
.A(n_2143),
.B(n_2144),
.Y(n_2794)
);

OR2x6_ASAP7_75t_L g2795 ( 
.A(n_2050),
.B(n_2134),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2077),
.B(n_2080),
.Y(n_2796)
);

AOI21xp5_ASAP7_75t_L g2797 ( 
.A1(n_2470),
.A2(n_2493),
.B(n_2027),
.Y(n_2797)
);

OAI21x1_ASAP7_75t_L g2798 ( 
.A1(n_2514),
.A2(n_2523),
.B(n_2522),
.Y(n_2798)
);

OR2x2_ASAP7_75t_L g2799 ( 
.A(n_2309),
.B(n_2057),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_L g2800 ( 
.A(n_2077),
.B(n_2080),
.Y(n_2800)
);

AOI21xp5_ASAP7_75t_L g2801 ( 
.A1(n_2027),
.A2(n_2214),
.B(n_2419),
.Y(n_2801)
);

A2O1A1Ixp33_ASAP7_75t_L g2802 ( 
.A1(n_2163),
.A2(n_2334),
.B(n_2176),
.C(n_2416),
.Y(n_2802)
);

AO31x2_ASAP7_75t_L g2803 ( 
.A1(n_2285),
.A2(n_2328),
.A3(n_2251),
.B(n_2244),
.Y(n_2803)
);

AOI21x1_ASAP7_75t_L g2804 ( 
.A1(n_2280),
.A2(n_2134),
.B(n_2420),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2153),
.B(n_2185),
.Y(n_2805)
);

OAI22xp5_ASAP7_75t_L g2806 ( 
.A1(n_2176),
.A2(n_2380),
.B1(n_2570),
.B2(n_2563),
.Y(n_2806)
);

AOI21xp5_ASAP7_75t_L g2807 ( 
.A1(n_2419),
.A2(n_2041),
.B(n_2121),
.Y(n_2807)
);

INVx3_ASAP7_75t_SL g2808 ( 
.A(n_2441),
.Y(n_2808)
);

AOI211x1_ASAP7_75t_L g2809 ( 
.A1(n_2219),
.A2(n_2338),
.B(n_2244),
.C(n_2224),
.Y(n_2809)
);

OAI22xp5_ASAP7_75t_L g2810 ( 
.A1(n_2418),
.A2(n_2183),
.B1(n_2327),
.B2(n_2052),
.Y(n_2810)
);

AND2x2_ASAP7_75t_L g2811 ( 
.A(n_2153),
.B(n_2185),
.Y(n_2811)
);

AND2x2_ASAP7_75t_L g2812 ( 
.A(n_2240),
.B(n_2091),
.Y(n_2812)
);

OAI21x1_ASAP7_75t_L g2813 ( 
.A1(n_2522),
.A2(n_2502),
.B(n_2046),
.Y(n_2813)
);

OAI22xp5_ASAP7_75t_L g2814 ( 
.A1(n_2418),
.A2(n_2327),
.B1(n_2347),
.B2(n_2104),
.Y(n_2814)
);

OAI21xp5_ASAP7_75t_L g2815 ( 
.A1(n_2402),
.A2(n_2386),
.B(n_2358),
.Y(n_2815)
);

AOI21xp5_ASAP7_75t_SL g2816 ( 
.A1(n_2361),
.A2(n_2565),
.B(n_2025),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_L g2817 ( 
.A(n_2348),
.B(n_2270),
.Y(n_2817)
);

INVx2_ASAP7_75t_L g2818 ( 
.A(n_2038),
.Y(n_2818)
);

OAI22xp5_ASAP7_75t_L g2819 ( 
.A1(n_2347),
.A2(n_2104),
.B1(n_2417),
.B2(n_2386),
.Y(n_2819)
);

OAI21x1_ASAP7_75t_L g2820 ( 
.A1(n_2522),
.A2(n_2568),
.B(n_2046),
.Y(n_2820)
);

OAI21x1_ASAP7_75t_SL g2821 ( 
.A1(n_2462),
.A2(n_2224),
.B(n_2222),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2125),
.Y(n_2822)
);

OAI21x1_ASAP7_75t_L g2823 ( 
.A1(n_2046),
.A2(n_2568),
.B(n_2264),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2348),
.B(n_2331),
.Y(n_2824)
);

A2O1A1Ixp33_ASAP7_75t_L g2825 ( 
.A1(n_2163),
.A2(n_2041),
.B(n_2120),
.C(n_2286),
.Y(n_2825)
);

AOI21xp5_ASAP7_75t_L g2826 ( 
.A1(n_2419),
.A2(n_2055),
.B(n_2447),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_L g2827 ( 
.A(n_2331),
.B(n_2079),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2125),
.Y(n_2828)
);

NOR2xp67_ASAP7_75t_L g2829 ( 
.A(n_2151),
.B(n_2420),
.Y(n_2829)
);

OA21x2_ASAP7_75t_L g2830 ( 
.A1(n_2289),
.A2(n_2397),
.B(n_2410),
.Y(n_2830)
);

OAI21xp33_ASAP7_75t_L g2831 ( 
.A1(n_2289),
.A2(n_2238),
.B(n_2222),
.Y(n_2831)
);

HB1xp67_ASAP7_75t_L g2832 ( 
.A(n_2079),
.Y(n_2832)
);

INVx2_ASAP7_75t_L g2833 ( 
.A(n_2038),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2148),
.Y(n_2834)
);

OAI21x1_ASAP7_75t_L g2835 ( 
.A1(n_2046),
.A2(n_2568),
.B(n_2264),
.Y(n_2835)
);

NOR2x1_ASAP7_75t_L g2836 ( 
.A(n_2390),
.B(n_2029),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_L g2837 ( 
.A(n_2576),
.B(n_2265),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2148),
.Y(n_2838)
);

BUFx2_ASAP7_75t_L g2839 ( 
.A(n_2576),
.Y(n_2839)
);

OAI21x1_ASAP7_75t_SL g2840 ( 
.A1(n_2238),
.A2(n_2249),
.B(n_2241),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_2240),
.B(n_2150),
.Y(n_2841)
);

OR2x2_ASAP7_75t_L g2842 ( 
.A(n_2122),
.B(n_2328),
.Y(n_2842)
);

AOI21xp5_ASAP7_75t_L g2843 ( 
.A1(n_2419),
.A2(n_2055),
.B(n_2447),
.Y(n_2843)
);

NOR2x1_ASAP7_75t_L g2844 ( 
.A(n_2390),
.B(n_2029),
.Y(n_2844)
);

INVx2_ASAP7_75t_L g2845 ( 
.A(n_2038),
.Y(n_2845)
);

AOI221xp5_ASAP7_75t_SL g2846 ( 
.A1(n_2417),
.A2(n_2434),
.B1(n_2332),
.B2(n_2150),
.C(n_2223),
.Y(n_2846)
);

OAI21x1_ASAP7_75t_SL g2847 ( 
.A1(n_2241),
.A2(n_2261),
.B(n_2249),
.Y(n_2847)
);

OAI21x1_ASAP7_75t_L g2848 ( 
.A1(n_2568),
.A2(n_2264),
.B(n_2200),
.Y(n_2848)
);

OAI22xp5_ASAP7_75t_L g2849 ( 
.A1(n_2358),
.A2(n_2412),
.B1(n_2147),
.B2(n_2178),
.Y(n_2849)
);

OAI21x1_ASAP7_75t_L g2850 ( 
.A1(n_2200),
.A2(n_2151),
.B(n_2565),
.Y(n_2850)
);

AOI221x1_ASAP7_75t_L g2851 ( 
.A1(n_2299),
.A2(n_2454),
.B1(n_2372),
.B2(n_2532),
.C(n_2457),
.Y(n_2851)
);

OAI21x1_ASAP7_75t_SL g2852 ( 
.A1(n_2261),
.A2(n_2263),
.B(n_2262),
.Y(n_2852)
);

A2O1A1Ixp33_ASAP7_75t_L g2853 ( 
.A1(n_2329),
.A2(n_2231),
.B(n_2228),
.C(n_2198),
.Y(n_2853)
);

OAI22xp5_ASAP7_75t_L g2854 ( 
.A1(n_2412),
.A2(n_2147),
.B1(n_2119),
.B2(n_2434),
.Y(n_2854)
);

OA22x2_ASAP7_75t_L g2855 ( 
.A1(n_2369),
.A2(n_2370),
.B1(n_2299),
.B2(n_2381),
.Y(n_2855)
);

BUFx6f_ASAP7_75t_L g2856 ( 
.A(n_2078),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2223),
.Y(n_2857)
);

AOI21x1_ASAP7_75t_L g2858 ( 
.A1(n_2280),
.A2(n_2345),
.B(n_2010),
.Y(n_2858)
);

OAI21xp5_ASAP7_75t_L g2859 ( 
.A1(n_2457),
.A2(n_2459),
.B(n_2308),
.Y(n_2859)
);

OAI21xp5_ASAP7_75t_L g2860 ( 
.A1(n_2459),
.A2(n_2055),
.B(n_2290),
.Y(n_2860)
);

AND2x2_ASAP7_75t_L g2861 ( 
.A(n_2254),
.B(n_2256),
.Y(n_2861)
);

INVxp67_ASAP7_75t_SL g2862 ( 
.A(n_2298),
.Y(n_2862)
);

BUFx3_ASAP7_75t_L g2863 ( 
.A(n_2094),
.Y(n_2863)
);

INVx3_ASAP7_75t_L g2864 ( 
.A(n_2151),
.Y(n_2864)
);

OAI21x1_ASAP7_75t_L g2865 ( 
.A1(n_2200),
.A2(n_2151),
.B(n_2565),
.Y(n_2865)
);

OAI21x1_ASAP7_75t_L g2866 ( 
.A1(n_2452),
.A2(n_2503),
.B(n_2010),
.Y(n_2866)
);

A2O1A1Ixp33_ASAP7_75t_L g2867 ( 
.A1(n_2132),
.A2(n_2179),
.B(n_2478),
.C(n_2517),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2254),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_L g2869 ( 
.A(n_2256),
.B(n_2350),
.Y(n_2869)
);

BUFx2_ASAP7_75t_L g2870 ( 
.A(n_2507),
.Y(n_2870)
);

AND3x4_ASAP7_75t_L g2871 ( 
.A(n_2094),
.B(n_2118),
.C(n_2107),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2350),
.B(n_2355),
.Y(n_2872)
);

AOI21xp5_ASAP7_75t_L g2873 ( 
.A1(n_2419),
.A2(n_2142),
.B(n_2137),
.Y(n_2873)
);

HB1xp67_ASAP7_75t_L g2874 ( 
.A(n_2122),
.Y(n_2874)
);

INVx3_ASAP7_75t_L g2875 ( 
.A(n_2351),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2397),
.Y(n_2876)
);

INVx2_ASAP7_75t_SL g2877 ( 
.A(n_2426),
.Y(n_2877)
);

OAI21x1_ASAP7_75t_L g2878 ( 
.A1(n_2452),
.A2(n_2503),
.B(n_2529),
.Y(n_2878)
);

AOI22xp33_ASAP7_75t_L g2879 ( 
.A1(n_2487),
.A2(n_2489),
.B1(n_2061),
.B2(n_2426),
.Y(n_2879)
);

INVxp67_ASAP7_75t_SL g2880 ( 
.A(n_2298),
.Y(n_2880)
);

AOI21xp5_ASAP7_75t_L g2881 ( 
.A1(n_2419),
.A2(n_2157),
.B(n_2149),
.Y(n_2881)
);

OAI22xp5_ASAP7_75t_L g2882 ( 
.A1(n_2489),
.A2(n_2294),
.B1(n_2262),
.B2(n_2263),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2355),
.B(n_2363),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2073),
.Y(n_2884)
);

OAI21x1_ASAP7_75t_L g2885 ( 
.A1(n_2452),
.A2(n_2503),
.B(n_2529),
.Y(n_2885)
);

BUFx2_ASAP7_75t_L g2886 ( 
.A(n_2507),
.Y(n_2886)
);

AND2x2_ASAP7_75t_L g2887 ( 
.A(n_2473),
.B(n_2520),
.Y(n_2887)
);

AO31x2_ASAP7_75t_L g2888 ( 
.A1(n_2532),
.A2(n_2454),
.A3(n_2258),
.B(n_2564),
.Y(n_2888)
);

AOI21xp5_ASAP7_75t_L g2889 ( 
.A1(n_2419),
.A2(n_2124),
.B(n_2287),
.Y(n_2889)
);

OAI21x1_ASAP7_75t_L g2890 ( 
.A1(n_2452),
.A2(n_2503),
.B(n_2529),
.Y(n_2890)
);

OAI21xp5_ASAP7_75t_L g2891 ( 
.A1(n_2492),
.A2(n_2439),
.B(n_2409),
.Y(n_2891)
);

INVx3_ASAP7_75t_L g2892 ( 
.A(n_2351),
.Y(n_2892)
);

OAI21x1_ASAP7_75t_L g2893 ( 
.A1(n_2529),
.A2(n_2501),
.B(n_2123),
.Y(n_2893)
);

NOR2xp67_ASAP7_75t_L g2894 ( 
.A(n_2025),
.B(n_2351),
.Y(n_2894)
);

BUFx6f_ASAP7_75t_L g2895 ( 
.A(n_2078),
.Y(n_2895)
);

AND2x4_ASAP7_75t_L g2896 ( 
.A(n_2310),
.B(n_2496),
.Y(n_2896)
);

OAI21x1_ASAP7_75t_L g2897 ( 
.A1(n_2501),
.A2(n_2123),
.B(n_2067),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_SL g2898 ( 
.A(n_2105),
.B(n_2393),
.Y(n_2898)
);

AND2x4_ASAP7_75t_L g2899 ( 
.A(n_2310),
.B(n_2496),
.Y(n_2899)
);

O2A1O1Ixp5_ASAP7_75t_L g2900 ( 
.A1(n_2320),
.A2(n_2283),
.B(n_2100),
.C(n_2103),
.Y(n_2900)
);

HB1xp67_ASAP7_75t_L g2901 ( 
.A(n_2473),
.Y(n_2901)
);

INVx5_ASAP7_75t_L g2902 ( 
.A(n_2025),
.Y(n_2902)
);

OR2x6_ASAP7_75t_L g2903 ( 
.A(n_2359),
.B(n_2384),
.Y(n_2903)
);

AOI21xp5_ASAP7_75t_L g2904 ( 
.A1(n_2482),
.A2(n_2439),
.B(n_2409),
.Y(n_2904)
);

AOI211x1_ASAP7_75t_L g2905 ( 
.A1(n_2272),
.A2(n_2279),
.B(n_2281),
.C(n_2292),
.Y(n_2905)
);

OAI22xp5_ASAP7_75t_L g2906 ( 
.A1(n_2272),
.A2(n_2292),
.B1(n_2281),
.B2(n_2279),
.Y(n_2906)
);

AOI21xp5_ASAP7_75t_L g2907 ( 
.A1(n_2482),
.A2(n_2439),
.B(n_2409),
.Y(n_2907)
);

AO32x2_ASAP7_75t_L g2908 ( 
.A1(n_2492),
.A2(n_2351),
.A3(n_2407),
.B1(n_2435),
.B2(n_2427),
.Y(n_2908)
);

OAI21xp5_ASAP7_75t_L g2909 ( 
.A1(n_2409),
.A2(n_2439),
.B(n_2449),
.Y(n_2909)
);

OR2x2_ASAP7_75t_L g2910 ( 
.A(n_2305),
.B(n_2311),
.Y(n_2910)
);

NOR2xp33_ASAP7_75t_L g2911 ( 
.A(n_2571),
.B(n_2088),
.Y(n_2911)
);

A2O1A1Ixp33_ASAP7_75t_L g2912 ( 
.A1(n_2179),
.A2(n_2517),
.B(n_2175),
.C(n_2160),
.Y(n_2912)
);

AOI21xp5_ASAP7_75t_L g2913 ( 
.A1(n_2482),
.A2(n_2518),
.B(n_2123),
.Y(n_2913)
);

NOR2xp33_ASAP7_75t_L g2914 ( 
.A(n_2109),
.B(n_2105),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2408),
.Y(n_2915)
);

OAI22x1_ASAP7_75t_L g2916 ( 
.A1(n_2268),
.A2(n_2472),
.B1(n_2229),
.B2(n_2406),
.Y(n_2916)
);

AO31x2_ASAP7_75t_L g2917 ( 
.A1(n_2073),
.A2(n_2303),
.A3(n_2258),
.B(n_2564),
.Y(n_2917)
);

OAI21xp5_ASAP7_75t_L g2918 ( 
.A1(n_2449),
.A2(n_2229),
.B(n_2543),
.Y(n_2918)
);

AOI21xp5_ASAP7_75t_L g2919 ( 
.A1(n_2482),
.A2(n_2518),
.B(n_2067),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2408),
.Y(n_2920)
);

AOI21xp5_ASAP7_75t_L g2921 ( 
.A1(n_2482),
.A2(n_2067),
.B(n_2359),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2073),
.Y(n_2922)
);

OAI21x1_ASAP7_75t_L g2923 ( 
.A1(n_2543),
.A2(n_2396),
.B(n_2301),
.Y(n_2923)
);

OAI21x1_ASAP7_75t_L g2924 ( 
.A1(n_2396),
.A2(n_2301),
.B(n_2410),
.Y(n_2924)
);

OAI21xp33_ASAP7_75t_L g2925 ( 
.A1(n_2374),
.A2(n_2379),
.B(n_2375),
.Y(n_2925)
);

OAI21x1_ASAP7_75t_L g2926 ( 
.A1(n_2422),
.A2(n_2450),
.B(n_2431),
.Y(n_2926)
);

OAI21x1_ASAP7_75t_L g2927 ( 
.A1(n_2422),
.A2(n_2450),
.B(n_2431),
.Y(n_2927)
);

AOI21xp5_ASAP7_75t_L g2928 ( 
.A1(n_2359),
.A2(n_2428),
.B(n_2384),
.Y(n_2928)
);

INVx2_ASAP7_75t_L g2929 ( 
.A(n_2110),
.Y(n_2929)
);

OAI22xp5_ASAP7_75t_L g2930 ( 
.A1(n_2268),
.A2(n_2584),
.B1(n_2247),
.B2(n_2169),
.Y(n_2930)
);

OAI21x1_ASAP7_75t_L g2931 ( 
.A1(n_2468),
.A2(n_2506),
.B(n_2504),
.Y(n_2931)
);

INVx6_ASAP7_75t_L g2932 ( 
.A(n_2451),
.Y(n_2932)
);

OAI21xp5_ASAP7_75t_L g2933 ( 
.A1(n_2411),
.A2(n_2445),
.B(n_2474),
.Y(n_2933)
);

OAI22x1_ASAP7_75t_L g2934 ( 
.A1(n_2472),
.A2(n_2520),
.B1(n_2498),
.B2(n_2516),
.Y(n_2934)
);

OAI21x1_ASAP7_75t_SL g2935 ( 
.A1(n_2025),
.A2(n_2527),
.B(n_2461),
.Y(n_2935)
);

OAI22xp5_ASAP7_75t_L g2936 ( 
.A1(n_2584),
.A2(n_2401),
.B1(n_2094),
.B2(n_2118),
.Y(n_2936)
);

BUFx10_ASAP7_75t_L g2937 ( 
.A(n_2312),
.Y(n_2937)
);

NAND2x1_ASAP7_75t_L g2938 ( 
.A(n_2461),
.B(n_2527),
.Y(n_2938)
);

HB1xp67_ASAP7_75t_L g2939 ( 
.A(n_2305),
.Y(n_2939)
);

AO31x2_ASAP7_75t_L g2940 ( 
.A1(n_2110),
.A2(n_2564),
.A3(n_2550),
.B(n_2549),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_L g2941 ( 
.A(n_2363),
.B(n_2365),
.Y(n_2941)
);

INVxp67_ASAP7_75t_L g2942 ( 
.A(n_2105),
.Y(n_2942)
);

OAI21x1_ASAP7_75t_L g2943 ( 
.A1(n_2468),
.A2(n_2504),
.B(n_2539),
.Y(n_2943)
);

AND2x4_ASAP7_75t_L g2944 ( 
.A(n_2310),
.B(n_2496),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2413),
.Y(n_2945)
);

BUFx3_ASAP7_75t_L g2946 ( 
.A(n_2107),
.Y(n_2946)
);

OA21x2_ASAP7_75t_L g2947 ( 
.A1(n_2479),
.A2(n_2526),
.B(n_2521),
.Y(n_2947)
);

OAI21x1_ASAP7_75t_L g2948 ( 
.A1(n_2479),
.A2(n_2521),
.B(n_2534),
.Y(n_2948)
);

OAI21x1_ASAP7_75t_L g2949 ( 
.A1(n_2506),
.A2(n_2526),
.B(n_2534),
.Y(n_2949)
);

OAI21xp5_ASAP7_75t_L g2950 ( 
.A1(n_2383),
.A2(n_2486),
.B(n_2496),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_L g2951 ( 
.A(n_2365),
.B(n_2373),
.Y(n_2951)
);

AOI21xp5_ASAP7_75t_L g2952 ( 
.A1(n_2359),
.A2(n_2428),
.B(n_2384),
.Y(n_2952)
);

AOI21xp5_ASAP7_75t_L g2953 ( 
.A1(n_2359),
.A2(n_2428),
.B(n_2384),
.Y(n_2953)
);

OA22x2_ASAP7_75t_L g2954 ( 
.A1(n_2429),
.A2(n_2442),
.B1(n_2384),
.B2(n_2428),
.Y(n_2954)
);

INVx2_ASAP7_75t_SL g2955 ( 
.A(n_2425),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2373),
.B(n_2376),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_L g2957 ( 
.A(n_2376),
.B(n_2382),
.Y(n_2957)
);

OAI21x1_ASAP7_75t_L g2958 ( 
.A1(n_2531),
.A2(n_2537),
.B(n_2539),
.Y(n_2958)
);

AO21x1_ASAP7_75t_L g2959 ( 
.A1(n_2382),
.A2(n_2387),
.B(n_2391),
.Y(n_2959)
);

OAI21x1_ASAP7_75t_L g2960 ( 
.A1(n_2531),
.A2(n_2538),
.B(n_2537),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_L g2961 ( 
.A(n_2387),
.B(n_2391),
.Y(n_2961)
);

OAI21x1_ASAP7_75t_L g2962 ( 
.A1(n_2538),
.A2(n_2394),
.B(n_2510),
.Y(n_2962)
);

OAI21xp5_ASAP7_75t_L g2963 ( 
.A1(n_2383),
.A2(n_2486),
.B(n_2037),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2413),
.Y(n_2964)
);

AOI22xp5_ASAP7_75t_L g2965 ( 
.A1(n_2487),
.A2(n_2061),
.B1(n_2345),
.B2(n_2312),
.Y(n_2965)
);

CKINVDCx5p33_ASAP7_75t_R g2966 ( 
.A(n_2061),
.Y(n_2966)
);

INVx2_ASAP7_75t_L g2967 ( 
.A(n_2110),
.Y(n_2967)
);

OAI21x1_ASAP7_75t_L g2968 ( 
.A1(n_2394),
.A2(n_2510),
.B(n_2549),
.Y(n_2968)
);

BUFx8_ASAP7_75t_SL g2969 ( 
.A(n_2312),
.Y(n_2969)
);

OAI21x1_ASAP7_75t_L g2970 ( 
.A1(n_2116),
.A2(n_2550),
.B(n_2549),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_L g2971 ( 
.A(n_2311),
.B(n_2116),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2443),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2116),
.B(n_2139),
.Y(n_2973)
);

OAI21xp5_ASAP7_75t_L g2974 ( 
.A1(n_2486),
.A2(n_2012),
.B(n_2037),
.Y(n_2974)
);

BUFx2_ASAP7_75t_L g2975 ( 
.A(n_2498),
.Y(n_2975)
);

INVx2_ASAP7_75t_L g2976 ( 
.A(n_2139),
.Y(n_2976)
);

AO22x2_ASAP7_75t_L g2977 ( 
.A1(n_2310),
.A2(n_2444),
.B1(n_2466),
.B2(n_2512),
.Y(n_2977)
);

OAI21xp5_ASAP7_75t_L g2978 ( 
.A1(n_2486),
.A2(n_2012),
.B(n_2037),
.Y(n_2978)
);

AND2x2_ASAP7_75t_L g2979 ( 
.A(n_2425),
.B(n_2012),
.Y(n_2979)
);

INVx3_ASAP7_75t_SL g2980 ( 
.A(n_2498),
.Y(n_2980)
);

OAI21x1_ASAP7_75t_L g2981 ( 
.A1(n_2139),
.A2(n_2550),
.B(n_2218),
.Y(n_2981)
);

NOR2x1_ASAP7_75t_SL g2982 ( 
.A(n_2428),
.B(n_2233),
.Y(n_2982)
);

OAI21x1_ASAP7_75t_L g2983 ( 
.A1(n_2145),
.A2(n_2154),
.B(n_2215),
.Y(n_2983)
);

INVxp67_ASAP7_75t_L g2984 ( 
.A(n_2012),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2145),
.B(n_2146),
.Y(n_2985)
);

AOI21xp5_ASAP7_75t_L g2986 ( 
.A1(n_2455),
.A2(n_2243),
.B(n_2078),
.Y(n_2986)
);

AOI21xp5_ASAP7_75t_L g2987 ( 
.A1(n_2455),
.A2(n_2440),
.B(n_2377),
.Y(n_2987)
);

OAI22xp5_ASAP7_75t_L g2988 ( 
.A1(n_2107),
.A2(n_2118),
.B1(n_2367),
.B2(n_2282),
.Y(n_2988)
);

AOI21xp5_ASAP7_75t_L g2989 ( 
.A1(n_2455),
.A2(n_2440),
.B(n_2377),
.Y(n_2989)
);

INVx1_ASAP7_75t_SL g2990 ( 
.A(n_2505),
.Y(n_2990)
);

OAI21x1_ASAP7_75t_L g2991 ( 
.A1(n_2145),
.A2(n_2303),
.B(n_2258),
.Y(n_2991)
);

AOI21xp5_ASAP7_75t_L g2992 ( 
.A1(n_2455),
.A2(n_2440),
.B(n_2377),
.Y(n_2992)
);

OAI21x1_ASAP7_75t_L g2993 ( 
.A1(n_2146),
.A2(n_2303),
.B(n_2232),
.Y(n_2993)
);

OAI21xp5_ASAP7_75t_L g2994 ( 
.A1(n_2037),
.A2(n_2101),
.B(n_2414),
.Y(n_2994)
);

AND2x2_ASAP7_75t_L g2995 ( 
.A(n_2101),
.B(n_2414),
.Y(n_2995)
);

OAI21x1_ASAP7_75t_L g2996 ( 
.A1(n_2146),
.A2(n_2245),
.B(n_2154),
.Y(n_2996)
);

INVx2_ASAP7_75t_L g2997 ( 
.A(n_2154),
.Y(n_2997)
);

NOR2xp33_ASAP7_75t_L g2998 ( 
.A(n_2481),
.B(n_2101),
.Y(n_2998)
);

OAI21xp5_ASAP7_75t_L g2999 ( 
.A1(n_2101),
.A2(n_2257),
.B(n_2174),
.Y(n_2999)
);

OAI21x1_ASAP7_75t_L g3000 ( 
.A1(n_2156),
.A2(n_2248),
.B(n_2232),
.Y(n_3000)
);

OAI21x1_ASAP7_75t_L g3001 ( 
.A1(n_2156),
.A2(n_2248),
.B(n_2232),
.Y(n_3001)
);

NAND2x1p5_ASAP7_75t_L g3002 ( 
.A(n_2407),
.B(n_2427),
.Y(n_3002)
);

INVxp67_ASAP7_75t_L g3003 ( 
.A(n_2174),
.Y(n_3003)
);

OA22x2_ASAP7_75t_L g3004 ( 
.A1(n_2174),
.A2(n_2257),
.B1(n_2205),
.B2(n_2414),
.Y(n_3004)
);

AOI21xp5_ASAP7_75t_L g3005 ( 
.A1(n_2213),
.A2(n_2246),
.B(n_2377),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_2156),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2215),
.B(n_2248),
.Y(n_3007)
);

NAND2xp5_ASAP7_75t_L g3008 ( 
.A(n_2215),
.B(n_2245),
.Y(n_3008)
);

BUFx3_ASAP7_75t_L g3009 ( 
.A(n_2233),
.Y(n_3009)
);

AO31x2_ASAP7_75t_L g3010 ( 
.A1(n_2216),
.A2(n_2245),
.A3(n_2218),
.B(n_2541),
.Y(n_3010)
);

O2A1O1Ixp5_ASAP7_75t_L g3011 ( 
.A1(n_2461),
.A2(n_2527),
.B(n_2427),
.C(n_2407),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_L g3012 ( 
.A(n_2216),
.B(n_2218),
.Y(n_3012)
);

AOI221xp5_ASAP7_75t_L g3013 ( 
.A1(n_2174),
.A2(n_2205),
.B1(n_2414),
.B2(n_2257),
.C(n_2512),
.Y(n_3013)
);

BUFx2_ASAP7_75t_SL g3014 ( 
.A(n_2407),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2466),
.Y(n_3015)
);

INVxp67_ASAP7_75t_SL g3016 ( 
.A(n_2530),
.Y(n_3016)
);

AOI21xp5_ASAP7_75t_L g3017 ( 
.A1(n_2213),
.A2(n_2440),
.B(n_2377),
.Y(n_3017)
);

AOI21xp33_ASAP7_75t_L g3018 ( 
.A1(n_2361),
.A2(n_2216),
.B(n_2541),
.Y(n_3018)
);

INVx1_ASAP7_75t_SL g3019 ( 
.A(n_2505),
.Y(n_3019)
);

AO31x2_ASAP7_75t_L g3020 ( 
.A1(n_2313),
.A2(n_2404),
.A3(n_2536),
.B(n_2524),
.Y(n_3020)
);

OAI21x1_ASAP7_75t_SL g3021 ( 
.A1(n_2461),
.A2(n_2527),
.B(n_2435),
.Y(n_3021)
);

NAND2x1_ASAP7_75t_L g3022 ( 
.A(n_2427),
.B(n_2435),
.Y(n_3022)
);

AOI21x1_ASAP7_75t_L g3023 ( 
.A1(n_2205),
.A2(n_2257),
.B(n_2536),
.Y(n_3023)
);

AO31x2_ASAP7_75t_L g3024 ( 
.A1(n_2313),
.A2(n_2403),
.A3(n_2536),
.B(n_2524),
.Y(n_3024)
);

OAI21x1_ASAP7_75t_L g3025 ( 
.A1(n_2313),
.A2(n_2399),
.B(n_2524),
.Y(n_3025)
);

BUFx6f_ASAP7_75t_L g3026 ( 
.A(n_2213),
.Y(n_3026)
);

OAI21x1_ASAP7_75t_L g3027 ( 
.A1(n_2315),
.A2(n_2399),
.B(n_2508),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2487),
.B(n_2205),
.Y(n_3028)
);

OAI21x1_ASAP7_75t_L g3029 ( 
.A1(n_2315),
.A2(n_2403),
.B(n_2508),
.Y(n_3029)
);

AND2x4_ASAP7_75t_L g3030 ( 
.A(n_2435),
.B(n_2213),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2487),
.B(n_2378),
.Y(n_3031)
);

OAI22xp5_ASAP7_75t_L g3032 ( 
.A1(n_2233),
.A2(n_2367),
.B1(n_2282),
.B2(n_2481),
.Y(n_3032)
);

OAI21x1_ASAP7_75t_L g3033 ( 
.A1(n_2315),
.A2(n_2399),
.B(n_2508),
.Y(n_3033)
);

OAI21xp33_ASAP7_75t_SL g3034 ( 
.A1(n_2456),
.A2(n_2541),
.B(n_2415),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_SL g3035 ( 
.A(n_2519),
.B(n_2213),
.Y(n_3035)
);

OAI21x1_ASAP7_75t_L g3036 ( 
.A1(n_2323),
.A2(n_2378),
.B(n_2403),
.Y(n_3036)
);

BUFx2_ASAP7_75t_L g3037 ( 
.A(n_2456),
.Y(n_3037)
);

BUFx3_ASAP7_75t_L g3038 ( 
.A(n_2282),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2323),
.B(n_2378),
.Y(n_3039)
);

O2A1O1Ixp5_ASAP7_75t_L g3040 ( 
.A1(n_2323),
.A2(n_2464),
.B(n_2404),
.C(n_2415),
.Y(n_3040)
);

OR2x2_ASAP7_75t_L g3041 ( 
.A(n_2326),
.B(n_2404),
.Y(n_3041)
);

AOI22xp5_ASAP7_75t_L g3042 ( 
.A1(n_2367),
.A2(n_2451),
.B1(n_2464),
.B2(n_2336),
.Y(n_3042)
);

OAI21x1_ASAP7_75t_L g3043 ( 
.A1(n_2326),
.A2(n_2415),
.B(n_2366),
.Y(n_3043)
);

OAI21xp5_ASAP7_75t_L g3044 ( 
.A1(n_2326),
.A2(n_2349),
.B(n_2464),
.Y(n_3044)
);

OAI21xp5_ASAP7_75t_L g3045 ( 
.A1(n_2333),
.A2(n_2349),
.B(n_2366),
.Y(n_3045)
);

OAI21xp5_ASAP7_75t_L g3046 ( 
.A1(n_2333),
.A2(n_2349),
.B(n_2366),
.Y(n_3046)
);

AND2x4_ASAP7_75t_L g3047 ( 
.A(n_2213),
.B(n_2243),
.Y(n_3047)
);

AOI21xp5_ASAP7_75t_L g3048 ( 
.A1(n_2243),
.A2(n_2246),
.B(n_2490),
.Y(n_3048)
);

OAI22xp5_ASAP7_75t_SL g3049 ( 
.A1(n_2456),
.A2(n_2243),
.B1(n_2246),
.B2(n_2490),
.Y(n_3049)
);

AOI21xp5_ASAP7_75t_L g3050 ( 
.A1(n_2243),
.A2(n_2246),
.B(n_2490),
.Y(n_3050)
);

A2O1A1Ixp33_ASAP7_75t_L g3051 ( 
.A1(n_2456),
.A2(n_2353),
.B(n_2336),
.C(n_2333),
.Y(n_3051)
);

INVx2_ASAP7_75t_SL g3052 ( 
.A(n_2243),
.Y(n_3052)
);

BUFx2_ASAP7_75t_L g3053 ( 
.A(n_2456),
.Y(n_3053)
);

OAI21xp5_ASAP7_75t_L g3054 ( 
.A1(n_2336),
.A2(n_2353),
.B(n_2456),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2353),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_2246),
.B(n_2377),
.Y(n_3056)
);

AOI21x1_ASAP7_75t_L g3057 ( 
.A1(n_2509),
.A2(n_2451),
.B(n_2440),
.Y(n_3057)
);

INVx4_ASAP7_75t_L g3058 ( 
.A(n_2246),
.Y(n_3058)
);

AOI21xp5_ASAP7_75t_L g3059 ( 
.A1(n_2440),
.A2(n_2476),
.B(n_2490),
.Y(n_3059)
);

AND2x2_ASAP7_75t_L g3060 ( 
.A(n_2476),
.B(n_2490),
.Y(n_3060)
);

AND2x2_ASAP7_75t_L g3061 ( 
.A(n_2476),
.B(n_2490),
.Y(n_3061)
);

OAI21x1_ASAP7_75t_L g3062 ( 
.A1(n_2509),
.A2(n_2476),
.B(n_2519),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2509),
.Y(n_3063)
);

AOI21xp5_ASAP7_75t_SL g3064 ( 
.A1(n_2519),
.A2(n_2476),
.B(n_2451),
.Y(n_3064)
);

OAI21x1_ASAP7_75t_L g3065 ( 
.A1(n_2509),
.A2(n_2476),
.B(n_2519),
.Y(n_3065)
);

AOI21xp33_ASAP7_75t_L g3066 ( 
.A1(n_2519),
.A2(n_2562),
.B(n_2548),
.Y(n_3066)
);

AO22x2_ASAP7_75t_L g3067 ( 
.A1(n_2509),
.A2(n_2562),
.B1(n_2574),
.B2(n_2548),
.Y(n_3067)
);

OAI22xp5_ASAP7_75t_L g3068 ( 
.A1(n_2519),
.A2(n_2559),
.B1(n_2588),
.B2(n_2562),
.Y(n_3068)
);

HB1xp67_ASAP7_75t_L g3069 ( 
.A(n_2509),
.Y(n_3069)
);

OAI21x1_ASAP7_75t_L g3070 ( 
.A1(n_2074),
.A2(n_2069),
.B(n_2098),
.Y(n_3070)
);

OAI21xp5_ASAP7_75t_L g3071 ( 
.A1(n_2014),
.A2(n_1054),
.B(n_2013),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_2040),
.B(n_2043),
.Y(n_3072)
);

OAI21x1_ASAP7_75t_L g3073 ( 
.A1(n_2074),
.A2(n_2069),
.B(n_2098),
.Y(n_3073)
);

A2O1A1Ixp33_ASAP7_75t_L g3074 ( 
.A1(n_2559),
.A2(n_1788),
.B(n_2588),
.C(n_2014),
.Y(n_3074)
);

A2O1A1Ixp33_ASAP7_75t_L g3075 ( 
.A1(n_2559),
.A2(n_1788),
.B(n_2588),
.C(n_2014),
.Y(n_3075)
);

NOR2xp33_ASAP7_75t_L g3076 ( 
.A(n_2087),
.B(n_666),
.Y(n_3076)
);

AND2x6_ASAP7_75t_L g3077 ( 
.A(n_2559),
.B(n_2588),
.Y(n_3077)
);

O2A1O1Ixp5_ASAP7_75t_L g3078 ( 
.A1(n_2026),
.A2(n_2548),
.B(n_2574),
.C(n_2562),
.Y(n_3078)
);

AO31x2_ASAP7_75t_L g3079 ( 
.A1(n_2026),
.A2(n_2074),
.A3(n_2300),
.B(n_2069),
.Y(n_3079)
);

AO32x2_ASAP7_75t_L g3080 ( 
.A1(n_2328),
.A2(n_2039),
.A3(n_2285),
.B1(n_2251),
.B2(n_2244),
.Y(n_3080)
);

INVx3_ASAP7_75t_L g3081 ( 
.A(n_2161),
.Y(n_3081)
);

AOI221x1_ASAP7_75t_L g3082 ( 
.A1(n_2002),
.A2(n_2082),
.B1(n_2013),
.B2(n_2562),
.C(n_2548),
.Y(n_3082)
);

OAI21x1_ASAP7_75t_L g3083 ( 
.A1(n_2074),
.A2(n_2069),
.B(n_2098),
.Y(n_3083)
);

O2A1O1Ixp33_ASAP7_75t_L g3084 ( 
.A1(n_2014),
.A2(n_2013),
.B(n_1989),
.C(n_1995),
.Y(n_3084)
);

AOI21x1_ASAP7_75t_L g3085 ( 
.A1(n_2058),
.A2(n_2210),
.B(n_2035),
.Y(n_3085)
);

AOI21xp5_ASAP7_75t_L g3086 ( 
.A1(n_1998),
.A2(n_1579),
.B(n_2555),
.Y(n_3086)
);

OAI21x1_ASAP7_75t_L g3087 ( 
.A1(n_2074),
.A2(n_2069),
.B(n_2098),
.Y(n_3087)
);

AO31x2_ASAP7_75t_L g3088 ( 
.A1(n_2026),
.A2(n_2074),
.A3(n_2300),
.B(n_2069),
.Y(n_3088)
);

INVx2_ASAP7_75t_L g3089 ( 
.A(n_2007),
.Y(n_3089)
);

OAI21xp5_ASAP7_75t_L g3090 ( 
.A1(n_2014),
.A2(n_1054),
.B(n_2013),
.Y(n_3090)
);

AO31x2_ASAP7_75t_L g3091 ( 
.A1(n_2026),
.A2(n_2074),
.A3(n_2300),
.B(n_2069),
.Y(n_3091)
);

NAND2x1p5_ASAP7_75t_L g3092 ( 
.A(n_2319),
.B(n_1415),
.Y(n_3092)
);

OAI21x1_ASAP7_75t_L g3093 ( 
.A1(n_2074),
.A2(n_2069),
.B(n_2098),
.Y(n_3093)
);

OAI21x1_ASAP7_75t_L g3094 ( 
.A1(n_2074),
.A2(n_2069),
.B(n_2098),
.Y(n_3094)
);

AO31x2_ASAP7_75t_L g3095 ( 
.A1(n_2026),
.A2(n_2074),
.A3(n_2300),
.B(n_2069),
.Y(n_3095)
);

OR2x2_ASAP7_75t_L g3096 ( 
.A(n_2551),
.B(n_2008),
.Y(n_3096)
);

AO21x1_ASAP7_75t_L g3097 ( 
.A1(n_2002),
.A2(n_2562),
.B(n_2548),
.Y(n_3097)
);

NAND2x1p5_ASAP7_75t_L g3098 ( 
.A(n_2319),
.B(n_1415),
.Y(n_3098)
);

AOI21xp5_ASAP7_75t_L g3099 ( 
.A1(n_1998),
.A2(n_1579),
.B(n_2555),
.Y(n_3099)
);

AND2x4_ASAP7_75t_L g3100 ( 
.A(n_2310),
.B(n_2085),
.Y(n_3100)
);

INVx1_ASAP7_75t_SL g3101 ( 
.A(n_2096),
.Y(n_3101)
);

AOI21xp5_ASAP7_75t_L g3102 ( 
.A1(n_1998),
.A2(n_1579),
.B(n_2555),
.Y(n_3102)
);

AND2x2_ASAP7_75t_L g3103 ( 
.A(n_1999),
.B(n_2083),
.Y(n_3103)
);

AOI21xp5_ASAP7_75t_L g3104 ( 
.A1(n_1998),
.A2(n_1579),
.B(n_2555),
.Y(n_3104)
);

OAI21x1_ASAP7_75t_L g3105 ( 
.A1(n_2074),
.A2(n_2069),
.B(n_2098),
.Y(n_3105)
);

OAI21x1_ASAP7_75t_L g3106 ( 
.A1(n_2074),
.A2(n_2069),
.B(n_2098),
.Y(n_3106)
);

AOI22xp5_ASAP7_75t_L g3107 ( 
.A1(n_2548),
.A2(n_2574),
.B1(n_2577),
.B2(n_2562),
.Y(n_3107)
);

AOI21xp5_ASAP7_75t_L g3108 ( 
.A1(n_1998),
.A2(n_1579),
.B(n_2555),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_2040),
.B(n_2043),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_2007),
.Y(n_3110)
);

BUFx6f_ASAP7_75t_L g3111 ( 
.A(n_2078),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_2040),
.B(n_2043),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_2040),
.B(n_2043),
.Y(n_3113)
);

OAI21x1_ASAP7_75t_L g3114 ( 
.A1(n_2074),
.A2(n_2069),
.B(n_2098),
.Y(n_3114)
);

OAI21xp5_ASAP7_75t_L g3115 ( 
.A1(n_2014),
.A2(n_1054),
.B(n_2013),
.Y(n_3115)
);

AOI21xp5_ASAP7_75t_L g3116 ( 
.A1(n_1998),
.A2(n_1579),
.B(n_2555),
.Y(n_3116)
);

OAI21x1_ASAP7_75t_L g3117 ( 
.A1(n_2074),
.A2(n_2069),
.B(n_2098),
.Y(n_3117)
);

AOI21xp5_ASAP7_75t_L g3118 ( 
.A1(n_1998),
.A2(n_1579),
.B(n_2555),
.Y(n_3118)
);

OAI21xp5_ASAP7_75t_L g3119 ( 
.A1(n_2014),
.A2(n_1054),
.B(n_2013),
.Y(n_3119)
);

AOI21x1_ASAP7_75t_SL g3120 ( 
.A1(n_2112),
.A2(n_1724),
.B(n_1722),
.Y(n_3120)
);

BUFx2_ASAP7_75t_L g3121 ( 
.A(n_2009),
.Y(n_3121)
);

AOI21xp5_ASAP7_75t_L g3122 ( 
.A1(n_1998),
.A2(n_1579),
.B(n_2555),
.Y(n_3122)
);

A2O1A1Ixp33_ASAP7_75t_L g3123 ( 
.A1(n_2559),
.A2(n_1788),
.B(n_2588),
.C(n_2014),
.Y(n_3123)
);

OAI21xp33_ASAP7_75t_L g3124 ( 
.A1(n_2002),
.A2(n_1788),
.B(n_2072),
.Y(n_3124)
);

OAI22xp33_ASAP7_75t_L g3125 ( 
.A1(n_2559),
.A2(n_2588),
.B1(n_2562),
.B2(n_2574),
.Y(n_3125)
);

INVx3_ASAP7_75t_L g3126 ( 
.A(n_2161),
.Y(n_3126)
);

AOI21xp5_ASAP7_75t_L g3127 ( 
.A1(n_1998),
.A2(n_1579),
.B(n_2555),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_SL g3128 ( 
.A(n_2003),
.B(n_2553),
.Y(n_3128)
);

OAI21x1_ASAP7_75t_SL g3129 ( 
.A1(n_2026),
.A2(n_2562),
.B(n_2548),
.Y(n_3129)
);

OAI21x1_ASAP7_75t_L g3130 ( 
.A1(n_2074),
.A2(n_2069),
.B(n_2098),
.Y(n_3130)
);

INVx2_ASAP7_75t_SL g3131 ( 
.A(n_2121),
.Y(n_3131)
);

NAND2x1p5_ASAP7_75t_L g3132 ( 
.A(n_2319),
.B(n_1415),
.Y(n_3132)
);

NAND2xp5_ASAP7_75t_SL g3133 ( 
.A(n_2003),
.B(n_2553),
.Y(n_3133)
);

NOR2xp33_ASAP7_75t_L g3134 ( 
.A(n_2087),
.B(n_666),
.Y(n_3134)
);

OAI21x1_ASAP7_75t_L g3135 ( 
.A1(n_2074),
.A2(n_2069),
.B(n_2098),
.Y(n_3135)
);

OAI21x1_ASAP7_75t_L g3136 ( 
.A1(n_2074),
.A2(n_2069),
.B(n_2098),
.Y(n_3136)
);

OAI21xp5_ASAP7_75t_L g3137 ( 
.A1(n_2014),
.A2(n_1054),
.B(n_2013),
.Y(n_3137)
);

AO21x2_ASAP7_75t_L g3138 ( 
.A1(n_2026),
.A2(n_2190),
.B(n_2181),
.Y(n_3138)
);

INVx3_ASAP7_75t_SL g3139 ( 
.A(n_2441),
.Y(n_3139)
);

AOI21xp5_ASAP7_75t_L g3140 ( 
.A1(n_1998),
.A2(n_1579),
.B(n_2555),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2321),
.Y(n_3141)
);

AO31x2_ASAP7_75t_L g3142 ( 
.A1(n_2026),
.A2(n_2074),
.A3(n_2300),
.B(n_2069),
.Y(n_3142)
);

OA22x2_ASAP7_75t_L g3143 ( 
.A1(n_2001),
.A2(n_2588),
.B1(n_2559),
.B2(n_2015),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_L g3144 ( 
.A(n_2040),
.B(n_2043),
.Y(n_3144)
);

OR2x2_ASAP7_75t_L g3145 ( 
.A(n_2756),
.B(n_2799),
.Y(n_3145)
);

O2A1O1Ixp33_ASAP7_75t_L g3146 ( 
.A1(n_2656),
.A2(n_3090),
.B(n_3115),
.C(n_3071),
.Y(n_3146)
);

AOI22xp5_ASAP7_75t_L g3147 ( 
.A1(n_3097),
.A2(n_2608),
.B1(n_2617),
.B2(n_3107),
.Y(n_3147)
);

INVx2_ASAP7_75t_SL g3148 ( 
.A(n_3004),
.Y(n_3148)
);

CKINVDCx20_ASAP7_75t_R g3149 ( 
.A(n_2785),
.Y(n_3149)
);

BUFx2_ASAP7_75t_L g3150 ( 
.A(n_3004),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_2609),
.B(n_2623),
.Y(n_3151)
);

CKINVDCx20_ASAP7_75t_R g3152 ( 
.A(n_2966),
.Y(n_3152)
);

AOI21xp5_ASAP7_75t_SL g3153 ( 
.A1(n_3082),
.A2(n_2734),
.B(n_2612),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_2647),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_2647),
.Y(n_3155)
);

AOI21xp5_ASAP7_75t_L g3156 ( 
.A1(n_3086),
.A2(n_3102),
.B(n_3099),
.Y(n_3156)
);

OR2x2_ASAP7_75t_SL g3157 ( 
.A(n_2591),
.B(n_2625),
.Y(n_3157)
);

AND2x4_ASAP7_75t_L g3158 ( 
.A(n_2622),
.B(n_2680),
.Y(n_3158)
);

BUFx2_ASAP7_75t_L g3159 ( 
.A(n_3004),
.Y(n_3159)
);

O2A1O1Ixp5_ASAP7_75t_L g3160 ( 
.A1(n_3097),
.A2(n_2608),
.B(n_3078),
.C(n_2605),
.Y(n_3160)
);

AND2x2_ASAP7_75t_L g3161 ( 
.A(n_2741),
.B(n_2794),
.Y(n_3161)
);

AOI21xp5_ASAP7_75t_L g3162 ( 
.A1(n_3086),
.A2(n_3102),
.B(n_3099),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_2686),
.Y(n_3163)
);

O2A1O1Ixp33_ASAP7_75t_L g3164 ( 
.A1(n_3071),
.A2(n_3090),
.B(n_3119),
.C(n_3115),
.Y(n_3164)
);

OAI22xp5_ASAP7_75t_L g3165 ( 
.A1(n_3107),
.A2(n_2617),
.B1(n_2661),
.B2(n_2605),
.Y(n_3165)
);

BUFx12f_ASAP7_75t_L g3166 ( 
.A(n_2707),
.Y(n_3166)
);

AND2x2_ASAP7_75t_L g3167 ( 
.A(n_2741),
.B(n_2794),
.Y(n_3167)
);

OR2x2_ASAP7_75t_L g3168 ( 
.A(n_2756),
.B(n_2799),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2686),
.Y(n_3169)
);

AOI21xp5_ASAP7_75t_L g3170 ( 
.A1(n_3104),
.A2(n_3116),
.B(n_3108),
.Y(n_3170)
);

INVx2_ASAP7_75t_L g3171 ( 
.A(n_2643),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_2643),
.Y(n_3172)
);

AND2x4_ASAP7_75t_L g3173 ( 
.A(n_2622),
.B(n_2680),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2716),
.Y(n_3174)
);

NOR2xp33_ASAP7_75t_SL g3175 ( 
.A(n_3124),
.B(n_3129),
.Y(n_3175)
);

INVx3_ASAP7_75t_L g3176 ( 
.A(n_3062),
.Y(n_3176)
);

A2O1A1Ixp33_ASAP7_75t_L g3177 ( 
.A1(n_3084),
.A2(n_2612),
.B(n_3124),
.C(n_2625),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_2716),
.Y(n_3178)
);

INVx3_ASAP7_75t_L g3179 ( 
.A(n_3062),
.Y(n_3179)
);

A2O1A1Ixp33_ASAP7_75t_L g3180 ( 
.A1(n_3084),
.A2(n_2591),
.B(n_3075),
.C(n_3074),
.Y(n_3180)
);

AOI22xp33_ASAP7_75t_L g3181 ( 
.A1(n_3143),
.A2(n_3077),
.B1(n_2606),
.B2(n_3125),
.Y(n_3181)
);

AND2x4_ASAP7_75t_L g3182 ( 
.A(n_2680),
.B(n_2896),
.Y(n_3182)
);

HB1xp67_ASAP7_75t_L g3183 ( 
.A(n_2832),
.Y(n_3183)
);

AOI21xp5_ASAP7_75t_L g3184 ( 
.A1(n_3104),
.A2(n_3116),
.B(n_3108),
.Y(n_3184)
);

CKINVDCx5p33_ASAP7_75t_R g3185 ( 
.A(n_2808),
.Y(n_3185)
);

AND2x4_ASAP7_75t_L g3186 ( 
.A(n_2680),
.B(n_2896),
.Y(n_3186)
);

OR2x6_ASAP7_75t_L g3187 ( 
.A(n_2807),
.B(n_2977),
.Y(n_3187)
);

AND2x4_ASAP7_75t_L g3188 ( 
.A(n_2680),
.B(n_2896),
.Y(n_3188)
);

INVx5_ASAP7_75t_L g3189 ( 
.A(n_2795),
.Y(n_3189)
);

OR2x2_ASAP7_75t_L g3190 ( 
.A(n_2837),
.B(n_2803),
.Y(n_3190)
);

BUFx6f_ASAP7_75t_L g3191 ( 
.A(n_2630),
.Y(n_3191)
);

A2O1A1Ixp33_ASAP7_75t_L g3192 ( 
.A1(n_3123),
.A2(n_2661),
.B(n_3137),
.C(n_3119),
.Y(n_3192)
);

INVx5_ASAP7_75t_L g3193 ( 
.A(n_2795),
.Y(n_3193)
);

AND2x4_ASAP7_75t_L g3194 ( 
.A(n_2680),
.B(n_2896),
.Y(n_3194)
);

AND2x2_ASAP7_75t_L g3195 ( 
.A(n_2805),
.B(n_2811),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_L g3196 ( 
.A(n_2609),
.B(n_2623),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_L g3197 ( 
.A(n_3072),
.B(n_3109),
.Y(n_3197)
);

INVx3_ASAP7_75t_L g3198 ( 
.A(n_3062),
.Y(n_3198)
);

BUFx2_ASAP7_75t_L g3199 ( 
.A(n_2908),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_2719),
.Y(n_3200)
);

AND2x4_ASAP7_75t_L g3201 ( 
.A(n_2680),
.B(n_2899),
.Y(n_3201)
);

A2O1A1Ixp33_ASAP7_75t_L g3202 ( 
.A1(n_3137),
.A2(n_2725),
.B(n_2675),
.C(n_2646),
.Y(n_3202)
);

AOI22xp5_ASAP7_75t_L g3203 ( 
.A1(n_2617),
.A2(n_2606),
.B1(n_3143),
.B2(n_2601),
.Y(n_3203)
);

BUFx4f_ASAP7_75t_L g3204 ( 
.A(n_3092),
.Y(n_3204)
);

NAND2x1p5_ASAP7_75t_L g3205 ( 
.A(n_2592),
.B(n_2902),
.Y(n_3205)
);

AOI22xp33_ASAP7_75t_L g3206 ( 
.A1(n_3143),
.A2(n_3077),
.B1(n_2607),
.B2(n_3129),
.Y(n_3206)
);

CKINVDCx5p33_ASAP7_75t_R g3207 ( 
.A(n_2808),
.Y(n_3207)
);

AND2x2_ASAP7_75t_L g3208 ( 
.A(n_2805),
.B(n_2811),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_2719),
.Y(n_3209)
);

INVx1_ASAP7_75t_SL g3210 ( 
.A(n_2604),
.Y(n_3210)
);

AO31x2_ASAP7_75t_L g3211 ( 
.A1(n_2670),
.A2(n_2676),
.A3(n_3053),
.B(n_3037),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_2759),
.Y(n_3212)
);

OR2x6_ASAP7_75t_L g3213 ( 
.A(n_2807),
.B(n_2977),
.Y(n_3213)
);

INVx2_ASAP7_75t_L g3214 ( 
.A(n_2643),
.Y(n_3214)
);

CKINVDCx11_ASAP7_75t_R g3215 ( 
.A(n_2808),
.Y(n_3215)
);

AOI21xp5_ASAP7_75t_L g3216 ( 
.A1(n_3118),
.A2(n_3127),
.B(n_3122),
.Y(n_3216)
);

BUFx3_ASAP7_75t_L g3217 ( 
.A(n_2969),
.Y(n_3217)
);

OAI22xp5_ASAP7_75t_L g3218 ( 
.A1(n_2687),
.A2(n_2601),
.B1(n_2662),
.B2(n_2815),
.Y(n_3218)
);

INVx2_ASAP7_75t_L g3219 ( 
.A(n_2678),
.Y(n_3219)
);

AOI21xp5_ASAP7_75t_L g3220 ( 
.A1(n_3118),
.A2(n_3127),
.B(n_3122),
.Y(n_3220)
);

INVx3_ASAP7_75t_L g3221 ( 
.A(n_3065),
.Y(n_3221)
);

INVx2_ASAP7_75t_L g3222 ( 
.A(n_2678),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_2759),
.Y(n_3223)
);

HB1xp67_ASAP7_75t_L g3224 ( 
.A(n_2839),
.Y(n_3224)
);

INVx2_ASAP7_75t_L g3225 ( 
.A(n_2678),
.Y(n_3225)
);

OAI21x1_ASAP7_75t_L g3226 ( 
.A1(n_2696),
.A2(n_2620),
.B(n_2590),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_2822),
.Y(n_3227)
);

AOI21xp5_ASAP7_75t_L g3228 ( 
.A1(n_3140),
.A2(n_2613),
.B(n_2602),
.Y(n_3228)
);

BUFx6f_ASAP7_75t_L g3229 ( 
.A(n_2630),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_2822),
.Y(n_3230)
);

INVx2_ASAP7_75t_SL g3231 ( 
.A(n_2665),
.Y(n_3231)
);

BUFx2_ASAP7_75t_SL g3232 ( 
.A(n_2747),
.Y(n_3232)
);

AND2x4_ASAP7_75t_L g3233 ( 
.A(n_2899),
.B(n_2944),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_2828),
.Y(n_3234)
);

OAI22xp5_ASAP7_75t_L g3235 ( 
.A1(n_2687),
.A2(n_2601),
.B1(n_2662),
.B2(n_2815),
.Y(n_3235)
);

INVx5_ASAP7_75t_L g3236 ( 
.A(n_2795),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_SL g3237 ( 
.A(n_2654),
.B(n_2747),
.Y(n_3237)
);

BUFx2_ASAP7_75t_L g3238 ( 
.A(n_2908),
.Y(n_3238)
);

A2O1A1Ixp33_ASAP7_75t_L g3239 ( 
.A1(n_2646),
.A2(n_2654),
.B(n_2710),
.C(n_2779),
.Y(n_3239)
);

OR2x2_ASAP7_75t_SL g3240 ( 
.A(n_2842),
.B(n_2758),
.Y(n_3240)
);

AOI21xp5_ASAP7_75t_L g3241 ( 
.A1(n_3140),
.A2(n_2613),
.B(n_2602),
.Y(n_3241)
);

BUFx2_ASAP7_75t_L g3242 ( 
.A(n_2908),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_SL g3243 ( 
.A(n_2724),
.B(n_2925),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2828),
.Y(n_3244)
);

AND2x4_ASAP7_75t_L g3245 ( 
.A(n_2899),
.B(n_2944),
.Y(n_3245)
);

AOI21xp5_ASAP7_75t_L g3246 ( 
.A1(n_2599),
.A2(n_2610),
.B(n_2626),
.Y(n_3246)
);

BUFx3_ASAP7_75t_L g3247 ( 
.A(n_2871),
.Y(n_3247)
);

AOI21xp5_ASAP7_75t_L g3248 ( 
.A1(n_2599),
.A2(n_2610),
.B(n_2626),
.Y(n_3248)
);

BUFx2_ASAP7_75t_R g3249 ( 
.A(n_3139),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_3072),
.B(n_3109),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_3112),
.B(n_3113),
.Y(n_3251)
);

OR2x2_ASAP7_75t_L g3252 ( 
.A(n_2837),
.B(n_2803),
.Y(n_3252)
);

AND2x2_ASAP7_75t_L g3253 ( 
.A(n_2664),
.B(n_2682),
.Y(n_3253)
);

NOR2xp33_ASAP7_75t_L g3254 ( 
.A(n_3076),
.B(n_3134),
.Y(n_3254)
);

OR2x2_ASAP7_75t_L g3255 ( 
.A(n_2803),
.B(n_2827),
.Y(n_3255)
);

NAND2xp5_ASAP7_75t_L g3256 ( 
.A(n_3112),
.B(n_3113),
.Y(n_3256)
);

AOI21xp5_ASAP7_75t_L g3257 ( 
.A1(n_2649),
.A2(n_2629),
.B(n_2645),
.Y(n_3257)
);

BUFx6f_ASAP7_75t_L g3258 ( 
.A(n_2630),
.Y(n_3258)
);

INVx2_ASAP7_75t_SL g3259 ( 
.A(n_2665),
.Y(n_3259)
);

INVxp67_ASAP7_75t_SL g3260 ( 
.A(n_2959),
.Y(n_3260)
);

OAI22xp5_ASAP7_75t_SL g3261 ( 
.A1(n_2689),
.A2(n_2782),
.B1(n_3049),
.B2(n_2607),
.Y(n_3261)
);

INVx2_ASAP7_75t_L g3262 ( 
.A(n_2818),
.Y(n_3262)
);

BUFx6f_ASAP7_75t_L g3263 ( 
.A(n_2630),
.Y(n_3263)
);

HB1xp67_ASAP7_75t_L g3264 ( 
.A(n_2839),
.Y(n_3264)
);

CKINVDCx20_ASAP7_75t_R g3265 ( 
.A(n_3139),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_2834),
.Y(n_3266)
);

AND2x4_ASAP7_75t_L g3267 ( 
.A(n_2899),
.B(n_2944),
.Y(n_3267)
);

OAI21xp33_ASAP7_75t_L g3268 ( 
.A1(n_2689),
.A2(n_2700),
.B(n_2683),
.Y(n_3268)
);

OAI22xp5_ASAP7_75t_L g3269 ( 
.A1(n_2683),
.A2(n_3067),
.B1(n_2787),
.B2(n_2782),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_3144),
.B(n_2959),
.Y(n_3270)
);

INVx3_ASAP7_75t_L g3271 ( 
.A(n_3065),
.Y(n_3271)
);

BUFx6f_ASAP7_75t_L g3272 ( 
.A(n_2630),
.Y(n_3272)
);

NAND2xp5_ASAP7_75t_L g3273 ( 
.A(n_3144),
.B(n_2905),
.Y(n_3273)
);

BUFx3_ASAP7_75t_L g3274 ( 
.A(n_2871),
.Y(n_3274)
);

BUFx2_ASAP7_75t_L g3275 ( 
.A(n_2908),
.Y(n_3275)
);

OAI22xp5_ASAP7_75t_L g3276 ( 
.A1(n_3067),
.A2(n_2787),
.B1(n_2859),
.B2(n_2819),
.Y(n_3276)
);

AND2x2_ASAP7_75t_L g3277 ( 
.A(n_2664),
.B(n_2682),
.Y(n_3277)
);

OAI22xp5_ASAP7_75t_L g3278 ( 
.A1(n_3067),
.A2(n_2859),
.B1(n_2819),
.B2(n_2641),
.Y(n_3278)
);

NOR2xp67_ASAP7_75t_SL g3279 ( 
.A(n_2816),
.B(n_3064),
.Y(n_3279)
);

INVxp67_ASAP7_75t_SL g3280 ( 
.A(n_2710),
.Y(n_3280)
);

OR2x2_ASAP7_75t_L g3281 ( 
.A(n_2803),
.B(n_2827),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_L g3282 ( 
.A(n_2905),
.B(n_2708),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_2834),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_2838),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_2838),
.Y(n_3285)
);

AND2x4_ASAP7_75t_L g3286 ( 
.A(n_2944),
.B(n_2903),
.Y(n_3286)
);

AOI22xp33_ASAP7_75t_L g3287 ( 
.A1(n_3077),
.A2(n_2670),
.B1(n_3067),
.B2(n_2635),
.Y(n_3287)
);

INVx2_ASAP7_75t_L g3288 ( 
.A(n_2818),
.Y(n_3288)
);

BUFx6f_ASAP7_75t_L g3289 ( 
.A(n_2630),
.Y(n_3289)
);

AOI21xp5_ASAP7_75t_L g3290 ( 
.A1(n_2649),
.A2(n_2629),
.B(n_2645),
.Y(n_3290)
);

AOI21xp5_ASAP7_75t_L g3291 ( 
.A1(n_2666),
.A2(n_2843),
.B(n_2826),
.Y(n_3291)
);

INVx1_ASAP7_75t_SL g3292 ( 
.A(n_2604),
.Y(n_3292)
);

AND2x2_ASAP7_75t_L g3293 ( 
.A(n_2887),
.B(n_2812),
.Y(n_3293)
);

AOI21xp5_ASAP7_75t_L g3294 ( 
.A1(n_2666),
.A2(n_2843),
.B(n_2826),
.Y(n_3294)
);

AND2x2_ASAP7_75t_L g3295 ( 
.A(n_2887),
.B(n_2812),
.Y(n_3295)
);

BUFx2_ASAP7_75t_L g3296 ( 
.A(n_2908),
.Y(n_3296)
);

HB1xp67_ASAP7_75t_L g3297 ( 
.A(n_2874),
.Y(n_3297)
);

OAI22xp5_ASAP7_75t_L g3298 ( 
.A1(n_3067),
.A2(n_3068),
.B1(n_2739),
.B2(n_2810),
.Y(n_3298)
);

AND2x4_ASAP7_75t_L g3299 ( 
.A(n_2903),
.B(n_2589),
.Y(n_3299)
);

CKINVDCx6p67_ASAP7_75t_R g3300 ( 
.A(n_3139),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_L g3301 ( 
.A(n_2708),
.B(n_2723),
.Y(n_3301)
);

AND2x2_ASAP7_75t_L g3302 ( 
.A(n_2628),
.B(n_2653),
.Y(n_3302)
);

AOI21x1_ASAP7_75t_L g3303 ( 
.A1(n_2590),
.A2(n_3085),
.B(n_2620),
.Y(n_3303)
);

INVx2_ASAP7_75t_SL g3304 ( 
.A(n_2665),
.Y(n_3304)
);

OAI21xp5_ASAP7_75t_L g3305 ( 
.A1(n_3082),
.A2(n_2627),
.B(n_2731),
.Y(n_3305)
);

A2O1A1Ixp33_ASAP7_75t_SL g3306 ( 
.A1(n_2700),
.A2(n_2739),
.B(n_2942),
.C(n_2676),
.Y(n_3306)
);

BUFx3_ASAP7_75t_L g3307 ( 
.A(n_2871),
.Y(n_3307)
);

BUFx2_ASAP7_75t_L g3308 ( 
.A(n_2908),
.Y(n_3308)
);

INVx2_ASAP7_75t_L g3309 ( 
.A(n_2833),
.Y(n_3309)
);

OR2x6_ASAP7_75t_SL g3310 ( 
.A(n_2930),
.B(n_2806),
.Y(n_3310)
);

NOR2xp33_ASAP7_75t_L g3311 ( 
.A(n_2674),
.B(n_2618),
.Y(n_3311)
);

OR2x6_ASAP7_75t_L g3312 ( 
.A(n_2977),
.B(n_2795),
.Y(n_3312)
);

OR2x2_ASAP7_75t_SL g3313 ( 
.A(n_2842),
.B(n_2758),
.Y(n_3313)
);

BUFx2_ASAP7_75t_L g3314 ( 
.A(n_2908),
.Y(n_3314)
);

AOI21xp5_ASAP7_75t_L g3315 ( 
.A1(n_2596),
.A2(n_3049),
.B(n_2597),
.Y(n_3315)
);

OAI22xp5_ASAP7_75t_L g3316 ( 
.A1(n_3068),
.A2(n_2810),
.B1(n_2802),
.B2(n_2748),
.Y(n_3316)
);

INVxp67_ASAP7_75t_L g3317 ( 
.A(n_2821),
.Y(n_3317)
);

NOR2xp33_ASAP7_75t_L g3318 ( 
.A(n_2598),
.B(n_3128),
.Y(n_3318)
);

INVxp67_ASAP7_75t_SL g3319 ( 
.A(n_2830),
.Y(n_3319)
);

A2O1A1Ixp33_ASAP7_75t_SL g3320 ( 
.A1(n_2748),
.A2(n_2911),
.B(n_2740),
.C(n_2728),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_2723),
.B(n_2726),
.Y(n_3321)
);

O2A1O1Ixp33_ASAP7_75t_L g3322 ( 
.A1(n_2635),
.A2(n_2672),
.B(n_3066),
.C(n_3133),
.Y(n_3322)
);

BUFx5_ASAP7_75t_L g3323 ( 
.A(n_3077),
.Y(n_3323)
);

INVx3_ASAP7_75t_L g3324 ( 
.A(n_3065),
.Y(n_3324)
);

AND2x4_ASAP7_75t_L g3325 ( 
.A(n_2903),
.B(n_2589),
.Y(n_3325)
);

CKINVDCx5p33_ASAP7_75t_R g3326 ( 
.A(n_2707),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_2857),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_2857),
.Y(n_3328)
);

AND2x2_ASAP7_75t_L g3329 ( 
.A(n_2628),
.B(n_2653),
.Y(n_3329)
);

OAI22xp5_ASAP7_75t_L g3330 ( 
.A1(n_2849),
.A2(n_2814),
.B1(n_2854),
.B2(n_2809),
.Y(n_3330)
);

CKINVDCx8_ASAP7_75t_R g3331 ( 
.A(n_3014),
.Y(n_3331)
);

BUFx2_ASAP7_75t_L g3332 ( 
.A(n_2762),
.Y(n_3332)
);

AND2x2_ASAP7_75t_L g3333 ( 
.A(n_3103),
.B(n_3080),
.Y(n_3333)
);

A2O1A1Ixp33_ASAP7_75t_L g3334 ( 
.A1(n_2779),
.A2(n_2667),
.B(n_2783),
.C(n_2688),
.Y(n_3334)
);

BUFx2_ASAP7_75t_L g3335 ( 
.A(n_2762),
.Y(n_3335)
);

INVx2_ASAP7_75t_L g3336 ( 
.A(n_2833),
.Y(n_3336)
);

OAI22xp5_ASAP7_75t_L g3337 ( 
.A1(n_2849),
.A2(n_2814),
.B1(n_2854),
.B2(n_2809),
.Y(n_3337)
);

NOR2xp33_ASAP7_75t_SL g3338 ( 
.A(n_2672),
.B(n_2771),
.Y(n_3338)
);

CKINVDCx20_ASAP7_75t_R g3339 ( 
.A(n_2901),
.Y(n_3339)
);

AOI21xp5_ASAP7_75t_L g3340 ( 
.A1(n_2596),
.A2(n_2597),
.B(n_2600),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_L g3341 ( 
.A(n_2726),
.B(n_2730),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_2868),
.Y(n_3342)
);

INVx2_ASAP7_75t_L g3343 ( 
.A(n_2845),
.Y(n_3343)
);

INVx2_ASAP7_75t_SL g3344 ( 
.A(n_2762),
.Y(n_3344)
);

OAI22xp5_ASAP7_75t_L g3345 ( 
.A1(n_2806),
.A2(n_2667),
.B1(n_3066),
.B2(n_3053),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_2868),
.Y(n_3346)
);

OAI21xp33_ASAP7_75t_SL g3347 ( 
.A1(n_2855),
.A2(n_2877),
.B(n_2702),
.Y(n_3347)
);

O2A1O1Ixp5_ASAP7_75t_L g3348 ( 
.A1(n_2783),
.A2(n_2688),
.B(n_2740),
.C(n_2786),
.Y(n_3348)
);

INVx2_ASAP7_75t_L g3349 ( 
.A(n_2845),
.Y(n_3349)
);

BUFx3_ASAP7_75t_L g3350 ( 
.A(n_2744),
.Y(n_3350)
);

INVx3_ASAP7_75t_L g3351 ( 
.A(n_2630),
.Y(n_3351)
);

BUFx6f_ASAP7_75t_L g3352 ( 
.A(n_2633),
.Y(n_3352)
);

AND2x4_ASAP7_75t_L g3353 ( 
.A(n_2903),
.B(n_2589),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_L g3354 ( 
.A(n_2730),
.B(n_2733),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_2733),
.B(n_2736),
.Y(n_3355)
);

INVx2_ASAP7_75t_L g3356 ( 
.A(n_2845),
.Y(n_3356)
);

NAND2xp5_ASAP7_75t_SL g3357 ( 
.A(n_2925),
.B(n_2853),
.Y(n_3357)
);

BUFx10_ASAP7_75t_L g3358 ( 
.A(n_2932),
.Y(n_3358)
);

INVx2_ASAP7_75t_L g3359 ( 
.A(n_2884),
.Y(n_3359)
);

INVx3_ASAP7_75t_L g3360 ( 
.A(n_2633),
.Y(n_3360)
);

A2O1A1Ixp33_ASAP7_75t_L g3361 ( 
.A1(n_2846),
.A2(n_3034),
.B(n_2801),
.C(n_2766),
.Y(n_3361)
);

INVx2_ASAP7_75t_SL g3362 ( 
.A(n_2863),
.Y(n_3362)
);

NAND2x1p5_ASAP7_75t_L g3363 ( 
.A(n_2592),
.B(n_2902),
.Y(n_3363)
);

NOR2x1_ASAP7_75t_SL g3364 ( 
.A(n_2795),
.B(n_2930),
.Y(n_3364)
);

INVx8_ASAP7_75t_L g3365 ( 
.A(n_2902),
.Y(n_3365)
);

INVxp67_ASAP7_75t_SL g3366 ( 
.A(n_2830),
.Y(n_3366)
);

AND2x4_ASAP7_75t_L g3367 ( 
.A(n_2903),
.B(n_2589),
.Y(n_3367)
);

AND2x2_ASAP7_75t_L g3368 ( 
.A(n_3103),
.B(n_3080),
.Y(n_3368)
);

OAI22xp5_ASAP7_75t_L g3369 ( 
.A1(n_3037),
.A2(n_2879),
.B1(n_2882),
.B2(n_2855),
.Y(n_3369)
);

OAI22xp5_ASAP7_75t_L g3370 ( 
.A1(n_2882),
.A2(n_2855),
.B1(n_3028),
.B2(n_2758),
.Y(n_3370)
);

OAI21x1_ASAP7_75t_L g3371 ( 
.A1(n_2696),
.A2(n_3085),
.B(n_2673),
.Y(n_3371)
);

NOR2xp33_ASAP7_75t_L g3372 ( 
.A(n_2639),
.B(n_2713),
.Y(n_3372)
);

INVx1_ASAP7_75t_L g3373 ( 
.A(n_2611),
.Y(n_3373)
);

AND2x2_ASAP7_75t_L g3374 ( 
.A(n_3080),
.B(n_2803),
.Y(n_3374)
);

OR2x2_ASAP7_75t_L g3375 ( 
.A(n_2803),
.B(n_2684),
.Y(n_3375)
);

AOI21x1_ASAP7_75t_L g3376 ( 
.A1(n_2655),
.A2(n_2781),
.B(n_3057),
.Y(n_3376)
);

NOR2xp33_ASAP7_75t_L g3377 ( 
.A(n_2715),
.B(n_2914),
.Y(n_3377)
);

AOI21xp33_ASAP7_75t_SL g3378 ( 
.A1(n_3032),
.A2(n_2998),
.B(n_2751),
.Y(n_3378)
);

BUFx2_ASAP7_75t_L g3379 ( 
.A(n_2863),
.Y(n_3379)
);

NAND2xp5_ASAP7_75t_L g3380 ( 
.A(n_2736),
.B(n_2743),
.Y(n_3380)
);

AND2x2_ASAP7_75t_L g3381 ( 
.A(n_3080),
.B(n_2803),
.Y(n_3381)
);

AOI21xp5_ASAP7_75t_L g3382 ( 
.A1(n_2596),
.A2(n_2597),
.B(n_2600),
.Y(n_3382)
);

AND2x4_ASAP7_75t_SL g3383 ( 
.A(n_2795),
.B(n_2937),
.Y(n_3383)
);

CKINVDCx5p33_ASAP7_75t_R g3384 ( 
.A(n_2707),
.Y(n_3384)
);

INVxp67_ASAP7_75t_SL g3385 ( 
.A(n_2830),
.Y(n_3385)
);

AOI21xp5_ASAP7_75t_L g3386 ( 
.A1(n_2600),
.A2(n_2595),
.B(n_3138),
.Y(n_3386)
);

AOI21xp5_ASAP7_75t_L g3387 ( 
.A1(n_2595),
.A2(n_3138),
.B(n_2669),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_2611),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_2619),
.Y(n_3389)
);

BUFx12f_ASAP7_75t_L g3390 ( 
.A(n_2707),
.Y(n_3390)
);

AOI21xp5_ASAP7_75t_L g3391 ( 
.A1(n_2595),
.A2(n_3138),
.B(n_2669),
.Y(n_3391)
);

INVx2_ASAP7_75t_L g3392 ( 
.A(n_2884),
.Y(n_3392)
);

AOI21xp5_ASAP7_75t_L g3393 ( 
.A1(n_3138),
.A2(n_2669),
.B(n_2660),
.Y(n_3393)
);

AND2x4_ASAP7_75t_L g3394 ( 
.A(n_2903),
.B(n_3100),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_L g3395 ( 
.A(n_2743),
.B(n_2745),
.Y(n_3395)
);

HB1xp67_ASAP7_75t_L g3396 ( 
.A(n_2648),
.Y(n_3396)
);

AND2x4_ASAP7_75t_L g3397 ( 
.A(n_3100),
.B(n_2829),
.Y(n_3397)
);

NOR2xp33_ASAP7_75t_L g3398 ( 
.A(n_2657),
.B(n_2659),
.Y(n_3398)
);

NAND2xp33_ASAP7_75t_L g3399 ( 
.A(n_3032),
.B(n_3077),
.Y(n_3399)
);

INVx3_ASAP7_75t_L g3400 ( 
.A(n_2633),
.Y(n_3400)
);

BUFx3_ASAP7_75t_L g3401 ( 
.A(n_2744),
.Y(n_3401)
);

BUFx3_ASAP7_75t_L g3402 ( 
.A(n_2744),
.Y(n_3402)
);

AND2x4_ASAP7_75t_L g3403 ( 
.A(n_3100),
.B(n_2829),
.Y(n_3403)
);

OR2x2_ASAP7_75t_L g3404 ( 
.A(n_2684),
.B(n_2693),
.Y(n_3404)
);

AND2x4_ASAP7_75t_L g3405 ( 
.A(n_3100),
.B(n_2877),
.Y(n_3405)
);

AOI22xp33_ASAP7_75t_L g3406 ( 
.A1(n_3077),
.A2(n_2751),
.B1(n_2737),
.B2(n_2877),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_2745),
.B(n_2746),
.Y(n_3407)
);

INVx4_ASAP7_75t_L g3408 ( 
.A(n_2902),
.Y(n_3408)
);

AOI21xp5_ASAP7_75t_L g3409 ( 
.A1(n_2660),
.A2(n_2638),
.B(n_2640),
.Y(n_3409)
);

AOI21xp5_ASAP7_75t_L g3410 ( 
.A1(n_2660),
.A2(n_2638),
.B(n_2640),
.Y(n_3410)
);

INVx5_ASAP7_75t_L g3411 ( 
.A(n_2699),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_L g3412 ( 
.A(n_2746),
.B(n_2749),
.Y(n_3412)
);

INVx3_ASAP7_75t_SL g3413 ( 
.A(n_2980),
.Y(n_3413)
);

INVx2_ASAP7_75t_L g3414 ( 
.A(n_2884),
.Y(n_3414)
);

OR2x6_ASAP7_75t_L g3415 ( 
.A(n_2977),
.B(n_2954),
.Y(n_3415)
);

INVx3_ASAP7_75t_L g3416 ( 
.A(n_2633),
.Y(n_3416)
);

INVx5_ASAP7_75t_L g3417 ( 
.A(n_2699),
.Y(n_3417)
);

AND2x4_ASAP7_75t_L g3418 ( 
.A(n_2921),
.B(n_2928),
.Y(n_3418)
);

OAI22xp5_ASAP7_75t_L g3419 ( 
.A1(n_3028),
.A2(n_2758),
.B1(n_2831),
.B2(n_2659),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_2749),
.B(n_2750),
.Y(n_3420)
);

AOI21xp5_ASAP7_75t_L g3421 ( 
.A1(n_2638),
.A2(n_2640),
.B(n_2644),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_L g3422 ( 
.A(n_2750),
.B(n_2757),
.Y(n_3422)
);

CKINVDCx16_ASAP7_75t_R g3423 ( 
.A(n_2671),
.Y(n_3423)
);

AOI22xp5_ASAP7_75t_L g3424 ( 
.A1(n_3077),
.A2(n_2846),
.B1(n_2737),
.B2(n_2758),
.Y(n_3424)
);

AOI21xp5_ASAP7_75t_L g3425 ( 
.A1(n_2644),
.A2(n_2658),
.B(n_3070),
.Y(n_3425)
);

OAI22xp5_ASAP7_75t_L g3426 ( 
.A1(n_2831),
.A2(n_2657),
.B1(n_2768),
.B2(n_2757),
.Y(n_3426)
);

INVx5_ASAP7_75t_L g3427 ( 
.A(n_2699),
.Y(n_3427)
);

A2O1A1Ixp33_ASAP7_75t_L g3428 ( 
.A1(n_3034),
.A2(n_2801),
.B(n_2766),
.C(n_2753),
.Y(n_3428)
);

BUFx3_ASAP7_75t_L g3429 ( 
.A(n_2744),
.Y(n_3429)
);

AO21x2_ASAP7_75t_L g3430 ( 
.A1(n_2753),
.A2(n_2786),
.B(n_3063),
.Y(n_3430)
);

BUFx2_ASAP7_75t_L g3431 ( 
.A(n_2863),
.Y(n_3431)
);

INVx4_ASAP7_75t_L g3432 ( 
.A(n_2902),
.Y(n_3432)
);

INVx2_ASAP7_75t_L g3433 ( 
.A(n_2922),
.Y(n_3433)
);

BUFx2_ASAP7_75t_L g3434 ( 
.A(n_2946),
.Y(n_3434)
);

AND2x4_ASAP7_75t_L g3435 ( 
.A(n_2921),
.B(n_2928),
.Y(n_3435)
);

OR2x6_ASAP7_75t_L g3436 ( 
.A(n_2977),
.B(n_2954),
.Y(n_3436)
);

INVxp67_ASAP7_75t_SL g3437 ( 
.A(n_2830),
.Y(n_3437)
);

INVx2_ASAP7_75t_L g3438 ( 
.A(n_2922),
.Y(n_3438)
);

INVx2_ASAP7_75t_SL g3439 ( 
.A(n_2946),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_2768),
.B(n_2769),
.Y(n_3440)
);

AND2x4_ASAP7_75t_L g3441 ( 
.A(n_2952),
.B(n_2953),
.Y(n_3441)
);

INVx2_ASAP7_75t_SL g3442 ( 
.A(n_2946),
.Y(n_3442)
);

INVx2_ASAP7_75t_L g3443 ( 
.A(n_2922),
.Y(n_3443)
);

O2A1O1Ixp33_ASAP7_75t_L g3444 ( 
.A1(n_2771),
.A2(n_2821),
.B(n_2860),
.C(n_2627),
.Y(n_3444)
);

AND2x4_ASAP7_75t_L g3445 ( 
.A(n_2952),
.B(n_2953),
.Y(n_3445)
);

INVx2_ASAP7_75t_L g3446 ( 
.A(n_2929),
.Y(n_3446)
);

CKINVDCx6p67_ASAP7_75t_R g3447 ( 
.A(n_2980),
.Y(n_3447)
);

AND2x2_ASAP7_75t_L g3448 ( 
.A(n_3080),
.B(n_2995),
.Y(n_3448)
);

OR2x6_ASAP7_75t_L g3449 ( 
.A(n_2954),
.B(n_2721),
.Y(n_3449)
);

AO21x1_ASAP7_75t_L g3450 ( 
.A1(n_2860),
.A2(n_3031),
.B(n_2906),
.Y(n_3450)
);

INVx1_ASAP7_75t_SL g3451 ( 
.A(n_2648),
.Y(n_3451)
);

BUFx2_ASAP7_75t_L g3452 ( 
.A(n_2671),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_2769),
.B(n_2817),
.Y(n_3453)
);

NOR2xp33_ASAP7_75t_L g3454 ( 
.A(n_2668),
.B(n_2685),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_3141),
.Y(n_3455)
);

INVx5_ASAP7_75t_L g3456 ( 
.A(n_2699),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_SL g3457 ( 
.A(n_2825),
.B(n_2965),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_2861),
.Y(n_3458)
);

INVx3_ASAP7_75t_L g3459 ( 
.A(n_2633),
.Y(n_3459)
);

INVx2_ASAP7_75t_L g3460 ( 
.A(n_2929),
.Y(n_3460)
);

OAI22xp5_ASAP7_75t_L g3461 ( 
.A1(n_2668),
.A2(n_2685),
.B1(n_2778),
.B2(n_2777),
.Y(n_3461)
);

NOR2xp33_ASAP7_75t_L g3462 ( 
.A(n_2651),
.B(n_2652),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_2861),
.Y(n_3463)
);

HB1xp67_ASAP7_75t_L g3464 ( 
.A(n_3101),
.Y(n_3464)
);

A2O1A1Ixp33_ASAP7_75t_L g3465 ( 
.A1(n_2965),
.A2(n_2764),
.B(n_2711),
.C(n_2867),
.Y(n_3465)
);

AOI21xp5_ASAP7_75t_L g3466 ( 
.A1(n_2644),
.A2(n_2658),
.B(n_3070),
.Y(n_3466)
);

BUFx3_ASAP7_75t_L g3467 ( 
.A(n_2671),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_2945),
.Y(n_3468)
);

CKINVDCx5p33_ASAP7_75t_R g3469 ( 
.A(n_3101),
.Y(n_3469)
);

AND2x4_ASAP7_75t_L g3470 ( 
.A(n_2594),
.B(n_2709),
.Y(n_3470)
);

NAND2x1p5_ASAP7_75t_L g3471 ( 
.A(n_2592),
.B(n_2902),
.Y(n_3471)
);

OAI31xp33_ASAP7_75t_L g3472 ( 
.A1(n_2912),
.A2(n_3031),
.A3(n_3077),
.B(n_2731),
.Y(n_3472)
);

NOR2xp33_ASAP7_75t_L g3473 ( 
.A(n_2651),
.B(n_2652),
.Y(n_3473)
);

AOI21xp5_ASAP7_75t_L g3474 ( 
.A1(n_2658),
.A2(n_3073),
.B(n_3070),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_L g3475 ( 
.A(n_2817),
.B(n_2777),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_2945),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_2778),
.B(n_2790),
.Y(n_3477)
);

BUFx6f_ASAP7_75t_L g3478 ( 
.A(n_2633),
.Y(n_3478)
);

O2A1O1Ixp33_ASAP7_75t_L g3479 ( 
.A1(n_2706),
.A2(n_2691),
.B(n_2764),
.C(n_2906),
.Y(n_3479)
);

BUFx3_ASAP7_75t_L g3480 ( 
.A(n_2694),
.Y(n_3480)
);

CKINVDCx8_ASAP7_75t_R g3481 ( 
.A(n_3014),
.Y(n_3481)
);

OAI21x1_ASAP7_75t_L g3482 ( 
.A1(n_2696),
.A2(n_2673),
.B(n_2655),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_L g3483 ( 
.A(n_2790),
.B(n_2793),
.Y(n_3483)
);

BUFx2_ASAP7_75t_L g3484 ( 
.A(n_2694),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_L g3485 ( 
.A(n_2793),
.B(n_2796),
.Y(n_3485)
);

NOR2xp67_ASAP7_75t_SL g3486 ( 
.A(n_2694),
.B(n_2902),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_2964),
.Y(n_3487)
);

BUFx6f_ASAP7_75t_L g3488 ( 
.A(n_2663),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_L g3489 ( 
.A(n_2796),
.B(n_2800),
.Y(n_3489)
);

CKINVDCx20_ASAP7_75t_R g3490 ( 
.A(n_3009),
.Y(n_3490)
);

CKINVDCx16_ASAP7_75t_R g3491 ( 
.A(n_3009),
.Y(n_3491)
);

OA21x2_ASAP7_75t_L g3492 ( 
.A1(n_2636),
.A2(n_2673),
.B(n_2624),
.Y(n_3492)
);

AOI21xp5_ASAP7_75t_L g3493 ( 
.A1(n_3073),
.A2(n_3087),
.B(n_3083),
.Y(n_3493)
);

AND2x2_ASAP7_75t_L g3494 ( 
.A(n_3080),
.B(n_2995),
.Y(n_3494)
);

AND2x4_ASAP7_75t_L g3495 ( 
.A(n_2594),
.B(n_2709),
.Y(n_3495)
);

AND2x2_ASAP7_75t_L g3496 ( 
.A(n_3080),
.B(n_2979),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_2800),
.B(n_2701),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_2701),
.B(n_2703),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_SL g3499 ( 
.A(n_2936),
.B(n_2898),
.Y(n_3499)
);

BUFx2_ASAP7_75t_L g3500 ( 
.A(n_2975),
.Y(n_3500)
);

AND2x2_ASAP7_75t_L g3501 ( 
.A(n_2979),
.B(n_2754),
.Y(n_3501)
);

AND2x2_ASAP7_75t_L g3502 ( 
.A(n_2754),
.B(n_2974),
.Y(n_3502)
);

OR2x2_ASAP7_75t_L g3503 ( 
.A(n_2693),
.B(n_3096),
.Y(n_3503)
);

BUFx2_ASAP7_75t_L g3504 ( 
.A(n_2975),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_2703),
.B(n_2729),
.Y(n_3505)
);

OAI22xp33_ASAP7_75t_L g3506 ( 
.A1(n_2851),
.A2(n_2990),
.B1(n_3019),
.B2(n_2592),
.Y(n_3506)
);

AND2x4_ASAP7_75t_L g3507 ( 
.A(n_2594),
.B(n_2709),
.Y(n_3507)
);

OAI22xp5_ASAP7_75t_L g3508 ( 
.A1(n_2695),
.A2(n_2697),
.B1(n_2634),
.B2(n_2642),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_L g3509 ( 
.A(n_2775),
.B(n_2872),
.Y(n_3509)
);

INVx2_ASAP7_75t_SL g3510 ( 
.A(n_2732),
.Y(n_3510)
);

INVx6_ASAP7_75t_L g3511 ( 
.A(n_2937),
.Y(n_3511)
);

AND2x4_ASAP7_75t_L g3512 ( 
.A(n_3131),
.B(n_3047),
.Y(n_3512)
);

BUFx4_ASAP7_75t_SL g3513 ( 
.A(n_3009),
.Y(n_3513)
);

NAND2x1p5_ASAP7_75t_L g3514 ( 
.A(n_2858),
.B(n_2721),
.Y(n_3514)
);

HB1xp67_ASAP7_75t_L g3515 ( 
.A(n_2870),
.Y(n_3515)
);

INVx3_ASAP7_75t_L g3516 ( 
.A(n_2663),
.Y(n_3516)
);

CKINVDCx20_ASAP7_75t_R g3517 ( 
.A(n_3038),
.Y(n_3517)
);

BUFx3_ASAP7_75t_L g3518 ( 
.A(n_2732),
.Y(n_3518)
);

OR2x6_ASAP7_75t_L g3519 ( 
.A(n_2637),
.B(n_2720),
.Y(n_3519)
);

INVx1_ASAP7_75t_SL g3520 ( 
.A(n_2742),
.Y(n_3520)
);

OAI22xp5_ASAP7_75t_L g3521 ( 
.A1(n_2695),
.A2(n_2697),
.B1(n_2634),
.B2(n_2642),
.Y(n_3521)
);

NOR2xp67_ASAP7_75t_SL g3522 ( 
.A(n_3038),
.B(n_2932),
.Y(n_3522)
);

O2A1O1Ixp33_ASAP7_75t_L g3523 ( 
.A1(n_2706),
.A2(n_2691),
.B(n_2900),
.C(n_2847),
.Y(n_3523)
);

NAND2xp5_ASAP7_75t_SL g3524 ( 
.A(n_2936),
.B(n_2836),
.Y(n_3524)
);

AND2x2_ASAP7_75t_L g3525 ( 
.A(n_2754),
.B(n_2974),
.Y(n_3525)
);

OAI22xp5_ASAP7_75t_L g3526 ( 
.A1(n_2631),
.A2(n_2650),
.B1(n_2891),
.B2(n_2841),
.Y(n_3526)
);

OR2x2_ASAP7_75t_L g3527 ( 
.A(n_3096),
.B(n_2910),
.Y(n_3527)
);

INVx2_ASAP7_75t_L g3528 ( 
.A(n_2967),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_2872),
.B(n_2883),
.Y(n_3529)
);

INVx2_ASAP7_75t_SL g3530 ( 
.A(n_2742),
.Y(n_3530)
);

AOI22xp33_ASAP7_75t_L g3531 ( 
.A1(n_3077),
.A2(n_2990),
.B1(n_3019),
.B2(n_2692),
.Y(n_3531)
);

AOI22xp33_ASAP7_75t_L g3532 ( 
.A1(n_2692),
.A2(n_2637),
.B1(n_3121),
.B2(n_2720),
.Y(n_3532)
);

OAI22xp5_ASAP7_75t_L g3533 ( 
.A1(n_2631),
.A2(n_2650),
.B1(n_2891),
.B2(n_2841),
.Y(n_3533)
);

AOI21xp5_ASAP7_75t_L g3534 ( 
.A1(n_3073),
.A2(n_3087),
.B(n_3083),
.Y(n_3534)
);

INVx3_ASAP7_75t_L g3535 ( 
.A(n_2663),
.Y(n_3535)
);

INVx2_ASAP7_75t_L g3536 ( 
.A(n_2967),
.Y(n_3536)
);

AND2x2_ASAP7_75t_L g3537 ( 
.A(n_2754),
.B(n_2978),
.Y(n_3537)
);

OAI22xp5_ASAP7_75t_L g3538 ( 
.A1(n_2824),
.A2(n_3013),
.B1(n_2704),
.B2(n_2705),
.Y(n_3538)
);

INVxp67_ASAP7_75t_L g3539 ( 
.A(n_2761),
.Y(n_3539)
);

BUFx6f_ASAP7_75t_L g3540 ( 
.A(n_2663),
.Y(n_3540)
);

INVx2_ASAP7_75t_L g3541 ( 
.A(n_2967),
.Y(n_3541)
);

NOR2x1_ASAP7_75t_SL g3542 ( 
.A(n_2988),
.B(n_2858),
.Y(n_3542)
);

AND2x2_ASAP7_75t_L g3543 ( 
.A(n_2754),
.B(n_2978),
.Y(n_3543)
);

NOR2xp67_ASAP7_75t_L g3544 ( 
.A(n_2916),
.B(n_3057),
.Y(n_3544)
);

OR2x6_ASAP7_75t_L g3545 ( 
.A(n_3121),
.B(n_2621),
.Y(n_3545)
);

BUFx12f_ASAP7_75t_L g3546 ( 
.A(n_2937),
.Y(n_3546)
);

AOI21xp5_ASAP7_75t_L g3547 ( 
.A1(n_3083),
.A2(n_3093),
.B(n_3087),
.Y(n_3547)
);

INVx6_ASAP7_75t_L g3548 ( 
.A(n_2937),
.Y(n_3548)
);

AND2x2_ASAP7_75t_L g3549 ( 
.A(n_2754),
.B(n_2994),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_2883),
.B(n_2941),
.Y(n_3550)
);

AND2x2_ASAP7_75t_L g3551 ( 
.A(n_2754),
.B(n_2994),
.Y(n_3551)
);

HB1xp67_ASAP7_75t_L g3552 ( 
.A(n_2870),
.Y(n_3552)
);

HB1xp67_ASAP7_75t_L g3553 ( 
.A(n_2886),
.Y(n_3553)
);

INVx1_ASAP7_75t_SL g3554 ( 
.A(n_2761),
.Y(n_3554)
);

HB1xp67_ASAP7_75t_L g3555 ( 
.A(n_2886),
.Y(n_3555)
);

OR2x2_ASAP7_75t_L g3556 ( 
.A(n_2910),
.B(n_2939),
.Y(n_3556)
);

O2A1O1Ixp5_ASAP7_75t_L g3557 ( 
.A1(n_2760),
.A2(n_2752),
.B(n_2918),
.C(n_2797),
.Y(n_3557)
);

AND2x2_ASAP7_75t_L g3558 ( 
.A(n_2999),
.B(n_2763),
.Y(n_3558)
);

INVx5_ASAP7_75t_L g3559 ( 
.A(n_2663),
.Y(n_3559)
);

AND2x2_ASAP7_75t_L g3560 ( 
.A(n_2999),
.B(n_2763),
.Y(n_3560)
);

BUFx3_ASAP7_75t_L g3561 ( 
.A(n_2776),
.Y(n_3561)
);

BUFx12f_ASAP7_75t_L g3562 ( 
.A(n_3038),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_2972),
.Y(n_3563)
);

AND2x4_ASAP7_75t_L g3564 ( 
.A(n_3131),
.B(n_3047),
.Y(n_3564)
);

A2O1A1Ixp33_ASAP7_75t_L g3565 ( 
.A1(n_2711),
.A2(n_2760),
.B(n_2712),
.C(n_2788),
.Y(n_3565)
);

OAI22xp5_ASAP7_75t_L g3566 ( 
.A1(n_2824),
.A2(n_3013),
.B1(n_2704),
.B2(n_2705),
.Y(n_3566)
);

OR2x6_ASAP7_75t_L g3567 ( 
.A(n_2621),
.B(n_2752),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_2941),
.B(n_2951),
.Y(n_3568)
);

AND2x2_ASAP7_75t_L g3569 ( 
.A(n_2776),
.B(n_2792),
.Y(n_3569)
);

INVx3_ASAP7_75t_SL g3570 ( 
.A(n_2980),
.Y(n_3570)
);

AOI21xp5_ASAP7_75t_L g3571 ( 
.A1(n_3093),
.A2(n_3105),
.B(n_3094),
.Y(n_3571)
);

AND2x4_ASAP7_75t_L g3572 ( 
.A(n_3131),
.B(n_3047),
.Y(n_3572)
);

INVx6_ASAP7_75t_L g3573 ( 
.A(n_2932),
.Y(n_3573)
);

INVx2_ASAP7_75t_L g3574 ( 
.A(n_2976),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_L g3575 ( 
.A(n_2951),
.B(n_2956),
.Y(n_3575)
);

AND2x2_ASAP7_75t_L g3576 ( 
.A(n_2792),
.B(n_2962),
.Y(n_3576)
);

AND2x4_ASAP7_75t_L g3577 ( 
.A(n_3047),
.B(n_2955),
.Y(n_3577)
);

BUFx10_ASAP7_75t_L g3578 ( 
.A(n_2932),
.Y(n_3578)
);

AO21x1_ASAP7_75t_L g3579 ( 
.A1(n_2711),
.A2(n_3063),
.B(n_3069),
.Y(n_3579)
);

AOI21xp5_ASAP7_75t_L g3580 ( 
.A1(n_3093),
.A2(n_3105),
.B(n_3094),
.Y(n_3580)
);

INVx2_ASAP7_75t_L g3581 ( 
.A(n_2976),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_2956),
.B(n_2957),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_2957),
.B(n_2961),
.Y(n_3583)
);

AND2x4_ASAP7_75t_L g3584 ( 
.A(n_2955),
.B(n_3030),
.Y(n_3584)
);

NAND2xp5_ASAP7_75t_SL g3585 ( 
.A(n_2836),
.B(n_2844),
.Y(n_3585)
);

AOI21xp5_ASAP7_75t_L g3586 ( 
.A1(n_3094),
.A2(n_3106),
.B(n_3105),
.Y(n_3586)
);

AOI22xp33_ASAP7_75t_L g3587 ( 
.A1(n_2692),
.A2(n_2789),
.B1(n_2955),
.B2(n_2916),
.Y(n_3587)
);

AND2x4_ASAP7_75t_L g3588 ( 
.A(n_3030),
.B(n_2950),
.Y(n_3588)
);

INVx3_ASAP7_75t_L g3589 ( 
.A(n_2663),
.Y(n_3589)
);

AND2x4_ASAP7_75t_L g3590 ( 
.A(n_3030),
.B(n_2950),
.Y(n_3590)
);

INVx2_ASAP7_75t_L g3591 ( 
.A(n_2976),
.Y(n_3591)
);

INVx2_ASAP7_75t_SL g3592 ( 
.A(n_2844),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_2961),
.B(n_2869),
.Y(n_3593)
);

BUFx3_ASAP7_75t_L g3594 ( 
.A(n_2934),
.Y(n_3594)
);

BUFx2_ASAP7_75t_L g3595 ( 
.A(n_2856),
.Y(n_3595)
);

AND2x4_ASAP7_75t_L g3596 ( 
.A(n_3030),
.B(n_3060),
.Y(n_3596)
);

INVx5_ASAP7_75t_L g3597 ( 
.A(n_2856),
.Y(n_3597)
);

AOI21xp5_ASAP7_75t_L g3598 ( 
.A1(n_3106),
.A2(n_3117),
.B(n_3114),
.Y(n_3598)
);

INVx2_ASAP7_75t_L g3599 ( 
.A(n_2997),
.Y(n_3599)
);

BUFx4_ASAP7_75t_SL g3600 ( 
.A(n_2876),
.Y(n_3600)
);

CKINVDCx20_ASAP7_75t_R g3601 ( 
.A(n_2933),
.Y(n_3601)
);

INVx3_ASAP7_75t_L g3602 ( 
.A(n_2856),
.Y(n_3602)
);

CKINVDCx11_ASAP7_75t_R g3603 ( 
.A(n_2856),
.Y(n_3603)
);

BUFx2_ASAP7_75t_L g3604 ( 
.A(n_2856),
.Y(n_3604)
);

NOR2xp33_ASAP7_75t_L g3605 ( 
.A(n_2933),
.B(n_2984),
.Y(n_3605)
);

BUFx6f_ASAP7_75t_L g3606 ( 
.A(n_2856),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_2869),
.B(n_2876),
.Y(n_3607)
);

INVx2_ASAP7_75t_SL g3608 ( 
.A(n_2895),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3015),
.Y(n_3609)
);

OR2x2_ASAP7_75t_L g3610 ( 
.A(n_2962),
.B(n_2971),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_2840),
.Y(n_3611)
);

AND2x2_ASAP7_75t_L g3612 ( 
.A(n_3060),
.B(n_3061),
.Y(n_3612)
);

BUFx12f_ASAP7_75t_L g3613 ( 
.A(n_2932),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_L g3614 ( 
.A(n_2915),
.B(n_2920),
.Y(n_3614)
);

AOI221xp5_ASAP7_75t_L g3615 ( 
.A1(n_2692),
.A2(n_2840),
.B1(n_2852),
.B2(n_2847),
.C(n_3054),
.Y(n_3615)
);

NAND2xp5_ASAP7_75t_L g3616 ( 
.A(n_2915),
.B(n_2920),
.Y(n_3616)
);

INVx2_ASAP7_75t_SL g3617 ( 
.A(n_2934),
.Y(n_3617)
);

INVx2_ASAP7_75t_L g3618 ( 
.A(n_2997),
.Y(n_3618)
);

CKINVDCx5p33_ASAP7_75t_R g3619 ( 
.A(n_2988),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_2852),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_2862),
.B(n_2880),
.Y(n_3621)
);

OR2x6_ASAP7_75t_L g3622 ( 
.A(n_2621),
.B(n_3092),
.Y(n_3622)
);

O2A1O1Ixp5_ASAP7_75t_L g3623 ( 
.A1(n_2918),
.A2(n_2797),
.B(n_2889),
.C(n_3018),
.Y(n_3623)
);

OR2x6_ASAP7_75t_L g3624 ( 
.A(n_2621),
.B(n_3092),
.Y(n_3624)
);

OAI21xp5_ASAP7_75t_L g3625 ( 
.A1(n_2851),
.A2(n_3114),
.B(n_3106),
.Y(n_3625)
);

NOR2xp33_ASAP7_75t_L g3626 ( 
.A(n_3003),
.B(n_2909),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3055),
.Y(n_3627)
);

CKINVDCx5p33_ASAP7_75t_R g3628 ( 
.A(n_3061),
.Y(n_3628)
);

BUFx2_ASAP7_75t_L g3629 ( 
.A(n_2895),
.Y(n_3629)
);

INVx2_ASAP7_75t_L g3630 ( 
.A(n_2997),
.Y(n_3630)
);

NOR2xp33_ASAP7_75t_L g3631 ( 
.A(n_2909),
.B(n_2904),
.Y(n_3631)
);

INVx2_ASAP7_75t_SL g3632 ( 
.A(n_3022),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_2830),
.B(n_2923),
.Y(n_3633)
);

INVx1_ASAP7_75t_SL g3634 ( 
.A(n_2895),
.Y(n_3634)
);

BUFx12f_ASAP7_75t_L g3635 ( 
.A(n_3092),
.Y(n_3635)
);

NAND2x1p5_ASAP7_75t_L g3636 ( 
.A(n_2897),
.B(n_2804),
.Y(n_3636)
);

BUFx6f_ASAP7_75t_L g3637 ( 
.A(n_2895),
.Y(n_3637)
);

AND2x2_ASAP7_75t_L g3638 ( 
.A(n_2968),
.B(n_2963),
.Y(n_3638)
);

AND2x4_ASAP7_75t_L g3639 ( 
.A(n_2963),
.B(n_2850),
.Y(n_3639)
);

AND2x4_ASAP7_75t_L g3640 ( 
.A(n_2850),
.B(n_2865),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3055),
.Y(n_3641)
);

AOI22xp5_ASAP7_75t_L g3642 ( 
.A1(n_2692),
.A2(n_3098),
.B1(n_3132),
.B2(n_3016),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_2971),
.Y(n_3643)
);

OAI22xp5_ASAP7_75t_L g3644 ( 
.A1(n_2904),
.A2(n_2907),
.B1(n_3132),
.B2(n_3098),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_2968),
.Y(n_3645)
);

NOR2xp33_ASAP7_75t_L g3646 ( 
.A(n_2907),
.B(n_3058),
.Y(n_3646)
);

BUFx2_ASAP7_75t_L g3647 ( 
.A(n_2895),
.Y(n_3647)
);

BUFx2_ASAP7_75t_L g3648 ( 
.A(n_2895),
.Y(n_3648)
);

AND2x2_ASAP7_75t_L g3649 ( 
.A(n_2789),
.B(n_2717),
.Y(n_3649)
);

HB1xp67_ASAP7_75t_L g3650 ( 
.A(n_2923),
.Y(n_3650)
);

O2A1O1Ixp33_ASAP7_75t_L g3651 ( 
.A1(n_3035),
.A2(n_3120),
.B(n_3018),
.C(n_3054),
.Y(n_3651)
);

BUFx12f_ASAP7_75t_L g3652 ( 
.A(n_3098),
.Y(n_3652)
);

AND2x4_ASAP7_75t_L g3653 ( 
.A(n_2850),
.B(n_2865),
.Y(n_3653)
);

A2O1A1Ixp33_ASAP7_75t_L g3654 ( 
.A1(n_2712),
.A2(n_2788),
.B(n_2889),
.C(n_2873),
.Y(n_3654)
);

A2O1A1Ixp33_ASAP7_75t_L g3655 ( 
.A1(n_2712),
.A2(n_2788),
.B(n_2873),
.C(n_2881),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_L g3656 ( 
.A(n_2923),
.B(n_2924),
.Y(n_3656)
);

AND2x2_ASAP7_75t_L g3657 ( 
.A(n_2789),
.B(n_2717),
.Y(n_3657)
);

AOI21xp33_ASAP7_75t_L g3658 ( 
.A1(n_2718),
.A2(n_2727),
.B(n_2679),
.Y(n_3658)
);

AOI21xp5_ASAP7_75t_L g3659 ( 
.A1(n_3114),
.A2(n_3130),
.B(n_3117),
.Y(n_3659)
);

AND2x4_ASAP7_75t_L g3660 ( 
.A(n_2865),
.B(n_2603),
.Y(n_3660)
);

AOI21xp5_ASAP7_75t_L g3661 ( 
.A1(n_3117),
.A2(n_3135),
.B(n_3130),
.Y(n_3661)
);

BUFx3_ASAP7_75t_L g3662 ( 
.A(n_2895),
.Y(n_3662)
);

INVx2_ASAP7_75t_L g3663 ( 
.A(n_3006),
.Y(n_3663)
);

OAI22xp5_ASAP7_75t_L g3664 ( 
.A1(n_3098),
.A2(n_3132),
.B1(n_3042),
.B2(n_3126),
.Y(n_3664)
);

INVx2_ASAP7_75t_L g3665 ( 
.A(n_3006),
.Y(n_3665)
);

BUFx10_ASAP7_75t_L g3666 ( 
.A(n_3026),
.Y(n_3666)
);

OR2x2_ASAP7_75t_L g3667 ( 
.A(n_2924),
.B(n_2947),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_2924),
.B(n_2947),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_L g3669 ( 
.A(n_2947),
.B(n_2614),
.Y(n_3669)
);

HB1xp67_ASAP7_75t_L g3670 ( 
.A(n_2614),
.Y(n_3670)
);

AND2x4_ASAP7_75t_L g3671 ( 
.A(n_2603),
.B(n_2632),
.Y(n_3671)
);

AND2x4_ASAP7_75t_SL g3672 ( 
.A(n_3042),
.B(n_2603),
.Y(n_3672)
);

A2O1A1Ixp33_ASAP7_75t_SL g3673 ( 
.A1(n_2875),
.A2(n_2892),
.B(n_2791),
.C(n_2864),
.Y(n_3673)
);

AO32x2_ASAP7_75t_L g3674 ( 
.A1(n_3052),
.A2(n_3058),
.A3(n_3051),
.B1(n_3040),
.B2(n_3023),
.Y(n_3674)
);

BUFx3_ASAP7_75t_L g3675 ( 
.A(n_3026),
.Y(n_3675)
);

INVx3_ASAP7_75t_L g3676 ( 
.A(n_3026),
.Y(n_3676)
);

BUFx12f_ASAP7_75t_L g3677 ( 
.A(n_3132),
.Y(n_3677)
);

AOI22xp33_ASAP7_75t_SL g3678 ( 
.A1(n_3218),
.A2(n_2789),
.B1(n_2614),
.B2(n_2982),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_L g3679 ( 
.A(n_3270),
.B(n_2614),
.Y(n_3679)
);

AOI22xp33_ASAP7_75t_SL g3680 ( 
.A1(n_3218),
.A2(n_2789),
.B1(n_2614),
.B2(n_2982),
.Y(n_3680)
);

AOI22xp33_ASAP7_75t_L g3681 ( 
.A1(n_3305),
.A2(n_2789),
.B1(n_2881),
.B2(n_2947),
.Y(n_3681)
);

OAI22xp5_ASAP7_75t_L g3682 ( 
.A1(n_3147),
.A2(n_3126),
.B1(n_2603),
.B2(n_2690),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3154),
.Y(n_3683)
);

INVx2_ASAP7_75t_L g3684 ( 
.A(n_3667),
.Y(n_3684)
);

AOI22xp33_ASAP7_75t_L g3685 ( 
.A1(n_3305),
.A2(n_2789),
.B1(n_2947),
.B2(n_3110),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3154),
.Y(n_3686)
);

CKINVDCx11_ASAP7_75t_R g3687 ( 
.A(n_3149),
.Y(n_3687)
);

BUFx8_ASAP7_75t_L g3688 ( 
.A(n_3217),
.Y(n_3688)
);

BUFx4_ASAP7_75t_SL g3689 ( 
.A(n_3265),
.Y(n_3689)
);

AOI22xp5_ASAP7_75t_L g3690 ( 
.A1(n_3165),
.A2(n_2789),
.B1(n_2718),
.B2(n_3081),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3155),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3155),
.Y(n_3692)
);

INVx1_ASAP7_75t_SL g3693 ( 
.A(n_3520),
.Y(n_3693)
);

AOI22xp33_ASAP7_75t_L g3694 ( 
.A1(n_3235),
.A2(n_3276),
.B1(n_3261),
.B2(n_3165),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3163),
.Y(n_3695)
);

INVx6_ASAP7_75t_L g3696 ( 
.A(n_3189),
.Y(n_3696)
);

AND2x2_ASAP7_75t_L g3697 ( 
.A(n_3448),
.B(n_2789),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_L g3698 ( 
.A(n_3270),
.B(n_2614),
.Y(n_3698)
);

NOR2xp33_ASAP7_75t_L g3699 ( 
.A(n_3254),
.B(n_3058),
.Y(n_3699)
);

AOI22xp33_ASAP7_75t_L g3700 ( 
.A1(n_3235),
.A2(n_2789),
.B1(n_3006),
.B2(n_3110),
.Y(n_3700)
);

INVx1_ASAP7_75t_L g3701 ( 
.A(n_3163),
.Y(n_3701)
);

OAI22xp5_ASAP7_75t_L g3702 ( 
.A1(n_3147),
.A2(n_3126),
.B1(n_2690),
.B2(n_2632),
.Y(n_3702)
);

OAI21xp5_ASAP7_75t_SL g3703 ( 
.A1(n_3164),
.A2(n_2781),
.B(n_3126),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3169),
.Y(n_3704)
);

NAND2x1p5_ASAP7_75t_L g3705 ( 
.A(n_3486),
.B(n_2804),
.Y(n_3705)
);

BUFx12f_ASAP7_75t_L g3706 ( 
.A(n_3215),
.Y(n_3706)
);

INVx6_ASAP7_75t_L g3707 ( 
.A(n_3189),
.Y(n_3707)
);

BUFx6f_ASAP7_75t_L g3708 ( 
.A(n_3191),
.Y(n_3708)
);

INVx1_ASAP7_75t_L g3709 ( 
.A(n_3169),
.Y(n_3709)
);

AOI22xp33_ASAP7_75t_L g3710 ( 
.A1(n_3276),
.A2(n_2789),
.B1(n_3089),
.B2(n_3110),
.Y(n_3710)
);

CKINVDCx20_ASAP7_75t_R g3711 ( 
.A(n_3152),
.Y(n_3711)
);

BUFx4f_ASAP7_75t_L g3712 ( 
.A(n_3365),
.Y(n_3712)
);

AOI22xp33_ASAP7_75t_L g3713 ( 
.A1(n_3261),
.A2(n_3089),
.B1(n_3081),
.B2(n_2690),
.Y(n_3713)
);

AOI22xp5_ASAP7_75t_L g3714 ( 
.A1(n_3203),
.A2(n_3316),
.B1(n_3181),
.B2(n_3177),
.Y(n_3714)
);

INVx1_ASAP7_75t_L g3715 ( 
.A(n_3174),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3174),
.Y(n_3716)
);

INVx6_ASAP7_75t_L g3717 ( 
.A(n_3189),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3178),
.Y(n_3718)
);

AOI22xp33_ASAP7_75t_SL g3719 ( 
.A1(n_3232),
.A2(n_2614),
.B1(n_2717),
.B2(n_2718),
.Y(n_3719)
);

BUFx12f_ASAP7_75t_L g3720 ( 
.A(n_3157),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_3178),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_3200),
.Y(n_3722)
);

OAI22xp5_ASAP7_75t_L g3723 ( 
.A1(n_3192),
.A2(n_2690),
.B1(n_3081),
.B2(n_2632),
.Y(n_3723)
);

OAI22xp33_ASAP7_75t_L g3724 ( 
.A1(n_3203),
.A2(n_3175),
.B1(n_3316),
.B2(n_3424),
.Y(n_3724)
);

INVx1_ASAP7_75t_SL g3725 ( 
.A(n_3520),
.Y(n_3725)
);

OAI22xp5_ASAP7_75t_L g3726 ( 
.A1(n_3239),
.A2(n_2632),
.B1(n_3081),
.B2(n_3056),
.Y(n_3726)
);

INVx5_ASAP7_75t_L g3727 ( 
.A(n_3187),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_L g3728 ( 
.A(n_3461),
.B(n_3374),
.Y(n_3728)
);

INVx2_ASAP7_75t_L g3729 ( 
.A(n_3667),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_L g3730 ( 
.A(n_3461),
.B(n_2593),
.Y(n_3730)
);

AOI22xp33_ASAP7_75t_SL g3731 ( 
.A1(n_3232),
.A2(n_2717),
.B1(n_2755),
.B2(n_2727),
.Y(n_3731)
);

AOI22xp33_ASAP7_75t_L g3732 ( 
.A1(n_3278),
.A2(n_3089),
.B1(n_3041),
.B2(n_3045),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_L g3733 ( 
.A(n_3374),
.B(n_2593),
.Y(n_3733)
);

AOI22xp33_ASAP7_75t_L g3734 ( 
.A1(n_3278),
.A2(n_3041),
.B1(n_3045),
.B2(n_3044),
.Y(n_3734)
);

BUFx2_ASAP7_75t_L g3735 ( 
.A(n_3247),
.Y(n_3735)
);

CKINVDCx11_ASAP7_75t_R g3736 ( 
.A(n_3490),
.Y(n_3736)
);

INVx1_ASAP7_75t_L g3737 ( 
.A(n_3209),
.Y(n_3737)
);

INVx1_ASAP7_75t_SL g3738 ( 
.A(n_3554),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3212),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3212),
.Y(n_3740)
);

INVx2_ASAP7_75t_L g3741 ( 
.A(n_3171),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3223),
.Y(n_3742)
);

BUFx4f_ASAP7_75t_L g3743 ( 
.A(n_3365),
.Y(n_3743)
);

BUFx3_ASAP7_75t_L g3744 ( 
.A(n_3217),
.Y(n_3744)
);

INVx2_ASAP7_75t_L g3745 ( 
.A(n_3171),
.Y(n_3745)
);

OAI22xp5_ASAP7_75t_L g3746 ( 
.A1(n_3157),
.A2(n_3056),
.B1(n_2773),
.B2(n_2791),
.Y(n_3746)
);

OAI22xp5_ASAP7_75t_L g3747 ( 
.A1(n_3202),
.A2(n_2864),
.B1(n_2773),
.B2(n_2791),
.Y(n_3747)
);

OAI22xp5_ASAP7_75t_L g3748 ( 
.A1(n_3164),
.A2(n_2864),
.B1(n_2773),
.B2(n_2791),
.Y(n_3748)
);

AOI22xp33_ASAP7_75t_L g3749 ( 
.A1(n_3269),
.A2(n_3044),
.B1(n_3046),
.B2(n_2773),
.Y(n_3749)
);

OAI22xp5_ASAP7_75t_L g3750 ( 
.A1(n_3180),
.A2(n_2864),
.B1(n_2722),
.B2(n_2894),
.Y(n_3750)
);

BUFx12f_ASAP7_75t_L g3751 ( 
.A(n_3185),
.Y(n_3751)
);

AOI22xp33_ASAP7_75t_L g3752 ( 
.A1(n_3269),
.A2(n_3046),
.B1(n_2722),
.B2(n_3012),
.Y(n_3752)
);

OAI22xp33_ASAP7_75t_L g3753 ( 
.A1(n_3175),
.A2(n_2913),
.B1(n_2919),
.B2(n_2722),
.Y(n_3753)
);

CKINVDCx11_ASAP7_75t_R g3754 ( 
.A(n_3517),
.Y(n_3754)
);

BUFx2_ASAP7_75t_L g3755 ( 
.A(n_3247),
.Y(n_3755)
);

AOI22xp33_ASAP7_75t_L g3756 ( 
.A1(n_3381),
.A2(n_2722),
.B1(n_3012),
.B2(n_3008),
.Y(n_3756)
);

BUFx12f_ASAP7_75t_L g3757 ( 
.A(n_3207),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_3223),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3227),
.Y(n_3759)
);

OR2x2_ASAP7_75t_L g3760 ( 
.A(n_3145),
.B(n_2717),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3227),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3230),
.Y(n_3762)
);

INVx2_ASAP7_75t_L g3763 ( 
.A(n_3171),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3230),
.Y(n_3764)
);

INVx4_ASAP7_75t_L g3765 ( 
.A(n_3300),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_3234),
.Y(n_3766)
);

INVx4_ASAP7_75t_L g3767 ( 
.A(n_3300),
.Y(n_3767)
);

INVx2_ASAP7_75t_SL g3768 ( 
.A(n_3559),
.Y(n_3768)
);

CKINVDCx20_ASAP7_75t_R g3769 ( 
.A(n_3217),
.Y(n_3769)
);

OAI22xp33_ASAP7_75t_L g3770 ( 
.A1(n_3424),
.A2(n_2913),
.B1(n_2919),
.B2(n_2894),
.Y(n_3770)
);

INVx1_ASAP7_75t_SL g3771 ( 
.A(n_3554),
.Y(n_3771)
);

OAI22xp5_ASAP7_75t_L g3772 ( 
.A1(n_3153),
.A2(n_3052),
.B1(n_2717),
.B2(n_3111),
.Y(n_3772)
);

CKINVDCx20_ASAP7_75t_R g3773 ( 
.A(n_3300),
.Y(n_3773)
);

INVx1_ASAP7_75t_SL g3774 ( 
.A(n_3600),
.Y(n_3774)
);

INVx1_ASAP7_75t_L g3775 ( 
.A(n_3234),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_L g3776 ( 
.A(n_3381),
.B(n_2593),
.Y(n_3776)
);

INVx3_ASAP7_75t_L g3777 ( 
.A(n_3176),
.Y(n_3777)
);

BUFx3_ASAP7_75t_L g3778 ( 
.A(n_3166),
.Y(n_3778)
);

INVx1_ASAP7_75t_L g3779 ( 
.A(n_3244),
.Y(n_3779)
);

BUFx6f_ASAP7_75t_L g3780 ( 
.A(n_3191),
.Y(n_3780)
);

AOI22xp5_ASAP7_75t_L g3781 ( 
.A1(n_3237),
.A2(n_2897),
.B1(n_2813),
.B2(n_2985),
.Y(n_3781)
);

INVx1_ASAP7_75t_L g3782 ( 
.A(n_3244),
.Y(n_3782)
);

INVx3_ASAP7_75t_L g3783 ( 
.A(n_3176),
.Y(n_3783)
);

BUFx10_ASAP7_75t_L g3784 ( 
.A(n_3511),
.Y(n_3784)
);

OAI22xp33_ASAP7_75t_L g3785 ( 
.A1(n_3330),
.A2(n_3111),
.B1(n_3026),
.B2(n_3023),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_3266),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3266),
.Y(n_3787)
);

AND2x2_ASAP7_75t_L g3788 ( 
.A(n_3448),
.B(n_2717),
.Y(n_3788)
);

BUFx8_ASAP7_75t_L g3789 ( 
.A(n_3166),
.Y(n_3789)
);

BUFx12f_ASAP7_75t_L g3790 ( 
.A(n_3326),
.Y(n_3790)
);

AOI22xp33_ASAP7_75t_L g3791 ( 
.A1(n_3298),
.A2(n_3039),
.B1(n_3008),
.B2(n_3007),
.Y(n_3791)
);

AOI22xp33_ASAP7_75t_SL g3792 ( 
.A1(n_3298),
.A2(n_2755),
.B1(n_2727),
.B2(n_3120),
.Y(n_3792)
);

BUFx4f_ASAP7_75t_SL g3793 ( 
.A(n_3562),
.Y(n_3793)
);

AOI22xp33_ASAP7_75t_L g3794 ( 
.A1(n_3369),
.A2(n_3039),
.B1(n_3007),
.B2(n_2985),
.Y(n_3794)
);

CKINVDCx14_ASAP7_75t_R g3795 ( 
.A(n_3339),
.Y(n_3795)
);

HB1xp67_ASAP7_75t_L g3796 ( 
.A(n_3650),
.Y(n_3796)
);

AOI22xp33_ASAP7_75t_L g3797 ( 
.A1(n_3369),
.A2(n_2973),
.B1(n_2813),
.B2(n_2927),
.Y(n_3797)
);

BUFx10_ASAP7_75t_L g3798 ( 
.A(n_3511),
.Y(n_3798)
);

INVx5_ASAP7_75t_L g3799 ( 
.A(n_3187),
.Y(n_3799)
);

AOI22xp33_ASAP7_75t_L g3800 ( 
.A1(n_3472),
.A2(n_2973),
.B1(n_2813),
.B2(n_2927),
.Y(n_3800)
);

INVx1_ASAP7_75t_L g3801 ( 
.A(n_3283),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3283),
.Y(n_3802)
);

OAI22xp33_ASAP7_75t_L g3803 ( 
.A1(n_3330),
.A2(n_3111),
.B1(n_3026),
.B2(n_3058),
.Y(n_3803)
);

CKINVDCx14_ASAP7_75t_R g3804 ( 
.A(n_3302),
.Y(n_3804)
);

CKINVDCx20_ASAP7_75t_R g3805 ( 
.A(n_3491),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_3284),
.Y(n_3806)
);

AOI22xp33_ASAP7_75t_L g3807 ( 
.A1(n_3472),
.A2(n_2949),
.B1(n_2960),
.B2(n_2958),
.Y(n_3807)
);

CKINVDCx5p33_ASAP7_75t_R g3808 ( 
.A(n_3469),
.Y(n_3808)
);

OAI22x1_ASAP7_75t_L g3809 ( 
.A1(n_3150),
.A2(n_3052),
.B1(n_3002),
.B2(n_3142),
.Y(n_3809)
);

BUFx12f_ASAP7_75t_L g3810 ( 
.A(n_3384),
.Y(n_3810)
);

INVx2_ASAP7_75t_L g3811 ( 
.A(n_3172),
.Y(n_3811)
);

INVx1_ASAP7_75t_L g3812 ( 
.A(n_3284),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3285),
.Y(n_3813)
);

OAI21xp5_ASAP7_75t_SL g3814 ( 
.A1(n_3146),
.A2(n_3002),
.B(n_2986),
.Y(n_3814)
);

AOI22xp33_ASAP7_75t_L g3815 ( 
.A1(n_3268),
.A2(n_2949),
.B1(n_2960),
.B2(n_2958),
.Y(n_3815)
);

INVx2_ASAP7_75t_L g3816 ( 
.A(n_3172),
.Y(n_3816)
);

AOI22xp33_ASAP7_75t_SL g3817 ( 
.A1(n_3337),
.A2(n_2755),
.B1(n_2784),
.B2(n_3130),
.Y(n_3817)
);

INVx1_ASAP7_75t_L g3818 ( 
.A(n_3285),
.Y(n_3818)
);

AOI22xp33_ASAP7_75t_L g3819 ( 
.A1(n_3268),
.A2(n_2949),
.B1(n_2960),
.B2(n_2958),
.Y(n_3819)
);

OAI22xp5_ASAP7_75t_L g3820 ( 
.A1(n_3153),
.A2(n_3111),
.B1(n_3026),
.B2(n_3002),
.Y(n_3820)
);

BUFx8_ASAP7_75t_SL g3821 ( 
.A(n_3562),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3327),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_L g3823 ( 
.A(n_3508),
.B(n_2593),
.Y(n_3823)
);

INVx1_ASAP7_75t_L g3824 ( 
.A(n_3327),
.Y(n_3824)
);

INVx6_ASAP7_75t_L g3825 ( 
.A(n_3189),
.Y(n_3825)
);

INVx3_ASAP7_75t_SL g3826 ( 
.A(n_3447),
.Y(n_3826)
);

OAI22xp33_ASAP7_75t_L g3827 ( 
.A1(n_3337),
.A2(n_3111),
.B1(n_3026),
.B2(n_3050),
.Y(n_3827)
);

AOI22xp33_ASAP7_75t_L g3828 ( 
.A1(n_3406),
.A2(n_2943),
.B1(n_2948),
.B2(n_2931),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_3328),
.Y(n_3829)
);

INVx2_ASAP7_75t_L g3830 ( 
.A(n_3172),
.Y(n_3830)
);

AOI22xp33_ASAP7_75t_SL g3831 ( 
.A1(n_3347),
.A2(n_2784),
.B1(n_3135),
.B2(n_3136),
.Y(n_3831)
);

AOI22xp33_ASAP7_75t_L g3832 ( 
.A1(n_3206),
.A2(n_2943),
.B1(n_2948),
.B2(n_2931),
.Y(n_3832)
);

CKINVDCx20_ASAP7_75t_R g3833 ( 
.A(n_3491),
.Y(n_3833)
);

INVx1_ASAP7_75t_SL g3834 ( 
.A(n_3500),
.Y(n_3834)
);

AOI22xp33_ASAP7_75t_SL g3835 ( 
.A1(n_3347),
.A2(n_2784),
.B1(n_3135),
.B2(n_3136),
.Y(n_3835)
);

AOI22xp33_ASAP7_75t_SL g3836 ( 
.A1(n_3370),
.A2(n_3551),
.B1(n_3549),
.B2(n_3502),
.Y(n_3836)
);

BUFx8_ASAP7_75t_L g3837 ( 
.A(n_3166),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_3328),
.Y(n_3838)
);

BUFx2_ASAP7_75t_L g3839 ( 
.A(n_3247),
.Y(n_3839)
);

AOI22xp33_ASAP7_75t_L g3840 ( 
.A1(n_3287),
.A2(n_2943),
.B1(n_2948),
.B2(n_2931),
.Y(n_3840)
);

AOI22xp33_ASAP7_75t_SL g3841 ( 
.A1(n_3370),
.A2(n_3136),
.B1(n_2679),
.B2(n_2681),
.Y(n_3841)
);

INVx2_ASAP7_75t_SL g3842 ( 
.A(n_3559),
.Y(n_3842)
);

OAI21xp5_ASAP7_75t_SL g3843 ( 
.A1(n_3146),
.A2(n_3002),
.B(n_2986),
.Y(n_3843)
);

AOI22xp33_ASAP7_75t_L g3844 ( 
.A1(n_3323),
.A2(n_2926),
.B1(n_2927),
.B2(n_2897),
.Y(n_3844)
);

AOI22xp33_ASAP7_75t_L g3845 ( 
.A1(n_3323),
.A2(n_2926),
.B1(n_3027),
.B2(n_3029),
.Y(n_3845)
);

AOI22xp33_ASAP7_75t_SL g3846 ( 
.A1(n_3549),
.A2(n_2679),
.B1(n_2681),
.B2(n_2772),
.Y(n_3846)
);

INVx4_ASAP7_75t_SL g3847 ( 
.A(n_3415),
.Y(n_3847)
);

OAI22xp5_ASAP7_75t_L g3848 ( 
.A1(n_3357),
.A2(n_3280),
.B1(n_3310),
.B2(n_3601),
.Y(n_3848)
);

AOI22xp33_ASAP7_75t_SL g3849 ( 
.A1(n_3551),
.A2(n_2681),
.B1(n_2772),
.B2(n_2738),
.Y(n_3849)
);

INVx3_ASAP7_75t_L g3850 ( 
.A(n_3176),
.Y(n_3850)
);

AOI22xp33_ASAP7_75t_L g3851 ( 
.A1(n_3323),
.A2(n_2926),
.B1(n_3025),
.B2(n_2993),
.Y(n_3851)
);

INVx6_ASAP7_75t_L g3852 ( 
.A(n_3189),
.Y(n_3852)
);

CKINVDCx20_ASAP7_75t_R g3853 ( 
.A(n_3628),
.Y(n_3853)
);

INVx2_ASAP7_75t_L g3854 ( 
.A(n_3214),
.Y(n_3854)
);

INVx6_ASAP7_75t_L g3855 ( 
.A(n_3189),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3342),
.Y(n_3856)
);

INVx1_ASAP7_75t_SL g3857 ( 
.A(n_3500),
.Y(n_3857)
);

INVx1_ASAP7_75t_L g3858 ( 
.A(n_3342),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_3346),
.Y(n_3859)
);

CKINVDCx20_ASAP7_75t_R g3860 ( 
.A(n_3423),
.Y(n_3860)
);

AOI22xp33_ASAP7_75t_L g3861 ( 
.A1(n_3323),
.A2(n_2970),
.B1(n_3027),
.B2(n_3029),
.Y(n_3861)
);

BUFx2_ASAP7_75t_SL g3862 ( 
.A(n_3331),
.Y(n_3862)
);

BUFx2_ASAP7_75t_L g3863 ( 
.A(n_3274),
.Y(n_3863)
);

CKINVDCx6p67_ASAP7_75t_R g3864 ( 
.A(n_3274),
.Y(n_3864)
);

OAI22xp5_ASAP7_75t_L g3865 ( 
.A1(n_3310),
.A2(n_3111),
.B1(n_3059),
.B2(n_3050),
.Y(n_3865)
);

INVx3_ASAP7_75t_L g3866 ( 
.A(n_3176),
.Y(n_3866)
);

AOI22xp33_ASAP7_75t_SL g3867 ( 
.A1(n_3502),
.A2(n_2772),
.B1(n_2738),
.B2(n_2735),
.Y(n_3867)
);

OAI22xp33_ASAP7_75t_L g3868 ( 
.A1(n_3338),
.A2(n_3111),
.B1(n_3059),
.B2(n_3048),
.Y(n_3868)
);

AOI22xp33_ASAP7_75t_L g3869 ( 
.A1(n_3323),
.A2(n_3450),
.B1(n_3415),
.B2(n_3436),
.Y(n_3869)
);

AOI22xp33_ASAP7_75t_L g3870 ( 
.A1(n_3323),
.A2(n_2993),
.B1(n_3000),
.B2(n_3043),
.Y(n_3870)
);

AOI22xp33_ASAP7_75t_L g3871 ( 
.A1(n_3323),
.A2(n_2993),
.B1(n_3000),
.B2(n_3043),
.Y(n_3871)
);

INVx1_ASAP7_75t_L g3872 ( 
.A(n_3346),
.Y(n_3872)
);

BUFx3_ASAP7_75t_L g3873 ( 
.A(n_3390),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_3373),
.Y(n_3874)
);

INVx2_ASAP7_75t_L g3875 ( 
.A(n_3214),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_L g3876 ( 
.A(n_3508),
.B(n_3521),
.Y(n_3876)
);

AOI22xp33_ASAP7_75t_L g3877 ( 
.A1(n_3323),
.A2(n_2991),
.B1(n_2983),
.B2(n_3043),
.Y(n_3877)
);

OAI22xp5_ASAP7_75t_L g3878 ( 
.A1(n_3243),
.A2(n_3274),
.B1(n_3307),
.B2(n_3334),
.Y(n_3878)
);

INVx2_ASAP7_75t_L g3879 ( 
.A(n_3214),
.Y(n_3879)
);

BUFx10_ASAP7_75t_L g3880 ( 
.A(n_3511),
.Y(n_3880)
);

AOI21xp5_ASAP7_75t_L g3881 ( 
.A1(n_3257),
.A2(n_3290),
.B(n_3162),
.Y(n_3881)
);

BUFx2_ASAP7_75t_L g3882 ( 
.A(n_3307),
.Y(n_3882)
);

OAI22xp5_ASAP7_75t_L g3883 ( 
.A1(n_3307),
.A2(n_3048),
.B1(n_3017),
.B2(n_3005),
.Y(n_3883)
);

BUFx6f_ASAP7_75t_L g3884 ( 
.A(n_3229),
.Y(n_3884)
);

CKINVDCx11_ASAP7_75t_R g3885 ( 
.A(n_3562),
.Y(n_3885)
);

BUFx8_ASAP7_75t_L g3886 ( 
.A(n_3390),
.Y(n_3886)
);

OAI22xp33_ASAP7_75t_R g3887 ( 
.A1(n_3311),
.A2(n_2593),
.B1(n_3095),
.B2(n_3091),
.Y(n_3887)
);

OAI22xp5_ASAP7_75t_L g3888 ( 
.A1(n_3444),
.A2(n_3017),
.B1(n_3005),
.B2(n_2938),
.Y(n_3888)
);

BUFx12f_ASAP7_75t_L g3889 ( 
.A(n_3390),
.Y(n_3889)
);

CKINVDCx11_ASAP7_75t_R g3890 ( 
.A(n_3210),
.Y(n_3890)
);

BUFx2_ASAP7_75t_L g3891 ( 
.A(n_3518),
.Y(n_3891)
);

INVx1_ASAP7_75t_SL g3892 ( 
.A(n_3504),
.Y(n_3892)
);

OAI22xp5_ASAP7_75t_L g3893 ( 
.A1(n_3444),
.A2(n_2938),
.B1(n_2992),
.B2(n_2989),
.Y(n_3893)
);

INVx6_ASAP7_75t_L g3894 ( 
.A(n_3189),
.Y(n_3894)
);

INVx4_ASAP7_75t_L g3895 ( 
.A(n_3365),
.Y(n_3895)
);

AOI22xp33_ASAP7_75t_L g3896 ( 
.A1(n_3450),
.A2(n_3000),
.B1(n_3036),
.B2(n_3033),
.Y(n_3896)
);

INVx2_ASAP7_75t_L g3897 ( 
.A(n_3219),
.Y(n_3897)
);

INVx2_ASAP7_75t_L g3898 ( 
.A(n_3219),
.Y(n_3898)
);

INVx2_ASAP7_75t_SL g3899 ( 
.A(n_3559),
.Y(n_3899)
);

BUFx2_ASAP7_75t_L g3900 ( 
.A(n_3518),
.Y(n_3900)
);

BUFx3_ASAP7_75t_L g3901 ( 
.A(n_3332),
.Y(n_3901)
);

INVx2_ASAP7_75t_L g3902 ( 
.A(n_3219),
.Y(n_3902)
);

OAI22xp5_ASAP7_75t_L g3903 ( 
.A1(n_3538),
.A2(n_2992),
.B1(n_2989),
.B2(n_2987),
.Y(n_3903)
);

INVx3_ASAP7_75t_L g3904 ( 
.A(n_3179),
.Y(n_3904)
);

AOI22xp33_ASAP7_75t_L g3905 ( 
.A1(n_3415),
.A2(n_2996),
.B1(n_3036),
.B2(n_3033),
.Y(n_3905)
);

OAI22x1_ASAP7_75t_L g3906 ( 
.A1(n_3150),
.A2(n_2593),
.B1(n_3095),
.B2(n_3091),
.Y(n_3906)
);

BUFx2_ASAP7_75t_SL g3907 ( 
.A(n_3331),
.Y(n_3907)
);

AND2x2_ASAP7_75t_L g3908 ( 
.A(n_3494),
.B(n_2593),
.Y(n_3908)
);

CKINVDCx5p33_ASAP7_75t_R g3909 ( 
.A(n_3513),
.Y(n_3909)
);

INVx4_ASAP7_75t_L g3910 ( 
.A(n_3365),
.Y(n_3910)
);

AND2x2_ASAP7_75t_L g3911 ( 
.A(n_3494),
.B(n_3142),
.Y(n_3911)
);

AOI22xp33_ASAP7_75t_L g3912 ( 
.A1(n_3415),
.A2(n_2996),
.B1(n_3033),
.B2(n_2991),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3373),
.Y(n_3913)
);

BUFx12f_ASAP7_75t_L g3914 ( 
.A(n_3619),
.Y(n_3914)
);

INVx2_ASAP7_75t_L g3915 ( 
.A(n_3222),
.Y(n_3915)
);

OR2x2_ASAP7_75t_L g3916 ( 
.A(n_3145),
.B(n_3142),
.Y(n_3916)
);

NAND2x1p5_ASAP7_75t_L g3917 ( 
.A(n_3486),
.B(n_2848),
.Y(n_3917)
);

CKINVDCx5p33_ASAP7_75t_R g3918 ( 
.A(n_3249),
.Y(n_3918)
);

HB1xp67_ASAP7_75t_L g3919 ( 
.A(n_3224),
.Y(n_3919)
);

INVx2_ASAP7_75t_L g3920 ( 
.A(n_3222),
.Y(n_3920)
);

BUFx2_ASAP7_75t_L g3921 ( 
.A(n_3518),
.Y(n_3921)
);

INVx1_ASAP7_75t_SL g3922 ( 
.A(n_3504),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3388),
.Y(n_3923)
);

OAI22xp5_ASAP7_75t_L g3924 ( 
.A1(n_3538),
.A2(n_2987),
.B1(n_2892),
.B2(n_2875),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3388),
.Y(n_3925)
);

INVx2_ASAP7_75t_L g3926 ( 
.A(n_3222),
.Y(n_3926)
);

INVx6_ASAP7_75t_L g3927 ( 
.A(n_3193),
.Y(n_3927)
);

INVx2_ASAP7_75t_L g3928 ( 
.A(n_3225),
.Y(n_3928)
);

AOI22xp33_ASAP7_75t_SL g3929 ( 
.A1(n_3525),
.A2(n_2738),
.B1(n_2735),
.B2(n_2624),
.Y(n_3929)
);

BUFx3_ASAP7_75t_L g3930 ( 
.A(n_3332),
.Y(n_3930)
);

BUFx8_ASAP7_75t_L g3931 ( 
.A(n_3546),
.Y(n_3931)
);

OAI22xp5_ASAP7_75t_L g3932 ( 
.A1(n_3566),
.A2(n_2875),
.B1(n_2892),
.B2(n_3022),
.Y(n_3932)
);

OAI22xp33_ASAP7_75t_L g3933 ( 
.A1(n_3338),
.A2(n_2875),
.B1(n_2892),
.B2(n_3095),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_3521),
.B(n_3426),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3389),
.Y(n_3935)
);

AOI22xp33_ASAP7_75t_SL g3936 ( 
.A1(n_3525),
.A2(n_2735),
.B1(n_2624),
.B2(n_2698),
.Y(n_3936)
);

OAI22xp5_ASAP7_75t_L g3937 ( 
.A1(n_3566),
.A2(n_3142),
.B1(n_3095),
.B2(n_3091),
.Y(n_3937)
);

INVx3_ASAP7_75t_L g3938 ( 
.A(n_3179),
.Y(n_3938)
);

AOI22xp33_ASAP7_75t_L g3939 ( 
.A1(n_3415),
.A2(n_2983),
.B1(n_3025),
.B2(n_2981),
.Y(n_3939)
);

AOI22xp5_ASAP7_75t_L g3940 ( 
.A1(n_3399),
.A2(n_2893),
.B1(n_2848),
.B2(n_2698),
.Y(n_3940)
);

BUFx8_ASAP7_75t_L g3941 ( 
.A(n_3546),
.Y(n_3941)
);

AOI22xp5_ASAP7_75t_L g3942 ( 
.A1(n_3345),
.A2(n_2893),
.B1(n_2848),
.B2(n_2698),
.Y(n_3942)
);

OAI21xp5_ASAP7_75t_SL g3943 ( 
.A1(n_3322),
.A2(n_3142),
.B(n_3095),
.Y(n_3943)
);

AOI22xp33_ASAP7_75t_SL g3944 ( 
.A1(n_3537),
.A2(n_3142),
.B1(n_3079),
.B2(n_3088),
.Y(n_3944)
);

BUFx2_ASAP7_75t_L g3945 ( 
.A(n_3561),
.Y(n_3945)
);

AOI22xp33_ASAP7_75t_L g3946 ( 
.A1(n_3436),
.A2(n_2981),
.B1(n_3025),
.B2(n_2970),
.Y(n_3946)
);

AOI22xp5_ASAP7_75t_SL g3947 ( 
.A1(n_3159),
.A2(n_3142),
.B1(n_3095),
.B2(n_3091),
.Y(n_3947)
);

BUFx8_ASAP7_75t_L g3948 ( 
.A(n_3546),
.Y(n_3948)
);

AOI22xp33_ASAP7_75t_L g3949 ( 
.A1(n_3436),
.A2(n_2981),
.B1(n_2996),
.B2(n_3001),
.Y(n_3949)
);

AOI22xp33_ASAP7_75t_L g3950 ( 
.A1(n_3436),
.A2(n_3001),
.B1(n_2991),
.B2(n_2893),
.Y(n_3950)
);

INVx3_ASAP7_75t_L g3951 ( 
.A(n_3179),
.Y(n_3951)
);

INVx5_ASAP7_75t_L g3952 ( 
.A(n_3187),
.Y(n_3952)
);

INVx3_ASAP7_75t_L g3953 ( 
.A(n_3179),
.Y(n_3953)
);

AOI22xp33_ASAP7_75t_L g3954 ( 
.A1(n_3436),
.A2(n_3531),
.B1(n_3506),
.B2(n_3345),
.Y(n_3954)
);

BUFx12f_ASAP7_75t_L g3955 ( 
.A(n_3358),
.Y(n_3955)
);

OAI22xp33_ASAP7_75t_R g3956 ( 
.A1(n_3190),
.A2(n_3095),
.B1(n_3091),
.B2(n_3088),
.Y(n_3956)
);

CKINVDCx11_ASAP7_75t_R g3957 ( 
.A(n_3210),
.Y(n_3957)
);

OAI22xp33_ASAP7_75t_L g3958 ( 
.A1(n_3378),
.A2(n_3091),
.B1(n_3088),
.B2(n_3079),
.Y(n_3958)
);

BUFx3_ASAP7_75t_L g3959 ( 
.A(n_3335),
.Y(n_3959)
);

NAND2x1p5_ASAP7_75t_L g3960 ( 
.A(n_3522),
.B(n_2835),
.Y(n_3960)
);

BUFx2_ASAP7_75t_SL g3961 ( 
.A(n_3331),
.Y(n_3961)
);

INVx3_ASAP7_75t_L g3962 ( 
.A(n_3198),
.Y(n_3962)
);

CKINVDCx14_ASAP7_75t_R g3963 ( 
.A(n_3302),
.Y(n_3963)
);

AOI22xp33_ASAP7_75t_L g3964 ( 
.A1(n_3537),
.A2(n_2935),
.B1(n_2780),
.B2(n_2798),
.Y(n_3964)
);

AND2x2_ASAP7_75t_L g3965 ( 
.A(n_3333),
.B(n_3091),
.Y(n_3965)
);

BUFx12f_ASAP7_75t_L g3966 ( 
.A(n_3358),
.Y(n_3966)
);

AND2x4_ASAP7_75t_L g3967 ( 
.A(n_3397),
.B(n_2823),
.Y(n_3967)
);

AOI22xp33_ASAP7_75t_L g3968 ( 
.A1(n_3543),
.A2(n_2935),
.B1(n_2780),
.B2(n_2798),
.Y(n_3968)
);

CKINVDCx20_ASAP7_75t_R g3969 ( 
.A(n_3423),
.Y(n_3969)
);

NAND2xp5_ASAP7_75t_L g3970 ( 
.A(n_3426),
.B(n_3088),
.Y(n_3970)
);

INVx11_ASAP7_75t_L g3971 ( 
.A(n_3613),
.Y(n_3971)
);

OAI22xp33_ASAP7_75t_R g3972 ( 
.A1(n_3190),
.A2(n_3088),
.B1(n_3079),
.B2(n_2616),
.Y(n_3972)
);

AOI22xp33_ASAP7_75t_SL g3973 ( 
.A1(n_3543),
.A2(n_3088),
.B1(n_3079),
.B2(n_2636),
.Y(n_3973)
);

INVx6_ASAP7_75t_L g3974 ( 
.A(n_3193),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_L g3975 ( 
.A(n_3273),
.B(n_3088),
.Y(n_3975)
);

INVx2_ASAP7_75t_L g3976 ( 
.A(n_3225),
.Y(n_3976)
);

INVxp33_ASAP7_75t_L g3977 ( 
.A(n_3372),
.Y(n_3977)
);

AOI22xp5_ASAP7_75t_L g3978 ( 
.A1(n_3457),
.A2(n_2780),
.B1(n_2636),
.B2(n_2767),
.Y(n_3978)
);

CKINVDCx11_ASAP7_75t_R g3979 ( 
.A(n_3292),
.Y(n_3979)
);

AOI22xp33_ASAP7_75t_SL g3980 ( 
.A1(n_3501),
.A2(n_3375),
.B1(n_3159),
.B2(n_3368),
.Y(n_3980)
);

AND2x2_ASAP7_75t_L g3981 ( 
.A(n_3333),
.B(n_3079),
.Y(n_3981)
);

INVx6_ASAP7_75t_L g3982 ( 
.A(n_3193),
.Y(n_3982)
);

INVx2_ASAP7_75t_SL g3983 ( 
.A(n_3559),
.Y(n_3983)
);

AOI22xp33_ASAP7_75t_L g3984 ( 
.A1(n_3375),
.A2(n_2798),
.B1(n_2767),
.B2(n_2677),
.Y(n_3984)
);

OAI21xp5_ASAP7_75t_L g3985 ( 
.A1(n_3160),
.A2(n_2677),
.B(n_2714),
.Y(n_3985)
);

CKINVDCx11_ASAP7_75t_R g3986 ( 
.A(n_3292),
.Y(n_3986)
);

INVx6_ASAP7_75t_L g3987 ( 
.A(n_3193),
.Y(n_3987)
);

INVx6_ASAP7_75t_L g3988 ( 
.A(n_3193),
.Y(n_3988)
);

AOI22xp33_ASAP7_75t_SL g3989 ( 
.A1(n_3501),
.A2(n_3079),
.B1(n_2677),
.B2(n_2714),
.Y(n_3989)
);

OR2x2_ASAP7_75t_L g3990 ( 
.A(n_3168),
.B(n_3079),
.Y(n_3990)
);

INVx2_ASAP7_75t_SL g3991 ( 
.A(n_3559),
.Y(n_3991)
);

AOI22xp33_ASAP7_75t_L g3992 ( 
.A1(n_3649),
.A2(n_2767),
.B1(n_3021),
.B2(n_2714),
.Y(n_3992)
);

OR2x2_ASAP7_75t_L g3993 ( 
.A(n_3168),
.B(n_2615),
.Y(n_3993)
);

BUFx2_ASAP7_75t_SL g3994 ( 
.A(n_3481),
.Y(n_3994)
);

CKINVDCx20_ASAP7_75t_R g3995 ( 
.A(n_3396),
.Y(n_3995)
);

INVx4_ASAP7_75t_L g3996 ( 
.A(n_3408),
.Y(n_3996)
);

HB1xp67_ASAP7_75t_L g3997 ( 
.A(n_3264),
.Y(n_3997)
);

CKINVDCx6p67_ASAP7_75t_R g3998 ( 
.A(n_3350),
.Y(n_3998)
);

BUFx2_ASAP7_75t_L g3999 ( 
.A(n_3561),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_L g4000 ( 
.A(n_3273),
.B(n_3151),
.Y(n_4000)
);

BUFx3_ASAP7_75t_L g4001 ( 
.A(n_3335),
.Y(n_4001)
);

AOI22xp33_ASAP7_75t_L g4002 ( 
.A1(n_3649),
.A2(n_3021),
.B1(n_2866),
.B2(n_2823),
.Y(n_4002)
);

OAI22xp5_ASAP7_75t_L g4003 ( 
.A1(n_3361),
.A2(n_2616),
.B1(n_2615),
.B2(n_3011),
.Y(n_4003)
);

AOI22xp33_ASAP7_75t_L g4004 ( 
.A1(n_3657),
.A2(n_2866),
.B1(n_2823),
.B2(n_2835),
.Y(n_4004)
);

AOI22xp5_ASAP7_75t_L g4005 ( 
.A1(n_3318),
.A2(n_2835),
.B1(n_2820),
.B2(n_2878),
.Y(n_4005)
);

INVx6_ASAP7_75t_L g4006 ( 
.A(n_3193),
.Y(n_4006)
);

BUFx12f_ASAP7_75t_L g4007 ( 
.A(n_3358),
.Y(n_4007)
);

OAI21xp5_ASAP7_75t_SL g4008 ( 
.A1(n_3322),
.A2(n_2616),
.B(n_2615),
.Y(n_4008)
);

INVx1_ASAP7_75t_SL g4009 ( 
.A(n_3451),
.Y(n_4009)
);

AND2x4_ASAP7_75t_L g4010 ( 
.A(n_3397),
.B(n_2866),
.Y(n_4010)
);

BUFx4_ASAP7_75t_SL g4011 ( 
.A(n_3249),
.Y(n_4011)
);

BUFx3_ASAP7_75t_L g4012 ( 
.A(n_3379),
.Y(n_4012)
);

BUFx6f_ASAP7_75t_L g4013 ( 
.A(n_3229),
.Y(n_4013)
);

AOI22xp33_ASAP7_75t_SL g4014 ( 
.A1(n_3368),
.A2(n_2616),
.B1(n_2765),
.B2(n_2774),
.Y(n_4014)
);

INVx1_ASAP7_75t_L g4015 ( 
.A(n_3455),
.Y(n_4015)
);

CKINVDCx6p67_ASAP7_75t_R g4016 ( 
.A(n_3350),
.Y(n_4016)
);

AOI22xp33_ASAP7_75t_SL g4017 ( 
.A1(n_3496),
.A2(n_2616),
.B1(n_2765),
.B2(n_2774),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_3468),
.Y(n_4018)
);

INVx8_ASAP7_75t_L g4019 ( 
.A(n_3635),
.Y(n_4019)
);

INVx1_ASAP7_75t_SL g4020 ( 
.A(n_3451),
.Y(n_4020)
);

BUFx2_ASAP7_75t_L g4021 ( 
.A(n_3561),
.Y(n_4021)
);

INVx1_ASAP7_75t_SL g4022 ( 
.A(n_3379),
.Y(n_4022)
);

INVx1_ASAP7_75t_L g4023 ( 
.A(n_3468),
.Y(n_4023)
);

BUFx12f_ASAP7_75t_L g4024 ( 
.A(n_3358),
.Y(n_4024)
);

OAI22xp33_ASAP7_75t_L g4025 ( 
.A1(n_3378),
.A2(n_2616),
.B1(n_2615),
.B2(n_2888),
.Y(n_4025)
);

INVx3_ASAP7_75t_SL g4026 ( 
.A(n_3447),
.Y(n_4026)
);

INVx1_ASAP7_75t_L g4027 ( 
.A(n_3476),
.Y(n_4027)
);

INVx6_ASAP7_75t_L g4028 ( 
.A(n_3193),
.Y(n_4028)
);

INVx6_ASAP7_75t_L g4029 ( 
.A(n_3236),
.Y(n_4029)
);

AOI22xp33_ASAP7_75t_SL g4030 ( 
.A1(n_3496),
.A2(n_2616),
.B1(n_2765),
.B2(n_2774),
.Y(n_4030)
);

HB1xp67_ASAP7_75t_L g4031 ( 
.A(n_3610),
.Y(n_4031)
);

INVx2_ASAP7_75t_L g4032 ( 
.A(n_3262),
.Y(n_4032)
);

INVx4_ASAP7_75t_L g4033 ( 
.A(n_3408),
.Y(n_4033)
);

CKINVDCx20_ASAP7_75t_R g4034 ( 
.A(n_3464),
.Y(n_4034)
);

CKINVDCx20_ASAP7_75t_R g4035 ( 
.A(n_3183),
.Y(n_4035)
);

AOI22xp33_ASAP7_75t_L g4036 ( 
.A1(n_3657),
.A2(n_2820),
.B1(n_2890),
.B2(n_2878),
.Y(n_4036)
);

AOI22xp33_ASAP7_75t_L g4037 ( 
.A1(n_3312),
.A2(n_2820),
.B1(n_2890),
.B2(n_2878),
.Y(n_4037)
);

CKINVDCx6p67_ASAP7_75t_R g4038 ( 
.A(n_3350),
.Y(n_4038)
);

BUFx2_ASAP7_75t_L g4039 ( 
.A(n_3452),
.Y(n_4039)
);

AOI22xp33_ASAP7_75t_L g4040 ( 
.A1(n_3312),
.A2(n_2890),
.B1(n_2885),
.B2(n_2770),
.Y(n_4040)
);

BUFx6f_ASAP7_75t_L g4041 ( 
.A(n_3229),
.Y(n_4041)
);

INVx2_ASAP7_75t_L g4042 ( 
.A(n_3262),
.Y(n_4042)
);

BUFx2_ASAP7_75t_L g4043 ( 
.A(n_3452),
.Y(n_4043)
);

NAND2x1p5_ASAP7_75t_L g4044 ( 
.A(n_3522),
.B(n_2885),
.Y(n_4044)
);

INVx6_ASAP7_75t_L g4045 ( 
.A(n_3236),
.Y(n_4045)
);

INVx2_ASAP7_75t_L g4046 ( 
.A(n_3288),
.Y(n_4046)
);

AOI22xp5_ASAP7_75t_L g4047 ( 
.A1(n_3260),
.A2(n_2885),
.B1(n_2770),
.B2(n_2888),
.Y(n_4047)
);

OAI22xp33_ASAP7_75t_L g4048 ( 
.A1(n_3255),
.A2(n_3281),
.B1(n_3312),
.B2(n_3213),
.Y(n_4048)
);

BUFx2_ASAP7_75t_SL g4049 ( 
.A(n_3481),
.Y(n_4049)
);

INVx1_ASAP7_75t_SL g4050 ( 
.A(n_3431),
.Y(n_4050)
);

INVx6_ASAP7_75t_L g4051 ( 
.A(n_3236),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_3487),
.Y(n_4052)
);

AOI22xp33_ASAP7_75t_L g4053 ( 
.A1(n_3312),
.A2(n_3148),
.B1(n_3213),
.B2(n_3187),
.Y(n_4053)
);

AOI22xp33_ASAP7_75t_L g4054 ( 
.A1(n_3312),
.A2(n_2770),
.B1(n_2888),
.B2(n_2940),
.Y(n_4054)
);

AOI22xp33_ASAP7_75t_SL g4055 ( 
.A1(n_3419),
.A2(n_2615),
.B1(n_2888),
.B2(n_2917),
.Y(n_4055)
);

INVx6_ASAP7_75t_L g4056 ( 
.A(n_3236),
.Y(n_4056)
);

INVxp67_ASAP7_75t_L g4057 ( 
.A(n_3515),
.Y(n_4057)
);

AOI22xp33_ASAP7_75t_SL g4058 ( 
.A1(n_3419),
.A2(n_2615),
.B1(n_2888),
.B2(n_2917),
.Y(n_4058)
);

BUFx4f_ASAP7_75t_L g4059 ( 
.A(n_3205),
.Y(n_4059)
);

BUFx8_ASAP7_75t_SL g4060 ( 
.A(n_3484),
.Y(n_4060)
);

INVx1_ASAP7_75t_SL g4061 ( 
.A(n_3431),
.Y(n_4061)
);

AOI22xp33_ASAP7_75t_L g4062 ( 
.A1(n_3148),
.A2(n_2888),
.B1(n_3024),
.B2(n_2917),
.Y(n_4062)
);

AOI22xp5_ASAP7_75t_SL g4063 ( 
.A1(n_3199),
.A2(n_2615),
.B1(n_2888),
.B2(n_2917),
.Y(n_4063)
);

BUFx6f_ASAP7_75t_SL g4064 ( 
.A(n_3567),
.Y(n_4064)
);

AOI22xp33_ASAP7_75t_L g4065 ( 
.A1(n_3187),
.A2(n_3024),
.B1(n_2940),
.B2(n_3010),
.Y(n_4065)
);

AOI22xp33_ASAP7_75t_L g4066 ( 
.A1(n_3213),
.A2(n_3024),
.B1(n_2940),
.B2(n_3010),
.Y(n_4066)
);

INVx2_ASAP7_75t_SL g4067 ( 
.A(n_3559),
.Y(n_4067)
);

AOI22xp33_ASAP7_75t_L g4068 ( 
.A1(n_3213),
.A2(n_3024),
.B1(n_2940),
.B2(n_3010),
.Y(n_4068)
);

INVx2_ASAP7_75t_SL g4069 ( 
.A(n_3559),
.Y(n_4069)
);

INVx6_ASAP7_75t_L g4070 ( 
.A(n_3236),
.Y(n_4070)
);

BUFx2_ASAP7_75t_L g4071 ( 
.A(n_3484),
.Y(n_4071)
);

HB1xp67_ASAP7_75t_L g4072 ( 
.A(n_3610),
.Y(n_4072)
);

AOI22xp33_ASAP7_75t_L g4073 ( 
.A1(n_3213),
.A2(n_3024),
.B1(n_2940),
.B2(n_3010),
.Y(n_4073)
);

AND2x2_ASAP7_75t_L g4074 ( 
.A(n_3293),
.B(n_2917),
.Y(n_4074)
);

OAI22xp33_ASAP7_75t_L g4075 ( 
.A1(n_3255),
.A2(n_2917),
.B1(n_2940),
.B2(n_3010),
.Y(n_4075)
);

NAND2xp5_ASAP7_75t_L g4076 ( 
.A(n_3151),
.B(n_2917),
.Y(n_4076)
);

INVx6_ASAP7_75t_L g4077 ( 
.A(n_3236),
.Y(n_4077)
);

INVx2_ASAP7_75t_L g4078 ( 
.A(n_3288),
.Y(n_4078)
);

OAI22xp5_ASAP7_75t_L g4079 ( 
.A1(n_3281),
.A2(n_2940),
.B1(n_3010),
.B2(n_3020),
.Y(n_4079)
);

OAI22xp5_ASAP7_75t_L g4080 ( 
.A1(n_3252),
.A2(n_3010),
.B1(n_3020),
.B2(n_3024),
.Y(n_4080)
);

OAI22xp5_ASAP7_75t_L g4081 ( 
.A1(n_3252),
.A2(n_3020),
.B1(n_3024),
.B2(n_3240),
.Y(n_4081)
);

INVx3_ASAP7_75t_L g4082 ( 
.A(n_3198),
.Y(n_4082)
);

INVx2_ASAP7_75t_SL g4083 ( 
.A(n_3597),
.Y(n_4083)
);

CKINVDCx6p67_ASAP7_75t_R g4084 ( 
.A(n_3401),
.Y(n_4084)
);

INVx1_ASAP7_75t_SL g4085 ( 
.A(n_3434),
.Y(n_4085)
);

AOI22xp5_ASAP7_75t_L g4086 ( 
.A1(n_3526),
.A2(n_3020),
.B1(n_3533),
.B2(n_3454),
.Y(n_4086)
);

AND2x2_ASAP7_75t_L g4087 ( 
.A(n_3293),
.B(n_3020),
.Y(n_4087)
);

AOI22xp33_ASAP7_75t_L g4088 ( 
.A1(n_3594),
.A2(n_3020),
.B1(n_3532),
.B2(n_3587),
.Y(n_4088)
);

AOI22xp33_ASAP7_75t_SL g4089 ( 
.A1(n_3199),
.A2(n_3020),
.B1(n_3242),
.B2(n_3238),
.Y(n_4089)
);

CKINVDCx11_ASAP7_75t_R g4090 ( 
.A(n_3413),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_3563),
.Y(n_4091)
);

CKINVDCx6p67_ASAP7_75t_R g4092 ( 
.A(n_3401),
.Y(n_4092)
);

INVx1_ASAP7_75t_L g4093 ( 
.A(n_3563),
.Y(n_4093)
);

CKINVDCx11_ASAP7_75t_R g4094 ( 
.A(n_3413),
.Y(n_4094)
);

AOI22xp33_ASAP7_75t_L g4095 ( 
.A1(n_3594),
.A2(n_3617),
.B1(n_3670),
.B2(n_3282),
.Y(n_4095)
);

AOI22xp33_ASAP7_75t_SL g4096 ( 
.A1(n_3238),
.A2(n_3275),
.B1(n_3296),
.B2(n_3242),
.Y(n_4096)
);

AOI22xp33_ASAP7_75t_SL g4097 ( 
.A1(n_3275),
.A2(n_3308),
.B1(n_3314),
.B2(n_3296),
.Y(n_4097)
);

AOI22xp33_ASAP7_75t_L g4098 ( 
.A1(n_3594),
.A2(n_3617),
.B1(n_3282),
.B2(n_3449),
.Y(n_4098)
);

AOI22xp33_ASAP7_75t_L g4099 ( 
.A1(n_3449),
.A2(n_3631),
.B1(n_3405),
.B2(n_3533),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_L g4100 ( 
.A(n_3196),
.B(n_3197),
.Y(n_4100)
);

AOI22xp33_ASAP7_75t_SL g4101 ( 
.A1(n_3308),
.A2(n_3314),
.B1(n_3364),
.B2(n_3526),
.Y(n_4101)
);

AOI22xp33_ASAP7_75t_L g4102 ( 
.A1(n_3449),
.A2(n_3405),
.B1(n_3509),
.B2(n_3505),
.Y(n_4102)
);

INVx4_ASAP7_75t_L g4103 ( 
.A(n_3408),
.Y(n_4103)
);

BUFx8_ASAP7_75t_L g4104 ( 
.A(n_3613),
.Y(n_4104)
);

OAI22xp5_ASAP7_75t_L g4105 ( 
.A1(n_3240),
.A2(n_3313),
.B1(n_3465),
.B2(n_3290),
.Y(n_4105)
);

BUFx2_ASAP7_75t_L g4106 ( 
.A(n_3434),
.Y(n_4106)
);

INVx6_ASAP7_75t_L g4107 ( 
.A(n_3578),
.Y(n_4107)
);

INVx6_ASAP7_75t_L g4108 ( 
.A(n_3578),
.Y(n_4108)
);

OAI21xp5_ASAP7_75t_L g4109 ( 
.A1(n_3160),
.A2(n_3257),
.B(n_3479),
.Y(n_4109)
);

AOI22xp33_ASAP7_75t_L g4110 ( 
.A1(n_3449),
.A2(n_3405),
.B1(n_3509),
.B2(n_3505),
.Y(n_4110)
);

INVx2_ASAP7_75t_L g4111 ( 
.A(n_3288),
.Y(n_4111)
);

AOI22xp33_ASAP7_75t_SL g4112 ( 
.A1(n_3364),
.A2(n_3542),
.B1(n_3366),
.B2(n_3385),
.Y(n_4112)
);

CKINVDCx20_ASAP7_75t_R g4113 ( 
.A(n_3297),
.Y(n_4113)
);

INVx4_ASAP7_75t_L g4114 ( 
.A(n_3408),
.Y(n_4114)
);

OAI22xp5_ASAP7_75t_L g4115 ( 
.A1(n_3313),
.A2(n_3428),
.B1(n_3605),
.B2(n_3317),
.Y(n_4115)
);

BUFx4f_ASAP7_75t_SL g4116 ( 
.A(n_3613),
.Y(n_4116)
);

AOI22xp33_ASAP7_75t_L g4117 ( 
.A1(n_3449),
.A2(n_3405),
.B1(n_3398),
.B2(n_3462),
.Y(n_4117)
);

AOI22xp33_ASAP7_75t_L g4118 ( 
.A1(n_3473),
.A2(n_3626),
.B1(n_3503),
.B2(n_3404),
.Y(n_4118)
);

OAI21xp5_ASAP7_75t_SL g4119 ( 
.A1(n_3479),
.A2(n_3523),
.B(n_3317),
.Y(n_4119)
);

INVx4_ASAP7_75t_L g4120 ( 
.A(n_3432),
.Y(n_4120)
);

CKINVDCx5p33_ASAP7_75t_R g4121 ( 
.A(n_3377),
.Y(n_4121)
);

BUFx12f_ASAP7_75t_L g4122 ( 
.A(n_3578),
.Y(n_4122)
);

AOI22xp33_ASAP7_75t_L g4123 ( 
.A1(n_3404),
.A2(n_3503),
.B1(n_3430),
.B2(n_3635),
.Y(n_4123)
);

INVx1_ASAP7_75t_L g4124 ( 
.A(n_3609),
.Y(n_4124)
);

BUFx2_ASAP7_75t_SL g4125 ( 
.A(n_3481),
.Y(n_4125)
);

CKINVDCx5p33_ASAP7_75t_R g4126 ( 
.A(n_3447),
.Y(n_4126)
);

INVx1_ASAP7_75t_L g4127 ( 
.A(n_3627),
.Y(n_4127)
);

OAI22xp5_ASAP7_75t_L g4128 ( 
.A1(n_3156),
.A2(n_3162),
.B1(n_3184),
.B2(n_3170),
.Y(n_4128)
);

CKINVDCx5p33_ASAP7_75t_R g4129 ( 
.A(n_3301),
.Y(n_4129)
);

BUFx2_ASAP7_75t_L g4130 ( 
.A(n_3539),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_3627),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_3641),
.Y(n_4132)
);

AOI22xp33_ASAP7_75t_SL g4133 ( 
.A1(n_3542),
.A2(n_3437),
.B1(n_3319),
.B2(n_3294),
.Y(n_4133)
);

CKINVDCx5p33_ASAP7_75t_R g4134 ( 
.A(n_3301),
.Y(n_4134)
);

BUFx2_ASAP7_75t_L g4135 ( 
.A(n_3539),
.Y(n_4135)
);

CKINVDCx11_ASAP7_75t_R g4136 ( 
.A(n_3413),
.Y(n_4136)
);

AOI22xp33_ASAP7_75t_L g4137 ( 
.A1(n_3430),
.A2(n_3652),
.B1(n_3677),
.B2(n_3635),
.Y(n_4137)
);

AOI22xp33_ASAP7_75t_L g4138 ( 
.A1(n_3430),
.A2(n_3677),
.B1(n_3652),
.B2(n_3435),
.Y(n_4138)
);

INVx1_ASAP7_75t_L g4139 ( 
.A(n_3641),
.Y(n_4139)
);

AOI22xp33_ASAP7_75t_SL g4140 ( 
.A1(n_3291),
.A2(n_3294),
.B1(n_3669),
.B2(n_3625),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_3621),
.Y(n_4141)
);

OAI22x1_ASAP7_75t_L g4142 ( 
.A1(n_3642),
.A2(n_3639),
.B1(n_3173),
.B2(n_3158),
.Y(n_4142)
);

BUFx2_ASAP7_75t_L g4143 ( 
.A(n_3552),
.Y(n_4143)
);

AOI22xp5_ASAP7_75t_SL g4144 ( 
.A1(n_3467),
.A2(n_3480),
.B1(n_3245),
.B2(n_3267),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_3621),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_3458),
.Y(n_4146)
);

INVx6_ASAP7_75t_L g4147 ( 
.A(n_3578),
.Y(n_4147)
);

AOI22xp33_ASAP7_75t_L g4148 ( 
.A1(n_3430),
.A2(n_3677),
.B1(n_3652),
.B2(n_3435),
.Y(n_4148)
);

OAI22xp5_ASAP7_75t_L g4149 ( 
.A1(n_3156),
.A2(n_3184),
.B1(n_3216),
.B2(n_3170),
.Y(n_4149)
);

INVx1_ASAP7_75t_L g4150 ( 
.A(n_3458),
.Y(n_4150)
);

INVx8_ASAP7_75t_L g4151 ( 
.A(n_3622),
.Y(n_4151)
);

BUFx12f_ASAP7_75t_L g4152 ( 
.A(n_3603),
.Y(n_4152)
);

NAND2xp5_ASAP7_75t_L g4153 ( 
.A(n_3196),
.B(n_3197),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_3463),
.Y(n_4154)
);

AOI21xp33_ASAP7_75t_L g4155 ( 
.A1(n_3306),
.A2(n_3320),
.B(n_3348),
.Y(n_4155)
);

AOI22xp33_ASAP7_75t_L g4156 ( 
.A1(n_3418),
.A2(n_3435),
.B1(n_3251),
.B2(n_3256),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_3463),
.Y(n_4157)
);

BUFx12f_ASAP7_75t_L g4158 ( 
.A(n_3573),
.Y(n_4158)
);

CKINVDCx20_ASAP7_75t_R g4159 ( 
.A(n_3556),
.Y(n_4159)
);

INVx2_ASAP7_75t_SL g4160 ( 
.A(n_3597),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_3614),
.Y(n_4161)
);

NAND2xp5_ASAP7_75t_L g4162 ( 
.A(n_3250),
.B(n_3251),
.Y(n_4162)
);

NAND2x1p5_ASAP7_75t_L g4163 ( 
.A(n_3279),
.B(n_3432),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_3614),
.Y(n_4164)
);

CKINVDCx20_ASAP7_75t_R g4165 ( 
.A(n_3556),
.Y(n_4165)
);

CKINVDCx11_ASAP7_75t_R g4166 ( 
.A(n_3570),
.Y(n_4166)
);

AOI22xp33_ASAP7_75t_SL g4167 ( 
.A1(n_3291),
.A2(n_3669),
.B1(n_3625),
.B2(n_3638),
.Y(n_4167)
);

INVx3_ASAP7_75t_L g4168 ( 
.A(n_3198),
.Y(n_4168)
);

AOI22xp33_ASAP7_75t_L g4169 ( 
.A1(n_3418),
.A2(n_3435),
.B1(n_3256),
.B2(n_3250),
.Y(n_4169)
);

AOI22xp33_ASAP7_75t_SL g4170 ( 
.A1(n_3638),
.A2(n_3639),
.B1(n_3418),
.B2(n_3383),
.Y(n_4170)
);

AOI22xp5_ASAP7_75t_L g4171 ( 
.A1(n_3615),
.A2(n_3341),
.B1(n_3354),
.B2(n_3321),
.Y(n_4171)
);

INVx1_ASAP7_75t_SL g4172 ( 
.A(n_3569),
.Y(n_4172)
);

AOI22xp33_ASAP7_75t_L g4173 ( 
.A1(n_3418),
.A2(n_3475),
.B1(n_3453),
.B2(n_3642),
.Y(n_4173)
);

CKINVDCx20_ASAP7_75t_R g4174 ( 
.A(n_3527),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_3616),
.Y(n_4175)
);

BUFx12f_ASAP7_75t_L g4176 ( 
.A(n_3573),
.Y(n_4176)
);

AND2x2_ASAP7_75t_L g4177 ( 
.A(n_3295),
.B(n_3161),
.Y(n_4177)
);

BUFx2_ASAP7_75t_SL g4178 ( 
.A(n_3544),
.Y(n_4178)
);

AOI22xp33_ASAP7_75t_L g4179 ( 
.A1(n_3453),
.A2(n_3475),
.B1(n_3615),
.B2(n_3519),
.Y(n_4179)
);

AND2x4_ASAP7_75t_L g4180 ( 
.A(n_3967),
.B(n_3544),
.Y(n_4180)
);

AND2x2_ASAP7_75t_L g4181 ( 
.A(n_3804),
.B(n_3253),
.Y(n_4181)
);

AOI21x1_ASAP7_75t_SL g4182 ( 
.A1(n_3934),
.A2(n_3576),
.B(n_3656),
.Y(n_4182)
);

OAI22xp5_ASAP7_75t_L g4183 ( 
.A1(n_3694),
.A2(n_3329),
.B1(n_3277),
.B2(n_3253),
.Y(n_4183)
);

AOI21x1_ASAP7_75t_SL g4184 ( 
.A1(n_3934),
.A2(n_3576),
.B(n_3656),
.Y(n_4184)
);

O2A1O1Ixp33_ASAP7_75t_L g4185 ( 
.A1(n_4155),
.A2(n_3348),
.B(n_3523),
.C(n_3557),
.Y(n_4185)
);

AND2x2_ASAP7_75t_L g4186 ( 
.A(n_3963),
.B(n_4177),
.Y(n_4186)
);

AND2x2_ASAP7_75t_L g4187 ( 
.A(n_4177),
.B(n_3277),
.Y(n_4187)
);

OA21x2_ASAP7_75t_L g4188 ( 
.A1(n_3881),
.A2(n_3226),
.B(n_3315),
.Y(n_4188)
);

AND2x2_ASAP7_75t_L g4189 ( 
.A(n_4074),
.B(n_3161),
.Y(n_4189)
);

AND2x2_ASAP7_75t_L g4190 ( 
.A(n_4074),
.B(n_3167),
.Y(n_4190)
);

OR2x2_ASAP7_75t_L g4191 ( 
.A(n_3728),
.B(n_3211),
.Y(n_4191)
);

AND2x2_ASAP7_75t_L g4192 ( 
.A(n_4087),
.B(n_3167),
.Y(n_4192)
);

NAND2xp5_ASAP7_75t_L g4193 ( 
.A(n_3876),
.B(n_3668),
.Y(n_4193)
);

AND2x2_ASAP7_75t_L g4194 ( 
.A(n_4087),
.B(n_3195),
.Y(n_4194)
);

INVx3_ASAP7_75t_L g4195 ( 
.A(n_4010),
.Y(n_4195)
);

AOI21x1_ASAP7_75t_SL g4196 ( 
.A1(n_3876),
.A2(n_3975),
.B(n_3970),
.Y(n_4196)
);

O2A1O1Ixp33_ASAP7_75t_L g4197 ( 
.A1(n_4155),
.A2(n_3557),
.B(n_3524),
.C(n_3220),
.Y(n_4197)
);

AND2x4_ASAP7_75t_SL g4198 ( 
.A(n_3864),
.B(n_3233),
.Y(n_4198)
);

NAND2xp5_ASAP7_75t_L g4199 ( 
.A(n_4086),
.B(n_3668),
.Y(n_4199)
);

OAI22xp5_ASAP7_75t_L g4200 ( 
.A1(n_3714),
.A2(n_3848),
.B1(n_4086),
.B2(n_3728),
.Y(n_4200)
);

AND2x2_ASAP7_75t_L g4201 ( 
.A(n_4096),
.B(n_3195),
.Y(n_4201)
);

AOI21xp5_ASAP7_75t_L g4202 ( 
.A1(n_3881),
.A2(n_3220),
.B(n_3216),
.Y(n_4202)
);

AND2x2_ASAP7_75t_L g4203 ( 
.A(n_4096),
.B(n_3208),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_4127),
.Y(n_4204)
);

AND2x2_ASAP7_75t_L g4205 ( 
.A(n_4097),
.B(n_3788),
.Y(n_4205)
);

AND2x2_ASAP7_75t_L g4206 ( 
.A(n_4097),
.B(n_3788),
.Y(n_4206)
);

AND2x2_ASAP7_75t_L g4207 ( 
.A(n_3697),
.B(n_3208),
.Y(n_4207)
);

OA21x2_ASAP7_75t_L g4208 ( 
.A1(n_3943),
.A2(n_3226),
.B(n_3315),
.Y(n_4208)
);

AND2x4_ASAP7_75t_L g4209 ( 
.A(n_3967),
.B(n_3397),
.Y(n_4209)
);

OAI22xp5_ASAP7_75t_L g4210 ( 
.A1(n_3714),
.A2(n_3329),
.B1(n_3499),
.B2(n_3295),
.Y(n_4210)
);

HB1xp67_ASAP7_75t_L g4211 ( 
.A(n_3919),
.Y(n_4211)
);

INVx1_ASAP7_75t_SL g4212 ( 
.A(n_3890),
.Y(n_4212)
);

OR2x2_ASAP7_75t_L g4213 ( 
.A(n_3733),
.B(n_3211),
.Y(n_4213)
);

NAND2xp5_ASAP7_75t_L g4214 ( 
.A(n_3975),
.B(n_3211),
.Y(n_4214)
);

AND2x2_ASAP7_75t_L g4215 ( 
.A(n_3697),
.B(n_3612),
.Y(n_4215)
);

A2O1A1Ixp33_ASAP7_75t_SL g4216 ( 
.A1(n_4109),
.A2(n_3620),
.B(n_3611),
.C(n_3248),
.Y(n_4216)
);

O2A1O1Ixp33_ASAP7_75t_L g4217 ( 
.A1(n_3848),
.A2(n_3565),
.B(n_3241),
.C(n_3228),
.Y(n_4217)
);

CKINVDCx5p33_ASAP7_75t_R g4218 ( 
.A(n_3687),
.Y(n_4218)
);

INVxp67_ASAP7_75t_L g4219 ( 
.A(n_3997),
.Y(n_4219)
);

CKINVDCx6p67_ASAP7_75t_R g4220 ( 
.A(n_3706),
.Y(n_4220)
);

OAI22xp5_ASAP7_75t_L g4221 ( 
.A1(n_3713),
.A2(n_3228),
.B1(n_3241),
.B2(n_3321),
.Y(n_4221)
);

AND2x2_ASAP7_75t_L g4222 ( 
.A(n_3965),
.B(n_3612),
.Y(n_4222)
);

AND2x2_ASAP7_75t_L g4223 ( 
.A(n_3965),
.B(n_3558),
.Y(n_4223)
);

AND2x4_ASAP7_75t_L g4224 ( 
.A(n_3967),
.B(n_3397),
.Y(n_4224)
);

HB1xp67_ASAP7_75t_L g4225 ( 
.A(n_4143),
.Y(n_4225)
);

AND2x2_ASAP7_75t_L g4226 ( 
.A(n_3981),
.B(n_3558),
.Y(n_4226)
);

INVx2_ASAP7_75t_L g4227 ( 
.A(n_3741),
.Y(n_4227)
);

AOI21xp5_ASAP7_75t_L g4228 ( 
.A1(n_4128),
.A2(n_4149),
.B(n_4105),
.Y(n_4228)
);

OA21x2_ASAP7_75t_L g4229 ( 
.A1(n_3943),
.A2(n_3226),
.B(n_3246),
.Y(n_4229)
);

INVx2_ASAP7_75t_L g4230 ( 
.A(n_3741),
.Y(n_4230)
);

OAI22xp5_ASAP7_75t_L g4231 ( 
.A1(n_3878),
.A2(n_3354),
.B1(n_3355),
.B2(n_3341),
.Y(n_4231)
);

NOR2xp67_ASAP7_75t_L g4232 ( 
.A(n_3809),
.B(n_3633),
.Y(n_4232)
);

AOI21x1_ASAP7_75t_SL g4233 ( 
.A1(n_3970),
.A2(n_3555),
.B(n_3553),
.Y(n_4233)
);

OR2x2_ASAP7_75t_L g4234 ( 
.A(n_3733),
.B(n_3211),
.Y(n_4234)
);

OAI22xp5_ASAP7_75t_L g4235 ( 
.A1(n_3878),
.A2(n_3380),
.B1(n_3395),
.B2(n_3355),
.Y(n_4235)
);

AO21x1_ASAP7_75t_L g4236 ( 
.A1(n_4105),
.A2(n_3651),
.B(n_3633),
.Y(n_4236)
);

INVxp33_ASAP7_75t_SL g4237 ( 
.A(n_4011),
.Y(n_4237)
);

A2O1A1Ixp33_ASAP7_75t_L g4238 ( 
.A1(n_3836),
.A2(n_3623),
.B(n_3651),
.C(n_3248),
.Y(n_4238)
);

INVx2_ASAP7_75t_L g4239 ( 
.A(n_3741),
.Y(n_4239)
);

OR2x2_ASAP7_75t_L g4240 ( 
.A(n_3776),
.B(n_3211),
.Y(n_4240)
);

OA22x2_ASAP7_75t_L g4241 ( 
.A1(n_4115),
.A2(n_3519),
.B1(n_3286),
.B2(n_3639),
.Y(n_4241)
);

AND2x2_ASAP7_75t_L g4242 ( 
.A(n_3981),
.B(n_3560),
.Y(n_4242)
);

O2A1O1Ixp5_ASAP7_75t_L g4243 ( 
.A1(n_4115),
.A2(n_3585),
.B(n_3623),
.C(n_3620),
.Y(n_4243)
);

OAI22xp5_ASAP7_75t_L g4244 ( 
.A1(n_3980),
.A2(n_3380),
.B1(n_3407),
.B2(n_3395),
.Y(n_4244)
);

NAND2xp5_ASAP7_75t_L g4245 ( 
.A(n_3730),
.B(n_3211),
.Y(n_4245)
);

OAI22xp5_ASAP7_75t_L g4246 ( 
.A1(n_3980),
.A2(n_3407),
.B1(n_3420),
.B2(n_3412),
.Y(n_4246)
);

OR2x2_ASAP7_75t_L g4247 ( 
.A(n_3776),
.B(n_3527),
.Y(n_4247)
);

NAND2xp5_ASAP7_75t_L g4248 ( 
.A(n_3730),
.B(n_3643),
.Y(n_4248)
);

CKINVDCx5p33_ASAP7_75t_R g4249 ( 
.A(n_3711),
.Y(n_4249)
);

BUFx3_ASAP7_75t_L g4250 ( 
.A(n_3706),
.Y(n_4250)
);

INVx2_ASAP7_75t_L g4251 ( 
.A(n_3745),
.Y(n_4251)
);

BUFx2_ASAP7_75t_L g4252 ( 
.A(n_4152),
.Y(n_4252)
);

AOI21xp5_ASAP7_75t_SL g4253 ( 
.A1(n_4109),
.A2(n_3772),
.B(n_3937),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_L g4254 ( 
.A(n_3823),
.B(n_3643),
.Y(n_4254)
);

NAND2xp5_ASAP7_75t_L g4255 ( 
.A(n_3823),
.B(n_3593),
.Y(n_4255)
);

AOI21xp5_ASAP7_75t_SL g4256 ( 
.A1(n_3772),
.A2(n_3654),
.B(n_3655),
.Y(n_4256)
);

NAND2xp5_ASAP7_75t_L g4257 ( 
.A(n_4141),
.B(n_3593),
.Y(n_4257)
);

BUFx6f_ASAP7_75t_L g4258 ( 
.A(n_3720),
.Y(n_4258)
);

HB1xp67_ASAP7_75t_L g4259 ( 
.A(n_4143),
.Y(n_4259)
);

INVx2_ASAP7_75t_L g4260 ( 
.A(n_3745),
.Y(n_4260)
);

OR2x2_ASAP7_75t_L g4261 ( 
.A(n_3760),
.B(n_3412),
.Y(n_4261)
);

A2O1A1Ixp33_ASAP7_75t_SL g4262 ( 
.A1(n_3985),
.A2(n_3611),
.B(n_3246),
.C(n_3646),
.Y(n_4262)
);

INVx2_ASAP7_75t_L g4263 ( 
.A(n_3745),
.Y(n_4263)
);

AOI21xp5_ASAP7_75t_L g4264 ( 
.A1(n_4128),
.A2(n_3386),
.B(n_3387),
.Y(n_4264)
);

OA21x2_ASAP7_75t_L g4265 ( 
.A1(n_4008),
.A2(n_3703),
.B(n_4047),
.Y(n_4265)
);

AOI21xp5_ASAP7_75t_SL g4266 ( 
.A1(n_3937),
.A2(n_3402),
.B(n_3401),
.Y(n_4266)
);

OR2x2_ASAP7_75t_L g4267 ( 
.A(n_3760),
.B(n_3916),
.Y(n_4267)
);

AND2x4_ASAP7_75t_L g4268 ( 
.A(n_3967),
.B(n_3403),
.Y(n_4268)
);

AOI21xp5_ASAP7_75t_SL g4269 ( 
.A1(n_3865),
.A2(n_3429),
.B(n_3402),
.Y(n_4269)
);

OA21x2_ASAP7_75t_L g4270 ( 
.A1(n_4008),
.A2(n_3371),
.B(n_3482),
.Y(n_4270)
);

NOR2xp67_ASAP7_75t_L g4271 ( 
.A(n_3809),
.B(n_4142),
.Y(n_4271)
);

OR2x2_ASAP7_75t_L g4272 ( 
.A(n_3916),
.B(n_3420),
.Y(n_4272)
);

OA21x2_ASAP7_75t_L g4273 ( 
.A1(n_3703),
.A2(n_3371),
.B(n_3482),
.Y(n_4273)
);

OA21x2_ASAP7_75t_L g4274 ( 
.A1(n_4047),
.A2(n_3371),
.B(n_3482),
.Y(n_4274)
);

O2A1O1Ixp33_ASAP7_75t_L g4275 ( 
.A1(n_3724),
.A2(n_3489),
.B(n_3422),
.C(n_3477),
.Y(n_4275)
);

CKINVDCx9p33_ASAP7_75t_R g4276 ( 
.A(n_4011),
.Y(n_4276)
);

INVx2_ASAP7_75t_L g4277 ( 
.A(n_3763),
.Y(n_4277)
);

INVx1_ASAP7_75t_L g4278 ( 
.A(n_4127),
.Y(n_4278)
);

AND2x2_ASAP7_75t_L g4279 ( 
.A(n_3908),
.B(n_3560),
.Y(n_4279)
);

INVx2_ASAP7_75t_L g4280 ( 
.A(n_3763),
.Y(n_4280)
);

INVx1_ASAP7_75t_L g4281 ( 
.A(n_4131),
.Y(n_4281)
);

INVx2_ASAP7_75t_L g4282 ( 
.A(n_3763),
.Y(n_4282)
);

OA21x2_ASAP7_75t_L g4283 ( 
.A1(n_3985),
.A2(n_3386),
.B(n_3393),
.Y(n_4283)
);

AND2x2_ASAP7_75t_L g4284 ( 
.A(n_3908),
.B(n_3596),
.Y(n_4284)
);

O2A1O1Ixp5_ASAP7_75t_L g4285 ( 
.A1(n_3865),
.A2(n_3679),
.B(n_3698),
.C(n_3958),
.Y(n_4285)
);

OAI22xp5_ASAP7_75t_L g4286 ( 
.A1(n_3836),
.A2(n_3489),
.B1(n_3550),
.B2(n_3485),
.Y(n_4286)
);

OAI22xp5_ASAP7_75t_L g4287 ( 
.A1(n_3720),
.A2(n_3440),
.B1(n_3550),
.B2(n_3583),
.Y(n_4287)
);

OR2x2_ASAP7_75t_L g4288 ( 
.A(n_3990),
.B(n_3422),
.Y(n_4288)
);

AOI21xp5_ASAP7_75t_L g4289 ( 
.A1(n_4149),
.A2(n_3391),
.B(n_3387),
.Y(n_4289)
);

INVx2_ASAP7_75t_L g4290 ( 
.A(n_3811),
.Y(n_4290)
);

AOI21xp5_ASAP7_75t_L g4291 ( 
.A1(n_3887),
.A2(n_3391),
.B(n_3393),
.Y(n_4291)
);

A2O1A1Ixp33_ASAP7_75t_L g4292 ( 
.A1(n_3947),
.A2(n_3639),
.B(n_3441),
.C(n_3445),
.Y(n_4292)
);

O2A1O1Ixp33_ASAP7_75t_L g4293 ( 
.A1(n_4119),
.A2(n_3575),
.B(n_3497),
.C(n_3568),
.Y(n_4293)
);

O2A1O1Ixp33_ASAP7_75t_L g4294 ( 
.A1(n_4119),
.A2(n_3582),
.B(n_3483),
.C(n_3497),
.Y(n_4294)
);

NAND2xp5_ASAP7_75t_L g4295 ( 
.A(n_4141),
.B(n_3440),
.Y(n_4295)
);

OA21x2_ASAP7_75t_L g4296 ( 
.A1(n_3679),
.A2(n_3382),
.B(n_3340),
.Y(n_4296)
);

AND2x2_ASAP7_75t_L g4297 ( 
.A(n_3911),
.B(n_3596),
.Y(n_4297)
);

O2A1O1Ixp33_ASAP7_75t_L g4298 ( 
.A1(n_3698),
.A2(n_3583),
.B(n_3485),
.C(n_3568),
.Y(n_4298)
);

NAND2xp5_ASAP7_75t_L g4299 ( 
.A(n_4145),
.B(n_3477),
.Y(n_4299)
);

NOR2xp67_ASAP7_75t_L g4300 ( 
.A(n_4142),
.B(n_3198),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_4131),
.Y(n_4301)
);

AND2x6_ASAP7_75t_L g4302 ( 
.A(n_4010),
.B(n_3233),
.Y(n_4302)
);

AND2x4_ASAP7_75t_SL g4303 ( 
.A(n_3864),
.B(n_3233),
.Y(n_4303)
);

OAI22xp5_ASAP7_75t_L g4304 ( 
.A1(n_3720),
.A2(n_3582),
.B1(n_3529),
.B2(n_3483),
.Y(n_4304)
);

BUFx12f_ASAP7_75t_L g4305 ( 
.A(n_3706),
.Y(n_4305)
);

OAI22xp5_ASAP7_75t_L g4306 ( 
.A1(n_4171),
.A2(n_3575),
.B1(n_3529),
.B2(n_3498),
.Y(n_4306)
);

AOI21xp5_ASAP7_75t_L g4307 ( 
.A1(n_3887),
.A2(n_3972),
.B(n_3956),
.Y(n_4307)
);

HB1xp67_ASAP7_75t_L g4308 ( 
.A(n_4057),
.Y(n_4308)
);

BUFx3_ASAP7_75t_L g4309 ( 
.A(n_3688),
.Y(n_4309)
);

AND2x4_ASAP7_75t_L g4310 ( 
.A(n_4144),
.B(n_3403),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_L g4311 ( 
.A(n_4145),
.B(n_3498),
.Y(n_4311)
);

OAI22xp5_ASAP7_75t_L g4312 ( 
.A1(n_4171),
.A2(n_3573),
.B1(n_3530),
.B2(n_3510),
.Y(n_4312)
);

AND2x2_ASAP7_75t_L g4313 ( 
.A(n_3911),
.B(n_4172),
.Y(n_4313)
);

OAI211xp5_ASAP7_75t_L g4314 ( 
.A1(n_4167),
.A2(n_3658),
.B(n_3382),
.C(n_3340),
.Y(n_4314)
);

OR2x2_ASAP7_75t_L g4315 ( 
.A(n_3990),
.B(n_3510),
.Y(n_4315)
);

O2A1O1Ixp5_ASAP7_75t_L g4316 ( 
.A1(n_4000),
.A2(n_3607),
.B(n_3616),
.C(n_3579),
.Y(n_4316)
);

OA21x2_ASAP7_75t_L g4317 ( 
.A1(n_4054),
.A2(n_3410),
.B(n_3409),
.Y(n_4317)
);

OAI22xp5_ASAP7_75t_L g4318 ( 
.A1(n_3719),
.A2(n_3573),
.B1(n_3530),
.B2(n_3607),
.Y(n_4318)
);

CKINVDCx5p33_ASAP7_75t_R g4319 ( 
.A(n_3736),
.Y(n_4319)
);

AND2x2_ASAP7_75t_L g4320 ( 
.A(n_4172),
.B(n_3596),
.Y(n_4320)
);

OAI22xp5_ASAP7_75t_L g4321 ( 
.A1(n_3719),
.A2(n_3573),
.B1(n_3672),
.B2(n_3467),
.Y(n_4321)
);

NAND2xp5_ASAP7_75t_L g4322 ( 
.A(n_4000),
.B(n_3645),
.Y(n_4322)
);

OA21x2_ASAP7_75t_L g4323 ( 
.A1(n_4040),
.A2(n_3843),
.B(n_3814),
.Y(n_4323)
);

AND2x2_ASAP7_75t_L g4324 ( 
.A(n_4144),
.B(n_3596),
.Y(n_4324)
);

AND2x2_ASAP7_75t_L g4325 ( 
.A(n_3735),
.B(n_3755),
.Y(n_4325)
);

INVx2_ASAP7_75t_L g4326 ( 
.A(n_3811),
.Y(n_4326)
);

O2A1O1Ixp5_ASAP7_75t_L g4327 ( 
.A1(n_4003),
.A2(n_3579),
.B(n_3660),
.C(n_3645),
.Y(n_4327)
);

CKINVDCx5p33_ASAP7_75t_R g4328 ( 
.A(n_3754),
.Y(n_4328)
);

INVxp67_ASAP7_75t_SL g4329 ( 
.A(n_4031),
.Y(n_4329)
);

O2A1O1Ixp5_ASAP7_75t_L g4330 ( 
.A1(n_4003),
.A2(n_3660),
.B(n_3590),
.C(n_3588),
.Y(n_4330)
);

NAND2xp5_ASAP7_75t_L g4331 ( 
.A(n_4161),
.B(n_3569),
.Y(n_4331)
);

OA21x2_ASAP7_75t_L g4332 ( 
.A1(n_3814),
.A2(n_3410),
.B(n_3409),
.Y(n_4332)
);

OA21x2_ASAP7_75t_L g4333 ( 
.A1(n_3843),
.A2(n_3421),
.B(n_3425),
.Y(n_4333)
);

AND2x2_ASAP7_75t_L g4334 ( 
.A(n_3735),
.B(n_3588),
.Y(n_4334)
);

NAND2xp5_ASAP7_75t_L g4335 ( 
.A(n_4161),
.B(n_3592),
.Y(n_4335)
);

OAI22xp5_ASAP7_75t_L g4336 ( 
.A1(n_4167),
.A2(n_4179),
.B1(n_4089),
.B2(n_3690),
.Y(n_4336)
);

OAI22xp5_ASAP7_75t_L g4337 ( 
.A1(n_4089),
.A2(n_3672),
.B1(n_3480),
.B2(n_3467),
.Y(n_4337)
);

CKINVDCx11_ASAP7_75t_R g4338 ( 
.A(n_3769),
.Y(n_4338)
);

HB1xp67_ASAP7_75t_L g4339 ( 
.A(n_4057),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_SL g4340 ( 
.A(n_4126),
.B(n_3233),
.Y(n_4340)
);

NAND2xp5_ASAP7_75t_L g4341 ( 
.A(n_4164),
.B(n_3592),
.Y(n_4341)
);

INVx1_ASAP7_75t_L g4342 ( 
.A(n_4132),
.Y(n_4342)
);

AOI21xp5_ASAP7_75t_SL g4343 ( 
.A1(n_4163),
.A2(n_3429),
.B(n_3402),
.Y(n_4343)
);

AND2x2_ASAP7_75t_L g4344 ( 
.A(n_3755),
.B(n_3588),
.Y(n_4344)
);

OAI22xp5_ASAP7_75t_L g4345 ( 
.A1(n_3690),
.A2(n_3672),
.B1(n_3480),
.B2(n_3429),
.Y(n_4345)
);

AOI21xp5_ASAP7_75t_L g4346 ( 
.A1(n_3972),
.A2(n_3466),
.B(n_3425),
.Y(n_4346)
);

OAI22xp5_ASAP7_75t_L g4347 ( 
.A1(n_4174),
.A2(n_4118),
.B1(n_4101),
.B2(n_3954),
.Y(n_4347)
);

AND2x4_ASAP7_75t_L g4348 ( 
.A(n_4010),
.B(n_3727),
.Y(n_4348)
);

AOI211xp5_ASAP7_75t_L g4349 ( 
.A1(n_3956),
.A2(n_3658),
.B(n_3644),
.C(n_3271),
.Y(n_4349)
);

O2A1O1Ixp33_ASAP7_75t_L g4350 ( 
.A1(n_4025),
.A2(n_3673),
.B(n_3324),
.C(n_3221),
.Y(n_4350)
);

A2O1A1Ixp33_ASAP7_75t_L g4351 ( 
.A1(n_3947),
.A2(n_3441),
.B(n_3445),
.C(n_3279),
.Y(n_4351)
);

AOI21xp5_ASAP7_75t_L g4352 ( 
.A1(n_3831),
.A2(n_3474),
.B(n_3466),
.Y(n_4352)
);

AOI221xp5_ASAP7_75t_L g4353 ( 
.A1(n_4081),
.A2(n_3441),
.B1(n_3445),
.B2(n_3324),
.C(n_3271),
.Y(n_4353)
);

NAND2xp5_ASAP7_75t_L g4354 ( 
.A(n_4164),
.B(n_3221),
.Y(n_4354)
);

OR2x2_ASAP7_75t_L g4355 ( 
.A(n_3993),
.B(n_3344),
.Y(n_4355)
);

INVx2_ASAP7_75t_L g4356 ( 
.A(n_3811),
.Y(n_4356)
);

AOI21xp5_ASAP7_75t_SL g4357 ( 
.A1(n_4163),
.A2(n_3906),
.B(n_3820),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_4132),
.Y(n_4358)
);

OA21x2_ASAP7_75t_L g4359 ( 
.A1(n_4065),
.A2(n_3421),
.B(n_3474),
.Y(n_4359)
);

BUFx2_ASAP7_75t_L g4360 ( 
.A(n_4152),
.Y(n_4360)
);

OAI22xp5_ASAP7_75t_L g4361 ( 
.A1(n_4101),
.A2(n_3231),
.B1(n_3259),
.B2(n_3304),
.Y(n_4361)
);

OAI22xp5_ASAP7_75t_L g4362 ( 
.A1(n_3792),
.A2(n_3231),
.B1(n_3259),
.B2(n_3304),
.Y(n_4362)
);

OR2x2_ASAP7_75t_L g4363 ( 
.A(n_3993),
.B(n_3344),
.Y(n_4363)
);

INVx1_ASAP7_75t_L g4364 ( 
.A(n_4139),
.Y(n_4364)
);

A2O1A1Ixp33_ASAP7_75t_L g4365 ( 
.A1(n_4081),
.A2(n_3441),
.B(n_3445),
.C(n_3158),
.Y(n_4365)
);

AOI21xp5_ASAP7_75t_SL g4366 ( 
.A1(n_4163),
.A2(n_3567),
.B(n_3514),
.Y(n_4366)
);

O2A1O1Ixp33_ASAP7_75t_L g4367 ( 
.A1(n_3726),
.A2(n_3644),
.B(n_3324),
.C(n_3271),
.Y(n_4367)
);

NOR2xp67_ASAP7_75t_L g4368 ( 
.A(n_3727),
.B(n_3221),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_4139),
.Y(n_4369)
);

AOI21x1_ASAP7_75t_SL g4370 ( 
.A1(n_4031),
.A2(n_3671),
.B(n_3660),
.Y(n_4370)
);

HB1xp67_ASAP7_75t_L g4371 ( 
.A(n_4130),
.Y(n_4371)
);

OAI31xp33_ASAP7_75t_L g4372 ( 
.A1(n_3770),
.A2(n_3664),
.A3(n_3383),
.B(n_3514),
.Y(n_4372)
);

NOR2x1_ASAP7_75t_SL g4373 ( 
.A(n_4178),
.B(n_3862),
.Y(n_4373)
);

AND2x2_ASAP7_75t_L g4374 ( 
.A(n_3839),
.B(n_3588),
.Y(n_4374)
);

AND2x2_ASAP7_75t_L g4375 ( 
.A(n_3839),
.B(n_3590),
.Y(n_4375)
);

OR2x2_ASAP7_75t_L g4376 ( 
.A(n_4076),
.B(n_3362),
.Y(n_4376)
);

AOI21xp5_ASAP7_75t_L g4377 ( 
.A1(n_3831),
.A2(n_3534),
.B(n_3493),
.Y(n_4377)
);

INVx4_ASAP7_75t_L g4378 ( 
.A(n_3889),
.Y(n_4378)
);

OA21x2_ASAP7_75t_L g4379 ( 
.A1(n_4066),
.A2(n_3534),
.B(n_3493),
.Y(n_4379)
);

AOI21xp5_ASAP7_75t_L g4380 ( 
.A1(n_3835),
.A2(n_3906),
.B(n_4140),
.Y(n_4380)
);

NAND2xp5_ASAP7_75t_L g4381 ( 
.A(n_4175),
.B(n_3221),
.Y(n_4381)
);

NAND2xp5_ASAP7_75t_L g4382 ( 
.A(n_4175),
.B(n_3271),
.Y(n_4382)
);

OA21x2_ASAP7_75t_L g4383 ( 
.A1(n_4068),
.A2(n_3547),
.B(n_3586),
.Y(n_4383)
);

OR2x2_ASAP7_75t_L g4384 ( 
.A(n_4076),
.B(n_3362),
.Y(n_4384)
);

OR2x2_ASAP7_75t_L g4385 ( 
.A(n_4072),
.B(n_3439),
.Y(n_4385)
);

AND2x2_ASAP7_75t_L g4386 ( 
.A(n_3863),
.B(n_3882),
.Y(n_4386)
);

OAI22xp5_ASAP7_75t_L g4387 ( 
.A1(n_3792),
.A2(n_3590),
.B1(n_3519),
.B2(n_3570),
.Y(n_4387)
);

BUFx2_ASAP7_75t_L g4388 ( 
.A(n_4152),
.Y(n_4388)
);

AND2x4_ASAP7_75t_L g4389 ( 
.A(n_4010),
.B(n_3727),
.Y(n_4389)
);

AOI21x1_ASAP7_75t_SL g4390 ( 
.A1(n_4072),
.A2(n_3671),
.B(n_3660),
.Y(n_4390)
);

AOI21xp5_ASAP7_75t_SL g4391 ( 
.A1(n_3820),
.A2(n_3567),
.B(n_3514),
.Y(n_4391)
);

O2A1O1Ixp5_ASAP7_75t_L g4392 ( 
.A1(n_3746),
.A2(n_3590),
.B(n_3664),
.C(n_3470),
.Y(n_4392)
);

OAI22xp5_ASAP7_75t_L g4393 ( 
.A1(n_3835),
.A2(n_3519),
.B1(n_3570),
.B2(n_3584),
.Y(n_4393)
);

AND2x2_ASAP7_75t_L g4394 ( 
.A(n_3863),
.B(n_3584),
.Y(n_4394)
);

CKINVDCx20_ASAP7_75t_R g4395 ( 
.A(n_3805),
.Y(n_4395)
);

BUFx3_ASAP7_75t_L g4396 ( 
.A(n_3688),
.Y(n_4396)
);

NAND2xp5_ASAP7_75t_L g4397 ( 
.A(n_4100),
.B(n_3324),
.Y(n_4397)
);

AOI21xp5_ASAP7_75t_L g4398 ( 
.A1(n_4140),
.A2(n_3903),
.B(n_3731),
.Y(n_4398)
);

INVx5_ASAP7_75t_L g4399 ( 
.A(n_3696),
.Y(n_4399)
);

A2O1A1Ixp33_ASAP7_75t_SL g4400 ( 
.A1(n_3777),
.A2(n_3676),
.B(n_3459),
.C(n_3416),
.Y(n_4400)
);

O2A1O1Ixp33_ASAP7_75t_L g4401 ( 
.A1(n_3726),
.A2(n_3598),
.B(n_3586),
.C(n_3580),
.Y(n_4401)
);

A2O1A1Ixp33_ASAP7_75t_L g4402 ( 
.A1(n_4063),
.A2(n_3158),
.B(n_3173),
.C(n_3403),
.Y(n_4402)
);

AND2x2_ASAP7_75t_L g4403 ( 
.A(n_3882),
.B(n_3584),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_3683),
.Y(n_4404)
);

AOI21xp5_ASAP7_75t_L g4405 ( 
.A1(n_3903),
.A2(n_3571),
.B(n_3661),
.Y(n_4405)
);

O2A1O1Ixp5_ASAP7_75t_L g4406 ( 
.A1(n_3746),
.A2(n_3470),
.B(n_3507),
.C(n_3495),
.Y(n_4406)
);

AND2x4_ASAP7_75t_L g4407 ( 
.A(n_3727),
.B(n_3403),
.Y(n_4407)
);

AND2x4_ASAP7_75t_L g4408 ( 
.A(n_3727),
.B(n_3245),
.Y(n_4408)
);

O2A1O1Ixp5_ASAP7_75t_L g4409 ( 
.A1(n_3785),
.A2(n_3507),
.B(n_3470),
.C(n_3495),
.Y(n_4409)
);

INVx2_ASAP7_75t_L g4410 ( 
.A(n_3816),
.Y(n_4410)
);

O2A1O1Ixp33_ASAP7_75t_L g4411 ( 
.A1(n_3747),
.A2(n_3598),
.B(n_3580),
.C(n_3571),
.Y(n_4411)
);

NOR2xp67_ASAP7_75t_L g4412 ( 
.A(n_3727),
.B(n_3597),
.Y(n_4412)
);

NAND2xp5_ASAP7_75t_L g4413 ( 
.A(n_4100),
.B(n_3439),
.Y(n_4413)
);

OR2x2_ASAP7_75t_L g4414 ( 
.A(n_4153),
.B(n_3442),
.Y(n_4414)
);

OA21x2_ASAP7_75t_L g4415 ( 
.A1(n_4073),
.A2(n_3547),
.B(n_3659),
.Y(n_4415)
);

OA21x2_ASAP7_75t_L g4416 ( 
.A1(n_3896),
.A2(n_3661),
.B(n_3659),
.Y(n_4416)
);

OA21x2_ASAP7_75t_L g4417 ( 
.A1(n_3942),
.A2(n_3303),
.B(n_3376),
.Y(n_4417)
);

O2A1O1Ixp33_ASAP7_75t_L g4418 ( 
.A1(n_3747),
.A2(n_3636),
.B(n_3442),
.C(n_3608),
.Y(n_4418)
);

INVx2_ASAP7_75t_L g4419 ( 
.A(n_3816),
.Y(n_4419)
);

OAI22xp5_ASAP7_75t_L g4420 ( 
.A1(n_4129),
.A2(n_3519),
.B1(n_3584),
.B2(n_3577),
.Y(n_4420)
);

AOI21xp5_ASAP7_75t_SL g4421 ( 
.A1(n_3705),
.A2(n_3567),
.B(n_3158),
.Y(n_4421)
);

OAI211xp5_ASAP7_75t_L g4422 ( 
.A1(n_4133),
.A2(n_3492),
.B(n_3376),
.C(n_3629),
.Y(n_4422)
);

INVxp67_ASAP7_75t_L g4423 ( 
.A(n_3699),
.Y(n_4423)
);

O2A1O1Ixp5_ASAP7_75t_L g4424 ( 
.A1(n_3977),
.A2(n_3932),
.B(n_3750),
.C(n_3924),
.Y(n_4424)
);

AOI21xp5_ASAP7_75t_L g4425 ( 
.A1(n_3731),
.A2(n_3567),
.B(n_3492),
.Y(n_4425)
);

BUFx2_ASAP7_75t_L g4426 ( 
.A(n_3860),
.Y(n_4426)
);

AND2x2_ASAP7_75t_L g4427 ( 
.A(n_4039),
.B(n_3512),
.Y(n_4427)
);

AND2x2_ASAP7_75t_L g4428 ( 
.A(n_4039),
.B(n_3512),
.Y(n_4428)
);

AOI21xp5_ASAP7_75t_SL g4429 ( 
.A1(n_3705),
.A2(n_3173),
.B(n_3640),
.Y(n_4429)
);

BUFx6f_ASAP7_75t_L g4430 ( 
.A(n_3708),
.Y(n_4430)
);

OR2x2_ASAP7_75t_L g4431 ( 
.A(n_4153),
.B(n_3595),
.Y(n_4431)
);

NAND2xp5_ASAP7_75t_L g4432 ( 
.A(n_4162),
.B(n_3632),
.Y(n_4432)
);

BUFx3_ASAP7_75t_L g4433 ( 
.A(n_3688),
.Y(n_4433)
);

AOI21xp5_ASAP7_75t_SL g4434 ( 
.A1(n_3705),
.A2(n_3173),
.B(n_3640),
.Y(n_4434)
);

AND2x2_ASAP7_75t_L g4435 ( 
.A(n_4043),
.B(n_3512),
.Y(n_4435)
);

AND2x2_ASAP7_75t_L g4436 ( 
.A(n_4043),
.B(n_3564),
.Y(n_4436)
);

HB1xp67_ASAP7_75t_L g4437 ( 
.A(n_4130),
.Y(n_4437)
);

OA21x2_ASAP7_75t_L g4438 ( 
.A1(n_3942),
.A2(n_3303),
.B(n_3653),
.Y(n_4438)
);

AND2x4_ASAP7_75t_L g4439 ( 
.A(n_3727),
.B(n_3245),
.Y(n_4439)
);

OAI22xp5_ASAP7_75t_L g4440 ( 
.A1(n_4134),
.A2(n_3944),
.B1(n_4165),
.B2(n_4159),
.Y(n_4440)
);

O2A1O1Ixp5_ASAP7_75t_L g4441 ( 
.A1(n_3932),
.A2(n_3470),
.B(n_3507),
.C(n_3495),
.Y(n_4441)
);

BUFx6f_ASAP7_75t_L g4442 ( 
.A(n_3708),
.Y(n_4442)
);

BUFx2_ASAP7_75t_R g4443 ( 
.A(n_3821),
.Y(n_4443)
);

OA21x2_ASAP7_75t_L g4444 ( 
.A1(n_4037),
.A2(n_3640),
.B(n_3653),
.Y(n_4444)
);

AOI21xp5_ASAP7_75t_L g4445 ( 
.A1(n_3944),
.A2(n_3753),
.B(n_3933),
.Y(n_4445)
);

OA21x2_ASAP7_75t_L g4446 ( 
.A1(n_4062),
.A2(n_3640),
.B(n_3653),
.Y(n_4446)
);

OR2x2_ASAP7_75t_L g4447 ( 
.A(n_4162),
.B(n_3595),
.Y(n_4447)
);

INVx1_ASAP7_75t_L g4448 ( 
.A(n_3683),
.Y(n_4448)
);

INVx1_ASAP7_75t_L g4449 ( 
.A(n_3686),
.Y(n_4449)
);

OR2x2_ASAP7_75t_L g4450 ( 
.A(n_4009),
.B(n_4020),
.Y(n_4450)
);

OAI22xp5_ASAP7_75t_L g4451 ( 
.A1(n_3752),
.A2(n_3577),
.B1(n_3204),
.B2(n_3411),
.Y(n_4451)
);

OAI22xp5_ASAP7_75t_L g4452 ( 
.A1(n_4099),
.A2(n_3577),
.B1(n_3204),
.B2(n_3411),
.Y(n_4452)
);

AND2x2_ASAP7_75t_L g4453 ( 
.A(n_4071),
.B(n_4106),
.Y(n_4453)
);

OR2x2_ASAP7_75t_L g4454 ( 
.A(n_4009),
.B(n_3604),
.Y(n_4454)
);

INVx3_ASAP7_75t_L g4455 ( 
.A(n_3777),
.Y(n_4455)
);

INVx1_ASAP7_75t_L g4456 ( 
.A(n_3686),
.Y(n_4456)
);

OA21x2_ASAP7_75t_L g4457 ( 
.A1(n_4036),
.A2(n_3653),
.B(n_3629),
.Y(n_4457)
);

INVx1_ASAP7_75t_L g4458 ( 
.A(n_3691),
.Y(n_4458)
);

AND2x2_ASAP7_75t_L g4459 ( 
.A(n_4071),
.B(n_3564),
.Y(n_4459)
);

HB1xp67_ASAP7_75t_L g4460 ( 
.A(n_4135),
.Y(n_4460)
);

OA21x2_ASAP7_75t_L g4461 ( 
.A1(n_3978),
.A2(n_3604),
.B(n_3647),
.Y(n_4461)
);

OAI22xp5_ASAP7_75t_L g4462 ( 
.A1(n_3794),
.A2(n_3577),
.B1(n_3204),
.B2(n_3456),
.Y(n_4462)
);

AND2x2_ASAP7_75t_L g4463 ( 
.A(n_4106),
.B(n_3564),
.Y(n_4463)
);

O2A1O1Ixp5_ASAP7_75t_L g4464 ( 
.A1(n_3750),
.A2(n_3495),
.B(n_3507),
.C(n_3572),
.Y(n_4464)
);

AND2x2_ASAP7_75t_L g4465 ( 
.A(n_3891),
.B(n_3572),
.Y(n_4465)
);

AOI21xp5_ASAP7_75t_SL g4466 ( 
.A1(n_3960),
.A2(n_3432),
.B(n_3267),
.Y(n_4466)
);

OAI22xp5_ASAP7_75t_L g4467 ( 
.A1(n_3791),
.A2(n_3732),
.B1(n_3973),
.B2(n_3678),
.Y(n_4467)
);

NAND2xp5_ASAP7_75t_L g4468 ( 
.A(n_3684),
.B(n_3632),
.Y(n_4468)
);

OA22x2_ASAP7_75t_L g4469 ( 
.A1(n_3918),
.A2(n_3286),
.B1(n_3325),
.B2(n_3394),
.Y(n_4469)
);

NAND2xp5_ASAP7_75t_L g4470 ( 
.A(n_3684),
.B(n_3647),
.Y(n_4470)
);

O2A1O1Ixp5_ASAP7_75t_L g4471 ( 
.A1(n_3924),
.A2(n_3572),
.B(n_3602),
.C(n_3589),
.Y(n_4471)
);

O2A1O1Ixp5_ASAP7_75t_L g4472 ( 
.A1(n_3827),
.A2(n_3572),
.B(n_3602),
.C(n_3589),
.Y(n_4472)
);

O2A1O1Ixp5_ASAP7_75t_L g4473 ( 
.A1(n_3723),
.A2(n_3676),
.B(n_3602),
.C(n_3589),
.Y(n_4473)
);

OA21x2_ASAP7_75t_L g4474 ( 
.A1(n_3978),
.A2(n_3648),
.B(n_3665),
.Y(n_4474)
);

CKINVDCx5p33_ASAP7_75t_R g4475 ( 
.A(n_3689),
.Y(n_4475)
);

OAI22xp5_ASAP7_75t_L g4476 ( 
.A1(n_3973),
.A2(n_3678),
.B1(n_3680),
.B2(n_3797),
.Y(n_4476)
);

A2O1A1Ixp33_ASAP7_75t_L g4477 ( 
.A1(n_4063),
.A2(n_3383),
.B(n_3286),
.C(n_3267),
.Y(n_4477)
);

INVx2_ASAP7_75t_L g4478 ( 
.A(n_3816),
.Y(n_4478)
);

INVxp33_ASAP7_75t_L g4479 ( 
.A(n_4060),
.Y(n_4479)
);

AND2x2_ASAP7_75t_L g4480 ( 
.A(n_3891),
.B(n_3648),
.Y(n_4480)
);

OR2x2_ASAP7_75t_L g4481 ( 
.A(n_4020),
.B(n_3608),
.Y(n_4481)
);

OR2x2_ASAP7_75t_L g4482 ( 
.A(n_3693),
.B(n_3608),
.Y(n_4482)
);

BUFx3_ASAP7_75t_L g4483 ( 
.A(n_3688),
.Y(n_4483)
);

INVx1_ASAP7_75t_L g4484 ( 
.A(n_3691),
.Y(n_4484)
);

INVx2_ASAP7_75t_L g4485 ( 
.A(n_3830),
.Y(n_4485)
);

BUFx2_ASAP7_75t_L g4486 ( 
.A(n_3969),
.Y(n_4486)
);

INVx2_ASAP7_75t_L g4487 ( 
.A(n_3830),
.Y(n_4487)
);

AND2x2_ASAP7_75t_L g4488 ( 
.A(n_3900),
.B(n_3245),
.Y(n_4488)
);

AND2x2_ASAP7_75t_L g4489 ( 
.A(n_3900),
.B(n_3267),
.Y(n_4489)
);

AOI221xp5_ASAP7_75t_L g4490 ( 
.A1(n_4055),
.A2(n_3541),
.B1(n_3536),
.B2(n_3574),
.C(n_3528),
.Y(n_4490)
);

O2A1O1Ixp5_ASAP7_75t_L g4491 ( 
.A1(n_3723),
.A2(n_3676),
.B(n_3602),
.C(n_3589),
.Y(n_4491)
);

OR2x2_ASAP7_75t_L g4492 ( 
.A(n_3693),
.B(n_3634),
.Y(n_4492)
);

OAI22xp5_ASAP7_75t_L g4493 ( 
.A1(n_3680),
.A2(n_3204),
.B1(n_3411),
.B2(n_3427),
.Y(n_4493)
);

AND2x2_ASAP7_75t_L g4494 ( 
.A(n_3921),
.B(n_3662),
.Y(n_4494)
);

INVx1_ASAP7_75t_L g4495 ( 
.A(n_3692),
.Y(n_4495)
);

OA21x2_ASAP7_75t_L g4496 ( 
.A1(n_3984),
.A2(n_3446),
.B(n_3665),
.Y(n_4496)
);

AND2x2_ASAP7_75t_L g4497 ( 
.A(n_3921),
.B(n_3662),
.Y(n_4497)
);

O2A1O1Ixp5_ASAP7_75t_L g4498 ( 
.A1(n_3682),
.A2(n_3676),
.B(n_3535),
.C(n_3516),
.Y(n_4498)
);

INVx3_ASAP7_75t_L g4499 ( 
.A(n_3777),
.Y(n_4499)
);

OA21x2_ASAP7_75t_L g4500 ( 
.A1(n_3992),
.A2(n_3446),
.B(n_3665),
.Y(n_4500)
);

O2A1O1Ixp33_ASAP7_75t_L g4501 ( 
.A1(n_3803),
.A2(n_3636),
.B(n_3634),
.C(n_3351),
.Y(n_4501)
);

OR2x2_ASAP7_75t_L g4502 ( 
.A(n_3725),
.B(n_3738),
.Y(n_4502)
);

OAI22xp5_ASAP7_75t_L g4503 ( 
.A1(n_3817),
.A2(n_3417),
.B1(n_3427),
.B2(n_3411),
.Y(n_4503)
);

INVx1_ASAP7_75t_L g4504 ( 
.A(n_3692),
.Y(n_4504)
);

AOI21x1_ASAP7_75t_L g4505 ( 
.A1(n_3796),
.A2(n_3492),
.B(n_3663),
.Y(n_4505)
);

NAND2xp5_ASAP7_75t_L g4506 ( 
.A(n_3684),
.B(n_3309),
.Y(n_4506)
);

BUFx3_ASAP7_75t_L g4507 ( 
.A(n_3909),
.Y(n_4507)
);

OAI22xp5_ASAP7_75t_L g4508 ( 
.A1(n_3817),
.A2(n_3417),
.B1(n_3427),
.B2(n_3411),
.Y(n_4508)
);

AND2x2_ASAP7_75t_L g4509 ( 
.A(n_3945),
.B(n_3662),
.Y(n_4509)
);

A2O1A1Ixp33_ASAP7_75t_L g4510 ( 
.A1(n_4055),
.A2(n_3286),
.B(n_3299),
.C(n_3367),
.Y(n_4510)
);

AND2x2_ASAP7_75t_L g4511 ( 
.A(n_3945),
.B(n_3675),
.Y(n_4511)
);

AND2x2_ASAP7_75t_L g4512 ( 
.A(n_3999),
.B(n_3675),
.Y(n_4512)
);

INVx1_ASAP7_75t_L g4513 ( 
.A(n_3695),
.Y(n_4513)
);

AOI21xp5_ASAP7_75t_L g4514 ( 
.A1(n_4133),
.A2(n_3492),
.B(n_3636),
.Y(n_4514)
);

NOR2xp33_ASAP7_75t_R g4515 ( 
.A(n_3795),
.B(n_3548),
.Y(n_4515)
);

OAI22xp5_ASAP7_75t_L g4516 ( 
.A1(n_3869),
.A2(n_3710),
.B1(n_4034),
.B2(n_3995),
.Y(n_4516)
);

BUFx2_ASAP7_75t_L g4517 ( 
.A(n_3833),
.Y(n_4517)
);

AND2x4_ASAP7_75t_L g4518 ( 
.A(n_3799),
.B(n_3299),
.Y(n_4518)
);

INVx2_ASAP7_75t_L g4519 ( 
.A(n_3830),
.Y(n_4519)
);

OAI22xp5_ASAP7_75t_L g4520 ( 
.A1(n_3989),
.A2(n_3417),
.B1(n_3411),
.B2(n_3427),
.Y(n_4520)
);

CKINVDCx14_ASAP7_75t_R g4521 ( 
.A(n_3853),
.Y(n_4521)
);

NAND2xp5_ASAP7_75t_L g4522 ( 
.A(n_3729),
.B(n_3725),
.Y(n_4522)
);

AOI221xp5_ASAP7_75t_L g4523 ( 
.A1(n_4058),
.A2(n_3438),
.B1(n_3433),
.B2(n_3663),
.C(n_3630),
.Y(n_4523)
);

OAI22xp5_ASAP7_75t_L g4524 ( 
.A1(n_3989),
.A2(n_3417),
.B1(n_3411),
.B2(n_3427),
.Y(n_4524)
);

INVx2_ASAP7_75t_L g4525 ( 
.A(n_3854),
.Y(n_4525)
);

OR2x2_ASAP7_75t_L g4526 ( 
.A(n_3738),
.B(n_3351),
.Y(n_4526)
);

INVx3_ASAP7_75t_L g4527 ( 
.A(n_3777),
.Y(n_4527)
);

AND2x4_ASAP7_75t_L g4528 ( 
.A(n_3799),
.B(n_3299),
.Y(n_4528)
);

NOR2xp67_ASAP7_75t_R g4529 ( 
.A(n_3914),
.B(n_3417),
.Y(n_4529)
);

AND2x4_ASAP7_75t_L g4530 ( 
.A(n_3799),
.B(n_3299),
.Y(n_4530)
);

INVx1_ASAP7_75t_L g4531 ( 
.A(n_3695),
.Y(n_4531)
);

AND2x4_ASAP7_75t_L g4532 ( 
.A(n_3799),
.B(n_3325),
.Y(n_4532)
);

OA21x2_ASAP7_75t_L g4533 ( 
.A1(n_4004),
.A2(n_3443),
.B(n_3663),
.Y(n_4533)
);

OR2x2_ASAP7_75t_L g4534 ( 
.A(n_3771),
.B(n_3351),
.Y(n_4534)
);

INVx1_ASAP7_75t_L g4535 ( 
.A(n_3701),
.Y(n_4535)
);

AOI21xp5_ASAP7_75t_L g4536 ( 
.A1(n_3883),
.A2(n_3427),
.B(n_3417),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_3701),
.Y(n_4537)
);

INVx2_ASAP7_75t_L g4538 ( 
.A(n_3854),
.Y(n_4538)
);

O2A1O1Ixp33_ASAP7_75t_L g4539 ( 
.A1(n_3748),
.A2(n_4048),
.B(n_3868),
.C(n_3682),
.Y(n_4539)
);

AND2x4_ASAP7_75t_L g4540 ( 
.A(n_3799),
.B(n_3325),
.Y(n_4540)
);

AND2x2_ASAP7_75t_L g4541 ( 
.A(n_3999),
.B(n_4021),
.Y(n_4541)
);

O2A1O1Ixp33_ASAP7_75t_L g4542 ( 
.A1(n_3702),
.A2(n_3351),
.B(n_3360),
.C(n_3400),
.Y(n_4542)
);

CKINVDCx5p33_ASAP7_75t_R g4543 ( 
.A(n_3689),
.Y(n_4543)
);

OA21x2_ASAP7_75t_L g4544 ( 
.A1(n_3815),
.A2(n_3443),
.B(n_3630),
.Y(n_4544)
);

AND2x2_ASAP7_75t_L g4545 ( 
.A(n_4021),
.B(n_3675),
.Y(n_4545)
);

O2A1O1Ixp33_ASAP7_75t_L g4546 ( 
.A1(n_3748),
.A2(n_3360),
.B(n_3400),
.C(n_3535),
.Y(n_4546)
);

AOI21xp5_ASAP7_75t_SL g4547 ( 
.A1(n_3960),
.A2(n_3432),
.B(n_3186),
.Y(n_4547)
);

INVx2_ASAP7_75t_L g4548 ( 
.A(n_3854),
.Y(n_4548)
);

HB1xp67_ASAP7_75t_L g4549 ( 
.A(n_4135),
.Y(n_4549)
);

BUFx6f_ASAP7_75t_L g4550 ( 
.A(n_3708),
.Y(n_4550)
);

OA21x2_ASAP7_75t_L g4551 ( 
.A1(n_3819),
.A2(n_3443),
.B(n_3630),
.Y(n_4551)
);

AND2x4_ASAP7_75t_L g4552 ( 
.A(n_3799),
.B(n_3353),
.Y(n_4552)
);

AND2x2_ASAP7_75t_L g4553 ( 
.A(n_3834),
.B(n_3857),
.Y(n_4553)
);

INVx1_ASAP7_75t_L g4554 ( 
.A(n_3704),
.Y(n_4554)
);

AND2x2_ASAP7_75t_L g4555 ( 
.A(n_3834),
.B(n_3597),
.Y(n_4555)
);

BUFx3_ASAP7_75t_L g4556 ( 
.A(n_3751),
.Y(n_4556)
);

O2A1O1Ixp33_ASAP7_75t_L g4557 ( 
.A1(n_3702),
.A2(n_3459),
.B(n_3360),
.C(n_3535),
.Y(n_4557)
);

BUFx6f_ASAP7_75t_L g4558 ( 
.A(n_3708),
.Y(n_4558)
);

NAND2xp5_ASAP7_75t_L g4559 ( 
.A(n_3729),
.B(n_3438),
.Y(n_4559)
);

AND2x2_ASAP7_75t_L g4560 ( 
.A(n_3857),
.B(n_3597),
.Y(n_4560)
);

OAI22xp5_ASAP7_75t_L g4561 ( 
.A1(n_3914),
.A2(n_4017),
.B1(n_4030),
.B2(n_3864),
.Y(n_4561)
);

O2A1O1Ixp33_ASAP7_75t_L g4562 ( 
.A1(n_4080),
.A2(n_3459),
.B(n_3360),
.C(n_3535),
.Y(n_4562)
);

OA21x2_ASAP7_75t_L g4563 ( 
.A1(n_4138),
.A2(n_3438),
.B(n_3618),
.Y(n_4563)
);

NAND2xp5_ASAP7_75t_L g4564 ( 
.A(n_3729),
.B(n_3446),
.Y(n_4564)
);

A2O1A1Ixp33_ASAP7_75t_SL g4565 ( 
.A1(n_3783),
.A2(n_3400),
.B(n_3416),
.C(n_3459),
.Y(n_4565)
);

OR2x2_ASAP7_75t_L g4566 ( 
.A(n_3771),
.B(n_3516),
.Y(n_4566)
);

O2A1O1Ixp33_ASAP7_75t_L g4567 ( 
.A1(n_4080),
.A2(n_3516),
.B(n_3400),
.C(n_3416),
.Y(n_4567)
);

AOI211xp5_ASAP7_75t_L g4568 ( 
.A1(n_3883),
.A2(n_3888),
.B(n_3893),
.C(n_4075),
.Y(n_4568)
);

AND2x2_ASAP7_75t_L g4569 ( 
.A(n_3892),
.B(n_3597),
.Y(n_4569)
);

AND2x2_ASAP7_75t_L g4570 ( 
.A(n_3892),
.B(n_3597),
.Y(n_4570)
);

AND2x6_ASAP7_75t_L g4571 ( 
.A(n_3778),
.B(n_3182),
.Y(n_4571)
);

O2A1O1Ixp33_ASAP7_75t_L g4572 ( 
.A1(n_4079),
.A2(n_3416),
.B(n_3516),
.C(n_3363),
.Y(n_4572)
);

AOI21xp5_ASAP7_75t_SL g4573 ( 
.A1(n_3960),
.A2(n_3188),
.B(n_3194),
.Y(n_4573)
);

OA21x2_ASAP7_75t_L g4574 ( 
.A1(n_4148),
.A2(n_3433),
.B(n_3618),
.Y(n_4574)
);

CKINVDCx20_ASAP7_75t_R g4575 ( 
.A(n_3885),
.Y(n_4575)
);

AND2x2_ASAP7_75t_L g4576 ( 
.A(n_3922),
.B(n_3901),
.Y(n_4576)
);

AND2x2_ASAP7_75t_L g4577 ( 
.A(n_3922),
.B(n_3666),
.Y(n_4577)
);

NAND2xp5_ASAP7_75t_L g4578 ( 
.A(n_3704),
.B(n_3709),
.Y(n_4578)
);

BUFx2_ASAP7_75t_L g4579 ( 
.A(n_3901),
.Y(n_4579)
);

OA22x2_ASAP7_75t_L g4580 ( 
.A1(n_3774),
.A2(n_3325),
.B1(n_3353),
.B2(n_3367),
.Y(n_4580)
);

NAND2xp5_ASAP7_75t_L g4581 ( 
.A(n_3709),
.B(n_3715),
.Y(n_4581)
);

NAND2xp5_ASAP7_75t_L g4582 ( 
.A(n_3715),
.B(n_3414),
.Y(n_4582)
);

INVx1_ASAP7_75t_L g4583 ( 
.A(n_3716),
.Y(n_4583)
);

AOI21xp5_ASAP7_75t_L g4584 ( 
.A1(n_4058),
.A2(n_3456),
.B(n_3427),
.Y(n_4584)
);

AOI21xp5_ASAP7_75t_L g4585 ( 
.A1(n_3841),
.A2(n_3456),
.B(n_3417),
.Y(n_4585)
);

NAND2xp5_ASAP7_75t_L g4586 ( 
.A(n_3716),
.B(n_3460),
.Y(n_4586)
);

AOI211xp5_ASAP7_75t_L g4587 ( 
.A1(n_3888),
.A2(n_3893),
.B(n_4079),
.C(n_4005),
.Y(n_4587)
);

OAI22xp5_ASAP7_75t_L g4588 ( 
.A1(n_3914),
.A2(n_3456),
.B1(n_3548),
.B2(n_3205),
.Y(n_4588)
);

OAI22xp5_ASAP7_75t_L g4589 ( 
.A1(n_4017),
.A2(n_3456),
.B1(n_3363),
.B2(n_3471),
.Y(n_4589)
);

NAND2xp5_ASAP7_75t_L g4590 ( 
.A(n_3718),
.B(n_3392),
.Y(n_4590)
);

AOI21x1_ASAP7_75t_SL g4591 ( 
.A1(n_4090),
.A2(n_3188),
.B(n_3194),
.Y(n_4591)
);

AND2x2_ASAP7_75t_L g4592 ( 
.A(n_3901),
.B(n_3666),
.Y(n_4592)
);

INVx1_ASAP7_75t_SL g4593 ( 
.A(n_3957),
.Y(n_4593)
);

AND2x2_ASAP7_75t_L g4594 ( 
.A(n_3930),
.B(n_3666),
.Y(n_4594)
);

OAI22xp5_ASAP7_75t_L g4595 ( 
.A1(n_4030),
.A2(n_3456),
.B1(n_3363),
.B2(n_3471),
.Y(n_4595)
);

BUFx6f_ASAP7_75t_L g4596 ( 
.A(n_3708),
.Y(n_4596)
);

AOI21x1_ASAP7_75t_SL g4597 ( 
.A1(n_4094),
.A2(n_3188),
.B(n_3194),
.Y(n_4597)
);

O2A1O1Ixp33_ASAP7_75t_L g4598 ( 
.A1(n_4173),
.A2(n_3471),
.B(n_3205),
.C(n_3545),
.Y(n_4598)
);

BUFx3_ASAP7_75t_L g4599 ( 
.A(n_3751),
.Y(n_4599)
);

AND2x2_ASAP7_75t_L g4600 ( 
.A(n_3930),
.B(n_3666),
.Y(n_4600)
);

CKINVDCx5p33_ASAP7_75t_R g4601 ( 
.A(n_3751),
.Y(n_4601)
);

AND2x2_ASAP7_75t_L g4602 ( 
.A(n_3930),
.B(n_3540),
.Y(n_4602)
);

INVx2_ASAP7_75t_L g4603 ( 
.A(n_3875),
.Y(n_4603)
);

AOI21xp5_ASAP7_75t_L g4604 ( 
.A1(n_3841),
.A2(n_3456),
.B(n_3545),
.Y(n_4604)
);

AOI21xp5_ASAP7_75t_L g4605 ( 
.A1(n_3846),
.A2(n_3849),
.B(n_3867),
.Y(n_4605)
);

BUFx2_ASAP7_75t_L g4606 ( 
.A(n_3959),
.Y(n_4606)
);

INVx1_ASAP7_75t_L g4607 ( 
.A(n_3721),
.Y(n_4607)
);

INVx1_ASAP7_75t_L g4608 ( 
.A(n_3722),
.Y(n_4608)
);

AND2x2_ASAP7_75t_L g4609 ( 
.A(n_3959),
.B(n_3540),
.Y(n_4609)
);

INVxp67_ASAP7_75t_L g4610 ( 
.A(n_3744),
.Y(n_4610)
);

OR2x2_ASAP7_75t_L g4611 ( 
.A(n_4146),
.B(n_4150),
.Y(n_4611)
);

INVx1_ASAP7_75t_L g4612 ( 
.A(n_3722),
.Y(n_4612)
);

OAI22xp5_ASAP7_75t_L g4613 ( 
.A1(n_4014),
.A2(n_3545),
.B1(n_3367),
.B2(n_3394),
.Y(n_4613)
);

OAI22xp5_ASAP7_75t_L g4614 ( 
.A1(n_4014),
.A2(n_3756),
.B1(n_3800),
.B2(n_4035),
.Y(n_4614)
);

OAI22xp5_ASAP7_75t_L g4615 ( 
.A1(n_4113),
.A2(n_3545),
.B1(n_3367),
.B2(n_3394),
.Y(n_4615)
);

O2A1O1Ixp33_ASAP7_75t_L g4616 ( 
.A1(n_3685),
.A2(n_3545),
.B(n_3624),
.C(n_3622),
.Y(n_4616)
);

OAI22xp5_ASAP7_75t_L g4617 ( 
.A1(n_3681),
.A2(n_3353),
.B1(n_3637),
.B2(n_3606),
.Y(n_4617)
);

AND2x2_ASAP7_75t_L g4618 ( 
.A(n_3959),
.B(n_3478),
.Y(n_4618)
);

CKINVDCx20_ASAP7_75t_R g4619 ( 
.A(n_3979),
.Y(n_4619)
);

AND2x4_ASAP7_75t_L g4620 ( 
.A(n_3952),
.B(n_3353),
.Y(n_4620)
);

AND2x2_ASAP7_75t_L g4621 ( 
.A(n_4001),
.B(n_3478),
.Y(n_4621)
);

O2A1O1Ixp5_ASAP7_75t_L g4622 ( 
.A1(n_3783),
.A2(n_3188),
.B(n_3194),
.C(n_3201),
.Y(n_4622)
);

INVx2_ASAP7_75t_SL g4623 ( 
.A(n_4001),
.Y(n_4623)
);

NOR2xp33_ASAP7_75t_L g4624 ( 
.A(n_3757),
.B(n_3488),
.Y(n_4624)
);

BUFx2_ASAP7_75t_L g4625 ( 
.A(n_4001),
.Y(n_4625)
);

OA21x2_ASAP7_75t_L g4626 ( 
.A1(n_3964),
.A2(n_3349),
.B(n_3618),
.Y(n_4626)
);

INVx2_ASAP7_75t_L g4627 ( 
.A(n_3875),
.Y(n_4627)
);

AOI21xp5_ASAP7_75t_L g4628 ( 
.A1(n_3846),
.A2(n_3622),
.B(n_3624),
.Y(n_4628)
);

AND2x2_ASAP7_75t_L g4629 ( 
.A(n_4012),
.B(n_3488),
.Y(n_4629)
);

NAND2x1p5_ASAP7_75t_L g4630 ( 
.A(n_4059),
.B(n_3201),
.Y(n_4630)
);

AND2x2_ASAP7_75t_L g4631 ( 
.A(n_4012),
.B(n_3488),
.Y(n_4631)
);

O2A1O1Ixp33_ASAP7_75t_L g4632 ( 
.A1(n_4095),
.A2(n_3674),
.B(n_3349),
.C(n_3581),
.Y(n_4632)
);

OAI22xp5_ASAP7_75t_L g4633 ( 
.A1(n_3700),
.A2(n_3488),
.B1(n_3258),
.B2(n_3263),
.Y(n_4633)
);

INVx1_ASAP7_75t_L g4634 ( 
.A(n_3737),
.Y(n_4634)
);

AND2x2_ASAP7_75t_L g4635 ( 
.A(n_4012),
.B(n_3488),
.Y(n_4635)
);

O2A1O1Ixp5_ASAP7_75t_L g4636 ( 
.A1(n_3783),
.A2(n_3201),
.B(n_3599),
.C(n_3591),
.Y(n_4636)
);

AND2x2_ASAP7_75t_L g4637 ( 
.A(n_4022),
.B(n_3488),
.Y(n_4637)
);

O2A1O1Ixp33_ASAP7_75t_L g4638 ( 
.A1(n_3774),
.A2(n_3622),
.B(n_3624),
.C(n_3349),
.Y(n_4638)
);

CKINVDCx12_ASAP7_75t_R g4639 ( 
.A(n_3793),
.Y(n_4639)
);

O2A1O1Ixp5_ASAP7_75t_L g4640 ( 
.A1(n_3783),
.A2(n_3201),
.B(n_3599),
.C(n_3591),
.Y(n_4640)
);

INVx1_ASAP7_75t_L g4641 ( 
.A(n_3739),
.Y(n_4641)
);

AOI21xp5_ASAP7_75t_L g4642 ( 
.A1(n_3849),
.A2(n_3624),
.B(n_3622),
.Y(n_4642)
);

NAND2xp5_ASAP7_75t_L g4643 ( 
.A(n_3739),
.B(n_3740),
.Y(n_4643)
);

AND2x2_ASAP7_75t_L g4644 ( 
.A(n_4022),
.B(n_4050),
.Y(n_4644)
);

AND2x2_ASAP7_75t_L g4645 ( 
.A(n_4050),
.B(n_3258),
.Y(n_4645)
);

BUFx6f_ASAP7_75t_L g4646 ( 
.A(n_3708),
.Y(n_4646)
);

NOR2xp67_ASAP7_75t_L g4647 ( 
.A(n_3952),
.B(n_3591),
.Y(n_4647)
);

NOR2xp67_ASAP7_75t_L g4648 ( 
.A(n_3952),
.B(n_3581),
.Y(n_4648)
);

AND2x2_ASAP7_75t_L g4649 ( 
.A(n_4061),
.B(n_3258),
.Y(n_4649)
);

AND2x2_ASAP7_75t_L g4650 ( 
.A(n_4061),
.B(n_3258),
.Y(n_4650)
);

AND2x2_ASAP7_75t_L g4651 ( 
.A(n_4085),
.B(n_3258),
.Y(n_4651)
);

BUFx5_ASAP7_75t_L g4652 ( 
.A(n_3955),
.Y(n_4652)
);

AND2x2_ASAP7_75t_L g4653 ( 
.A(n_4085),
.B(n_3263),
.Y(n_4653)
);

O2A1O1Ixp5_ASAP7_75t_L g4654 ( 
.A1(n_3850),
.A2(n_3343),
.B(n_3574),
.C(n_3541),
.Y(n_4654)
);

NAND2xp5_ASAP7_75t_L g4655 ( 
.A(n_3742),
.B(n_3758),
.Y(n_4655)
);

CKINVDCx20_ASAP7_75t_R g4656 ( 
.A(n_3986),
.Y(n_4656)
);

O2A1O1Ixp33_ASAP7_75t_L g4657 ( 
.A1(n_3807),
.A2(n_3624),
.B(n_3541),
.C(n_3574),
.Y(n_4657)
);

INVx1_ASAP7_75t_L g4658 ( 
.A(n_3742),
.Y(n_4658)
);

INVx1_ASAP7_75t_L g4659 ( 
.A(n_3758),
.Y(n_4659)
);

AOI21x1_ASAP7_75t_SL g4660 ( 
.A1(n_4136),
.A2(n_3674),
.B(n_3272),
.Y(n_4660)
);

BUFx6f_ASAP7_75t_L g4661 ( 
.A(n_3780),
.Y(n_4661)
);

AND2x2_ASAP7_75t_SL g4662 ( 
.A(n_4059),
.B(n_3263),
.Y(n_4662)
);

INVx1_ASAP7_75t_L g4663 ( 
.A(n_3759),
.Y(n_4663)
);

OAI22xp5_ASAP7_75t_L g4664 ( 
.A1(n_3749),
.A2(n_4121),
.B1(n_4169),
.B2(n_4156),
.Y(n_4664)
);

AND2x2_ASAP7_75t_L g4665 ( 
.A(n_4170),
.B(n_3263),
.Y(n_4665)
);

INVx2_ASAP7_75t_L g4666 ( 
.A(n_3875),
.Y(n_4666)
);

AOI21xp5_ASAP7_75t_L g4667 ( 
.A1(n_3867),
.A2(n_3263),
.B(n_3272),
.Y(n_4667)
);

OA21x2_ASAP7_75t_L g4668 ( 
.A1(n_3968),
.A2(n_3336),
.B(n_3536),
.Y(n_4668)
);

AND2x2_ASAP7_75t_L g4669 ( 
.A(n_4170),
.B(n_3263),
.Y(n_4669)
);

INVxp33_ASAP7_75t_SL g4670 ( 
.A(n_3808),
.Y(n_4670)
);

AND2x4_ASAP7_75t_SL g4671 ( 
.A(n_3998),
.B(n_3272),
.Y(n_4671)
);

O2A1O1Ixp33_ASAP7_75t_L g4672 ( 
.A1(n_4123),
.A2(n_3744),
.B(n_3832),
.C(n_3828),
.Y(n_4672)
);

AND2x2_ASAP7_75t_L g4673 ( 
.A(n_4112),
.B(n_3272),
.Y(n_4673)
);

AND2x4_ASAP7_75t_L g4674 ( 
.A(n_3952),
.B(n_3272),
.Y(n_4674)
);

AND2x2_ASAP7_75t_L g4675 ( 
.A(n_4112),
.B(n_3272),
.Y(n_4675)
);

AOI21x1_ASAP7_75t_SL g4676 ( 
.A1(n_4166),
.A2(n_3674),
.B(n_3289),
.Y(n_4676)
);

AOI21xp5_ASAP7_75t_L g4677 ( 
.A1(n_3936),
.A2(n_3289),
.B(n_3637),
.Y(n_4677)
);

AOI21xp5_ASAP7_75t_SL g4678 ( 
.A1(n_3917),
.A2(n_3289),
.B(n_3637),
.Y(n_4678)
);

O2A1O1Ixp33_ASAP7_75t_L g4679 ( 
.A1(n_3744),
.A2(n_3674),
.B(n_3309),
.C(n_3336),
.Y(n_4679)
);

AND2x2_ASAP7_75t_SL g4680 ( 
.A(n_4059),
.B(n_3289),
.Y(n_4680)
);

AND2x2_ASAP7_75t_L g4681 ( 
.A(n_4154),
.B(n_3289),
.Y(n_4681)
);

AND2x2_ASAP7_75t_L g4682 ( 
.A(n_4157),
.B(n_3289),
.Y(n_4682)
);

INVx1_ASAP7_75t_L g4683 ( 
.A(n_3761),
.Y(n_4683)
);

INVx1_ASAP7_75t_L g4684 ( 
.A(n_3762),
.Y(n_4684)
);

AOI21xp5_ASAP7_75t_L g4685 ( 
.A1(n_3936),
.A2(n_3478),
.B(n_3637),
.Y(n_4685)
);

O2A1O1Ixp5_ASAP7_75t_L g4686 ( 
.A1(n_3850),
.A2(n_3309),
.B(n_3336),
.C(n_3343),
.Y(n_4686)
);

CKINVDCx20_ASAP7_75t_R g4687 ( 
.A(n_3773),
.Y(n_4687)
);

OR2x2_ASAP7_75t_L g4688 ( 
.A(n_4157),
.B(n_3762),
.Y(n_4688)
);

CKINVDCx5p33_ASAP7_75t_R g4689 ( 
.A(n_3757),
.Y(n_4689)
);

BUFx3_ASAP7_75t_L g4690 ( 
.A(n_3757),
.Y(n_4690)
);

NOR2x1_ASAP7_75t_SL g4691 ( 
.A(n_4178),
.B(n_3862),
.Y(n_4691)
);

CKINVDCx20_ASAP7_75t_R g4692 ( 
.A(n_3790),
.Y(n_4692)
);

O2A1O1Ixp5_ASAP7_75t_L g4693 ( 
.A1(n_3850),
.A2(n_3356),
.B(n_3359),
.C(n_3414),
.Y(n_4693)
);

AND2x4_ASAP7_75t_L g4694 ( 
.A(n_3952),
.B(n_3768),
.Y(n_4694)
);

AOI21xp5_ASAP7_75t_L g4695 ( 
.A1(n_3929),
.A2(n_3352),
.B(n_3637),
.Y(n_4695)
);

NAND2xp5_ASAP7_75t_L g4696 ( 
.A(n_3764),
.B(n_3528),
.Y(n_4696)
);

AND2x2_ASAP7_75t_L g4697 ( 
.A(n_4044),
.B(n_3352),
.Y(n_4697)
);

INVx1_ASAP7_75t_L g4698 ( 
.A(n_3766),
.Y(n_4698)
);

OR2x6_ASAP7_75t_L g4699 ( 
.A(n_4151),
.B(n_3352),
.Y(n_4699)
);

INVx1_ASAP7_75t_L g4700 ( 
.A(n_3766),
.Y(n_4700)
);

NAND2xp5_ASAP7_75t_L g4701 ( 
.A(n_3775),
.B(n_3359),
.Y(n_4701)
);

AND2x2_ASAP7_75t_L g4702 ( 
.A(n_4044),
.B(n_3352),
.Y(n_4702)
);

AND2x2_ASAP7_75t_L g4703 ( 
.A(n_4044),
.B(n_3352),
.Y(n_4703)
);

NOR3xp33_ASAP7_75t_SL g4704 ( 
.A(n_4561),
.B(n_3837),
.C(n_3789),
.Y(n_4704)
);

AND2x2_ASAP7_75t_L g4705 ( 
.A(n_4324),
.B(n_3996),
.Y(n_4705)
);

OAI22xp5_ASAP7_75t_L g4706 ( 
.A1(n_4200),
.A2(n_4088),
.B1(n_4098),
.B2(n_4117),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4688),
.Y(n_4707)
);

NAND3xp33_ASAP7_75t_SL g4708 ( 
.A(n_4307),
.B(n_3929),
.C(n_4005),
.Y(n_4708)
);

INVx1_ASAP7_75t_L g4709 ( 
.A(n_4688),
.Y(n_4709)
);

INVx2_ASAP7_75t_L g4710 ( 
.A(n_4505),
.Y(n_4710)
);

OR2x2_ASAP7_75t_L g4711 ( 
.A(n_4191),
.B(n_3779),
.Y(n_4711)
);

AOI222xp33_ASAP7_75t_L g4712 ( 
.A1(n_4286),
.A2(n_3734),
.B1(n_4053),
.B2(n_3847),
.C1(n_3840),
.C2(n_3952),
.Y(n_4712)
);

INVx1_ASAP7_75t_L g4713 ( 
.A(n_4611),
.Y(n_4713)
);

INVx1_ASAP7_75t_L g4714 ( 
.A(n_4611),
.Y(n_4714)
);

CKINVDCx16_ASAP7_75t_R g4715 ( 
.A(n_4305),
.Y(n_4715)
);

AO31x2_ASAP7_75t_L g4716 ( 
.A1(n_4236),
.A2(n_3897),
.A3(n_3898),
.B(n_3879),
.Y(n_4716)
);

XOR2x2_ASAP7_75t_SL g4717 ( 
.A(n_4200),
.B(n_3781),
.Y(n_4717)
);

CKINVDCx5p33_ASAP7_75t_R g4718 ( 
.A(n_4249),
.Y(n_4718)
);

CKINVDCx5p33_ASAP7_75t_R g4719 ( 
.A(n_4338),
.Y(n_4719)
);

NOR2xp33_ASAP7_75t_L g4720 ( 
.A(n_4237),
.B(n_3790),
.Y(n_4720)
);

AND2x2_ASAP7_75t_L g4721 ( 
.A(n_4324),
.B(n_3996),
.Y(n_4721)
);

AOI22xp33_ASAP7_75t_L g4722 ( 
.A1(n_4476),
.A2(n_3952),
.B1(n_4064),
.B2(n_4102),
.Y(n_4722)
);

NAND3xp33_ASAP7_75t_SL g4723 ( 
.A(n_4307),
.B(n_3940),
.C(n_3781),
.Y(n_4723)
);

INVx1_ASAP7_75t_L g4724 ( 
.A(n_4204),
.Y(n_4724)
);

BUFx3_ASAP7_75t_L g4725 ( 
.A(n_4305),
.Y(n_4725)
);

HB1xp67_ASAP7_75t_L g4726 ( 
.A(n_4225),
.Y(n_4726)
);

NOR2x1_ASAP7_75t_L g4727 ( 
.A(n_4253),
.B(n_3765),
.Y(n_4727)
);

NAND2x1p5_ASAP7_75t_L g4728 ( 
.A(n_4662),
.B(n_4059),
.Y(n_4728)
);

NAND2xp33_ASAP7_75t_SL g4729 ( 
.A(n_4515),
.B(n_3826),
.Y(n_4729)
);

CKINVDCx5p33_ASAP7_75t_R g4730 ( 
.A(n_4218),
.Y(n_4730)
);

NOR3xp33_ASAP7_75t_SL g4731 ( 
.A(n_4561),
.B(n_3837),
.C(n_3789),
.Y(n_4731)
);

INVx4_ASAP7_75t_L g4732 ( 
.A(n_4305),
.Y(n_4732)
);

BUFx3_ASAP7_75t_L g4733 ( 
.A(n_4250),
.Y(n_4733)
);

AND2x2_ASAP7_75t_L g4734 ( 
.A(n_4201),
.B(n_3996),
.Y(n_4734)
);

OR2x6_ASAP7_75t_L g4735 ( 
.A(n_4253),
.B(n_4151),
.Y(n_4735)
);

NOR2x1_ASAP7_75t_SL g4736 ( 
.A(n_4699),
.B(n_3907),
.Y(n_4736)
);

INVx2_ASAP7_75t_L g4737 ( 
.A(n_4505),
.Y(n_4737)
);

BUFx3_ASAP7_75t_L g4738 ( 
.A(n_4250),
.Y(n_4738)
);

CKINVDCx5p33_ASAP7_75t_R g4739 ( 
.A(n_4319),
.Y(n_4739)
);

NOR2xp33_ASAP7_75t_L g4740 ( 
.A(n_4220),
.B(n_3790),
.Y(n_4740)
);

CKINVDCx5p33_ASAP7_75t_R g4741 ( 
.A(n_4328),
.Y(n_4741)
);

INVx2_ASAP7_75t_L g4742 ( 
.A(n_4654),
.Y(n_4742)
);

INVx1_ASAP7_75t_L g4743 ( 
.A(n_4204),
.Y(n_4743)
);

AOI22xp33_ASAP7_75t_L g4744 ( 
.A1(n_4476),
.A2(n_4064),
.B1(n_4110),
.B2(n_4151),
.Y(n_4744)
);

HB1xp67_ASAP7_75t_L g4745 ( 
.A(n_4259),
.Y(n_4745)
);

BUFx4f_ASAP7_75t_SL g4746 ( 
.A(n_4575),
.Y(n_4746)
);

INVx1_ASAP7_75t_L g4747 ( 
.A(n_4278),
.Y(n_4747)
);

O2A1O1Ixp33_ASAP7_75t_L g4748 ( 
.A1(n_4238),
.A2(n_3850),
.B(n_3904),
.C(n_3866),
.Y(n_4748)
);

AND2x2_ASAP7_75t_L g4749 ( 
.A(n_4201),
.B(n_3996),
.Y(n_4749)
);

INVx2_ASAP7_75t_L g4750 ( 
.A(n_4686),
.Y(n_4750)
);

INVx1_ASAP7_75t_SL g4751 ( 
.A(n_4276),
.Y(n_4751)
);

NAND2xp33_ASAP7_75t_R g4752 ( 
.A(n_4265),
.B(n_3866),
.Y(n_4752)
);

NOR2xp33_ASAP7_75t_R g4753 ( 
.A(n_4521),
.B(n_3889),
.Y(n_4753)
);

AOI22xp33_ASAP7_75t_L g4754 ( 
.A1(n_4614),
.A2(n_4064),
.B1(n_4151),
.B2(n_3696),
.Y(n_4754)
);

HB1xp67_ASAP7_75t_L g4755 ( 
.A(n_4211),
.Y(n_4755)
);

CKINVDCx8_ASAP7_75t_R g4756 ( 
.A(n_4475),
.Y(n_4756)
);

AND2x4_ASAP7_75t_L g4757 ( 
.A(n_4310),
.B(n_3768),
.Y(n_4757)
);

NOR2xp33_ASAP7_75t_L g4758 ( 
.A(n_4220),
.B(n_3810),
.Y(n_4758)
);

BUFx6f_ASAP7_75t_L g4759 ( 
.A(n_4250),
.Y(n_4759)
);

NOR3xp33_ASAP7_75t_SL g4760 ( 
.A(n_4543),
.B(n_3837),
.C(n_3789),
.Y(n_4760)
);

INVx1_ASAP7_75t_SL g4761 ( 
.A(n_4212),
.Y(n_4761)
);

OAI22xp5_ASAP7_75t_L g4762 ( 
.A1(n_4440),
.A2(n_4002),
.B1(n_4016),
.B2(n_3998),
.Y(n_4762)
);

OAI21xp5_ASAP7_75t_L g4763 ( 
.A1(n_4228),
.A2(n_3940),
.B(n_3844),
.Y(n_4763)
);

CKINVDCx6p67_ASAP7_75t_R g4764 ( 
.A(n_4639),
.Y(n_4764)
);

CKINVDCx5p33_ASAP7_75t_R g4765 ( 
.A(n_4670),
.Y(n_4765)
);

INVx1_ASAP7_75t_L g4766 ( 
.A(n_4278),
.Y(n_4766)
);

NAND2xp33_ASAP7_75t_R g4767 ( 
.A(n_4265),
.B(n_3866),
.Y(n_4767)
);

HB1xp67_ASAP7_75t_L g4768 ( 
.A(n_4308),
.Y(n_4768)
);

AOI221xp5_ASAP7_75t_L g4769 ( 
.A1(n_4614),
.A2(n_4023),
.B1(n_4027),
.B2(n_4018),
.C(n_4015),
.Y(n_4769)
);

OAI22xp5_ASAP7_75t_L g4770 ( 
.A1(n_4440),
.A2(n_3998),
.B1(n_4038),
.B2(n_4016),
.Y(n_4770)
);

HB1xp67_ASAP7_75t_L g4771 ( 
.A(n_4339),
.Y(n_4771)
);

HB1xp67_ASAP7_75t_L g4772 ( 
.A(n_4450),
.Y(n_4772)
);

CKINVDCx16_ASAP7_75t_R g4773 ( 
.A(n_4619),
.Y(n_4773)
);

NOR3xp33_ASAP7_75t_SL g4774 ( 
.A(n_4314),
.B(n_3837),
.C(n_3789),
.Y(n_4774)
);

AOI22xp33_ASAP7_75t_L g4775 ( 
.A1(n_4336),
.A2(n_4064),
.B1(n_4151),
.B2(n_3696),
.Y(n_4775)
);

AOI221xp5_ASAP7_75t_L g4776 ( 
.A1(n_4336),
.A2(n_4027),
.B1(n_4023),
.B2(n_4018),
.C(n_4015),
.Y(n_4776)
);

AND2x2_ASAP7_75t_L g4777 ( 
.A(n_4203),
.B(n_4033),
.Y(n_4777)
);

HB1xp67_ASAP7_75t_L g4778 ( 
.A(n_4450),
.Y(n_4778)
);

INVx2_ASAP7_75t_L g4779 ( 
.A(n_4693),
.Y(n_4779)
);

HB1xp67_ASAP7_75t_L g4780 ( 
.A(n_4502),
.Y(n_4780)
);

INVx2_ASAP7_75t_L g4781 ( 
.A(n_4227),
.Y(n_4781)
);

AND2x2_ASAP7_75t_L g4782 ( 
.A(n_4203),
.B(n_4033),
.Y(n_4782)
);

CKINVDCx16_ASAP7_75t_R g4783 ( 
.A(n_4656),
.Y(n_4783)
);

AO31x2_ASAP7_75t_L g4784 ( 
.A1(n_4236),
.A2(n_3897),
.A3(n_3898),
.B(n_3879),
.Y(n_4784)
);

INVxp67_ASAP7_75t_L g4785 ( 
.A(n_4426),
.Y(n_4785)
);

NAND2xp33_ASAP7_75t_R g4786 ( 
.A(n_4265),
.B(n_3866),
.Y(n_4786)
);

INVx2_ASAP7_75t_L g4787 ( 
.A(n_4227),
.Y(n_4787)
);

CKINVDCx16_ASAP7_75t_R g4788 ( 
.A(n_4395),
.Y(n_4788)
);

INVx1_ASAP7_75t_L g4789 ( 
.A(n_4281),
.Y(n_4789)
);

NOR2x1_ASAP7_75t_L g4790 ( 
.A(n_4343),
.B(n_3765),
.Y(n_4790)
);

BUFx3_ASAP7_75t_L g4791 ( 
.A(n_4252),
.Y(n_4791)
);

OAI22xp5_ASAP7_75t_L g4792 ( 
.A1(n_4228),
.A2(n_4016),
.B1(n_4084),
.B2(n_4038),
.Y(n_4792)
);

AND2x2_ASAP7_75t_L g4793 ( 
.A(n_4189),
.B(n_4033),
.Y(n_4793)
);

NAND2xp33_ASAP7_75t_L g4794 ( 
.A(n_4601),
.B(n_3826),
.Y(n_4794)
);

OAI21x1_ASAP7_75t_L g4795 ( 
.A1(n_4660),
.A2(n_3938),
.B(n_3904),
.Y(n_4795)
);

NOR3xp33_ASAP7_75t_SL g4796 ( 
.A(n_4314),
.B(n_3886),
.C(n_3889),
.Y(n_4796)
);

BUFx3_ASAP7_75t_L g4797 ( 
.A(n_4252),
.Y(n_4797)
);

INVx1_ASAP7_75t_L g4798 ( 
.A(n_4281),
.Y(n_4798)
);

INVx2_ASAP7_75t_L g4799 ( 
.A(n_4227),
.Y(n_4799)
);

AND2x2_ASAP7_75t_L g4800 ( 
.A(n_4189),
.B(n_4033),
.Y(n_4800)
);

AND2x2_ASAP7_75t_L g4801 ( 
.A(n_4190),
.B(n_4103),
.Y(n_4801)
);

NOR2xp33_ASAP7_75t_R g4802 ( 
.A(n_4692),
.B(n_3810),
.Y(n_4802)
);

INVx1_ASAP7_75t_L g4803 ( 
.A(n_4301),
.Y(n_4803)
);

HB1xp67_ASAP7_75t_L g4804 ( 
.A(n_4502),
.Y(n_4804)
);

INVx1_ASAP7_75t_L g4805 ( 
.A(n_4301),
.Y(n_4805)
);

AND2x2_ASAP7_75t_L g4806 ( 
.A(n_4190),
.B(n_4103),
.Y(n_4806)
);

INVx2_ASAP7_75t_L g4807 ( 
.A(n_4230),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4342),
.Y(n_4808)
);

CKINVDCx5p33_ASAP7_75t_R g4809 ( 
.A(n_4687),
.Y(n_4809)
);

AOI22xp33_ASAP7_75t_L g4810 ( 
.A1(n_4467),
.A2(n_4151),
.B1(n_3696),
.B2(n_3717),
.Y(n_4810)
);

NAND2xp5_ASAP7_75t_L g4811 ( 
.A(n_4306),
.B(n_3779),
.Y(n_4811)
);

INVx1_ASAP7_75t_L g4812 ( 
.A(n_4342),
.Y(n_4812)
);

AND2x2_ASAP7_75t_L g4813 ( 
.A(n_4192),
.B(n_4103),
.Y(n_4813)
);

AND2x2_ASAP7_75t_L g4814 ( 
.A(n_4192),
.B(n_4103),
.Y(n_4814)
);

INVx2_ASAP7_75t_L g4815 ( 
.A(n_4230),
.Y(n_4815)
);

AOI22xp33_ASAP7_75t_L g4816 ( 
.A1(n_4467),
.A2(n_3696),
.B1(n_3717),
.B2(n_3707),
.Y(n_4816)
);

NOR2xp33_ASAP7_75t_R g4817 ( 
.A(n_4639),
.B(n_3810),
.Y(n_4817)
);

NAND2xp33_ASAP7_75t_R g4818 ( 
.A(n_4265),
.B(n_3904),
.Y(n_4818)
);

OAI22xp5_ASAP7_75t_L g4819 ( 
.A1(n_4605),
.A2(n_4084),
.B1(n_4092),
.B2(n_4038),
.Y(n_4819)
);

INVx1_ASAP7_75t_L g4820 ( 
.A(n_4358),
.Y(n_4820)
);

AND2x2_ASAP7_75t_SL g4821 ( 
.A(n_4323),
.B(n_4114),
.Y(n_4821)
);

AOI22xp33_ASAP7_75t_L g4822 ( 
.A1(n_4286),
.A2(n_3707),
.B1(n_3825),
.B2(n_3717),
.Y(n_4822)
);

INVx1_ASAP7_75t_L g4823 ( 
.A(n_4358),
.Y(n_4823)
);

NOR2xp33_ASAP7_75t_L g4824 ( 
.A(n_4443),
.B(n_3826),
.Y(n_4824)
);

HB1xp67_ASAP7_75t_L g4825 ( 
.A(n_4371),
.Y(n_4825)
);

A2O1A1Ixp33_ASAP7_75t_L g4826 ( 
.A1(n_4605),
.A2(n_4137),
.B(n_3950),
.C(n_3778),
.Y(n_4826)
);

NAND3xp33_ASAP7_75t_L g4827 ( 
.A(n_4398),
.B(n_3886),
.C(n_3786),
.Y(n_4827)
);

OAI22xp5_ASAP7_75t_L g4828 ( 
.A1(n_4398),
.A2(n_4084),
.B1(n_4092),
.B2(n_4026),
.Y(n_4828)
);

INVx1_ASAP7_75t_L g4829 ( 
.A(n_4364),
.Y(n_4829)
);

OR2x6_ASAP7_75t_L g4830 ( 
.A(n_4366),
.B(n_4019),
.Y(n_4830)
);

AND2x2_ASAP7_75t_L g4831 ( 
.A(n_4194),
.B(n_4114),
.Y(n_4831)
);

INVx5_ASAP7_75t_L g4832 ( 
.A(n_4258),
.Y(n_4832)
);

NAND2xp33_ASAP7_75t_SL g4833 ( 
.A(n_4186),
.B(n_4026),
.Y(n_4833)
);

AO21x2_ASAP7_75t_L g4834 ( 
.A1(n_4380),
.A2(n_3897),
.B(n_3879),
.Y(n_4834)
);

HB1xp67_ASAP7_75t_L g4835 ( 
.A(n_4437),
.Y(n_4835)
);

AOI22xp33_ASAP7_75t_L g4836 ( 
.A1(n_4347),
.A2(n_3707),
.B1(n_3825),
.B2(n_3717),
.Y(n_4836)
);

OR2x6_ASAP7_75t_L g4837 ( 
.A(n_4366),
.B(n_4019),
.Y(n_4837)
);

INVxp67_ASAP7_75t_L g4838 ( 
.A(n_4426),
.Y(n_4838)
);

INVx1_ASAP7_75t_L g4839 ( 
.A(n_4364),
.Y(n_4839)
);

CKINVDCx5p33_ASAP7_75t_R g4840 ( 
.A(n_4689),
.Y(n_4840)
);

NOR2xp33_ASAP7_75t_R g4841 ( 
.A(n_4507),
.B(n_3931),
.Y(n_4841)
);

AO31x2_ASAP7_75t_L g4842 ( 
.A1(n_4380),
.A2(n_3902),
.A3(n_3915),
.B(n_3898),
.Y(n_4842)
);

NOR2xp33_ASAP7_75t_R g4843 ( 
.A(n_4507),
.B(n_3931),
.Y(n_4843)
);

INVx2_ASAP7_75t_L g4844 ( 
.A(n_4230),
.Y(n_4844)
);

INVx2_ASAP7_75t_L g4845 ( 
.A(n_4239),
.Y(n_4845)
);

AND2x2_ASAP7_75t_L g4846 ( 
.A(n_4194),
.B(n_4114),
.Y(n_4846)
);

HB1xp67_ASAP7_75t_L g4847 ( 
.A(n_4460),
.Y(n_4847)
);

AO21x2_ASAP7_75t_L g4848 ( 
.A1(n_4245),
.A2(n_3915),
.B(n_3902),
.Y(n_4848)
);

CKINVDCx5p33_ASAP7_75t_R g4849 ( 
.A(n_4507),
.Y(n_4849)
);

INVxp67_ASAP7_75t_L g4850 ( 
.A(n_4486),
.Y(n_4850)
);

AND2x2_ASAP7_75t_L g4851 ( 
.A(n_4186),
.B(n_4114),
.Y(n_4851)
);

AND2x4_ASAP7_75t_L g4852 ( 
.A(n_4310),
.B(n_3768),
.Y(n_4852)
);

INVx2_ASAP7_75t_L g4853 ( 
.A(n_4239),
.Y(n_4853)
);

AND2x2_ASAP7_75t_L g4854 ( 
.A(n_4313),
.B(n_4222),
.Y(n_4854)
);

AOI22xp33_ASAP7_75t_L g4855 ( 
.A1(n_4347),
.A2(n_3707),
.B1(n_3825),
.B2(n_3717),
.Y(n_4855)
);

INVx2_ASAP7_75t_L g4856 ( 
.A(n_4239),
.Y(n_4856)
);

NAND2xp5_ASAP7_75t_L g4857 ( 
.A(n_4306),
.B(n_3782),
.Y(n_4857)
);

AND2x2_ASAP7_75t_L g4858 ( 
.A(n_4313),
.B(n_4120),
.Y(n_4858)
);

NOR3xp33_ASAP7_75t_SL g4859 ( 
.A(n_4362),
.B(n_4422),
.C(n_4387),
.Y(n_4859)
);

INVx1_ASAP7_75t_L g4860 ( 
.A(n_4369),
.Y(n_4860)
);

INVx1_ASAP7_75t_L g4861 ( 
.A(n_4369),
.Y(n_4861)
);

BUFx6f_ASAP7_75t_L g4862 ( 
.A(n_4258),
.Y(n_4862)
);

AO31x2_ASAP7_75t_L g4863 ( 
.A1(n_4291),
.A2(n_4362),
.A3(n_4245),
.B(n_4514),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4404),
.Y(n_4864)
);

INVx2_ASAP7_75t_L g4865 ( 
.A(n_4251),
.Y(n_4865)
);

INVx1_ASAP7_75t_L g4866 ( 
.A(n_4404),
.Y(n_4866)
);

INVx1_ASAP7_75t_L g4867 ( 
.A(n_4448),
.Y(n_4867)
);

BUFx5_ASAP7_75t_L g4868 ( 
.A(n_4571),
.Y(n_4868)
);

INVx6_ASAP7_75t_L g4869 ( 
.A(n_4258),
.Y(n_4869)
);

CKINVDCx20_ASAP7_75t_R g4870 ( 
.A(n_4486),
.Y(n_4870)
);

BUFx12f_ASAP7_75t_L g4871 ( 
.A(n_4378),
.Y(n_4871)
);

INVx1_ASAP7_75t_L g4872 ( 
.A(n_4448),
.Y(n_4872)
);

BUFx2_ASAP7_75t_L g4873 ( 
.A(n_4302),
.Y(n_4873)
);

NOR3xp33_ASAP7_75t_SL g4874 ( 
.A(n_4422),
.B(n_3886),
.C(n_3931),
.Y(n_4874)
);

AND2x2_ASAP7_75t_L g4875 ( 
.A(n_4222),
.B(n_4120),
.Y(n_4875)
);

CKINVDCx5p33_ASAP7_75t_R g4876 ( 
.A(n_4443),
.Y(n_4876)
);

OAI21xp5_ASAP7_75t_L g4877 ( 
.A1(n_4231),
.A2(n_3917),
.B(n_3786),
.Y(n_4877)
);

AND2x2_ASAP7_75t_L g4878 ( 
.A(n_4223),
.B(n_4120),
.Y(n_4878)
);

NAND2xp33_ASAP7_75t_L g4879 ( 
.A(n_4212),
.B(n_4026),
.Y(n_4879)
);

AO31x2_ASAP7_75t_L g4880 ( 
.A1(n_4291),
.A2(n_3915),
.A3(n_3920),
.B(n_3902),
.Y(n_4880)
);

OR2x6_ASAP7_75t_L g4881 ( 
.A(n_4357),
.B(n_4256),
.Y(n_4881)
);

HB1xp67_ASAP7_75t_L g4882 ( 
.A(n_4549),
.Y(n_4882)
);

OAI21xp5_ASAP7_75t_L g4883 ( 
.A1(n_4231),
.A2(n_3917),
.B(n_3787),
.Y(n_4883)
);

CKINVDCx5p33_ASAP7_75t_R g4884 ( 
.A(n_4593),
.Y(n_4884)
);

INVx2_ASAP7_75t_SL g4885 ( 
.A(n_4360),
.Y(n_4885)
);

NAND2xp5_ASAP7_75t_L g4886 ( 
.A(n_4293),
.B(n_4294),
.Y(n_4886)
);

AND2x2_ASAP7_75t_L g4887 ( 
.A(n_4223),
.B(n_4120),
.Y(n_4887)
);

NAND2xp5_ASAP7_75t_L g4888 ( 
.A(n_4293),
.B(n_3782),
.Y(n_4888)
);

CKINVDCx20_ASAP7_75t_R g4889 ( 
.A(n_4517),
.Y(n_4889)
);

AND2x4_ASAP7_75t_L g4890 ( 
.A(n_4310),
.B(n_3842),
.Y(n_4890)
);

INVx2_ASAP7_75t_L g4891 ( 
.A(n_4251),
.Y(n_4891)
);

NOR2xp33_ASAP7_75t_R g4892 ( 
.A(n_4360),
.B(n_3931),
.Y(n_4892)
);

AO31x2_ASAP7_75t_L g4893 ( 
.A1(n_4514),
.A2(n_3926),
.A3(n_3928),
.B(n_3920),
.Y(n_4893)
);

INVx2_ASAP7_75t_L g4894 ( 
.A(n_4251),
.Y(n_4894)
);

AND2x2_ASAP7_75t_L g4895 ( 
.A(n_4226),
.B(n_3907),
.Y(n_4895)
);

AOI22xp33_ASAP7_75t_L g4896 ( 
.A1(n_4244),
.A2(n_3707),
.B1(n_3852),
.B2(n_3825),
.Y(n_4896)
);

NOR2xp33_ASAP7_75t_L g4897 ( 
.A(n_4479),
.B(n_3765),
.Y(n_4897)
);

NAND2xp33_ASAP7_75t_R g4898 ( 
.A(n_4388),
.B(n_3904),
.Y(n_4898)
);

INVx2_ASAP7_75t_L g4899 ( 
.A(n_4260),
.Y(n_4899)
);

NOR3xp33_ASAP7_75t_SL g4900 ( 
.A(n_4387),
.B(n_3886),
.C(n_3941),
.Y(n_4900)
);

INVx1_ASAP7_75t_SL g4901 ( 
.A(n_4593),
.Y(n_4901)
);

O2A1O1Ixp33_ASAP7_75t_SL g4902 ( 
.A1(n_4235),
.A2(n_4210),
.B(n_4340),
.C(n_4183),
.Y(n_4902)
);

CKINVDCx12_ASAP7_75t_R g4903 ( 
.A(n_4181),
.Y(n_4903)
);

INVx2_ASAP7_75t_L g4904 ( 
.A(n_4260),
.Y(n_4904)
);

AO31x2_ASAP7_75t_L g4905 ( 
.A1(n_4445),
.A2(n_3976),
.A3(n_4046),
.B(n_4042),
.Y(n_4905)
);

INVx3_ASAP7_75t_L g4906 ( 
.A(n_4302),
.Y(n_4906)
);

INVx2_ASAP7_75t_L g4907 ( 
.A(n_4260),
.Y(n_4907)
);

INVx1_ASAP7_75t_L g4908 ( 
.A(n_4449),
.Y(n_4908)
);

AOI22xp5_ASAP7_75t_L g4909 ( 
.A1(n_4244),
.A2(n_3847),
.B1(n_4158),
.B2(n_4176),
.Y(n_4909)
);

AND2x2_ASAP7_75t_L g4910 ( 
.A(n_4226),
.B(n_3961),
.Y(n_4910)
);

HB1xp67_ASAP7_75t_L g4911 ( 
.A(n_4219),
.Y(n_4911)
);

NOR2xp33_ASAP7_75t_R g4912 ( 
.A(n_4388),
.B(n_3941),
.Y(n_4912)
);

CKINVDCx16_ASAP7_75t_R g4913 ( 
.A(n_4309),
.Y(n_4913)
);

HB1xp67_ASAP7_75t_L g4914 ( 
.A(n_4432),
.Y(n_4914)
);

AOI22xp33_ASAP7_75t_L g4915 ( 
.A1(n_4246),
.A2(n_3988),
.B1(n_3894),
.B2(n_3927),
.Y(n_4915)
);

CKINVDCx16_ASAP7_75t_R g4916 ( 
.A(n_4309),
.Y(n_4916)
);

NAND2xp5_ASAP7_75t_L g4917 ( 
.A(n_4298),
.B(n_3787),
.Y(n_4917)
);

AND2x2_ASAP7_75t_L g4918 ( 
.A(n_4242),
.B(n_3961),
.Y(n_4918)
);

HB1xp67_ASAP7_75t_L g4919 ( 
.A(n_4432),
.Y(n_4919)
);

BUFx2_ASAP7_75t_L g4920 ( 
.A(n_4302),
.Y(n_4920)
);

CKINVDCx5p33_ASAP7_75t_R g4921 ( 
.A(n_4556),
.Y(n_4921)
);

OR2x2_ASAP7_75t_SL g4922 ( 
.A(n_4323),
.B(n_4107),
.Y(n_4922)
);

BUFx12f_ASAP7_75t_L g4923 ( 
.A(n_4378),
.Y(n_4923)
);

INVx1_ASAP7_75t_L g4924 ( 
.A(n_4449),
.Y(n_4924)
);

OAI22xp33_ASAP7_75t_L g4925 ( 
.A1(n_4246),
.A2(n_4241),
.B1(n_4191),
.B2(n_4271),
.Y(n_4925)
);

AOI22xp33_ASAP7_75t_L g4926 ( 
.A1(n_4516),
.A2(n_3927),
.B1(n_3988),
.B2(n_4006),
.Y(n_4926)
);

AND2x2_ASAP7_75t_L g4927 ( 
.A(n_4242),
.B(n_3994),
.Y(n_4927)
);

INVx4_ASAP7_75t_L g4928 ( 
.A(n_4378),
.Y(n_4928)
);

INVx1_ASAP7_75t_L g4929 ( 
.A(n_4456),
.Y(n_4929)
);

NAND2xp33_ASAP7_75t_SL g4930 ( 
.A(n_4181),
.B(n_4325),
.Y(n_4930)
);

NOR2xp33_ASAP7_75t_R g4931 ( 
.A(n_4309),
.B(n_3941),
.Y(n_4931)
);

BUFx12f_ASAP7_75t_L g4932 ( 
.A(n_4378),
.Y(n_4932)
);

AOI22xp33_ASAP7_75t_SL g4933 ( 
.A1(n_4241),
.A2(n_4028),
.B1(n_3927),
.B2(n_3974),
.Y(n_4933)
);

BUFx3_ASAP7_75t_L g4934 ( 
.A(n_4396),
.Y(n_4934)
);

INVx2_ASAP7_75t_L g4935 ( 
.A(n_4263),
.Y(n_4935)
);

INVx2_ASAP7_75t_L g4936 ( 
.A(n_4263),
.Y(n_4936)
);

NAND2xp33_ASAP7_75t_R g4937 ( 
.A(n_4517),
.B(n_3938),
.Y(n_4937)
);

OR2x6_ASAP7_75t_L g4938 ( 
.A(n_4357),
.B(n_4256),
.Y(n_4938)
);

NAND2xp33_ASAP7_75t_R g4939 ( 
.A(n_4323),
.B(n_3938),
.Y(n_4939)
);

CKINVDCx16_ASAP7_75t_R g4940 ( 
.A(n_4396),
.Y(n_4940)
);

AOI22xp33_ASAP7_75t_L g4941 ( 
.A1(n_4516),
.A2(n_3927),
.B1(n_3988),
.B2(n_4006),
.Y(n_4941)
);

INVx2_ASAP7_75t_L g4942 ( 
.A(n_4263),
.Y(n_4942)
);

OAI22xp5_ASAP7_75t_L g4943 ( 
.A1(n_4235),
.A2(n_4092),
.B1(n_4108),
.B2(n_4147),
.Y(n_4943)
);

OAI22xp5_ASAP7_75t_L g4944 ( 
.A1(n_4587),
.A2(n_4107),
.B1(n_4108),
.B2(n_4147),
.Y(n_4944)
);

AND2x2_ASAP7_75t_L g4945 ( 
.A(n_4279),
.B(n_3994),
.Y(n_4945)
);

NOR3xp33_ASAP7_75t_SL g4946 ( 
.A(n_4393),
.B(n_3948),
.C(n_3941),
.Y(n_4946)
);

AOI22xp33_ASAP7_75t_L g4947 ( 
.A1(n_4205),
.A2(n_3927),
.B1(n_3988),
.B2(n_4006),
.Y(n_4947)
);

AND2x2_ASAP7_75t_L g4948 ( 
.A(n_4279),
.B(n_4049),
.Y(n_4948)
);

OR2x2_ASAP7_75t_L g4949 ( 
.A(n_4272),
.B(n_3801),
.Y(n_4949)
);

NAND2xp33_ASAP7_75t_SL g4950 ( 
.A(n_4325),
.B(n_3765),
.Y(n_4950)
);

HB1xp67_ASAP7_75t_L g4951 ( 
.A(n_4335),
.Y(n_4951)
);

BUFx3_ASAP7_75t_L g4952 ( 
.A(n_4396),
.Y(n_4952)
);

INVx1_ASAP7_75t_L g4953 ( 
.A(n_4456),
.Y(n_4953)
);

INVx1_ASAP7_75t_L g4954 ( 
.A(n_4458),
.Y(n_4954)
);

AOI22xp33_ASAP7_75t_SL g4955 ( 
.A1(n_4241),
.A2(n_4051),
.B1(n_3974),
.B2(n_3982),
.Y(n_4955)
);

CKINVDCx14_ASAP7_75t_R g4956 ( 
.A(n_4556),
.Y(n_4956)
);

INVx1_ASAP7_75t_L g4957 ( 
.A(n_4458),
.Y(n_4957)
);

CKINVDCx16_ASAP7_75t_R g4958 ( 
.A(n_4433),
.Y(n_4958)
);

NAND2xp5_ASAP7_75t_L g4959 ( 
.A(n_4298),
.B(n_3801),
.Y(n_4959)
);

INVx1_ASAP7_75t_L g4960 ( 
.A(n_4484),
.Y(n_4960)
);

CKINVDCx5p33_ASAP7_75t_R g4961 ( 
.A(n_4556),
.Y(n_4961)
);

AO21x2_ASAP7_75t_L g4962 ( 
.A1(n_4346),
.A2(n_4377),
.B(n_4352),
.Y(n_4962)
);

BUFx2_ASAP7_75t_L g4963 ( 
.A(n_4302),
.Y(n_4963)
);

NAND3xp33_ASAP7_75t_SL g4964 ( 
.A(n_4587),
.B(n_3851),
.C(n_3845),
.Y(n_4964)
);

NOR3xp33_ASAP7_75t_SL g4965 ( 
.A(n_4393),
.B(n_3948),
.C(n_3806),
.Y(n_4965)
);

AO21x2_ASAP7_75t_L g4966 ( 
.A1(n_4346),
.A2(n_3926),
.B(n_3920),
.Y(n_4966)
);

CKINVDCx16_ASAP7_75t_R g4967 ( 
.A(n_4433),
.Y(n_4967)
);

AND2x2_ASAP7_75t_L g4968 ( 
.A(n_4334),
.B(n_4049),
.Y(n_4968)
);

NOR2xp33_ASAP7_75t_R g4969 ( 
.A(n_4433),
.B(n_3948),
.Y(n_4969)
);

INVx2_ASAP7_75t_L g4970 ( 
.A(n_4277),
.Y(n_4970)
);

NAND2xp33_ASAP7_75t_R g4971 ( 
.A(n_4323),
.B(n_3938),
.Y(n_4971)
);

OAI21xp5_ASAP7_75t_SL g4972 ( 
.A1(n_4217),
.A2(n_3899),
.B(n_3842),
.Y(n_4972)
);

AND2x2_ASAP7_75t_L g4973 ( 
.A(n_4334),
.B(n_4125),
.Y(n_4973)
);

INVx1_ASAP7_75t_L g4974 ( 
.A(n_4484),
.Y(n_4974)
);

INVxp67_ASAP7_75t_SL g4975 ( 
.A(n_4232),
.Y(n_4975)
);

OAI21x1_ASAP7_75t_L g4976 ( 
.A1(n_4676),
.A2(n_3953),
.B(n_3951),
.Y(n_4976)
);

AND2x4_ASAP7_75t_L g4977 ( 
.A(n_4310),
.B(n_3842),
.Y(n_4977)
);

AND2x2_ASAP7_75t_L g4978 ( 
.A(n_4344),
.B(n_4125),
.Y(n_4978)
);

AND2x4_ASAP7_75t_L g4979 ( 
.A(n_4209),
.B(n_3899),
.Y(n_4979)
);

INVx1_ASAP7_75t_L g4980 ( 
.A(n_4495),
.Y(n_4980)
);

NAND2xp5_ASAP7_75t_L g4981 ( 
.A(n_4193),
.B(n_3802),
.Y(n_4981)
);

NOR2xp33_ASAP7_75t_R g4982 ( 
.A(n_4483),
.B(n_3948),
.Y(n_4982)
);

INVx2_ASAP7_75t_L g4983 ( 
.A(n_4277),
.Y(n_4983)
);

INVx2_ASAP7_75t_L g4984 ( 
.A(n_4277),
.Y(n_4984)
);

NAND2xp5_ASAP7_75t_L g4985 ( 
.A(n_4193),
.B(n_3802),
.Y(n_4985)
);

CKINVDCx5p33_ASAP7_75t_R g4986 ( 
.A(n_4599),
.Y(n_4986)
);

CKINVDCx5p33_ASAP7_75t_R g4987 ( 
.A(n_4599),
.Y(n_4987)
);

NAND3xp33_ASAP7_75t_SL g4988 ( 
.A(n_4568),
.B(n_3767),
.C(n_3806),
.Y(n_4988)
);

INVxp67_ASAP7_75t_L g4989 ( 
.A(n_4386),
.Y(n_4989)
);

CKINVDCx8_ASAP7_75t_R g4990 ( 
.A(n_4258),
.Y(n_4990)
);

INVx2_ASAP7_75t_L g4991 ( 
.A(n_4280),
.Y(n_4991)
);

HB1xp67_ASAP7_75t_L g4992 ( 
.A(n_4335),
.Y(n_4992)
);

BUFx3_ASAP7_75t_L g4993 ( 
.A(n_4483),
.Y(n_4993)
);

INVx2_ASAP7_75t_L g4994 ( 
.A(n_4280),
.Y(n_4994)
);

AND2x2_ASAP7_75t_L g4995 ( 
.A(n_4344),
.B(n_3899),
.Y(n_4995)
);

AND2x4_ASAP7_75t_SL g4996 ( 
.A(n_4258),
.B(n_3767),
.Y(n_4996)
);

NOR3xp33_ASAP7_75t_SL g4997 ( 
.A(n_4361),
.B(n_3813),
.C(n_3812),
.Y(n_4997)
);

INVx2_ASAP7_75t_L g4998 ( 
.A(n_4280),
.Y(n_4998)
);

INVx4_ASAP7_75t_L g4999 ( 
.A(n_4599),
.Y(n_4999)
);

OA21x2_ASAP7_75t_L g5000 ( 
.A1(n_4425),
.A2(n_3912),
.B(n_3905),
.Y(n_5000)
);

CKINVDCx11_ASAP7_75t_R g5001 ( 
.A(n_4690),
.Y(n_5001)
);

INVx3_ASAP7_75t_L g5002 ( 
.A(n_4302),
.Y(n_5002)
);

INVx1_ASAP7_75t_L g5003 ( 
.A(n_4495),
.Y(n_5003)
);

OR2x6_ASAP7_75t_L g5004 ( 
.A(n_4421),
.B(n_4019),
.Y(n_5004)
);

NOR2xp33_ASAP7_75t_R g5005 ( 
.A(n_4483),
.B(n_4116),
.Y(n_5005)
);

INVx2_ASAP7_75t_SL g5006 ( 
.A(n_4198),
.Y(n_5006)
);

INVx2_ASAP7_75t_L g5007 ( 
.A(n_4282),
.Y(n_5007)
);

CKINVDCx16_ASAP7_75t_R g5008 ( 
.A(n_4690),
.Y(n_5008)
);

INVx1_ASAP7_75t_L g5009 ( 
.A(n_4504),
.Y(n_5009)
);

NAND3xp33_ASAP7_75t_SL g5010 ( 
.A(n_4568),
.B(n_3767),
.C(n_3812),
.Y(n_5010)
);

A2O1A1Ixp33_ASAP7_75t_L g5011 ( 
.A1(n_4632),
.A2(n_3778),
.B(n_3873),
.C(n_3946),
.Y(n_5011)
);

AO32x2_ASAP7_75t_L g5012 ( 
.A1(n_4287),
.A2(n_4083),
.A3(n_4069),
.B1(n_3983),
.B2(n_3991),
.Y(n_5012)
);

BUFx3_ASAP7_75t_L g5013 ( 
.A(n_4690),
.Y(n_5013)
);

BUFx6f_ASAP7_75t_L g5014 ( 
.A(n_4258),
.Y(n_5014)
);

INVx2_ASAP7_75t_L g5015 ( 
.A(n_4282),
.Y(n_5015)
);

NAND2xp33_ASAP7_75t_R g5016 ( 
.A(n_4457),
.B(n_3951),
.Y(n_5016)
);

XNOR2xp5_ASAP7_75t_L g5017 ( 
.A(n_4210),
.B(n_3873),
.Y(n_5017)
);

BUFx10_ASAP7_75t_L g5018 ( 
.A(n_4662),
.Y(n_5018)
);

BUFx3_ASAP7_75t_L g5019 ( 
.A(n_4571),
.Y(n_5019)
);

BUFx2_ASAP7_75t_L g5020 ( 
.A(n_4302),
.Y(n_5020)
);

AND2x4_ASAP7_75t_L g5021 ( 
.A(n_4209),
.B(n_4224),
.Y(n_5021)
);

INVx4_ASAP7_75t_SL g5022 ( 
.A(n_4571),
.Y(n_5022)
);

BUFx2_ASAP7_75t_L g5023 ( 
.A(n_4302),
.Y(n_5023)
);

CKINVDCx5p33_ASAP7_75t_R g5024 ( 
.A(n_4610),
.Y(n_5024)
);

NOR2xp33_ASAP7_75t_R g5025 ( 
.A(n_4652),
.B(n_3873),
.Y(n_5025)
);

NAND2xp33_ASAP7_75t_R g5026 ( 
.A(n_4457),
.B(n_3951),
.Y(n_5026)
);

NAND2xp5_ASAP7_75t_L g5027 ( 
.A(n_4255),
.B(n_3813),
.Y(n_5027)
);

NOR2xp33_ASAP7_75t_R g5028 ( 
.A(n_4652),
.B(n_4104),
.Y(n_5028)
);

OAI21xp5_ASAP7_75t_L g5029 ( 
.A1(n_4285),
.A2(n_3822),
.B(n_3818),
.Y(n_5029)
);

AND2x2_ASAP7_75t_L g5030 ( 
.A(n_4374),
.B(n_3983),
.Y(n_5030)
);

INVx1_ASAP7_75t_SL g5031 ( 
.A(n_4386),
.Y(n_5031)
);

INVx2_ASAP7_75t_L g5032 ( 
.A(n_4282),
.Y(n_5032)
);

INVx2_ASAP7_75t_L g5033 ( 
.A(n_4290),
.Y(n_5033)
);

AND2x4_ASAP7_75t_L g5034 ( 
.A(n_4209),
.B(n_3983),
.Y(n_5034)
);

CKINVDCx16_ASAP7_75t_R g5035 ( 
.A(n_4183),
.Y(n_5035)
);

CKINVDCx5p33_ASAP7_75t_R g5036 ( 
.A(n_4624),
.Y(n_5036)
);

NAND2xp33_ASAP7_75t_R g5037 ( 
.A(n_4457),
.B(n_3951),
.Y(n_5037)
);

AND2x2_ASAP7_75t_L g5038 ( 
.A(n_4374),
.B(n_3991),
.Y(n_5038)
);

NOR3xp33_ASAP7_75t_SL g5039 ( 
.A(n_4361),
.B(n_3822),
.C(n_3818),
.Y(n_5039)
);

HB1xp67_ASAP7_75t_L g5040 ( 
.A(n_4341),
.Y(n_5040)
);

AND2x2_ASAP7_75t_L g5041 ( 
.A(n_4375),
.B(n_3991),
.Y(n_5041)
);

AND2x4_ASAP7_75t_SL g5042 ( 
.A(n_4209),
.B(n_3767),
.Y(n_5042)
);

INVx1_ASAP7_75t_L g5043 ( 
.A(n_4504),
.Y(n_5043)
);

AND2x2_ASAP7_75t_L g5044 ( 
.A(n_4375),
.B(n_4067),
.Y(n_5044)
);

NAND2xp5_ASAP7_75t_L g5045 ( 
.A(n_4255),
.B(n_3824),
.Y(n_5045)
);

AOI22xp33_ASAP7_75t_SL g5046 ( 
.A1(n_4205),
.A2(n_4070),
.B1(n_3974),
.B2(n_3982),
.Y(n_5046)
);

AOI22xp33_ASAP7_75t_SL g5047 ( 
.A1(n_4206),
.A2(n_4070),
.B1(n_3974),
.B2(n_3982),
.Y(n_5047)
);

AND2x4_ASAP7_75t_L g5048 ( 
.A(n_4224),
.B(n_4067),
.Y(n_5048)
);

O2A1O1Ixp5_ASAP7_75t_L g5049 ( 
.A1(n_4445),
.A2(n_3962),
.B(n_3953),
.C(n_4082),
.Y(n_5049)
);

NAND2xp33_ASAP7_75t_R g5050 ( 
.A(n_4457),
.B(n_3953),
.Y(n_5050)
);

INVx1_ASAP7_75t_L g5051 ( 
.A(n_4513),
.Y(n_5051)
);

O2A1O1Ixp33_ASAP7_75t_SL g5052 ( 
.A1(n_4199),
.A2(n_4067),
.B(n_4069),
.C(n_4083),
.Y(n_5052)
);

AND2x2_ASAP7_75t_SL g5053 ( 
.A(n_4206),
.B(n_3712),
.Y(n_5053)
);

AO32x2_ASAP7_75t_L g5054 ( 
.A1(n_4287),
.A2(n_4069),
.A3(n_4160),
.B1(n_4083),
.B2(n_3910),
.Y(n_5054)
);

NAND3xp33_ASAP7_75t_SL g5055 ( 
.A(n_4424),
.B(n_3829),
.C(n_3824),
.Y(n_5055)
);

INVx1_ASAP7_75t_L g5056 ( 
.A(n_4513),
.Y(n_5056)
);

CKINVDCx5p33_ASAP7_75t_R g5057 ( 
.A(n_4423),
.Y(n_5057)
);

OR2x6_ASAP7_75t_L g5058 ( 
.A(n_4421),
.B(n_4019),
.Y(n_5058)
);

INVx2_ASAP7_75t_L g5059 ( 
.A(n_4290),
.Y(n_5059)
);

INVx1_ASAP7_75t_L g5060 ( 
.A(n_4531),
.Y(n_5060)
);

CKINVDCx5p33_ASAP7_75t_R g5061 ( 
.A(n_4579),
.Y(n_5061)
);

INVx1_ASAP7_75t_L g5062 ( 
.A(n_4531),
.Y(n_5062)
);

CKINVDCx5p33_ASAP7_75t_R g5063 ( 
.A(n_4579),
.Y(n_5063)
);

AOI22xp33_ASAP7_75t_L g5064 ( 
.A1(n_4271),
.A2(n_3855),
.B1(n_3974),
.B2(n_3982),
.Y(n_5064)
);

NAND2xp33_ASAP7_75t_SL g5065 ( 
.A(n_4488),
.B(n_3895),
.Y(n_5065)
);

XOR2xp5_ASAP7_75t_L g5066 ( 
.A(n_4664),
.B(n_3829),
.Y(n_5066)
);

OR2x2_ASAP7_75t_L g5067 ( 
.A(n_4272),
.B(n_3838),
.Y(n_5067)
);

INVx2_ASAP7_75t_L g5068 ( 
.A(n_4290),
.Y(n_5068)
);

CKINVDCx5p33_ASAP7_75t_R g5069 ( 
.A(n_4606),
.Y(n_5069)
);

INVx4_ASAP7_75t_L g5070 ( 
.A(n_4571),
.Y(n_5070)
);

NOR2xp33_ASAP7_75t_L g5071 ( 
.A(n_4664),
.B(n_3971),
.Y(n_5071)
);

AND2x2_ASAP7_75t_L g5072 ( 
.A(n_4284),
.B(n_4160),
.Y(n_5072)
);

AND2x6_ASAP7_75t_SL g5073 ( 
.A(n_4199),
.B(n_3971),
.Y(n_5073)
);

CKINVDCx20_ASAP7_75t_R g5074 ( 
.A(n_4198),
.Y(n_5074)
);

AND2x2_ASAP7_75t_L g5075 ( 
.A(n_4284),
.B(n_4160),
.Y(n_5075)
);

INVx2_ASAP7_75t_L g5076 ( 
.A(n_4326),
.Y(n_5076)
);

AOI22xp33_ASAP7_75t_L g5077 ( 
.A1(n_4490),
.A2(n_4028),
.B1(n_3982),
.B2(n_3987),
.Y(n_5077)
);

AOI22xp33_ASAP7_75t_L g5078 ( 
.A1(n_4490),
.A2(n_3852),
.B1(n_4045),
.B2(n_3987),
.Y(n_5078)
);

NAND2xp5_ASAP7_75t_L g5079 ( 
.A(n_4295),
.B(n_3838),
.Y(n_5079)
);

NAND2xp33_ASAP7_75t_R g5080 ( 
.A(n_4673),
.B(n_3953),
.Y(n_5080)
);

NAND2xp5_ASAP7_75t_L g5081 ( 
.A(n_4295),
.B(n_3856),
.Y(n_5081)
);

INVx4_ASAP7_75t_SL g5082 ( 
.A(n_4571),
.Y(n_5082)
);

CKINVDCx5p33_ASAP7_75t_R g5083 ( 
.A(n_4606),
.Y(n_5083)
);

BUFx6f_ASAP7_75t_L g5084 ( 
.A(n_4430),
.Y(n_5084)
);

INVx1_ASAP7_75t_SL g5085 ( 
.A(n_4553),
.Y(n_5085)
);

AND2x4_ASAP7_75t_L g5086 ( 
.A(n_4224),
.B(n_4268),
.Y(n_5086)
);

AOI22xp33_ASAP7_75t_L g5087 ( 
.A1(n_4523),
.A2(n_4446),
.B1(n_4444),
.B2(n_4318),
.Y(n_5087)
);

AOI22xp33_ASAP7_75t_L g5088 ( 
.A1(n_4523),
.A2(n_4029),
.B1(n_3987),
.B2(n_3988),
.Y(n_5088)
);

NOR3xp33_ASAP7_75t_SL g5089 ( 
.A(n_4185),
.B(n_3858),
.C(n_3856),
.Y(n_5089)
);

NOR2xp33_ASAP7_75t_R g5090 ( 
.A(n_4652),
.B(n_4104),
.Y(n_5090)
);

BUFx6f_ASAP7_75t_L g5091 ( 
.A(n_4430),
.Y(n_5091)
);

NAND2xp5_ASAP7_75t_L g5092 ( 
.A(n_4299),
.B(n_4311),
.Y(n_5092)
);

AND2x2_ASAP7_75t_L g5093 ( 
.A(n_4297),
.B(n_3784),
.Y(n_5093)
);

INVx2_ASAP7_75t_L g5094 ( 
.A(n_4326),
.Y(n_5094)
);

HB1xp67_ASAP7_75t_SL g5095 ( 
.A(n_4652),
.Y(n_5095)
);

OR2x6_ASAP7_75t_L g5096 ( 
.A(n_4391),
.B(n_4019),
.Y(n_5096)
);

INVx1_ASAP7_75t_L g5097 ( 
.A(n_4535),
.Y(n_5097)
);

NAND2xp33_ASAP7_75t_R g5098 ( 
.A(n_4673),
.B(n_3962),
.Y(n_5098)
);

AND2x2_ASAP7_75t_L g5099 ( 
.A(n_4297),
.B(n_3784),
.Y(n_5099)
);

CKINVDCx5p33_ASAP7_75t_R g5100 ( 
.A(n_4625),
.Y(n_5100)
);

INVx2_ASAP7_75t_L g5101 ( 
.A(n_4326),
.Y(n_5101)
);

A2O1A1Ixp33_ASAP7_75t_L g5102 ( 
.A1(n_4275),
.A2(n_3939),
.B(n_3949),
.C(n_3743),
.Y(n_5102)
);

NOR2xp33_ASAP7_75t_R g5103 ( 
.A(n_4652),
.B(n_4104),
.Y(n_5103)
);

AND2x4_ASAP7_75t_L g5104 ( 
.A(n_4224),
.B(n_3962),
.Y(n_5104)
);

CKINVDCx5p33_ASAP7_75t_R g5105 ( 
.A(n_4625),
.Y(n_5105)
);

AND2x2_ASAP7_75t_SL g5106 ( 
.A(n_4662),
.B(n_3712),
.Y(n_5106)
);

AND2x2_ASAP7_75t_L g5107 ( 
.A(n_4207),
.B(n_3784),
.Y(n_5107)
);

NAND2xp5_ASAP7_75t_SL g5108 ( 
.A(n_4330),
.B(n_3712),
.Y(n_5108)
);

INVx2_ASAP7_75t_SL g5109 ( 
.A(n_4198),
.Y(n_5109)
);

INVx2_ASAP7_75t_L g5110 ( 
.A(n_4356),
.Y(n_5110)
);

NAND2xp5_ASAP7_75t_L g5111 ( 
.A(n_4299),
.B(n_3858),
.Y(n_5111)
);

NOR2x1_ASAP7_75t_L g5112 ( 
.A(n_4343),
.B(n_3962),
.Y(n_5112)
);

AND2x2_ASAP7_75t_L g5113 ( 
.A(n_4207),
.B(n_4187),
.Y(n_5113)
);

AOI21xp5_ASAP7_75t_L g5114 ( 
.A1(n_4266),
.A2(n_3743),
.B(n_3712),
.Y(n_5114)
);

INVxp67_ASAP7_75t_L g5115 ( 
.A(n_4311),
.Y(n_5115)
);

INVx1_ASAP7_75t_L g5116 ( 
.A(n_4535),
.Y(n_5116)
);

AND2x2_ASAP7_75t_L g5117 ( 
.A(n_4187),
.B(n_3784),
.Y(n_5117)
);

INVx2_ASAP7_75t_L g5118 ( 
.A(n_4356),
.Y(n_5118)
);

INVxp33_ASAP7_75t_SL g5119 ( 
.A(n_4529),
.Y(n_5119)
);

NAND2x1p5_ASAP7_75t_L g5120 ( 
.A(n_4680),
.B(n_3743),
.Y(n_5120)
);

AND2x2_ASAP7_75t_L g5121 ( 
.A(n_4215),
.B(n_4394),
.Y(n_5121)
);

CKINVDCx5p33_ASAP7_75t_R g5122 ( 
.A(n_4553),
.Y(n_5122)
);

HB1xp67_ASAP7_75t_L g5123 ( 
.A(n_4341),
.Y(n_5123)
);

OAI22xp5_ASAP7_75t_L g5124 ( 
.A1(n_4349),
.A2(n_4107),
.B1(n_4108),
.B2(n_4147),
.Y(n_5124)
);

NAND2xp5_ASAP7_75t_L g5125 ( 
.A(n_4257),
.B(n_3859),
.Y(n_5125)
);

NOR3xp33_ASAP7_75t_SL g5126 ( 
.A(n_4185),
.B(n_3872),
.C(n_3859),
.Y(n_5126)
);

INVx3_ASAP7_75t_L g5127 ( 
.A(n_4302),
.Y(n_5127)
);

AO31x2_ASAP7_75t_L g5128 ( 
.A1(n_4425),
.A2(n_4046),
.A3(n_4042),
.B(n_4032),
.Y(n_5128)
);

BUFx6f_ASAP7_75t_L g5129 ( 
.A(n_4430),
.Y(n_5129)
);

OAI22xp33_ASAP7_75t_L g5130 ( 
.A1(n_4213),
.A2(n_3852),
.B1(n_3987),
.B2(n_4006),
.Y(n_5130)
);

CKINVDCx16_ASAP7_75t_R g5131 ( 
.A(n_4304),
.Y(n_5131)
);

CKINVDCx20_ASAP7_75t_R g5132 ( 
.A(n_4303),
.Y(n_5132)
);

CKINVDCx5p33_ASAP7_75t_R g5133 ( 
.A(n_4304),
.Y(n_5133)
);

A2O1A1Ixp33_ASAP7_75t_L g5134 ( 
.A1(n_4275),
.A2(n_3743),
.B(n_4082),
.C(n_4168),
.Y(n_5134)
);

INVx1_ASAP7_75t_L g5135 ( 
.A(n_4537),
.Y(n_5135)
);

AO31x2_ASAP7_75t_L g5136 ( 
.A1(n_4318),
.A2(n_4214),
.A3(n_4377),
.B(n_4352),
.Y(n_5136)
);

OR2x6_ASAP7_75t_L g5137 ( 
.A(n_4391),
.B(n_4019),
.Y(n_5137)
);

NOR2xp33_ASAP7_75t_R g5138 ( 
.A(n_4652),
.B(n_4104),
.Y(n_5138)
);

AND2x2_ASAP7_75t_L g5139 ( 
.A(n_4215),
.B(n_3798),
.Y(n_5139)
);

OAI21x1_ASAP7_75t_L g5140 ( 
.A1(n_4498),
.A2(n_4168),
.B(n_4082),
.Y(n_5140)
);

INVx1_ASAP7_75t_L g5141 ( 
.A(n_4537),
.Y(n_5141)
);

NAND2xp5_ASAP7_75t_L g5142 ( 
.A(n_4257),
.B(n_3872),
.Y(n_5142)
);

AND2x2_ASAP7_75t_L g5143 ( 
.A(n_4394),
.B(n_3798),
.Y(n_5143)
);

INVx1_ASAP7_75t_L g5144 ( 
.A(n_4554),
.Y(n_5144)
);

NAND3xp33_ASAP7_75t_L g5145 ( 
.A(n_4197),
.B(n_3913),
.C(n_3874),
.Y(n_5145)
);

INVx6_ASAP7_75t_L g5146 ( 
.A(n_4399),
.Y(n_5146)
);

INVx2_ASAP7_75t_L g5147 ( 
.A(n_4356),
.Y(n_5147)
);

OAI222xp33_ASAP7_75t_L g5148 ( 
.A1(n_4469),
.A2(n_3847),
.B1(n_3877),
.B2(n_3871),
.C1(n_3870),
.C2(n_3861),
.Y(n_5148)
);

INVx2_ASAP7_75t_SL g5149 ( 
.A(n_4303),
.Y(n_5149)
);

INVx1_ASAP7_75t_L g5150 ( 
.A(n_4554),
.Y(n_5150)
);

AND2x2_ASAP7_75t_L g5151 ( 
.A(n_4403),
.B(n_3798),
.Y(n_5151)
);

INVx2_ASAP7_75t_L g5152 ( 
.A(n_4410),
.Y(n_5152)
);

HB1xp67_ASAP7_75t_L g5153 ( 
.A(n_4414),
.Y(n_5153)
);

NOR3xp33_ASAP7_75t_SL g5154 ( 
.A(n_4197),
.B(n_3913),
.C(n_3874),
.Y(n_5154)
);

BUFx3_ASAP7_75t_L g5155 ( 
.A(n_4571),
.Y(n_5155)
);

INVx1_ASAP7_75t_L g5156 ( 
.A(n_4583),
.Y(n_5156)
);

INVxp67_ASAP7_75t_L g5157 ( 
.A(n_4576),
.Y(n_5157)
);

AND2x4_ASAP7_75t_L g5158 ( 
.A(n_4268),
.B(n_4082),
.Y(n_5158)
);

NAND2xp5_ASAP7_75t_SL g5159 ( 
.A(n_4580),
.B(n_3798),
.Y(n_5159)
);

AO32x2_ASAP7_75t_L g5160 ( 
.A1(n_4312),
.A2(n_3910),
.A3(n_3895),
.B1(n_3847),
.B2(n_4124),
.Y(n_5160)
);

BUFx3_ASAP7_75t_L g5161 ( 
.A(n_4571),
.Y(n_5161)
);

INVx1_ASAP7_75t_L g5162 ( 
.A(n_4583),
.Y(n_5162)
);

INVx1_ASAP7_75t_L g5163 ( 
.A(n_4607),
.Y(n_5163)
);

CKINVDCx12_ASAP7_75t_R g5164 ( 
.A(n_4699),
.Y(n_5164)
);

BUFx6f_ASAP7_75t_L g5165 ( 
.A(n_4430),
.Y(n_5165)
);

HB1xp67_ASAP7_75t_L g5166 ( 
.A(n_4414),
.Y(n_5166)
);

OAI22xp5_ASAP7_75t_L g5167 ( 
.A1(n_4349),
.A2(n_4147),
.B1(n_4108),
.B2(n_4107),
.Y(n_5167)
);

AND2x4_ASAP7_75t_SL g5168 ( 
.A(n_4268),
.B(n_3880),
.Y(n_5168)
);

CKINVDCx12_ASAP7_75t_R g5169 ( 
.A(n_4699),
.Y(n_5169)
);

INVx1_ASAP7_75t_L g5170 ( 
.A(n_4607),
.Y(n_5170)
);

AND2x2_ASAP7_75t_L g5171 ( 
.A(n_4403),
.B(n_3880),
.Y(n_5171)
);

INVx2_ASAP7_75t_L g5172 ( 
.A(n_4410),
.Y(n_5172)
);

AOI22xp33_ASAP7_75t_L g5173 ( 
.A1(n_4446),
.A2(n_4077),
.B1(n_4070),
.B2(n_4056),
.Y(n_5173)
);

NOR2xp33_ASAP7_75t_L g5174 ( 
.A(n_4413),
.B(n_4288),
.Y(n_5174)
);

INVx1_ASAP7_75t_L g5175 ( 
.A(n_4608),
.Y(n_5175)
);

INVx1_ASAP7_75t_L g5176 ( 
.A(n_4608),
.Y(n_5176)
);

INVx1_ASAP7_75t_L g5177 ( 
.A(n_4612),
.Y(n_5177)
);

BUFx2_ASAP7_75t_L g5178 ( 
.A(n_4571),
.Y(n_5178)
);

INVx1_ASAP7_75t_L g5179 ( 
.A(n_4612),
.Y(n_5179)
);

CKINVDCx16_ASAP7_75t_R g5180 ( 
.A(n_4337),
.Y(n_5180)
);

INVx1_ASAP7_75t_L g5181 ( 
.A(n_4634),
.Y(n_5181)
);

NAND2xp5_ASAP7_75t_L g5182 ( 
.A(n_4413),
.B(n_3923),
.Y(n_5182)
);

INVx1_ASAP7_75t_L g5183 ( 
.A(n_4634),
.Y(n_5183)
);

BUFx2_ASAP7_75t_L g5184 ( 
.A(n_4665),
.Y(n_5184)
);

AOI22xp33_ASAP7_75t_L g5185 ( 
.A1(n_4446),
.A2(n_4077),
.B1(n_4070),
.B2(n_4056),
.Y(n_5185)
);

INVx2_ASAP7_75t_SL g5186 ( 
.A(n_4303),
.Y(n_5186)
);

NAND3xp33_ASAP7_75t_L g5187 ( 
.A(n_4202),
.B(n_4093),
.C(n_4091),
.Y(n_5187)
);

AND2x2_ASAP7_75t_L g5188 ( 
.A(n_4488),
.B(n_4489),
.Y(n_5188)
);

NAND2xp5_ASAP7_75t_L g5189 ( 
.A(n_4248),
.B(n_3923),
.Y(n_5189)
);

AO31x2_ASAP7_75t_L g5190 ( 
.A1(n_4214),
.A2(n_4111),
.A3(n_4078),
.B(n_4046),
.Y(n_5190)
);

INVx1_ASAP7_75t_L g5191 ( 
.A(n_4641),
.Y(n_5191)
);

NAND2xp5_ASAP7_75t_L g5192 ( 
.A(n_4248),
.B(n_3925),
.Y(n_5192)
);

CKINVDCx16_ASAP7_75t_R g5193 ( 
.A(n_4337),
.Y(n_5193)
);

BUFx2_ASAP7_75t_SL g5194 ( 
.A(n_4300),
.Y(n_5194)
);

INVx2_ASAP7_75t_L g5195 ( 
.A(n_4716),
.Y(n_5195)
);

INVx2_ASAP7_75t_L g5196 ( 
.A(n_4716),
.Y(n_5196)
);

AO21x2_ASAP7_75t_L g5197 ( 
.A1(n_4962),
.A2(n_4232),
.B(n_4679),
.Y(n_5197)
);

BUFx6f_ASAP7_75t_SL g5198 ( 
.A(n_4725),
.Y(n_5198)
);

OAI222xp33_ASAP7_75t_L g5199 ( 
.A1(n_5035),
.A2(n_4672),
.B1(n_4234),
.B2(n_4240),
.C1(n_4213),
.C2(n_4613),
.Y(n_5199)
);

INVx1_ASAP7_75t_L g5200 ( 
.A(n_4724),
.Y(n_5200)
);

INVxp67_ASAP7_75t_SL g5201 ( 
.A(n_4717),
.Y(n_5201)
);

INVx2_ASAP7_75t_L g5202 ( 
.A(n_4716),
.Y(n_5202)
);

INVx2_ASAP7_75t_L g5203 ( 
.A(n_4716),
.Y(n_5203)
);

INVxp67_ASAP7_75t_L g5204 ( 
.A(n_4885),
.Y(n_5204)
);

INVx1_ASAP7_75t_SL g5205 ( 
.A(n_4870),
.Y(n_5205)
);

AND2x2_ASAP7_75t_L g5206 ( 
.A(n_5113),
.B(n_4675),
.Y(n_5206)
);

AOI21xp5_ASAP7_75t_SL g5207 ( 
.A1(n_4881),
.A2(n_4493),
.B(n_4672),
.Y(n_5207)
);

AOI222xp33_ASAP7_75t_L g5208 ( 
.A1(n_4769),
.A2(n_4221),
.B1(n_4353),
.B2(n_4613),
.C1(n_4617),
.C2(n_4321),
.Y(n_5208)
);

INVx2_ASAP7_75t_L g5209 ( 
.A(n_4716),
.Y(n_5209)
);

AOI211x1_ASAP7_75t_L g5210 ( 
.A1(n_4925),
.A2(n_4221),
.B(n_4202),
.C(n_4312),
.Y(n_5210)
);

OA21x2_ASAP7_75t_L g5211 ( 
.A1(n_5087),
.A2(n_4289),
.B(n_4264),
.Y(n_5211)
);

INVx2_ASAP7_75t_L g5212 ( 
.A(n_4716),
.Y(n_5212)
);

OAI21xp5_ASAP7_75t_L g5213 ( 
.A1(n_4886),
.A2(n_4243),
.B(n_4316),
.Y(n_5213)
);

NAND2xp33_ASAP7_75t_R g5214 ( 
.A(n_4859),
.B(n_4675),
.Y(n_5214)
);

INVx2_ASAP7_75t_L g5215 ( 
.A(n_4784),
.Y(n_5215)
);

INVx1_ASAP7_75t_L g5216 ( 
.A(n_4724),
.Y(n_5216)
);

INVx2_ASAP7_75t_SL g5217 ( 
.A(n_5146),
.Y(n_5217)
);

HB1xp67_ASAP7_75t_L g5218 ( 
.A(n_4755),
.Y(n_5218)
);

INVx1_ASAP7_75t_L g5219 ( 
.A(n_4743),
.Y(n_5219)
);

BUFx6f_ASAP7_75t_L g5220 ( 
.A(n_4764),
.Y(n_5220)
);

INVx3_ASAP7_75t_L g5221 ( 
.A(n_4962),
.Y(n_5221)
);

AND2x2_ASAP7_75t_L g5222 ( 
.A(n_5113),
.B(n_4195),
.Y(n_5222)
);

INVx2_ASAP7_75t_L g5223 ( 
.A(n_4784),
.Y(n_5223)
);

NAND2xp5_ASAP7_75t_L g5224 ( 
.A(n_4776),
.B(n_4254),
.Y(n_5224)
);

AOI221xp5_ASAP7_75t_L g5225 ( 
.A1(n_4708),
.A2(n_4327),
.B1(n_4240),
.B2(n_4234),
.C(n_4353),
.Y(n_5225)
);

INVx4_ASAP7_75t_L g5226 ( 
.A(n_4764),
.Y(n_5226)
);

INVx2_ASAP7_75t_SL g5227 ( 
.A(n_5146),
.Y(n_5227)
);

INVx1_ASAP7_75t_L g5228 ( 
.A(n_4743),
.Y(n_5228)
);

BUFx3_ASAP7_75t_L g5229 ( 
.A(n_4876),
.Y(n_5229)
);

OR2x2_ASAP7_75t_L g5230 ( 
.A(n_5035),
.B(n_4254),
.Y(n_5230)
);

OR2x6_ASAP7_75t_L g5231 ( 
.A(n_4881),
.B(n_4266),
.Y(n_5231)
);

OR2x2_ASAP7_75t_L g5232 ( 
.A(n_4888),
.B(n_4397),
.Y(n_5232)
);

INVx4_ASAP7_75t_L g5233 ( 
.A(n_4732),
.Y(n_5233)
);

INVx1_ASAP7_75t_L g5234 ( 
.A(n_4747),
.Y(n_5234)
);

AND2x2_ASAP7_75t_L g5235 ( 
.A(n_5053),
.B(n_4195),
.Y(n_5235)
);

INVx3_ASAP7_75t_L g5236 ( 
.A(n_4962),
.Y(n_5236)
);

BUFx2_ASAP7_75t_L g5237 ( 
.A(n_4727),
.Y(n_5237)
);

AND2x2_ASAP7_75t_L g5238 ( 
.A(n_5053),
.B(n_4195),
.Y(n_5238)
);

INVx2_ASAP7_75t_L g5239 ( 
.A(n_4784),
.Y(n_5239)
);

INVx1_ASAP7_75t_L g5240 ( 
.A(n_4747),
.Y(n_5240)
);

AND2x2_ASAP7_75t_L g5241 ( 
.A(n_5053),
.B(n_4195),
.Y(n_5241)
);

AND2x2_ASAP7_75t_L g5242 ( 
.A(n_4727),
.B(n_4489),
.Y(n_5242)
);

AO21x2_ASAP7_75t_L g5243 ( 
.A1(n_4723),
.A2(n_4834),
.B(n_4737),
.Y(n_5243)
);

OR2x6_ASAP7_75t_L g5244 ( 
.A(n_4881),
.B(n_4429),
.Y(n_5244)
);

INVx2_ASAP7_75t_L g5245 ( 
.A(n_4784),
.Y(n_5245)
);

AND2x2_ASAP7_75t_L g5246 ( 
.A(n_4854),
.B(n_4665),
.Y(n_5246)
);

INVx1_ASAP7_75t_L g5247 ( 
.A(n_4766),
.Y(n_5247)
);

INVx1_ASAP7_75t_L g5248 ( 
.A(n_4766),
.Y(n_5248)
);

AND2x2_ASAP7_75t_L g5249 ( 
.A(n_4854),
.B(n_4669),
.Y(n_5249)
);

INVx1_ASAP7_75t_L g5250 ( 
.A(n_4789),
.Y(n_5250)
);

OA21x2_ASAP7_75t_L g5251 ( 
.A1(n_5140),
.A2(n_4289),
.B(n_4264),
.Y(n_5251)
);

OAI221xp5_ASAP7_75t_L g5252 ( 
.A1(n_4826),
.A2(n_4372),
.B1(n_4510),
.B2(n_4392),
.C(n_4657),
.Y(n_5252)
);

AO21x2_ASAP7_75t_L g5253 ( 
.A1(n_4834),
.A2(n_4405),
.B(n_4350),
.Y(n_5253)
);

INVx3_ASAP7_75t_L g5254 ( 
.A(n_5136),
.Y(n_5254)
);

AND2x2_ASAP7_75t_L g5255 ( 
.A(n_5121),
.B(n_4669),
.Y(n_5255)
);

INVx1_ASAP7_75t_L g5256 ( 
.A(n_4789),
.Y(n_5256)
);

INVx1_ASAP7_75t_L g5257 ( 
.A(n_4798),
.Y(n_5257)
);

OAI21xp5_ASAP7_75t_L g5258 ( 
.A1(n_5089),
.A2(n_4539),
.B(n_4409),
.Y(n_5258)
);

HB1xp67_ASAP7_75t_L g5259 ( 
.A(n_4726),
.Y(n_5259)
);

INVx1_ASAP7_75t_SL g5260 ( 
.A(n_4889),
.Y(n_5260)
);

INVx2_ASAP7_75t_L g5261 ( 
.A(n_4784),
.Y(n_5261)
);

BUFx2_ASAP7_75t_L g5262 ( 
.A(n_4833),
.Y(n_5262)
);

AOI222xp33_ASAP7_75t_L g5263 ( 
.A1(n_4964),
.A2(n_4617),
.B1(n_4321),
.B2(n_4493),
.C1(n_4451),
.C2(n_4300),
.Y(n_5263)
);

NOR2xp33_ASAP7_75t_L g5264 ( 
.A(n_4773),
.B(n_4288),
.Y(n_5264)
);

AND2x2_ASAP7_75t_L g5265 ( 
.A(n_5121),
.B(n_5042),
.Y(n_5265)
);

AO21x2_ASAP7_75t_L g5266 ( 
.A1(n_4834),
.A2(n_4405),
.B(n_4657),
.Y(n_5266)
);

AOI21xp5_ASAP7_75t_SL g5267 ( 
.A1(n_4881),
.A2(n_4418),
.B(n_4373),
.Y(n_5267)
);

NAND2xp5_ASAP7_75t_L g5268 ( 
.A(n_4917),
.B(n_4322),
.Y(n_5268)
);

INVx1_ASAP7_75t_L g5269 ( 
.A(n_4798),
.Y(n_5269)
);

AND2x2_ASAP7_75t_L g5270 ( 
.A(n_5042),
.B(n_4622),
.Y(n_5270)
);

AO21x2_ASAP7_75t_L g5271 ( 
.A1(n_4710),
.A2(n_4262),
.B(n_4401),
.Y(n_5271)
);

AOI21x1_ASAP7_75t_L g5272 ( 
.A1(n_4881),
.A2(n_4381),
.B(n_4354),
.Y(n_5272)
);

AND2x4_ASAP7_75t_L g5273 ( 
.A(n_5022),
.B(n_4348),
.Y(n_5273)
);

AO21x2_ASAP7_75t_L g5274 ( 
.A1(n_4710),
.A2(n_4401),
.B(n_4292),
.Y(n_5274)
);

INVx2_ASAP7_75t_SL g5275 ( 
.A(n_5146),
.Y(n_5275)
);

INVxp67_ASAP7_75t_SL g5276 ( 
.A(n_4717),
.Y(n_5276)
);

AND2x2_ASAP7_75t_L g5277 ( 
.A(n_5042),
.B(n_4268),
.Y(n_5277)
);

INVx1_ASAP7_75t_L g5278 ( 
.A(n_4803),
.Y(n_5278)
);

AO21x2_ASAP7_75t_L g5279 ( 
.A1(n_4710),
.A2(n_4411),
.B(n_4562),
.Y(n_5279)
);

AOI221xp5_ASAP7_75t_L g5280 ( 
.A1(n_4763),
.A2(n_4367),
.B1(n_4562),
.B2(n_4567),
.C(n_4572),
.Y(n_5280)
);

INVx2_ASAP7_75t_SL g5281 ( 
.A(n_5146),
.Y(n_5281)
);

AND2x2_ASAP7_75t_L g5282 ( 
.A(n_4821),
.B(n_4406),
.Y(n_5282)
);

INVx1_ASAP7_75t_L g5283 ( 
.A(n_4803),
.Y(n_5283)
);

INVx2_ASAP7_75t_L g5284 ( 
.A(n_4784),
.Y(n_5284)
);

AND2x2_ASAP7_75t_L g5285 ( 
.A(n_4821),
.B(n_4541),
.Y(n_5285)
);

INVx2_ASAP7_75t_SL g5286 ( 
.A(n_5112),
.Y(n_5286)
);

BUFx2_ASAP7_75t_L g5287 ( 
.A(n_4892),
.Y(n_5287)
);

AND2x2_ASAP7_75t_L g5288 ( 
.A(n_4821),
.B(n_4541),
.Y(n_5288)
);

AOI21x1_ASAP7_75t_L g5289 ( 
.A1(n_4938),
.A2(n_4381),
.B(n_4354),
.Y(n_5289)
);

AND2x2_ASAP7_75t_L g5290 ( 
.A(n_4757),
.B(n_4320),
.Y(n_5290)
);

AND2x2_ASAP7_75t_L g5291 ( 
.A(n_4757),
.B(n_4320),
.Y(n_5291)
);

INVx1_ASAP7_75t_L g5292 ( 
.A(n_4805),
.Y(n_5292)
);

INVx1_ASAP7_75t_L g5293 ( 
.A(n_4805),
.Y(n_5293)
);

INVx1_ASAP7_75t_L g5294 ( 
.A(n_4808),
.Y(n_5294)
);

HB1xp67_ASAP7_75t_L g5295 ( 
.A(n_4745),
.Y(n_5295)
);

AND2x2_ASAP7_75t_L g5296 ( 
.A(n_4757),
.B(n_4441),
.Y(n_5296)
);

AOI21x1_ASAP7_75t_L g5297 ( 
.A1(n_4938),
.A2(n_4382),
.B(n_4453),
.Y(n_5297)
);

INVx1_ASAP7_75t_L g5298 ( 
.A(n_4808),
.Y(n_5298)
);

AND2x4_ASAP7_75t_L g5299 ( 
.A(n_5022),
.B(n_4348),
.Y(n_5299)
);

AND2x2_ASAP7_75t_L g5300 ( 
.A(n_4757),
.B(n_4453),
.Y(n_5300)
);

BUFx6f_ASAP7_75t_L g5301 ( 
.A(n_4725),
.Y(n_5301)
);

INVx2_ASAP7_75t_L g5302 ( 
.A(n_4966),
.Y(n_5302)
);

BUFx2_ASAP7_75t_L g5303 ( 
.A(n_4912),
.Y(n_5303)
);

OA21x2_ASAP7_75t_L g5304 ( 
.A1(n_5140),
.A2(n_4491),
.B(n_4473),
.Y(n_5304)
);

INVx5_ASAP7_75t_SL g5305 ( 
.A(n_4759),
.Y(n_5305)
);

INVx2_ASAP7_75t_L g5306 ( 
.A(n_4966),
.Y(n_5306)
);

INVx1_ASAP7_75t_L g5307 ( 
.A(n_4812),
.Y(n_5307)
);

BUFx3_ASAP7_75t_L g5308 ( 
.A(n_4756),
.Y(n_5308)
);

AO21x2_ASAP7_75t_L g5309 ( 
.A1(n_4737),
.A2(n_4411),
.B(n_4567),
.Y(n_5309)
);

AND2x2_ASAP7_75t_L g5310 ( 
.A(n_4852),
.B(n_4464),
.Y(n_5310)
);

INVx1_ASAP7_75t_L g5311 ( 
.A(n_4812),
.Y(n_5311)
);

NOR2xp33_ASAP7_75t_L g5312 ( 
.A(n_4773),
.B(n_4623),
.Y(n_5312)
);

INVx1_ASAP7_75t_L g5313 ( 
.A(n_4820),
.Y(n_5313)
);

BUFx4f_ASAP7_75t_SL g5314 ( 
.A(n_4761),
.Y(n_5314)
);

INVx2_ASAP7_75t_L g5315 ( 
.A(n_4966),
.Y(n_5315)
);

INVxp67_ASAP7_75t_SL g5316 ( 
.A(n_5017),
.Y(n_5316)
);

INVx1_ASAP7_75t_L g5317 ( 
.A(n_4820),
.Y(n_5317)
);

OAI22xp5_ASAP7_75t_L g5318 ( 
.A1(n_5131),
.A2(n_4365),
.B1(n_4269),
.B2(n_4345),
.Y(n_5318)
);

INVxp67_ASAP7_75t_SL g5319 ( 
.A(n_5017),
.Y(n_5319)
);

OA21x2_ASAP7_75t_L g5320 ( 
.A1(n_5049),
.A2(n_4472),
.B(n_4471),
.Y(n_5320)
);

NAND2xp5_ASAP7_75t_L g5321 ( 
.A(n_4959),
.B(n_4322),
.Y(n_5321)
);

INVxp67_ASAP7_75t_SL g5322 ( 
.A(n_4785),
.Y(n_5322)
);

INVx1_ASAP7_75t_L g5323 ( 
.A(n_4823),
.Y(n_5323)
);

INVx1_ASAP7_75t_SL g5324 ( 
.A(n_4901),
.Y(n_5324)
);

AOI221xp5_ASAP7_75t_L g5325 ( 
.A1(n_5131),
.A2(n_5055),
.B1(n_4902),
.B2(n_5145),
.C(n_5187),
.Y(n_5325)
);

INVx5_ASAP7_75t_SL g5326 ( 
.A(n_4759),
.Y(n_5326)
);

BUFx2_ASAP7_75t_L g5327 ( 
.A(n_4753),
.Y(n_5327)
);

OR2x2_ASAP7_75t_L g5328 ( 
.A(n_4811),
.B(n_4397),
.Y(n_5328)
);

NAND2xp5_ASAP7_75t_L g5329 ( 
.A(n_5115),
.B(n_4329),
.Y(n_5329)
);

INVx2_ASAP7_75t_L g5330 ( 
.A(n_5128),
.Y(n_5330)
);

INVx1_ASAP7_75t_L g5331 ( 
.A(n_4823),
.Y(n_5331)
);

INVx1_ASAP7_75t_L g5332 ( 
.A(n_4829),
.Y(n_5332)
);

OA21x2_ASAP7_75t_L g5333 ( 
.A1(n_5187),
.A2(n_4640),
.B(n_4636),
.Y(n_5333)
);

INVx1_ASAP7_75t_L g5334 ( 
.A(n_4829),
.Y(n_5334)
);

NOR2xp33_ASAP7_75t_L g5335 ( 
.A(n_4783),
.B(n_4623),
.Y(n_5335)
);

INVx1_ASAP7_75t_L g5336 ( 
.A(n_4839),
.Y(n_5336)
);

OR2x2_ASAP7_75t_L g5337 ( 
.A(n_4857),
.B(n_4247),
.Y(n_5337)
);

INVx1_ASAP7_75t_L g5338 ( 
.A(n_4839),
.Y(n_5338)
);

HB1xp67_ASAP7_75t_L g5339 ( 
.A(n_4768),
.Y(n_5339)
);

AND2x4_ASAP7_75t_SL g5340 ( 
.A(n_5074),
.B(n_4694),
.Y(n_5340)
);

AND2x2_ASAP7_75t_L g5341 ( 
.A(n_4852),
.B(n_4576),
.Y(n_5341)
);

AOI22xp33_ASAP7_75t_L g5342 ( 
.A1(n_5000),
.A2(n_4446),
.B1(n_4444),
.B2(n_4533),
.Y(n_5342)
);

INVx1_ASAP7_75t_L g5343 ( 
.A(n_4860),
.Y(n_5343)
);

OR2x6_ASAP7_75t_L g5344 ( 
.A(n_4938),
.B(n_5194),
.Y(n_5344)
);

OAI222xp33_ASAP7_75t_L g5345 ( 
.A1(n_4938),
.A2(n_4267),
.B1(n_4469),
.B2(n_4580),
.C1(n_4616),
.C2(n_4604),
.Y(n_5345)
);

OA21x2_ASAP7_75t_L g5346 ( 
.A1(n_5145),
.A2(n_4695),
.B(n_4685),
.Y(n_5346)
);

INVx1_ASAP7_75t_L g5347 ( 
.A(n_4860),
.Y(n_5347)
);

NAND2xp5_ASAP7_75t_L g5348 ( 
.A(n_5092),
.B(n_4641),
.Y(n_5348)
);

NOR2xp33_ASAP7_75t_L g5349 ( 
.A(n_4783),
.B(n_4431),
.Y(n_5349)
);

NAND2xp5_ASAP7_75t_L g5350 ( 
.A(n_5126),
.B(n_4658),
.Y(n_5350)
);

NOR2x1p5_ASAP7_75t_L g5351 ( 
.A(n_4732),
.B(n_4455),
.Y(n_5351)
);

INVx2_ASAP7_75t_L g5352 ( 
.A(n_5128),
.Y(n_5352)
);

INVx1_ASAP7_75t_L g5353 ( 
.A(n_4861),
.Y(n_5353)
);

INVx3_ASAP7_75t_L g5354 ( 
.A(n_5136),
.Y(n_5354)
);

OA21x2_ASAP7_75t_L g5355 ( 
.A1(n_5148),
.A2(n_4695),
.B(n_4685),
.Y(n_5355)
);

INVx1_ASAP7_75t_L g5356 ( 
.A(n_4861),
.Y(n_5356)
);

AND2x2_ASAP7_75t_L g5357 ( 
.A(n_4852),
.B(n_4427),
.Y(n_5357)
);

AO21x2_ASAP7_75t_L g5358 ( 
.A1(n_4737),
.A2(n_4750),
.B(n_4742),
.Y(n_5358)
);

OAI221xp5_ASAP7_75t_L g5359 ( 
.A1(n_4754),
.A2(n_4372),
.B1(n_4474),
.B2(n_4438),
.C(n_4351),
.Y(n_5359)
);

NAND2xp5_ASAP7_75t_L g5360 ( 
.A(n_5154),
.B(n_4658),
.Y(n_5360)
);

INVx1_ASAP7_75t_L g5361 ( 
.A(n_4864),
.Y(n_5361)
);

INVx1_ASAP7_75t_L g5362 ( 
.A(n_4864),
.Y(n_5362)
);

AND2x2_ASAP7_75t_L g5363 ( 
.A(n_4852),
.B(n_4427),
.Y(n_5363)
);

AND2x2_ASAP7_75t_L g5364 ( 
.A(n_4890),
.B(n_4428),
.Y(n_5364)
);

AOI21x1_ASAP7_75t_L g5365 ( 
.A1(n_4938),
.A2(n_4382),
.B(n_4368),
.Y(n_5365)
);

OR2x2_ASAP7_75t_L g5366 ( 
.A(n_4981),
.B(n_4985),
.Y(n_5366)
);

AND2x2_ASAP7_75t_L g5367 ( 
.A(n_4890),
.B(n_4428),
.Y(n_5367)
);

NAND2xp5_ASAP7_75t_L g5368 ( 
.A(n_5174),
.B(n_4659),
.Y(n_5368)
);

AO21x2_ASAP7_75t_L g5369 ( 
.A1(n_4742),
.A2(n_4367),
.B(n_4677),
.Y(n_5369)
);

INVx2_ASAP7_75t_L g5370 ( 
.A(n_5128),
.Y(n_5370)
);

AND2x4_ASAP7_75t_L g5371 ( 
.A(n_5022),
.B(n_4348),
.Y(n_5371)
);

AND2x2_ASAP7_75t_L g5372 ( 
.A(n_4890),
.B(n_4435),
.Y(n_5372)
);

NAND2xp5_ASAP7_75t_L g5373 ( 
.A(n_4772),
.B(n_4659),
.Y(n_5373)
);

AOI22xp33_ASAP7_75t_SL g5374 ( 
.A1(n_5180),
.A2(n_4474),
.B1(n_4359),
.B2(n_4383),
.Y(n_5374)
);

OA21x2_ASAP7_75t_L g5375 ( 
.A1(n_5011),
.A2(n_4750),
.B(n_4742),
.Y(n_5375)
);

BUFx2_ASAP7_75t_L g5376 ( 
.A(n_4871),
.Y(n_5376)
);

AND2x2_ASAP7_75t_L g5377 ( 
.A(n_4890),
.B(n_4435),
.Y(n_5377)
);

AO21x2_ASAP7_75t_L g5378 ( 
.A1(n_4750),
.A2(n_4677),
.B(n_4667),
.Y(n_5378)
);

HB1xp67_ASAP7_75t_L g5379 ( 
.A(n_4771),
.Y(n_5379)
);

INVx1_ASAP7_75t_L g5380 ( 
.A(n_4866),
.Y(n_5380)
);

INVx2_ASAP7_75t_L g5381 ( 
.A(n_5128),
.Y(n_5381)
);

INVx1_ASAP7_75t_L g5382 ( 
.A(n_4866),
.Y(n_5382)
);

INVx2_ASAP7_75t_L g5383 ( 
.A(n_5128),
.Y(n_5383)
);

INVx2_ASAP7_75t_L g5384 ( 
.A(n_5128),
.Y(n_5384)
);

INVx1_ASAP7_75t_L g5385 ( 
.A(n_4867),
.Y(n_5385)
);

INVx1_ASAP7_75t_L g5386 ( 
.A(n_4867),
.Y(n_5386)
);

AOI21xp33_ASAP7_75t_SL g5387 ( 
.A1(n_4715),
.A2(n_4208),
.B(n_4520),
.Y(n_5387)
);

AO21x2_ASAP7_75t_L g5388 ( 
.A1(n_4779),
.A2(n_4667),
.B(n_4216),
.Y(n_5388)
);

INVx1_ASAP7_75t_L g5389 ( 
.A(n_4872),
.Y(n_5389)
);

INVx1_ASAP7_75t_L g5390 ( 
.A(n_4872),
.Y(n_5390)
);

OAI21xp5_ASAP7_75t_L g5391 ( 
.A1(n_4997),
.A2(n_4269),
.B(n_4418),
.Y(n_5391)
);

HB1xp67_ASAP7_75t_L g5392 ( 
.A(n_4911),
.Y(n_5392)
);

AO31x2_ASAP7_75t_L g5393 ( 
.A1(n_5102),
.A2(n_4477),
.A3(n_4508),
.B(n_4503),
.Y(n_5393)
);

INVx2_ASAP7_75t_L g5394 ( 
.A(n_4880),
.Y(n_5394)
);

AOI21xp5_ASAP7_75t_SL g5395 ( 
.A1(n_4988),
.A2(n_4691),
.B(n_4373),
.Y(n_5395)
);

INVx1_ASAP7_75t_L g5396 ( 
.A(n_4908),
.Y(n_5396)
);

OAI21xp5_ASAP7_75t_L g5397 ( 
.A1(n_5039),
.A2(n_4604),
.B(n_4229),
.Y(n_5397)
);

OR2x2_ASAP7_75t_L g5398 ( 
.A(n_4949),
.B(n_4247),
.Y(n_5398)
);

BUFx12f_ASAP7_75t_L g5399 ( 
.A(n_4732),
.Y(n_5399)
);

HB1xp67_ASAP7_75t_L g5400 ( 
.A(n_4778),
.Y(n_5400)
);

OAI21xp5_ASAP7_75t_L g5401 ( 
.A1(n_4827),
.A2(n_4229),
.B(n_4584),
.Y(n_5401)
);

AND2x4_ASAP7_75t_L g5402 ( 
.A(n_5022),
.B(n_4348),
.Y(n_5402)
);

AND2x2_ASAP7_75t_L g5403 ( 
.A(n_4977),
.B(n_4436),
.Y(n_5403)
);

AO21x2_ASAP7_75t_L g5404 ( 
.A1(n_4779),
.A2(n_4419),
.B(n_4410),
.Y(n_5404)
);

INVx1_ASAP7_75t_L g5405 ( 
.A(n_4908),
.Y(n_5405)
);

INVx1_ASAP7_75t_L g5406 ( 
.A(n_4924),
.Y(n_5406)
);

INVx2_ASAP7_75t_L g5407 ( 
.A(n_4880),
.Y(n_5407)
);

AOI221xp5_ASAP7_75t_L g5408 ( 
.A1(n_5066),
.A2(n_4572),
.B1(n_4589),
.B2(n_4595),
.C(n_4267),
.Y(n_5408)
);

INVx1_ASAP7_75t_L g5409 ( 
.A(n_4924),
.Y(n_5409)
);

INVx3_ASAP7_75t_L g5410 ( 
.A(n_5136),
.Y(n_5410)
);

INVx1_ASAP7_75t_L g5411 ( 
.A(n_4929),
.Y(n_5411)
);

AND2x2_ASAP7_75t_L g5412 ( 
.A(n_4977),
.B(n_4436),
.Y(n_5412)
);

AO21x2_ASAP7_75t_L g5413 ( 
.A1(n_4779),
.A2(n_4478),
.B(n_4419),
.Y(n_5413)
);

INVx2_ASAP7_75t_L g5414 ( 
.A(n_4880),
.Y(n_5414)
);

INVx2_ASAP7_75t_L g5415 ( 
.A(n_4880),
.Y(n_5415)
);

OA21x2_ASAP7_75t_L g5416 ( 
.A1(n_4795),
.A2(n_4536),
.B(n_4478),
.Y(n_5416)
);

INVx1_ASAP7_75t_L g5417 ( 
.A(n_4929),
.Y(n_5417)
);

AOI211xp5_ASAP7_75t_SL g5418 ( 
.A1(n_4762),
.A2(n_4524),
.B(n_4520),
.C(n_4508),
.Y(n_5418)
);

INVx1_ASAP7_75t_L g5419 ( 
.A(n_4953),
.Y(n_5419)
);

OR2x2_ASAP7_75t_L g5420 ( 
.A(n_4949),
.B(n_4431),
.Y(n_5420)
);

OAI221xp5_ASAP7_75t_L g5421 ( 
.A1(n_5066),
.A2(n_4474),
.B1(n_4438),
.B2(n_4208),
.C(n_4379),
.Y(n_5421)
);

INVx1_ASAP7_75t_L g5422 ( 
.A(n_4953),
.Y(n_5422)
);

AND2x2_ASAP7_75t_L g5423 ( 
.A(n_4977),
.B(n_4459),
.Y(n_5423)
);

NAND2xp5_ASAP7_75t_L g5424 ( 
.A(n_4780),
.B(n_4663),
.Y(n_5424)
);

AND2x4_ASAP7_75t_L g5425 ( 
.A(n_5022),
.B(n_4389),
.Y(n_5425)
);

INVx1_ASAP7_75t_L g5426 ( 
.A(n_4954),
.Y(n_5426)
);

INVx2_ASAP7_75t_L g5427 ( 
.A(n_4880),
.Y(n_5427)
);

INVx1_ASAP7_75t_L g5428 ( 
.A(n_4954),
.Y(n_5428)
);

INVx1_ASAP7_75t_L g5429 ( 
.A(n_4957),
.Y(n_5429)
);

AND2x2_ASAP7_75t_L g5430 ( 
.A(n_4977),
.B(n_4459),
.Y(n_5430)
);

INVx2_ASAP7_75t_L g5431 ( 
.A(n_4880),
.Y(n_5431)
);

INVx1_ASAP7_75t_L g5432 ( 
.A(n_4957),
.Y(n_5432)
);

NOR2xp33_ASAP7_75t_L g5433 ( 
.A(n_4715),
.B(n_4447),
.Y(n_5433)
);

INVx1_ASAP7_75t_L g5434 ( 
.A(n_4960),
.Y(n_5434)
);

INVx1_ASAP7_75t_L g5435 ( 
.A(n_4960),
.Y(n_5435)
);

INVx2_ASAP7_75t_L g5436 ( 
.A(n_4893),
.Y(n_5436)
);

INVx2_ASAP7_75t_L g5437 ( 
.A(n_4893),
.Y(n_5437)
);

NOR2xp33_ASAP7_75t_L g5438 ( 
.A(n_4751),
.B(n_4447),
.Y(n_5438)
);

INVx2_ASAP7_75t_SL g5439 ( 
.A(n_5112),
.Y(n_5439)
);

OAI33xp33_ASAP7_75t_L g5440 ( 
.A1(n_4706),
.A2(n_4503),
.A3(n_4524),
.B1(n_4522),
.B2(n_4595),
.B3(n_4589),
.Y(n_5440)
);

HB1xp67_ASAP7_75t_L g5441 ( 
.A(n_4804),
.Y(n_5441)
);

INVxp67_ASAP7_75t_L g5442 ( 
.A(n_4885),
.Y(n_5442)
);

INVx1_ASAP7_75t_L g5443 ( 
.A(n_4974),
.Y(n_5443)
);

INVx2_ASAP7_75t_L g5444 ( 
.A(n_4893),
.Y(n_5444)
);

INVx2_ASAP7_75t_L g5445 ( 
.A(n_4893),
.Y(n_5445)
);

AND2x2_ASAP7_75t_L g5446 ( 
.A(n_5021),
.B(n_4463),
.Y(n_5446)
);

INVx3_ASAP7_75t_L g5447 ( 
.A(n_5136),
.Y(n_5447)
);

OAI31xp33_ASAP7_75t_L g5448 ( 
.A1(n_4827),
.A2(n_4451),
.A3(n_4345),
.B(n_4462),
.Y(n_5448)
);

OA21x2_ASAP7_75t_L g5449 ( 
.A1(n_4795),
.A2(n_4536),
.B(n_4478),
.Y(n_5449)
);

AND2x2_ASAP7_75t_L g5450 ( 
.A(n_5021),
.B(n_4463),
.Y(n_5450)
);

AND2x2_ASAP7_75t_L g5451 ( 
.A(n_5021),
.B(n_4465),
.Y(n_5451)
);

NAND2xp5_ASAP7_75t_L g5452 ( 
.A(n_5153),
.B(n_4663),
.Y(n_5452)
);

AND2x4_ASAP7_75t_L g5453 ( 
.A(n_5082),
.B(n_4389),
.Y(n_5453)
);

AO21x2_ASAP7_75t_L g5454 ( 
.A1(n_4877),
.A2(n_4485),
.B(n_4419),
.Y(n_5454)
);

OAI22xp5_ASAP7_75t_SL g5455 ( 
.A1(n_5180),
.A2(n_4680),
.B1(n_4208),
.B2(n_4229),
.Y(n_5455)
);

AND2x2_ASAP7_75t_L g5456 ( 
.A(n_5021),
.B(n_4465),
.Y(n_5456)
);

INVx1_ASAP7_75t_L g5457 ( 
.A(n_4974),
.Y(n_5457)
);

OA21x2_ASAP7_75t_L g5458 ( 
.A1(n_4976),
.A2(n_4487),
.B(n_4485),
.Y(n_5458)
);

INVx3_ASAP7_75t_L g5459 ( 
.A(n_5136),
.Y(n_5459)
);

INVx2_ASAP7_75t_SL g5460 ( 
.A(n_4869),
.Y(n_5460)
);

AOI21xp5_ASAP7_75t_SL g5461 ( 
.A1(n_5010),
.A2(n_4691),
.B(n_4208),
.Y(n_5461)
);

INVx1_ASAP7_75t_L g5462 ( 
.A(n_4980),
.Y(n_5462)
);

BUFx2_ASAP7_75t_L g5463 ( 
.A(n_4871),
.Y(n_5463)
);

AND2x2_ASAP7_75t_L g5464 ( 
.A(n_5086),
.B(n_4644),
.Y(n_5464)
);

AOI22xp33_ASAP7_75t_L g5465 ( 
.A1(n_5000),
.A2(n_4444),
.B1(n_4533),
.B2(n_4626),
.Y(n_5465)
);

INVx1_ASAP7_75t_L g5466 ( 
.A(n_4980),
.Y(n_5466)
);

HB1xp67_ASAP7_75t_L g5467 ( 
.A(n_4825),
.Y(n_5467)
);

INVx1_ASAP7_75t_L g5468 ( 
.A(n_5003),
.Y(n_5468)
);

OAI21x1_ASAP7_75t_L g5469 ( 
.A1(n_4976),
.A2(n_4196),
.B(n_4233),
.Y(n_5469)
);

INVx2_ASAP7_75t_L g5470 ( 
.A(n_4893),
.Y(n_5470)
);

AND2x4_ASAP7_75t_L g5471 ( 
.A(n_5082),
.B(n_4389),
.Y(n_5471)
);

BUFx2_ASAP7_75t_L g5472 ( 
.A(n_4923),
.Y(n_5472)
);

AO21x2_ASAP7_75t_L g5473 ( 
.A1(n_4883),
.A2(n_4487),
.B(n_4485),
.Y(n_5473)
);

NAND2xp5_ASAP7_75t_L g5474 ( 
.A(n_5166),
.B(n_4683),
.Y(n_5474)
);

INVxp67_ASAP7_75t_L g5475 ( 
.A(n_4791),
.Y(n_5475)
);

INVx2_ASAP7_75t_L g5476 ( 
.A(n_4893),
.Y(n_5476)
);

INVx1_ASAP7_75t_L g5477 ( 
.A(n_5003),
.Y(n_5477)
);

OR2x2_ASAP7_75t_L g5478 ( 
.A(n_5067),
.B(n_4261),
.Y(n_5478)
);

AO21x2_ASAP7_75t_L g5479 ( 
.A1(n_4975),
.A2(n_4519),
.B(n_4487),
.Y(n_5479)
);

AND2x2_ASAP7_75t_L g5480 ( 
.A(n_5086),
.B(n_4644),
.Y(n_5480)
);

AOI21xp5_ASAP7_75t_SL g5481 ( 
.A1(n_4735),
.A2(n_4461),
.B(n_4229),
.Y(n_5481)
);

INVx1_ASAP7_75t_L g5482 ( 
.A(n_5009),
.Y(n_5482)
);

OR2x2_ASAP7_75t_L g5483 ( 
.A(n_5067),
.B(n_5027),
.Y(n_5483)
);

AND2x2_ASAP7_75t_L g5484 ( 
.A(n_5086),
.B(n_4480),
.Y(n_5484)
);

OR2x2_ASAP7_75t_L g5485 ( 
.A(n_5045),
.B(n_4707),
.Y(n_5485)
);

INVx2_ASAP7_75t_L g5486 ( 
.A(n_4842),
.Y(n_5486)
);

INVx3_ASAP7_75t_L g5487 ( 
.A(n_5136),
.Y(n_5487)
);

NOR2xp33_ASAP7_75t_R g5488 ( 
.A(n_4719),
.B(n_4652),
.Y(n_5488)
);

INVx2_ASAP7_75t_SL g5489 ( 
.A(n_4869),
.Y(n_5489)
);

OR2x2_ASAP7_75t_L g5490 ( 
.A(n_4707),
.B(n_4261),
.Y(n_5490)
);

INVx2_ASAP7_75t_SL g5491 ( 
.A(n_4869),
.Y(n_5491)
);

INVx1_ASAP7_75t_L g5492 ( 
.A(n_5009),
.Y(n_5492)
);

INVx1_ASAP7_75t_L g5493 ( 
.A(n_5043),
.Y(n_5493)
);

INVx1_ASAP7_75t_L g5494 ( 
.A(n_5043),
.Y(n_5494)
);

HB1xp67_ASAP7_75t_L g5495 ( 
.A(n_4835),
.Y(n_5495)
);

OR2x2_ASAP7_75t_L g5496 ( 
.A(n_4709),
.B(n_4331),
.Y(n_5496)
);

OR2x6_ASAP7_75t_L g5497 ( 
.A(n_5194),
.B(n_4735),
.Y(n_5497)
);

OR2x2_ASAP7_75t_L g5498 ( 
.A(n_4709),
.B(n_4331),
.Y(n_5498)
);

INVx2_ASAP7_75t_L g5499 ( 
.A(n_4842),
.Y(n_5499)
);

INVx2_ASAP7_75t_L g5500 ( 
.A(n_4842),
.Y(n_5500)
);

INVx1_ASAP7_75t_L g5501 ( 
.A(n_5051),
.Y(n_5501)
);

OR2x2_ASAP7_75t_L g5502 ( 
.A(n_4713),
.B(n_4376),
.Y(n_5502)
);

AOI21xp5_ASAP7_75t_L g5503 ( 
.A1(n_4735),
.A2(n_4584),
.B(n_4642),
.Y(n_5503)
);

INVx1_ASAP7_75t_L g5504 ( 
.A(n_5051),
.Y(n_5504)
);

INVx2_ASAP7_75t_L g5505 ( 
.A(n_4842),
.Y(n_5505)
);

OAI21xp5_ASAP7_75t_L g5506 ( 
.A1(n_5133),
.A2(n_4557),
.B(n_4542),
.Y(n_5506)
);

BUFx2_ASAP7_75t_L g5507 ( 
.A(n_4923),
.Y(n_5507)
);

INVx1_ASAP7_75t_L g5508 ( 
.A(n_5056),
.Y(n_5508)
);

AO21x2_ASAP7_75t_L g5509 ( 
.A1(n_4781),
.A2(n_4525),
.B(n_4519),
.Y(n_5509)
);

INVx1_ASAP7_75t_L g5510 ( 
.A(n_5056),
.Y(n_5510)
);

AND2x4_ASAP7_75t_L g5511 ( 
.A(n_5082),
.B(n_4389),
.Y(n_5511)
);

HB1xp67_ASAP7_75t_L g5512 ( 
.A(n_4847),
.Y(n_5512)
);

AOI21xp5_ASAP7_75t_SL g5513 ( 
.A1(n_4735),
.A2(n_4732),
.B(n_4736),
.Y(n_5513)
);

INVx2_ASAP7_75t_L g5514 ( 
.A(n_4842),
.Y(n_5514)
);

INVx1_ASAP7_75t_L g5515 ( 
.A(n_5060),
.Y(n_5515)
);

AOI22xp33_ASAP7_75t_L g5516 ( 
.A1(n_5000),
.A2(n_5193),
.B1(n_4712),
.B2(n_4722),
.Y(n_5516)
);

AND2x2_ASAP7_75t_L g5517 ( 
.A(n_5086),
.B(n_4480),
.Y(n_5517)
);

INVx1_ASAP7_75t_L g5518 ( 
.A(n_5060),
.Y(n_5518)
);

INVx1_ASAP7_75t_L g5519 ( 
.A(n_5062),
.Y(n_5519)
);

AND2x2_ASAP7_75t_L g5520 ( 
.A(n_5178),
.B(n_4734),
.Y(n_5520)
);

INVx2_ASAP7_75t_L g5521 ( 
.A(n_4842),
.Y(n_5521)
);

OAI21xp5_ASAP7_75t_L g5522 ( 
.A1(n_5071),
.A2(n_4731),
.B(n_4704),
.Y(n_5522)
);

OR2x6_ASAP7_75t_L g5523 ( 
.A(n_4735),
.B(n_4429),
.Y(n_5523)
);

INVx1_ASAP7_75t_L g5524 ( 
.A(n_5062),
.Y(n_5524)
);

INVx3_ASAP7_75t_L g5525 ( 
.A(n_5070),
.Y(n_5525)
);

OAI321xp33_ASAP7_75t_L g5526 ( 
.A1(n_4836),
.A2(n_4616),
.A3(n_4633),
.B1(n_4462),
.B2(n_4501),
.C(n_4452),
.Y(n_5526)
);

INVx2_ASAP7_75t_L g5527 ( 
.A(n_4905),
.Y(n_5527)
);

INVx1_ASAP7_75t_L g5528 ( 
.A(n_5097),
.Y(n_5528)
);

OR2x6_ASAP7_75t_L g5529 ( 
.A(n_5096),
.B(n_4434),
.Y(n_5529)
);

OA21x2_ASAP7_75t_L g5530 ( 
.A1(n_4972),
.A2(n_4525),
.B(n_4519),
.Y(n_5530)
);

INVx2_ASAP7_75t_L g5531 ( 
.A(n_4905),
.Y(n_5531)
);

AO21x2_ASAP7_75t_L g5532 ( 
.A1(n_4781),
.A2(n_4538),
.B(n_4525),
.Y(n_5532)
);

BUFx2_ASAP7_75t_L g5533 ( 
.A(n_4932),
.Y(n_5533)
);

AO21x2_ASAP7_75t_L g5534 ( 
.A1(n_4781),
.A2(n_4548),
.B(n_4538),
.Y(n_5534)
);

AND2x2_ASAP7_75t_L g5535 ( 
.A(n_5178),
.B(n_4494),
.Y(n_5535)
);

HB1xp67_ASAP7_75t_L g5536 ( 
.A(n_4882),
.Y(n_5536)
);

HB1xp67_ASAP7_75t_L g5537 ( 
.A(n_4838),
.Y(n_5537)
);

INVx2_ASAP7_75t_L g5538 ( 
.A(n_4905),
.Y(n_5538)
);

OA21x2_ASAP7_75t_L g5539 ( 
.A1(n_4787),
.A2(n_4807),
.B(n_4799),
.Y(n_5539)
);

INVxp67_ASAP7_75t_SL g5540 ( 
.A(n_4850),
.Y(n_5540)
);

INVx3_ASAP7_75t_L g5541 ( 
.A(n_5070),
.Y(n_5541)
);

OA21x2_ASAP7_75t_L g5542 ( 
.A1(n_4787),
.A2(n_4807),
.B(n_4799),
.Y(n_5542)
);

INVx2_ASAP7_75t_SL g5543 ( 
.A(n_4869),
.Y(n_5543)
);

INVx2_ASAP7_75t_L g5544 ( 
.A(n_4905),
.Y(n_5544)
);

INVx2_ASAP7_75t_L g5545 ( 
.A(n_4905),
.Y(n_5545)
);

AND2x2_ASAP7_75t_L g5546 ( 
.A(n_4734),
.B(n_4494),
.Y(n_5546)
);

INVx2_ASAP7_75t_L g5547 ( 
.A(n_4905),
.Y(n_5547)
);

OAI22xp5_ASAP7_75t_SL g5548 ( 
.A1(n_5193),
.A2(n_4680),
.B1(n_4461),
.B2(n_4529),
.Y(n_5548)
);

INVx1_ASAP7_75t_L g5549 ( 
.A(n_5097),
.Y(n_5549)
);

INVx1_ASAP7_75t_L g5550 ( 
.A(n_5116),
.Y(n_5550)
);

OA21x2_ASAP7_75t_L g5551 ( 
.A1(n_4787),
.A2(n_4548),
.B(n_4538),
.Y(n_5551)
);

AO21x2_ASAP7_75t_L g5552 ( 
.A1(n_4799),
.A2(n_4603),
.B(n_4548),
.Y(n_5552)
);

INVx3_ASAP7_75t_L g5553 ( 
.A(n_5070),
.Y(n_5553)
);

INVx1_ASAP7_75t_L g5554 ( 
.A(n_5116),
.Y(n_5554)
);

AND2x4_ASAP7_75t_L g5555 ( 
.A(n_5082),
.B(n_4399),
.Y(n_5555)
);

HB1xp67_ASAP7_75t_L g5556 ( 
.A(n_5029),
.Y(n_5556)
);

BUFx3_ASAP7_75t_L g5557 ( 
.A(n_4756),
.Y(n_5557)
);

INVx1_ASAP7_75t_L g5558 ( 
.A(n_5135),
.Y(n_5558)
);

INVx2_ASAP7_75t_L g5559 ( 
.A(n_4848),
.Y(n_5559)
);

NAND2x1_ASAP7_75t_L g5560 ( 
.A(n_4790),
.B(n_4434),
.Y(n_5560)
);

AND2x2_ASAP7_75t_L g5561 ( 
.A(n_4749),
.B(n_4497),
.Y(n_5561)
);

INVx1_ASAP7_75t_L g5562 ( 
.A(n_5135),
.Y(n_5562)
);

OA21x2_ASAP7_75t_L g5563 ( 
.A1(n_4807),
.A2(n_4627),
.B(n_4603),
.Y(n_5563)
);

AND2x2_ASAP7_75t_L g5564 ( 
.A(n_4749),
.B(n_4497),
.Y(n_5564)
);

INVx2_ASAP7_75t_L g5565 ( 
.A(n_4848),
.Y(n_5565)
);

AND2x2_ASAP7_75t_L g5566 ( 
.A(n_4777),
.B(n_4509),
.Y(n_5566)
);

AOI21xp33_ASAP7_75t_L g5567 ( 
.A1(n_4939),
.A2(n_4417),
.B(n_4438),
.Y(n_5567)
);

CKINVDCx20_ASAP7_75t_R g5568 ( 
.A(n_4746),
.Y(n_5568)
);

INVx1_ASAP7_75t_L g5569 ( 
.A(n_5141),
.Y(n_5569)
);

INVx1_ASAP7_75t_L g5570 ( 
.A(n_5141),
.Y(n_5570)
);

INVx1_ASAP7_75t_L g5571 ( 
.A(n_5144),
.Y(n_5571)
);

AND2x4_ASAP7_75t_L g5572 ( 
.A(n_5082),
.B(n_4399),
.Y(n_5572)
);

OAI221xp5_ASAP7_75t_SL g5573 ( 
.A1(n_5184),
.A2(n_4501),
.B1(n_4585),
.B2(n_4557),
.C(n_4542),
.Y(n_5573)
);

OR2x2_ASAP7_75t_L g5574 ( 
.A(n_4713),
.B(n_4714),
.Y(n_5574)
);

BUFx2_ASAP7_75t_L g5575 ( 
.A(n_4932),
.Y(n_5575)
);

INVx2_ASAP7_75t_L g5576 ( 
.A(n_4848),
.Y(n_5576)
);

AND2x4_ASAP7_75t_L g5577 ( 
.A(n_5019),
.B(n_4399),
.Y(n_5577)
);

BUFx2_ASAP7_75t_L g5578 ( 
.A(n_4791),
.Y(n_5578)
);

HB1xp67_ASAP7_75t_L g5579 ( 
.A(n_5157),
.Y(n_5579)
);

INVx1_ASAP7_75t_L g5580 ( 
.A(n_5144),
.Y(n_5580)
);

BUFx2_ASAP7_75t_L g5581 ( 
.A(n_4791),
.Y(n_5581)
);

INVx2_ASAP7_75t_L g5582 ( 
.A(n_5190),
.Y(n_5582)
);

AOI21xp5_ASAP7_75t_SL g5583 ( 
.A1(n_4736),
.A2(n_4461),
.B(n_4474),
.Y(n_5583)
);

INVx2_ASAP7_75t_L g5584 ( 
.A(n_5190),
.Y(n_5584)
);

AO21x2_ASAP7_75t_L g5585 ( 
.A1(n_4844),
.A2(n_4627),
.B(n_4603),
.Y(n_5585)
);

INVx3_ASAP7_75t_L g5586 ( 
.A(n_5070),
.Y(n_5586)
);

OR2x2_ASAP7_75t_L g5587 ( 
.A(n_4714),
.B(n_4376),
.Y(n_5587)
);

INVx2_ASAP7_75t_L g5588 ( 
.A(n_5190),
.Y(n_5588)
);

HB1xp67_ASAP7_75t_L g5589 ( 
.A(n_4951),
.Y(n_5589)
);

NAND2xp5_ASAP7_75t_L g5590 ( 
.A(n_4914),
.B(n_4683),
.Y(n_5590)
);

HB1xp67_ASAP7_75t_L g5591 ( 
.A(n_4992),
.Y(n_5591)
);

BUFx3_ASAP7_75t_L g5592 ( 
.A(n_4725),
.Y(n_5592)
);

BUFx3_ASAP7_75t_L g5593 ( 
.A(n_5001),
.Y(n_5593)
);

AND2x2_ASAP7_75t_L g5594 ( 
.A(n_4777),
.B(n_4509),
.Y(n_5594)
);

OA21x2_ASAP7_75t_L g5595 ( 
.A1(n_4844),
.A2(n_4666),
.B(n_4627),
.Y(n_5595)
);

INVx2_ASAP7_75t_L g5596 ( 
.A(n_5190),
.Y(n_5596)
);

INVx2_ASAP7_75t_L g5597 ( 
.A(n_5190),
.Y(n_5597)
);

AO21x2_ASAP7_75t_L g5598 ( 
.A1(n_4844),
.A2(n_4666),
.B(n_4628),
.Y(n_5598)
);

INVx1_ASAP7_75t_L g5599 ( 
.A(n_5150),
.Y(n_5599)
);

INVx2_ASAP7_75t_L g5600 ( 
.A(n_5195),
.Y(n_5600)
);

AND2x2_ASAP7_75t_L g5601 ( 
.A(n_5340),
.B(n_5282),
.Y(n_5601)
);

OR2x2_ASAP7_75t_L g5602 ( 
.A(n_5268),
.B(n_4711),
.Y(n_5602)
);

HB1xp67_ASAP7_75t_L g5603 ( 
.A(n_5324),
.Y(n_5603)
);

AND2x4_ASAP7_75t_L g5604 ( 
.A(n_5340),
.B(n_4797),
.Y(n_5604)
);

AND2x2_ASAP7_75t_L g5605 ( 
.A(n_5340),
.B(n_4797),
.Y(n_5605)
);

OR2x2_ASAP7_75t_L g5606 ( 
.A(n_5268),
.B(n_4711),
.Y(n_5606)
);

BUFx3_ASAP7_75t_L g5607 ( 
.A(n_5593),
.Y(n_5607)
);

AOI22xp33_ASAP7_75t_L g5608 ( 
.A1(n_5355),
.A2(n_5000),
.B1(n_4744),
.B2(n_4444),
.Y(n_5608)
);

AND2x2_ASAP7_75t_L g5609 ( 
.A(n_5282),
.B(n_4797),
.Y(n_5609)
);

BUFx3_ASAP7_75t_L g5610 ( 
.A(n_5593),
.Y(n_5610)
);

INVx2_ASAP7_75t_L g5611 ( 
.A(n_5195),
.Y(n_5611)
);

INVx1_ASAP7_75t_L g5612 ( 
.A(n_5200),
.Y(n_5612)
);

OAI22xp5_ASAP7_75t_L g5613 ( 
.A1(n_5210),
.A2(n_4922),
.B1(n_4770),
.B2(n_4855),
.Y(n_5613)
);

AND2x2_ASAP7_75t_L g5614 ( 
.A(n_5262),
.B(n_4999),
.Y(n_5614)
);

AOI222xp33_ASAP7_75t_L g5615 ( 
.A1(n_5201),
.A2(n_5184),
.B1(n_4775),
.B2(n_4819),
.C1(n_4810),
.C2(n_4816),
.Y(n_5615)
);

HB1xp67_ASAP7_75t_L g5616 ( 
.A(n_5324),
.Y(n_5616)
);

AND2x4_ASAP7_75t_L g5617 ( 
.A(n_5344),
.B(n_4733),
.Y(n_5617)
);

AND2x2_ASAP7_75t_L g5618 ( 
.A(n_5262),
.B(n_4999),
.Y(n_5618)
);

AND2x4_ASAP7_75t_L g5619 ( 
.A(n_5344),
.B(n_4733),
.Y(n_5619)
);

INVx1_ASAP7_75t_L g5620 ( 
.A(n_5200),
.Y(n_5620)
);

OAI221xp5_ASAP7_75t_SL g5621 ( 
.A1(n_5325),
.A2(n_4941),
.B1(n_4926),
.B2(n_4922),
.C(n_5077),
.Y(n_5621)
);

OR2x2_ASAP7_75t_L g5622 ( 
.A(n_5321),
.B(n_4863),
.Y(n_5622)
);

AND2x2_ASAP7_75t_L g5623 ( 
.A(n_5305),
.B(n_4999),
.Y(n_5623)
);

INVx2_ASAP7_75t_L g5624 ( 
.A(n_5195),
.Y(n_5624)
);

OAI22xp5_ASAP7_75t_L g5625 ( 
.A1(n_5210),
.A2(n_4874),
.B1(n_4965),
.B2(n_4774),
.Y(n_5625)
);

INVx1_ASAP7_75t_L g5626 ( 
.A(n_5400),
.Y(n_5626)
);

AND2x4_ASAP7_75t_L g5627 ( 
.A(n_5344),
.B(n_4733),
.Y(n_5627)
);

AND2x2_ASAP7_75t_L g5628 ( 
.A(n_5305),
.B(n_5326),
.Y(n_5628)
);

HB1xp67_ASAP7_75t_L g5629 ( 
.A(n_5392),
.Y(n_5629)
);

INVx1_ASAP7_75t_L g5630 ( 
.A(n_5441),
.Y(n_5630)
);

INVx1_ASAP7_75t_L g5631 ( 
.A(n_5216),
.Y(n_5631)
);

AND2x2_ASAP7_75t_L g5632 ( 
.A(n_5305),
.B(n_4999),
.Y(n_5632)
);

BUFx3_ASAP7_75t_L g5633 ( 
.A(n_5593),
.Y(n_5633)
);

AND2x2_ASAP7_75t_L g5634 ( 
.A(n_5305),
.B(n_5013),
.Y(n_5634)
);

NAND2xp5_ASAP7_75t_L g5635 ( 
.A(n_5213),
.B(n_5040),
.Y(n_5635)
);

INVx1_ASAP7_75t_L g5636 ( 
.A(n_5216),
.Y(n_5636)
);

AND2x2_ASAP7_75t_L g5637 ( 
.A(n_5305),
.B(n_5013),
.Y(n_5637)
);

INVx2_ASAP7_75t_L g5638 ( 
.A(n_5196),
.Y(n_5638)
);

OR2x2_ASAP7_75t_L g5639 ( 
.A(n_5321),
.B(n_4863),
.Y(n_5639)
);

NAND2xp5_ASAP7_75t_L g5640 ( 
.A(n_5213),
.B(n_5123),
.Y(n_5640)
);

OR2x6_ASAP7_75t_L g5641 ( 
.A(n_5207),
.B(n_4759),
.Y(n_5641)
);

INVx1_ASAP7_75t_L g5642 ( 
.A(n_5219),
.Y(n_5642)
);

HB1xp67_ASAP7_75t_L g5643 ( 
.A(n_5537),
.Y(n_5643)
);

AND2x2_ASAP7_75t_L g5644 ( 
.A(n_5326),
.B(n_5013),
.Y(n_5644)
);

INVx1_ASAP7_75t_L g5645 ( 
.A(n_5219),
.Y(n_5645)
);

OR2x2_ASAP7_75t_L g5646 ( 
.A(n_5337),
.B(n_4863),
.Y(n_5646)
);

OR2x2_ASAP7_75t_L g5647 ( 
.A(n_5337),
.B(n_4863),
.Y(n_5647)
);

CKINVDCx14_ASAP7_75t_R g5648 ( 
.A(n_5568),
.Y(n_5648)
);

NAND2xp5_ASAP7_75t_L g5649 ( 
.A(n_5322),
.B(n_5085),
.Y(n_5649)
);

INVx5_ASAP7_75t_L g5650 ( 
.A(n_5220),
.Y(n_5650)
);

INVx3_ASAP7_75t_SL g5651 ( 
.A(n_5226),
.Y(n_5651)
);

INVx3_ASAP7_75t_L g5652 ( 
.A(n_5346),
.Y(n_5652)
);

INVx2_ASAP7_75t_L g5653 ( 
.A(n_5196),
.Y(n_5653)
);

HB1xp67_ASAP7_75t_L g5654 ( 
.A(n_5218),
.Y(n_5654)
);

AND2x2_ASAP7_75t_L g5655 ( 
.A(n_5326),
.B(n_4738),
.Y(n_5655)
);

AND2x2_ASAP7_75t_L g5656 ( 
.A(n_5326),
.B(n_4738),
.Y(n_5656)
);

INVx2_ASAP7_75t_L g5657 ( 
.A(n_5196),
.Y(n_5657)
);

INVx1_ASAP7_75t_L g5658 ( 
.A(n_5228),
.Y(n_5658)
);

OAI222xp33_ASAP7_75t_L g5659 ( 
.A1(n_5421),
.A2(n_4955),
.B1(n_4933),
.B2(n_4469),
.C1(n_4580),
.C2(n_5108),
.Y(n_5659)
);

NOR2xp33_ASAP7_75t_L g5660 ( 
.A(n_5226),
.B(n_4788),
.Y(n_5660)
);

OR2x2_ASAP7_75t_L g5661 ( 
.A(n_5224),
.B(n_4863),
.Y(n_5661)
);

INVx1_ASAP7_75t_L g5662 ( 
.A(n_5228),
.Y(n_5662)
);

BUFx2_ASAP7_75t_L g5663 ( 
.A(n_5327),
.Y(n_5663)
);

AND2x4_ASAP7_75t_L g5664 ( 
.A(n_5344),
.B(n_4738),
.Y(n_5664)
);

NAND2xp5_ASAP7_75t_L g5665 ( 
.A(n_5540),
.B(n_4919),
.Y(n_5665)
);

BUFx2_ASAP7_75t_L g5666 ( 
.A(n_5327),
.Y(n_5666)
);

AND2x2_ASAP7_75t_L g5667 ( 
.A(n_5326),
.B(n_5008),
.Y(n_5667)
);

OR2x6_ASAP7_75t_L g5668 ( 
.A(n_5207),
.B(n_4759),
.Y(n_5668)
);

INVx2_ASAP7_75t_L g5669 ( 
.A(n_5202),
.Y(n_5669)
);

NAND2xp33_ASAP7_75t_L g5670 ( 
.A(n_5220),
.B(n_4817),
.Y(n_5670)
);

INVx2_ASAP7_75t_L g5671 ( 
.A(n_5202),
.Y(n_5671)
);

INVx1_ASAP7_75t_L g5672 ( 
.A(n_5234),
.Y(n_5672)
);

INVx1_ASAP7_75t_L g5673 ( 
.A(n_5234),
.Y(n_5673)
);

INVx2_ASAP7_75t_SL g5674 ( 
.A(n_5220),
.Y(n_5674)
);

AND2x2_ASAP7_75t_L g5675 ( 
.A(n_5265),
.B(n_5008),
.Y(n_5675)
);

INVx1_ASAP7_75t_L g5676 ( 
.A(n_5240),
.Y(n_5676)
);

INVx1_ASAP7_75t_L g5677 ( 
.A(n_5240),
.Y(n_5677)
);

AND2x2_ASAP7_75t_L g5678 ( 
.A(n_5265),
.B(n_5012),
.Y(n_5678)
);

OR2x2_ASAP7_75t_L g5679 ( 
.A(n_5224),
.B(n_4863),
.Y(n_5679)
);

AOI22xp33_ASAP7_75t_L g5680 ( 
.A1(n_5355),
.A2(n_4533),
.B1(n_4668),
.B2(n_4626),
.Y(n_5680)
);

NAND2xp5_ASAP7_75t_L g5681 ( 
.A(n_5339),
.B(n_5379),
.Y(n_5681)
);

AOI22xp33_ASAP7_75t_L g5682 ( 
.A1(n_5355),
.A2(n_4533),
.B1(n_4668),
.B2(n_4626),
.Y(n_5682)
);

INVx2_ASAP7_75t_L g5683 ( 
.A(n_5202),
.Y(n_5683)
);

NAND2xp5_ASAP7_75t_L g5684 ( 
.A(n_5259),
.B(n_5295),
.Y(n_5684)
);

OR2x2_ASAP7_75t_L g5685 ( 
.A(n_5232),
.B(n_5189),
.Y(n_5685)
);

NAND2xp5_ASAP7_75t_L g5686 ( 
.A(n_5467),
.B(n_5031),
.Y(n_5686)
);

INVx1_ASAP7_75t_L g5687 ( 
.A(n_5247),
.Y(n_5687)
);

INVx5_ASAP7_75t_L g5688 ( 
.A(n_5220),
.Y(n_5688)
);

OR2x2_ASAP7_75t_L g5689 ( 
.A(n_5232),
.B(n_5192),
.Y(n_5689)
);

INVx1_ASAP7_75t_L g5690 ( 
.A(n_5247),
.Y(n_5690)
);

AND2x4_ASAP7_75t_L g5691 ( 
.A(n_5344),
.B(n_5019),
.Y(n_5691)
);

INVx1_ASAP7_75t_L g5692 ( 
.A(n_5248),
.Y(n_5692)
);

INVx1_ASAP7_75t_L g5693 ( 
.A(n_5248),
.Y(n_5693)
);

HB1xp67_ASAP7_75t_L g5694 ( 
.A(n_5495),
.Y(n_5694)
);

NAND2xp5_ASAP7_75t_L g5695 ( 
.A(n_5512),
.B(n_4989),
.Y(n_5695)
);

AND2x2_ASAP7_75t_L g5696 ( 
.A(n_5341),
.B(n_5012),
.Y(n_5696)
);

BUFx2_ASAP7_75t_L g5697 ( 
.A(n_5229),
.Y(n_5697)
);

OAI22xp5_ASAP7_75t_L g5698 ( 
.A1(n_5325),
.A2(n_4796),
.B1(n_4916),
.B2(n_4913),
.Y(n_5698)
);

OAI22xp5_ASAP7_75t_L g5699 ( 
.A1(n_5455),
.A2(n_4916),
.B1(n_4940),
.B2(n_4913),
.Y(n_5699)
);

INVx1_ASAP7_75t_L g5700 ( 
.A(n_5250),
.Y(n_5700)
);

AND2x2_ASAP7_75t_L g5701 ( 
.A(n_5341),
.B(n_5012),
.Y(n_5701)
);

NAND2xp5_ASAP7_75t_L g5702 ( 
.A(n_5536),
.B(n_4940),
.Y(n_5702)
);

INVx2_ASAP7_75t_L g5703 ( 
.A(n_5203),
.Y(n_5703)
);

AND2x4_ASAP7_75t_L g5704 ( 
.A(n_5555),
.B(n_5019),
.Y(n_5704)
);

INVx2_ASAP7_75t_L g5705 ( 
.A(n_5203),
.Y(n_5705)
);

INVxp67_ASAP7_75t_L g5706 ( 
.A(n_5229),
.Y(n_5706)
);

OR2x2_ASAP7_75t_L g5707 ( 
.A(n_5483),
.B(n_5079),
.Y(n_5707)
);

INVx1_ASAP7_75t_L g5708 ( 
.A(n_5250),
.Y(n_5708)
);

INVx1_ASAP7_75t_L g5709 ( 
.A(n_5256),
.Y(n_5709)
);

INVx2_ASAP7_75t_L g5710 ( 
.A(n_5203),
.Y(n_5710)
);

AND2x2_ASAP7_75t_L g5711 ( 
.A(n_5300),
.B(n_5012),
.Y(n_5711)
);

AOI22xp33_ASAP7_75t_L g5712 ( 
.A1(n_5355),
.A2(n_4626),
.B1(n_4668),
.B2(n_4496),
.Y(n_5712)
);

INVx1_ASAP7_75t_L g5713 ( 
.A(n_5256),
.Y(n_5713)
);

AND2x2_ASAP7_75t_L g5714 ( 
.A(n_5300),
.B(n_5012),
.Y(n_5714)
);

INVx1_ASAP7_75t_L g5715 ( 
.A(n_5257),
.Y(n_5715)
);

INVx2_ASAP7_75t_L g5716 ( 
.A(n_5209),
.Y(n_5716)
);

AOI22xp5_ASAP7_75t_L g5717 ( 
.A1(n_5214),
.A2(n_4767),
.B1(n_4786),
.B2(n_4752),
.Y(n_5717)
);

INVx1_ASAP7_75t_L g5718 ( 
.A(n_5257),
.Y(n_5718)
);

INVx1_ASAP7_75t_L g5719 ( 
.A(n_5269),
.Y(n_5719)
);

AND2x2_ASAP7_75t_L g5720 ( 
.A(n_5285),
.B(n_5012),
.Y(n_5720)
);

INVxp67_ASAP7_75t_SL g5721 ( 
.A(n_5221),
.Y(n_5721)
);

INVx1_ASAP7_75t_L g5722 ( 
.A(n_5269),
.Y(n_5722)
);

OAI222xp33_ASAP7_75t_L g5723 ( 
.A1(n_5421),
.A2(n_5078),
.B1(n_5088),
.B2(n_4909),
.C1(n_5159),
.C2(n_4963),
.Y(n_5723)
);

NAND2xp5_ASAP7_75t_L g5724 ( 
.A(n_5589),
.B(n_4958),
.Y(n_5724)
);

OR2x2_ASAP7_75t_L g5725 ( 
.A(n_5483),
.B(n_5081),
.Y(n_5725)
);

AND2x2_ASAP7_75t_L g5726 ( 
.A(n_5285),
.B(n_4958),
.Y(n_5726)
);

NAND2xp5_ASAP7_75t_L g5727 ( 
.A(n_5591),
.B(n_5264),
.Y(n_5727)
);

AOI22xp33_ASAP7_75t_L g5728 ( 
.A1(n_5276),
.A2(n_5211),
.B1(n_5567),
.B2(n_5375),
.Y(n_5728)
);

NAND2xp5_ASAP7_75t_L g5729 ( 
.A(n_5579),
.B(n_4967),
.Y(n_5729)
);

HB1xp67_ASAP7_75t_L g5730 ( 
.A(n_5475),
.Y(n_5730)
);

INVx1_ASAP7_75t_L g5731 ( 
.A(n_5278),
.Y(n_5731)
);

INVx1_ASAP7_75t_L g5732 ( 
.A(n_5278),
.Y(n_5732)
);

BUFx3_ASAP7_75t_L g5733 ( 
.A(n_5229),
.Y(n_5733)
);

INVx1_ASAP7_75t_L g5734 ( 
.A(n_5283),
.Y(n_5734)
);

INVxp67_ASAP7_75t_L g5735 ( 
.A(n_5312),
.Y(n_5735)
);

NAND2xp5_ASAP7_75t_L g5736 ( 
.A(n_5578),
.B(n_4967),
.Y(n_5736)
);

INVx3_ASAP7_75t_L g5737 ( 
.A(n_5346),
.Y(n_5737)
);

AND2x2_ASAP7_75t_L g5738 ( 
.A(n_5288),
.B(n_4928),
.Y(n_5738)
);

NAND2xp5_ASAP7_75t_L g5739 ( 
.A(n_5578),
.B(n_5122),
.Y(n_5739)
);

OR2x2_ASAP7_75t_L g5740 ( 
.A(n_5398),
.B(n_5111),
.Y(n_5740)
);

OR2x2_ASAP7_75t_L g5741 ( 
.A(n_5398),
.B(n_5125),
.Y(n_5741)
);

INVx2_ASAP7_75t_L g5742 ( 
.A(n_5209),
.Y(n_5742)
);

INVx1_ASAP7_75t_L g5743 ( 
.A(n_5283),
.Y(n_5743)
);

AND2x2_ASAP7_75t_L g5744 ( 
.A(n_5288),
.B(n_4928),
.Y(n_5744)
);

AND2x4_ASAP7_75t_L g5745 ( 
.A(n_5555),
.B(n_5155),
.Y(n_5745)
);

INVxp67_ASAP7_75t_SL g5746 ( 
.A(n_5221),
.Y(n_5746)
);

AND2x2_ASAP7_75t_L g5747 ( 
.A(n_5246),
.B(n_4928),
.Y(n_5747)
);

BUFx6f_ASAP7_75t_L g5748 ( 
.A(n_5220),
.Y(n_5748)
);

INVx2_ASAP7_75t_SL g5749 ( 
.A(n_5220),
.Y(n_5749)
);

INVx2_ASAP7_75t_L g5750 ( 
.A(n_5209),
.Y(n_5750)
);

AND2x2_ASAP7_75t_L g5751 ( 
.A(n_5246),
.B(n_4928),
.Y(n_5751)
);

AND2x2_ASAP7_75t_L g5752 ( 
.A(n_5249),
.B(n_5054),
.Y(n_5752)
);

HB1xp67_ASAP7_75t_L g5753 ( 
.A(n_5475),
.Y(n_5753)
);

AND2x2_ASAP7_75t_L g5754 ( 
.A(n_5249),
.B(n_5054),
.Y(n_5754)
);

INVx1_ASAP7_75t_L g5755 ( 
.A(n_5292),
.Y(n_5755)
);

INVx3_ASAP7_75t_L g5756 ( 
.A(n_5346),
.Y(n_5756)
);

INVx2_ASAP7_75t_L g5757 ( 
.A(n_5212),
.Y(n_5757)
);

NAND2xp5_ASAP7_75t_L g5758 ( 
.A(n_5581),
.B(n_4759),
.Y(n_5758)
);

AND2x4_ASAP7_75t_L g5759 ( 
.A(n_5555),
.B(n_5155),
.Y(n_5759)
);

INVx1_ASAP7_75t_L g5760 ( 
.A(n_5292),
.Y(n_5760)
);

INVx1_ASAP7_75t_L g5761 ( 
.A(n_5293),
.Y(n_5761)
);

INVx1_ASAP7_75t_L g5762 ( 
.A(n_5293),
.Y(n_5762)
);

BUFx2_ASAP7_75t_L g5763 ( 
.A(n_5226),
.Y(n_5763)
);

INVx1_ASAP7_75t_L g5764 ( 
.A(n_5294),
.Y(n_5764)
);

AND2x2_ASAP7_75t_L g5765 ( 
.A(n_5464),
.B(n_5480),
.Y(n_5765)
);

OR2x2_ASAP7_75t_L g5766 ( 
.A(n_5574),
.B(n_5142),
.Y(n_5766)
);

AND2x2_ASAP7_75t_L g5767 ( 
.A(n_5464),
.B(n_5054),
.Y(n_5767)
);

AND2x2_ASAP7_75t_L g5768 ( 
.A(n_5480),
.B(n_5054),
.Y(n_5768)
);

INVx2_ASAP7_75t_L g5769 ( 
.A(n_5212),
.Y(n_5769)
);

INVx1_ASAP7_75t_L g5770 ( 
.A(n_5294),
.Y(n_5770)
);

INVx1_ASAP7_75t_L g5771 ( 
.A(n_5298),
.Y(n_5771)
);

AND2x2_ASAP7_75t_L g5772 ( 
.A(n_5235),
.B(n_5054),
.Y(n_5772)
);

INVxp67_ASAP7_75t_SL g5773 ( 
.A(n_5221),
.Y(n_5773)
);

AND2x2_ASAP7_75t_L g5774 ( 
.A(n_5235),
.B(n_5054),
.Y(n_5774)
);

NAND2xp5_ASAP7_75t_L g5775 ( 
.A(n_5581),
.B(n_5057),
.Y(n_5775)
);

INVx1_ASAP7_75t_L g5776 ( 
.A(n_5298),
.Y(n_5776)
);

AND2x2_ASAP7_75t_L g5777 ( 
.A(n_5238),
.B(n_4934),
.Y(n_5777)
);

INVx3_ASAP7_75t_L g5778 ( 
.A(n_5346),
.Y(n_5778)
);

NOR2x1_ASAP7_75t_L g5779 ( 
.A(n_5226),
.B(n_4879),
.Y(n_5779)
);

INVx1_ASAP7_75t_L g5780 ( 
.A(n_5307),
.Y(n_5780)
);

AND2x2_ASAP7_75t_L g5781 ( 
.A(n_5238),
.B(n_4934),
.Y(n_5781)
);

AOI22xp33_ASAP7_75t_L g5782 ( 
.A1(n_5211),
.A2(n_4668),
.B1(n_4496),
.B2(n_4551),
.Y(n_5782)
);

AOI222xp33_ASAP7_75t_L g5783 ( 
.A1(n_5199),
.A2(n_5167),
.B1(n_5124),
.B2(n_4828),
.C1(n_5064),
.C2(n_5173),
.Y(n_5783)
);

AND2x2_ASAP7_75t_L g5784 ( 
.A(n_5241),
.B(n_4934),
.Y(n_5784)
);

INVx1_ASAP7_75t_L g5785 ( 
.A(n_5307),
.Y(n_5785)
);

NAND2xp5_ASAP7_75t_L g5786 ( 
.A(n_5230),
.B(n_4952),
.Y(n_5786)
);

NAND2xp5_ASAP7_75t_L g5787 ( 
.A(n_5230),
.B(n_5556),
.Y(n_5787)
);

INVx1_ASAP7_75t_L g5788 ( 
.A(n_5311),
.Y(n_5788)
);

NAND2xp5_ASAP7_75t_L g5789 ( 
.A(n_5225),
.B(n_4952),
.Y(n_5789)
);

AND2x2_ASAP7_75t_L g5790 ( 
.A(n_5241),
.B(n_4952),
.Y(n_5790)
);

NAND2xp5_ASAP7_75t_L g5791 ( 
.A(n_5225),
.B(n_4993),
.Y(n_5791)
);

INVx1_ASAP7_75t_L g5792 ( 
.A(n_5311),
.Y(n_5792)
);

AND2x2_ASAP7_75t_L g5793 ( 
.A(n_5290),
.B(n_4993),
.Y(n_5793)
);

INVx2_ASAP7_75t_SL g5794 ( 
.A(n_5314),
.Y(n_5794)
);

INVx2_ASAP7_75t_L g5795 ( 
.A(n_5212),
.Y(n_5795)
);

INVx1_ASAP7_75t_L g5796 ( 
.A(n_5313),
.Y(n_5796)
);

OR2x2_ASAP7_75t_L g5797 ( 
.A(n_5574),
.B(n_5182),
.Y(n_5797)
);

HB1xp67_ASAP7_75t_L g5798 ( 
.A(n_5204),
.Y(n_5798)
);

INVx1_ASAP7_75t_L g5799 ( 
.A(n_5313),
.Y(n_5799)
);

INVx2_ASAP7_75t_SL g5800 ( 
.A(n_5205),
.Y(n_5800)
);

AOI22xp33_ASAP7_75t_L g5801 ( 
.A1(n_5211),
.A2(n_4496),
.B1(n_4551),
.B2(n_4544),
.Y(n_5801)
);

AND2x2_ASAP7_75t_L g5802 ( 
.A(n_5290),
.B(n_4993),
.Y(n_5802)
);

BUFx6f_ASAP7_75t_L g5803 ( 
.A(n_5308),
.Y(n_5803)
);

INVx3_ASAP7_75t_L g5804 ( 
.A(n_5560),
.Y(n_5804)
);

NAND2xp5_ASAP7_75t_L g5805 ( 
.A(n_5350),
.B(n_5061),
.Y(n_5805)
);

AND2x2_ASAP7_75t_L g5806 ( 
.A(n_5291),
.B(n_4782),
.Y(n_5806)
);

AND2x2_ASAP7_75t_L g5807 ( 
.A(n_5291),
.B(n_4782),
.Y(n_5807)
);

AND2x2_ASAP7_75t_L g5808 ( 
.A(n_5357),
.B(n_4705),
.Y(n_5808)
);

INVx1_ASAP7_75t_SL g5809 ( 
.A(n_5205),
.Y(n_5809)
);

OAI22xp5_ASAP7_75t_L g5810 ( 
.A1(n_5455),
.A2(n_4900),
.B1(n_4946),
.B2(n_4822),
.Y(n_5810)
);

INVx1_ASAP7_75t_L g5811 ( 
.A(n_5317),
.Y(n_5811)
);

INVx1_ASAP7_75t_L g5812 ( 
.A(n_5317),
.Y(n_5812)
);

INVx2_ASAP7_75t_L g5813 ( 
.A(n_5215),
.Y(n_5813)
);

INVx1_ASAP7_75t_L g5814 ( 
.A(n_5323),
.Y(n_5814)
);

INVx1_ASAP7_75t_L g5815 ( 
.A(n_5323),
.Y(n_5815)
);

OR2x2_ASAP7_75t_L g5816 ( 
.A(n_5485),
.B(n_5150),
.Y(n_5816)
);

AND2x2_ASAP7_75t_L g5817 ( 
.A(n_5357),
.B(n_5363),
.Y(n_5817)
);

NAND2xp5_ASAP7_75t_L g5818 ( 
.A(n_5350),
.B(n_5063),
.Y(n_5818)
);

INVx1_ASAP7_75t_L g5819 ( 
.A(n_5331),
.Y(n_5819)
);

HB1xp67_ASAP7_75t_L g5820 ( 
.A(n_5204),
.Y(n_5820)
);

NAND2xp5_ASAP7_75t_L g5821 ( 
.A(n_5316),
.B(n_5069),
.Y(n_5821)
);

AND2x2_ASAP7_75t_L g5822 ( 
.A(n_5363),
.B(n_4705),
.Y(n_5822)
);

INVx2_ASAP7_75t_L g5823 ( 
.A(n_5215),
.Y(n_5823)
);

NAND2xp5_ASAP7_75t_L g5824 ( 
.A(n_5319),
.B(n_5083),
.Y(n_5824)
);

INVx2_ASAP7_75t_L g5825 ( 
.A(n_5215),
.Y(n_5825)
);

HB1xp67_ASAP7_75t_L g5826 ( 
.A(n_5442),
.Y(n_5826)
);

AOI22xp33_ASAP7_75t_SL g5827 ( 
.A1(n_5211),
.A2(n_4317),
.B1(n_4383),
.B2(n_4379),
.Y(n_5827)
);

AND2x2_ASAP7_75t_L g5828 ( 
.A(n_5364),
.B(n_4721),
.Y(n_5828)
);

INVx1_ASAP7_75t_L g5829 ( 
.A(n_5331),
.Y(n_5829)
);

AND2x2_ASAP7_75t_L g5830 ( 
.A(n_5364),
.B(n_4721),
.Y(n_5830)
);

NAND2xp5_ASAP7_75t_L g5831 ( 
.A(n_5349),
.B(n_5100),
.Y(n_5831)
);

INVx1_ASAP7_75t_L g5832 ( 
.A(n_5332),
.Y(n_5832)
);

CKINVDCx5p33_ASAP7_75t_R g5833 ( 
.A(n_5308),
.Y(n_5833)
);

INVx2_ASAP7_75t_L g5834 ( 
.A(n_5223),
.Y(n_5834)
);

AND2x2_ASAP7_75t_L g5835 ( 
.A(n_5367),
.B(n_4873),
.Y(n_5835)
);

NAND3xp33_ASAP7_75t_L g5836 ( 
.A(n_5374),
.B(n_4971),
.C(n_4818),
.Y(n_5836)
);

INVx1_ASAP7_75t_L g5837 ( 
.A(n_5332),
.Y(n_5837)
);

NAND2xp5_ASAP7_75t_L g5838 ( 
.A(n_5442),
.B(n_5105),
.Y(n_5838)
);

INVx1_ASAP7_75t_L g5839 ( 
.A(n_5334),
.Y(n_5839)
);

INVx2_ASAP7_75t_L g5840 ( 
.A(n_5223),
.Y(n_5840)
);

AND2x2_ASAP7_75t_L g5841 ( 
.A(n_5367),
.B(n_4873),
.Y(n_5841)
);

INVx1_ASAP7_75t_L g5842 ( 
.A(n_5334),
.Y(n_5842)
);

INVx3_ASAP7_75t_L g5843 ( 
.A(n_5560),
.Y(n_5843)
);

INVx1_ASAP7_75t_L g5844 ( 
.A(n_5336),
.Y(n_5844)
);

INVx1_ASAP7_75t_L g5845 ( 
.A(n_5336),
.Y(n_5845)
);

NAND2xp5_ASAP7_75t_SL g5846 ( 
.A(n_5318),
.B(n_5119),
.Y(n_5846)
);

INVx1_ASAP7_75t_L g5847 ( 
.A(n_5338),
.Y(n_5847)
);

AND2x2_ASAP7_75t_L g5848 ( 
.A(n_5372),
.B(n_4920),
.Y(n_5848)
);

INVx1_ASAP7_75t_L g5849 ( 
.A(n_5338),
.Y(n_5849)
);

INVx1_ASAP7_75t_L g5850 ( 
.A(n_5343),
.Y(n_5850)
);

AOI22xp33_ASAP7_75t_SL g5851 ( 
.A1(n_5375),
.A2(n_4317),
.B1(n_4383),
.B2(n_4379),
.Y(n_5851)
);

OR2x2_ASAP7_75t_L g5852 ( 
.A(n_5485),
.B(n_5156),
.Y(n_5852)
);

INVx2_ASAP7_75t_L g5853 ( 
.A(n_5223),
.Y(n_5853)
);

CKINVDCx5p33_ASAP7_75t_R g5854 ( 
.A(n_5308),
.Y(n_5854)
);

INVx1_ASAP7_75t_L g5855 ( 
.A(n_5343),
.Y(n_5855)
);

OR2x2_ASAP7_75t_L g5856 ( 
.A(n_5366),
.B(n_5156),
.Y(n_5856)
);

NAND2xp5_ASAP7_75t_L g5857 ( 
.A(n_5438),
.B(n_5188),
.Y(n_5857)
);

INVx1_ASAP7_75t_L g5858 ( 
.A(n_5347),
.Y(n_5858)
);

AOI22xp33_ASAP7_75t_SL g5859 ( 
.A1(n_5375),
.A2(n_4317),
.B1(n_4383),
.B2(n_4379),
.Y(n_5859)
);

AND2x2_ASAP7_75t_L g5860 ( 
.A(n_5372),
.B(n_4920),
.Y(n_5860)
);

AND2x2_ASAP7_75t_L g5861 ( 
.A(n_5377),
.B(n_4963),
.Y(n_5861)
);

BUFx3_ASAP7_75t_L g5862 ( 
.A(n_5557),
.Y(n_5862)
);

INVx2_ASAP7_75t_L g5863 ( 
.A(n_5239),
.Y(n_5863)
);

NOR2xp67_ASAP7_75t_L g5864 ( 
.A(n_5387),
.B(n_4906),
.Y(n_5864)
);

NOR2xp67_ASAP7_75t_L g5865 ( 
.A(n_5387),
.B(n_4906),
.Y(n_5865)
);

INVx1_ASAP7_75t_L g5866 ( 
.A(n_5347),
.Y(n_5866)
);

INVx1_ASAP7_75t_L g5867 ( 
.A(n_5353),
.Y(n_5867)
);

INVx4_ASAP7_75t_L g5868 ( 
.A(n_5399),
.Y(n_5868)
);

NAND2xp5_ASAP7_75t_L g5869 ( 
.A(n_5254),
.B(n_5188),
.Y(n_5869)
);

INVx1_ASAP7_75t_L g5870 ( 
.A(n_5353),
.Y(n_5870)
);

AND2x2_ASAP7_75t_L g5871 ( 
.A(n_5377),
.B(n_5020),
.Y(n_5871)
);

INVx2_ASAP7_75t_L g5872 ( 
.A(n_5239),
.Y(n_5872)
);

INVx1_ASAP7_75t_L g5873 ( 
.A(n_5356),
.Y(n_5873)
);

INVx1_ASAP7_75t_L g5874 ( 
.A(n_5356),
.Y(n_5874)
);

AND2x2_ASAP7_75t_L g5875 ( 
.A(n_5403),
.B(n_5020),
.Y(n_5875)
);

AND2x2_ASAP7_75t_L g5876 ( 
.A(n_5403),
.B(n_5023),
.Y(n_5876)
);

INVx1_ASAP7_75t_L g5877 ( 
.A(n_5361),
.Y(n_5877)
);

AND2x2_ASAP7_75t_L g5878 ( 
.A(n_5412),
.B(n_5023),
.Y(n_5878)
);

HB1xp67_ASAP7_75t_L g5879 ( 
.A(n_5271),
.Y(n_5879)
);

AOI22xp33_ASAP7_75t_L g5880 ( 
.A1(n_5567),
.A2(n_4496),
.B1(n_4551),
.B2(n_4544),
.Y(n_5880)
);

NAND2xp5_ASAP7_75t_L g5881 ( 
.A(n_5254),
.B(n_5354),
.Y(n_5881)
);

AND2x4_ASAP7_75t_L g5882 ( 
.A(n_5555),
.B(n_5155),
.Y(n_5882)
);

AND2x2_ASAP7_75t_L g5883 ( 
.A(n_5412),
.B(n_5423),
.Y(n_5883)
);

AND2x2_ASAP7_75t_L g5884 ( 
.A(n_5423),
.B(n_4851),
.Y(n_5884)
);

INVx2_ASAP7_75t_L g5885 ( 
.A(n_5239),
.Y(n_5885)
);

INVx2_ASAP7_75t_SL g5886 ( 
.A(n_5260),
.Y(n_5886)
);

NAND2xp5_ASAP7_75t_L g5887 ( 
.A(n_5254),
.B(n_5162),
.Y(n_5887)
);

INVx4_ASAP7_75t_L g5888 ( 
.A(n_5399),
.Y(n_5888)
);

OR2x2_ASAP7_75t_L g5889 ( 
.A(n_5366),
.B(n_5478),
.Y(n_5889)
);

CKINVDCx5p33_ASAP7_75t_R g5890 ( 
.A(n_5557),
.Y(n_5890)
);

OR2x2_ASAP7_75t_L g5891 ( 
.A(n_5478),
.B(n_5162),
.Y(n_5891)
);

INVx1_ASAP7_75t_L g5892 ( 
.A(n_5361),
.Y(n_5892)
);

AND2x2_ASAP7_75t_L g5893 ( 
.A(n_5430),
.B(n_4851),
.Y(n_5893)
);

INVx2_ASAP7_75t_L g5894 ( 
.A(n_5245),
.Y(n_5894)
);

BUFx3_ASAP7_75t_L g5895 ( 
.A(n_5557),
.Y(n_5895)
);

INVx1_ASAP7_75t_L g5896 ( 
.A(n_5362),
.Y(n_5896)
);

AND2x2_ASAP7_75t_L g5897 ( 
.A(n_5430),
.B(n_5168),
.Y(n_5897)
);

AND2x2_ASAP7_75t_L g5898 ( 
.A(n_5255),
.B(n_5242),
.Y(n_5898)
);

OR2x2_ASAP7_75t_L g5899 ( 
.A(n_5490),
.B(n_5163),
.Y(n_5899)
);

NAND2xp5_ASAP7_75t_L g5900 ( 
.A(n_5254),
.B(n_5163),
.Y(n_5900)
);

NAND2xp5_ASAP7_75t_L g5901 ( 
.A(n_5354),
.B(n_5170),
.Y(n_5901)
);

AND2x2_ASAP7_75t_L g5902 ( 
.A(n_5255),
.B(n_5168),
.Y(n_5902)
);

AOI22xp33_ASAP7_75t_L g5903 ( 
.A1(n_5375),
.A2(n_4544),
.B1(n_4551),
.B2(n_4500),
.Y(n_5903)
);

AND2x2_ASAP7_75t_L g5904 ( 
.A(n_5242),
.B(n_5168),
.Y(n_5904)
);

NAND2xp5_ASAP7_75t_L g5905 ( 
.A(n_5354),
.B(n_5170),
.Y(n_5905)
);

NAND2xp5_ASAP7_75t_L g5906 ( 
.A(n_5354),
.B(n_5175),
.Y(n_5906)
);

INVx2_ASAP7_75t_L g5907 ( 
.A(n_5245),
.Y(n_5907)
);

AOI22xp33_ASAP7_75t_SL g5908 ( 
.A1(n_5252),
.A2(n_4317),
.B1(n_4415),
.B2(n_4359),
.Y(n_5908)
);

NAND2x1p5_ASAP7_75t_L g5909 ( 
.A(n_5237),
.B(n_4832),
.Y(n_5909)
);

HB1xp67_ASAP7_75t_L g5910 ( 
.A(n_5271),
.Y(n_5910)
);

INVx2_ASAP7_75t_L g5911 ( 
.A(n_5245),
.Y(n_5911)
);

INVx2_ASAP7_75t_L g5912 ( 
.A(n_5261),
.Y(n_5912)
);

INVx1_ASAP7_75t_L g5913 ( 
.A(n_5362),
.Y(n_5913)
);

AND2x2_ASAP7_75t_L g5914 ( 
.A(n_5296),
.B(n_4790),
.Y(n_5914)
);

INVx1_ASAP7_75t_L g5915 ( 
.A(n_5380),
.Y(n_5915)
);

INVx1_ASAP7_75t_L g5916 ( 
.A(n_5380),
.Y(n_5916)
);

NAND2xp5_ASAP7_75t_L g5917 ( 
.A(n_5410),
.B(n_5447),
.Y(n_5917)
);

INVx1_ASAP7_75t_L g5918 ( 
.A(n_5382),
.Y(n_5918)
);

AOI21xp33_ASAP7_75t_L g5919 ( 
.A1(n_5253),
.A2(n_5026),
.B(n_5016),
.Y(n_5919)
);

INVx8_ASAP7_75t_L g5920 ( 
.A(n_5399),
.Y(n_5920)
);

INVx1_ASAP7_75t_SL g5921 ( 
.A(n_5260),
.Y(n_5921)
);

AND2x2_ASAP7_75t_L g5922 ( 
.A(n_5296),
.B(n_4862),
.Y(n_5922)
);

INVx1_ASAP7_75t_L g5923 ( 
.A(n_5382),
.Y(n_5923)
);

INVx2_ASAP7_75t_L g5924 ( 
.A(n_5261),
.Y(n_5924)
);

OR2x2_ASAP7_75t_L g5925 ( 
.A(n_5490),
.B(n_5368),
.Y(n_5925)
);

AND2x2_ASAP7_75t_L g5926 ( 
.A(n_5310),
.B(n_4862),
.Y(n_5926)
);

AND2x2_ASAP7_75t_L g5927 ( 
.A(n_5310),
.B(n_4862),
.Y(n_5927)
);

INVx1_ASAP7_75t_L g5928 ( 
.A(n_5385),
.Y(n_5928)
);

AND2x2_ASAP7_75t_L g5929 ( 
.A(n_5451),
.B(n_4862),
.Y(n_5929)
);

INVx1_ASAP7_75t_L g5930 ( 
.A(n_5385),
.Y(n_5930)
);

INVx2_ASAP7_75t_L g5931 ( 
.A(n_5261),
.Y(n_5931)
);

HB1xp67_ASAP7_75t_L g5932 ( 
.A(n_5271),
.Y(n_5932)
);

NAND2xp5_ASAP7_75t_L g5933 ( 
.A(n_5410),
.B(n_5175),
.Y(n_5933)
);

INVx1_ASAP7_75t_L g5934 ( 
.A(n_5386),
.Y(n_5934)
);

INVx2_ASAP7_75t_L g5935 ( 
.A(n_5284),
.Y(n_5935)
);

INVx2_ASAP7_75t_L g5936 ( 
.A(n_5284),
.Y(n_5936)
);

INVx1_ASAP7_75t_L g5937 ( 
.A(n_5386),
.Y(n_5937)
);

INVx1_ASAP7_75t_L g5938 ( 
.A(n_5389),
.Y(n_5938)
);

AND2x4_ASAP7_75t_L g5939 ( 
.A(n_5572),
.B(n_5161),
.Y(n_5939)
);

AND2x4_ASAP7_75t_SL g5940 ( 
.A(n_5335),
.B(n_4760),
.Y(n_5940)
);

OAI21xp5_ASAP7_75t_L g5941 ( 
.A1(n_5836),
.A2(n_5374),
.B(n_5258),
.Y(n_5941)
);

INVx2_ASAP7_75t_L g5942 ( 
.A(n_5652),
.Y(n_5942)
);

AND2x2_ASAP7_75t_L g5943 ( 
.A(n_5726),
.B(n_5667),
.Y(n_5943)
);

OAI221xp5_ASAP7_75t_L g5944 ( 
.A1(n_5728),
.A2(n_5342),
.B1(n_5516),
.B2(n_5465),
.C(n_5397),
.Y(n_5944)
);

AOI222xp33_ASAP7_75t_L g5945 ( 
.A1(n_5608),
.A2(n_5199),
.B1(n_5791),
.B2(n_5789),
.C1(n_5440),
.C2(n_5680),
.Y(n_5945)
);

NOR2x1p5_ASAP7_75t_L g5946 ( 
.A(n_5607),
.B(n_5610),
.Y(n_5946)
);

AND2x2_ASAP7_75t_L g5947 ( 
.A(n_5697),
.B(n_5287),
.Y(n_5947)
);

OR2x2_ASAP7_75t_L g5948 ( 
.A(n_5603),
.B(n_5368),
.Y(n_5948)
);

NAND2xp5_ASAP7_75t_SL g5949 ( 
.A(n_5652),
.B(n_5237),
.Y(n_5949)
);

INVx2_ASAP7_75t_L g5950 ( 
.A(n_5652),
.Y(n_5950)
);

INVx4_ASAP7_75t_L g5951 ( 
.A(n_5803),
.Y(n_5951)
);

AOI221xp5_ASAP7_75t_L g5952 ( 
.A1(n_5919),
.A2(n_5440),
.B1(n_5236),
.B2(n_5221),
.C(n_5397),
.Y(n_5952)
);

AOI22xp5_ASAP7_75t_L g5953 ( 
.A1(n_5717),
.A2(n_5197),
.B1(n_5266),
.B2(n_5253),
.Y(n_5953)
);

INVx1_ASAP7_75t_L g5954 ( 
.A(n_5616),
.Y(n_5954)
);

HB1xp67_ASAP7_75t_L g5955 ( 
.A(n_5800),
.Y(n_5955)
);

INVx1_ASAP7_75t_L g5956 ( 
.A(n_5612),
.Y(n_5956)
);

INVx1_ASAP7_75t_L g5957 ( 
.A(n_5612),
.Y(n_5957)
);

INVxp67_ASAP7_75t_L g5958 ( 
.A(n_5794),
.Y(n_5958)
);

OAI21xp33_ASAP7_75t_L g5959 ( 
.A1(n_5908),
.A2(n_5258),
.B(n_5280),
.Y(n_5959)
);

AND2x2_ASAP7_75t_L g5960 ( 
.A(n_5726),
.B(n_5287),
.Y(n_5960)
);

INVx5_ASAP7_75t_SL g5961 ( 
.A(n_5803),
.Y(n_5961)
);

AOI22xp33_ASAP7_75t_L g5962 ( 
.A1(n_5661),
.A2(n_5197),
.B1(n_5236),
.B2(n_5253),
.Y(n_5962)
);

NAND2xp5_ASAP7_75t_L g5963 ( 
.A(n_5809),
.B(n_5410),
.Y(n_5963)
);

AOI32xp33_ASAP7_75t_L g5964 ( 
.A1(n_5827),
.A2(n_5236),
.A3(n_5408),
.B1(n_5447),
.B2(n_5410),
.Y(n_5964)
);

INVx2_ASAP7_75t_L g5965 ( 
.A(n_5737),
.Y(n_5965)
);

AND2x2_ASAP7_75t_L g5966 ( 
.A(n_5697),
.B(n_5667),
.Y(n_5966)
);

NOR4xp25_ASAP7_75t_SL g5967 ( 
.A(n_5621),
.B(n_5573),
.C(n_5037),
.D(n_5050),
.Y(n_5967)
);

OAI31xp33_ASAP7_75t_L g5968 ( 
.A1(n_5661),
.A2(n_5345),
.A3(n_5252),
.B(n_5359),
.Y(n_5968)
);

OR2x2_ASAP7_75t_L g5969 ( 
.A(n_5889),
.B(n_5420),
.Y(n_5969)
);

HB1xp67_ASAP7_75t_L g5970 ( 
.A(n_5800),
.Y(n_5970)
);

OAI22xp5_ASAP7_75t_L g5971 ( 
.A1(n_5641),
.A2(n_5408),
.B1(n_5318),
.B2(n_5573),
.Y(n_5971)
);

INVx2_ASAP7_75t_L g5972 ( 
.A(n_5737),
.Y(n_5972)
);

NAND3xp33_ASAP7_75t_L g5973 ( 
.A(n_5851),
.B(n_5236),
.C(n_5447),
.Y(n_5973)
);

INVx2_ASAP7_75t_L g5974 ( 
.A(n_5737),
.Y(n_5974)
);

INVx3_ASAP7_75t_L g5975 ( 
.A(n_5641),
.Y(n_5975)
);

INVx1_ASAP7_75t_L g5976 ( 
.A(n_5620),
.Y(n_5976)
);

INVxp67_ASAP7_75t_L g5977 ( 
.A(n_5794),
.Y(n_5977)
);

NAND3xp33_ASAP7_75t_L g5978 ( 
.A(n_5859),
.B(n_5459),
.C(n_5447),
.Y(n_5978)
);

AOI22xp5_ASAP7_75t_L g5979 ( 
.A1(n_5756),
.A2(n_5197),
.B1(n_5266),
.B2(n_5253),
.Y(n_5979)
);

INVx1_ASAP7_75t_L g5980 ( 
.A(n_5620),
.Y(n_5980)
);

NAND2xp5_ASAP7_75t_L g5981 ( 
.A(n_5921),
.B(n_5459),
.Y(n_5981)
);

OR2x2_ASAP7_75t_L g5982 ( 
.A(n_5889),
.B(n_5420),
.Y(n_5982)
);

BUFx3_ASAP7_75t_L g5983 ( 
.A(n_5607),
.Y(n_5983)
);

HB1xp67_ASAP7_75t_L g5984 ( 
.A(n_5886),
.Y(n_5984)
);

INVx2_ASAP7_75t_L g5985 ( 
.A(n_5756),
.Y(n_5985)
);

AND2x2_ASAP7_75t_L g5986 ( 
.A(n_5663),
.B(n_5303),
.Y(n_5986)
);

NAND2xp33_ASAP7_75t_R g5987 ( 
.A(n_5641),
.B(n_5231),
.Y(n_5987)
);

AOI22xp33_ASAP7_75t_L g5988 ( 
.A1(n_5679),
.A2(n_5756),
.B1(n_5778),
.B2(n_5932),
.Y(n_5988)
);

AOI22xp33_ASAP7_75t_L g5989 ( 
.A1(n_5679),
.A2(n_5197),
.B1(n_5243),
.B2(n_5266),
.Y(n_5989)
);

NAND3xp33_ASAP7_75t_L g5990 ( 
.A(n_5641),
.B(n_5487),
.C(n_5459),
.Y(n_5990)
);

INVx1_ASAP7_75t_SL g5991 ( 
.A(n_5663),
.Y(n_5991)
);

AND2x2_ASAP7_75t_L g5992 ( 
.A(n_5666),
.B(n_5303),
.Y(n_5992)
);

AOI22xp33_ASAP7_75t_L g5993 ( 
.A1(n_5778),
.A2(n_5243),
.B1(n_5266),
.B2(n_5459),
.Y(n_5993)
);

AND2x2_ASAP7_75t_L g5994 ( 
.A(n_5666),
.B(n_5675),
.Y(n_5994)
);

OAI221xp5_ASAP7_75t_L g5995 ( 
.A1(n_5668),
.A2(n_5401),
.B1(n_5359),
.B2(n_5391),
.C(n_5280),
.Y(n_5995)
);

OAI21xp5_ASAP7_75t_L g5996 ( 
.A1(n_5668),
.A2(n_5506),
.B(n_5487),
.Y(n_5996)
);

AOI221xp5_ASAP7_75t_L g5997 ( 
.A1(n_5778),
.A2(n_5487),
.B1(n_5481),
.B2(n_5401),
.C(n_5369),
.Y(n_5997)
);

INVx1_ASAP7_75t_L g5998 ( 
.A(n_5687),
.Y(n_5998)
);

NOR2xp33_ASAP7_75t_R g5999 ( 
.A(n_5648),
.B(n_4884),
.Y(n_5999)
);

AND2x4_ASAP7_75t_L g6000 ( 
.A(n_5886),
.B(n_5592),
.Y(n_6000)
);

OAI211xp5_ASAP7_75t_L g6001 ( 
.A1(n_5635),
.A2(n_5418),
.B(n_5506),
.C(n_5461),
.Y(n_6001)
);

AOI211xp5_ASAP7_75t_L g6002 ( 
.A1(n_5699),
.A2(n_5481),
.B(n_5548),
.C(n_5583),
.Y(n_6002)
);

AOI22xp33_ASAP7_75t_L g6003 ( 
.A1(n_5879),
.A2(n_5243),
.B1(n_5487),
.B2(n_5369),
.Y(n_6003)
);

OAI211xp5_ASAP7_75t_L g6004 ( 
.A1(n_5640),
.A2(n_5418),
.B(n_5461),
.C(n_5513),
.Y(n_6004)
);

NAND3xp33_ASAP7_75t_SL g6005 ( 
.A(n_5615),
.B(n_5263),
.C(n_5208),
.Y(n_6005)
);

AOI322xp5_ASAP7_75t_L g6006 ( 
.A1(n_5712),
.A2(n_5360),
.A3(n_5284),
.B1(n_5306),
.B2(n_5315),
.C1(n_5302),
.C2(n_5206),
.Y(n_6006)
);

AOI22xp33_ASAP7_75t_SL g6007 ( 
.A1(n_5720),
.A2(n_5378),
.B1(n_5548),
.B2(n_5243),
.Y(n_6007)
);

NAND2xp5_ASAP7_75t_L g6008 ( 
.A(n_5643),
.B(n_5360),
.Y(n_6008)
);

AOI22xp33_ASAP7_75t_SL g6009 ( 
.A1(n_5720),
.A2(n_5378),
.B1(n_5369),
.B2(n_5274),
.Y(n_6009)
);

INVx1_ASAP7_75t_L g6010 ( 
.A(n_5687),
.Y(n_6010)
);

AND2x4_ASAP7_75t_L g6011 ( 
.A(n_5675),
.B(n_5592),
.Y(n_6011)
);

INVx2_ASAP7_75t_L g6012 ( 
.A(n_5668),
.Y(n_6012)
);

BUFx6f_ASAP7_75t_L g6013 ( 
.A(n_5803),
.Y(n_6013)
);

NOR4xp25_ASAP7_75t_SL g6014 ( 
.A(n_5846),
.B(n_4937),
.C(n_4898),
.D(n_5080),
.Y(n_6014)
);

NAND2xp33_ASAP7_75t_SL g6015 ( 
.A(n_5803),
.B(n_4841),
.Y(n_6015)
);

AOI22xp5_ASAP7_75t_L g6016 ( 
.A1(n_5668),
.A2(n_5378),
.B1(n_5369),
.B2(n_5388),
.Y(n_6016)
);

AOI22xp5_ASAP7_75t_L g6017 ( 
.A1(n_5782),
.A2(n_5378),
.B1(n_5388),
.B2(n_5263),
.Y(n_6017)
);

INVx1_ASAP7_75t_L g6018 ( 
.A(n_5690),
.Y(n_6018)
);

OAI22xp5_ASAP7_75t_L g6019 ( 
.A1(n_5613),
.A2(n_5625),
.B1(n_5391),
.B2(n_5698),
.Y(n_6019)
);

INVx1_ASAP7_75t_L g6020 ( 
.A(n_5690),
.Y(n_6020)
);

AOI22xp5_ASAP7_75t_L g6021 ( 
.A1(n_5910),
.A2(n_5388),
.B1(n_5274),
.B2(n_5208),
.Y(n_6021)
);

INVx1_ASAP7_75t_L g6022 ( 
.A(n_5692),
.Y(n_6022)
);

AND2x2_ASAP7_75t_L g6023 ( 
.A(n_5765),
.B(n_5376),
.Y(n_6023)
);

OAI222xp33_ASAP7_75t_L g6024 ( 
.A1(n_5682),
.A2(n_5503),
.B1(n_5231),
.B2(n_5244),
.C1(n_5523),
.C2(n_5529),
.Y(n_6024)
);

AND2x2_ASAP7_75t_L g6025 ( 
.A(n_5765),
.B(n_5376),
.Y(n_6025)
);

INVx2_ASAP7_75t_L g6026 ( 
.A(n_5803),
.Y(n_6026)
);

AOI21xp33_ASAP7_75t_L g6027 ( 
.A1(n_5622),
.A2(n_5271),
.B(n_5388),
.Y(n_6027)
);

NAND2xp5_ASAP7_75t_L g6028 ( 
.A(n_5798),
.B(n_5433),
.Y(n_6028)
);

AOI22xp33_ASAP7_75t_L g6029 ( 
.A1(n_5622),
.A2(n_5358),
.B1(n_5274),
.B2(n_5404),
.Y(n_6029)
);

BUFx12f_ASAP7_75t_L g6030 ( 
.A(n_5833),
.Y(n_6030)
);

INVx2_ASAP7_75t_L g6031 ( 
.A(n_5862),
.Y(n_6031)
);

OAI31xp33_ASAP7_75t_L g6032 ( 
.A1(n_5659),
.A2(n_5345),
.A3(n_5503),
.B(n_5448),
.Y(n_6032)
);

HB1xp67_ASAP7_75t_L g6033 ( 
.A(n_5862),
.Y(n_6033)
);

INVx3_ASAP7_75t_L g6034 ( 
.A(n_5610),
.Y(n_6034)
);

AND2x4_ASAP7_75t_L g6035 ( 
.A(n_5604),
.B(n_5592),
.Y(n_6035)
);

AOI21xp33_ASAP7_75t_L g6036 ( 
.A1(n_5639),
.A2(n_5358),
.B(n_5274),
.Y(n_6036)
);

INVxp67_ASAP7_75t_SL g6037 ( 
.A(n_5633),
.Y(n_6037)
);

AND2x2_ASAP7_75t_L g6038 ( 
.A(n_5898),
.B(n_5463),
.Y(n_6038)
);

BUFx3_ASAP7_75t_L g6039 ( 
.A(n_5633),
.Y(n_6039)
);

OAI22xp33_ASAP7_75t_L g6040 ( 
.A1(n_5646),
.A2(n_5231),
.B1(n_5244),
.B2(n_5526),
.Y(n_6040)
);

INVx2_ASAP7_75t_L g6041 ( 
.A(n_5895),
.Y(n_6041)
);

INVx1_ASAP7_75t_L g6042 ( 
.A(n_5692),
.Y(n_6042)
);

CKINVDCx11_ASAP7_75t_R g6043 ( 
.A(n_5651),
.Y(n_6043)
);

NAND2xp5_ASAP7_75t_L g6044 ( 
.A(n_5820),
.B(n_5301),
.Y(n_6044)
);

INVx1_ASAP7_75t_L g6045 ( 
.A(n_5693),
.Y(n_6045)
);

INVx2_ASAP7_75t_L g6046 ( 
.A(n_5895),
.Y(n_6046)
);

NAND3xp33_ASAP7_75t_L g6047 ( 
.A(n_5639),
.B(n_5301),
.C(n_5231),
.Y(n_6047)
);

AOI22xp33_ASAP7_75t_L g6048 ( 
.A1(n_5646),
.A2(n_5358),
.B1(n_5413),
.B2(n_5404),
.Y(n_6048)
);

INVx2_ASAP7_75t_L g6049 ( 
.A(n_5733),
.Y(n_6049)
);

INVx2_ASAP7_75t_L g6050 ( 
.A(n_5733),
.Y(n_6050)
);

INVxp67_ASAP7_75t_L g6051 ( 
.A(n_5660),
.Y(n_6051)
);

INVx2_ASAP7_75t_L g6052 ( 
.A(n_5898),
.Y(n_6052)
);

OAI21x1_ASAP7_75t_L g6053 ( 
.A1(n_5804),
.A2(n_5297),
.B(n_5289),
.Y(n_6053)
);

AND2x2_ASAP7_75t_L g6054 ( 
.A(n_5793),
.B(n_5463),
.Y(n_6054)
);

AO21x2_ASAP7_75t_L g6055 ( 
.A1(n_5721),
.A2(n_5773),
.B(n_5746),
.Y(n_6055)
);

INVx1_ASAP7_75t_L g6056 ( 
.A(n_5693),
.Y(n_6056)
);

INVx2_ASAP7_75t_L g6057 ( 
.A(n_5647),
.Y(n_6057)
);

AND2x2_ASAP7_75t_L g6058 ( 
.A(n_5793),
.B(n_5472),
.Y(n_6058)
);

OA21x2_ASAP7_75t_L g6059 ( 
.A1(n_5903),
.A2(n_5306),
.B(n_5302),
.Y(n_6059)
);

INVx1_ASAP7_75t_L g6060 ( 
.A(n_5700),
.Y(n_6060)
);

BUFx2_ASAP7_75t_L g6061 ( 
.A(n_5706),
.Y(n_6061)
);

AOI22xp33_ASAP7_75t_L g6062 ( 
.A1(n_5647),
.A2(n_5358),
.B1(n_5413),
.B2(n_5404),
.Y(n_6062)
);

AOI221xp5_ASAP7_75t_L g6063 ( 
.A1(n_5787),
.A2(n_5583),
.B1(n_5526),
.B2(n_5413),
.C(n_5404),
.Y(n_6063)
);

OAI321xp33_ASAP7_75t_L g6064 ( 
.A1(n_5914),
.A2(n_5231),
.A3(n_5244),
.B1(n_5439),
.B2(n_5286),
.C(n_5297),
.Y(n_6064)
);

AND2x2_ASAP7_75t_L g6065 ( 
.A(n_5802),
.B(n_5472),
.Y(n_6065)
);

BUFx3_ASAP7_75t_L g6066 ( 
.A(n_5833),
.Y(n_6066)
);

NAND2xp5_ASAP7_75t_L g6067 ( 
.A(n_5826),
.B(n_5301),
.Y(n_6067)
);

AND2x2_ASAP7_75t_L g6068 ( 
.A(n_5802),
.B(n_5817),
.Y(n_6068)
);

NOR2xp33_ASAP7_75t_R g6069 ( 
.A(n_5854),
.B(n_4956),
.Y(n_6069)
);

INVxp67_ASAP7_75t_SL g6070 ( 
.A(n_5775),
.Y(n_6070)
);

AOI22xp33_ASAP7_75t_L g6071 ( 
.A1(n_5801),
.A2(n_5413),
.B1(n_5309),
.B2(n_5279),
.Y(n_6071)
);

NAND3xp33_ASAP7_75t_L g6072 ( 
.A(n_5854),
.B(n_5301),
.C(n_5233),
.Y(n_6072)
);

OAI221xp5_ASAP7_75t_L g6073 ( 
.A1(n_5880),
.A2(n_5448),
.B1(n_5244),
.B2(n_5267),
.C(n_5306),
.Y(n_6073)
);

NOR3xp33_ASAP7_75t_L g6074 ( 
.A(n_5868),
.B(n_5233),
.C(n_5507),
.Y(n_6074)
);

OAI22xp5_ASAP7_75t_L g6075 ( 
.A1(n_5864),
.A2(n_5244),
.B1(n_5267),
.B2(n_5497),
.Y(n_6075)
);

INVx2_ASAP7_75t_L g6076 ( 
.A(n_5922),
.Y(n_6076)
);

INVx2_ASAP7_75t_L g6077 ( 
.A(n_5922),
.Y(n_6077)
);

NAND3xp33_ASAP7_75t_L g6078 ( 
.A(n_5890),
.B(n_5301),
.C(n_5233),
.Y(n_6078)
);

INVx1_ASAP7_75t_L g6079 ( 
.A(n_5700),
.Y(n_6079)
);

NAND2xp33_ASAP7_75t_R g6080 ( 
.A(n_5890),
.B(n_5507),
.Y(n_6080)
);

HB1xp67_ASAP7_75t_L g6081 ( 
.A(n_5629),
.Y(n_6081)
);

INVx2_ASAP7_75t_L g6082 ( 
.A(n_5926),
.Y(n_6082)
);

NAND2xp5_ASAP7_75t_L g6083 ( 
.A(n_5730),
.B(n_5301),
.Y(n_6083)
);

BUFx2_ASAP7_75t_L g6084 ( 
.A(n_5604),
.Y(n_6084)
);

NAND2xp5_ASAP7_75t_L g6085 ( 
.A(n_5753),
.B(n_5206),
.Y(n_6085)
);

INVx1_ASAP7_75t_L g6086 ( 
.A(n_5708),
.Y(n_6086)
);

INVxp67_ASAP7_75t_L g6087 ( 
.A(n_5763),
.Y(n_6087)
);

INVxp67_ASAP7_75t_SL g6088 ( 
.A(n_5779),
.Y(n_6088)
);

OAI31xp33_ASAP7_75t_L g6089 ( 
.A1(n_5723),
.A2(n_5302),
.A3(n_5315),
.B(n_5286),
.Y(n_6089)
);

OA21x2_ASAP7_75t_L g6090 ( 
.A1(n_5881),
.A2(n_5315),
.B(n_5559),
.Y(n_6090)
);

AOI221xp5_ASAP7_75t_L g6091 ( 
.A1(n_5805),
.A2(n_5309),
.B1(n_5279),
.B2(n_5598),
.C(n_5473),
.Y(n_6091)
);

INVx1_ASAP7_75t_L g6092 ( 
.A(n_5708),
.Y(n_6092)
);

OAI22xp5_ASAP7_75t_L g6093 ( 
.A1(n_5865),
.A2(n_5497),
.B1(n_5523),
.B2(n_5134),
.Y(n_6093)
);

BUFx10_ASAP7_75t_L g6094 ( 
.A(n_5748),
.Y(n_6094)
);

AND2x2_ASAP7_75t_L g6095 ( 
.A(n_5817),
.B(n_5883),
.Y(n_6095)
);

AND2x2_ASAP7_75t_L g6096 ( 
.A(n_5883),
.B(n_5533),
.Y(n_6096)
);

AND2x2_ASAP7_75t_L g6097 ( 
.A(n_5634),
.B(n_5533),
.Y(n_6097)
);

INVxp67_ASAP7_75t_L g6098 ( 
.A(n_5763),
.Y(n_6098)
);

NAND2xp5_ASAP7_75t_L g6099 ( 
.A(n_5654),
.B(n_5328),
.Y(n_6099)
);

AOI22xp33_ASAP7_75t_L g6100 ( 
.A1(n_5818),
.A2(n_5309),
.B1(n_5279),
.B2(n_5598),
.Y(n_6100)
);

AOI22xp5_ASAP7_75t_L g6101 ( 
.A1(n_5914),
.A2(n_5598),
.B1(n_5473),
.B2(n_5454),
.Y(n_6101)
);

AOI22xp33_ASAP7_75t_L g6102 ( 
.A1(n_5727),
.A2(n_5309),
.B1(n_5279),
.B2(n_5598),
.Y(n_6102)
);

INVx1_ASAP7_75t_L g6103 ( 
.A(n_5709),
.Y(n_6103)
);

OAI22xp5_ASAP7_75t_L g6104 ( 
.A1(n_5810),
.A2(n_5857),
.B1(n_5497),
.B2(n_5843),
.Y(n_6104)
);

OR2x2_ASAP7_75t_L g6105 ( 
.A(n_5925),
.B(n_5502),
.Y(n_6105)
);

NOR3xp33_ASAP7_75t_L g6106 ( 
.A(n_5868),
.B(n_5233),
.C(n_5575),
.Y(n_6106)
);

AOI21xp33_ASAP7_75t_L g6107 ( 
.A1(n_5917),
.A2(n_5227),
.B(n_5217),
.Y(n_6107)
);

INVx2_ASAP7_75t_L g6108 ( 
.A(n_5926),
.Y(n_6108)
);

OR2x2_ASAP7_75t_L g6109 ( 
.A(n_5925),
.B(n_5502),
.Y(n_6109)
);

INVx3_ASAP7_75t_L g6110 ( 
.A(n_5804),
.Y(n_6110)
);

AOI22xp33_ASAP7_75t_SL g6111 ( 
.A1(n_5772),
.A2(n_5333),
.B1(n_5473),
.B2(n_5454),
.Y(n_6111)
);

CKINVDCx5p33_ASAP7_75t_R g6112 ( 
.A(n_5651),
.Y(n_6112)
);

INVxp67_ASAP7_75t_SL g6113 ( 
.A(n_5748),
.Y(n_6113)
);

OAI31xp33_ASAP7_75t_L g6114 ( 
.A1(n_5772),
.A2(n_5286),
.A3(n_5439),
.B(n_5407),
.Y(n_6114)
);

AOI221xp5_ASAP7_75t_L g6115 ( 
.A1(n_5752),
.A2(n_5473),
.B1(n_5454),
.B2(n_5479),
.C(n_5414),
.Y(n_6115)
);

AOI221xp5_ASAP7_75t_L g6116 ( 
.A1(n_5752),
.A2(n_5454),
.B1(n_5479),
.B2(n_5414),
.C(n_5415),
.Y(n_6116)
);

INVx1_ASAP7_75t_L g6117 ( 
.A(n_5709),
.Y(n_6117)
);

INVx1_ASAP7_75t_L g6118 ( 
.A(n_5713),
.Y(n_6118)
);

BUFx2_ASAP7_75t_L g6119 ( 
.A(n_5604),
.Y(n_6119)
);

INVx2_ASAP7_75t_L g6120 ( 
.A(n_5927),
.Y(n_6120)
);

AND2x4_ASAP7_75t_L g6121 ( 
.A(n_5605),
.B(n_5575),
.Y(n_6121)
);

INVx1_ASAP7_75t_SL g6122 ( 
.A(n_5605),
.Y(n_6122)
);

OAI22xp5_ASAP7_75t_L g6123 ( 
.A1(n_5804),
.A2(n_5497),
.B1(n_5523),
.B2(n_5529),
.Y(n_6123)
);

NAND3xp33_ASAP7_75t_L g6124 ( 
.A(n_5694),
.B(n_5333),
.C(n_5251),
.Y(n_6124)
);

INVx2_ASAP7_75t_L g6125 ( 
.A(n_5927),
.Y(n_6125)
);

INVx1_ASAP7_75t_L g6126 ( 
.A(n_5713),
.Y(n_6126)
);

HB1xp67_ASAP7_75t_L g6127 ( 
.A(n_5609),
.Y(n_6127)
);

NAND2xp5_ASAP7_75t_L g6128 ( 
.A(n_5626),
.B(n_5328),
.Y(n_6128)
);

OA211x2_ASAP7_75t_L g6129 ( 
.A1(n_5735),
.A2(n_5522),
.B(n_4824),
.C(n_4740),
.Y(n_6129)
);

OAI222xp33_ASAP7_75t_L g6130 ( 
.A1(n_5774),
.A2(n_5523),
.B1(n_5529),
.B2(n_5497),
.C1(n_5439),
.C2(n_5289),
.Y(n_6130)
);

AOI22xp33_ASAP7_75t_L g6131 ( 
.A1(n_5609),
.A2(n_5333),
.B1(n_5479),
.B2(n_4415),
.Y(n_6131)
);

INVx1_ASAP7_75t_L g6132 ( 
.A(n_5715),
.Y(n_6132)
);

AND2x2_ASAP7_75t_L g6133 ( 
.A(n_5634),
.B(n_5217),
.Y(n_6133)
);

AOI222xp33_ASAP7_75t_L g6134 ( 
.A1(n_5774),
.A2(n_5545),
.B1(n_5531),
.B2(n_5547),
.C1(n_5538),
.C2(n_5527),
.Y(n_6134)
);

OAI211xp5_ASAP7_75t_L g6135 ( 
.A1(n_5614),
.A2(n_5618),
.B(n_5783),
.C(n_5513),
.Y(n_6135)
);

HB1xp67_ASAP7_75t_L g6136 ( 
.A(n_5821),
.Y(n_6136)
);

AND2x4_ASAP7_75t_L g6137 ( 
.A(n_5777),
.B(n_5572),
.Y(n_6137)
);

INVx1_ASAP7_75t_L g6138 ( 
.A(n_5715),
.Y(n_6138)
);

AOI22xp33_ASAP7_75t_L g6139 ( 
.A1(n_5754),
.A2(n_5333),
.B1(n_5479),
.B2(n_4415),
.Y(n_6139)
);

INVx2_ASAP7_75t_L g6140 ( 
.A(n_5748),
.Y(n_6140)
);

INVx1_ASAP7_75t_L g6141 ( 
.A(n_5718),
.Y(n_6141)
);

NOR2xp33_ASAP7_75t_L g6142 ( 
.A(n_5868),
.B(n_4788),
.Y(n_6142)
);

INVx1_ASAP7_75t_L g6143 ( 
.A(n_5718),
.Y(n_6143)
);

AOI22xp33_ASAP7_75t_L g6144 ( 
.A1(n_5754),
.A2(n_4415),
.B1(n_4359),
.B2(n_5394),
.Y(n_6144)
);

AND2x2_ASAP7_75t_L g6145 ( 
.A(n_5601),
.B(n_5522),
.Y(n_6145)
);

OAI221xp5_ASAP7_75t_L g6146 ( 
.A1(n_5696),
.A2(n_5098),
.B1(n_5523),
.B2(n_5530),
.C(n_5529),
.Y(n_6146)
);

INVx2_ASAP7_75t_L g6147 ( 
.A(n_5748),
.Y(n_6147)
);

HB1xp67_ASAP7_75t_L g6148 ( 
.A(n_5824),
.Y(n_6148)
);

INVx1_ASAP7_75t_L g6149 ( 
.A(n_5719),
.Y(n_6149)
);

OR2x2_ASAP7_75t_L g6150 ( 
.A(n_5740),
.B(n_5587),
.Y(n_6150)
);

NAND4xp25_ASAP7_75t_L g6151 ( 
.A(n_5736),
.B(n_5525),
.C(n_5586),
.D(n_5541),
.Y(n_6151)
);

INVx2_ASAP7_75t_SL g6152 ( 
.A(n_5650),
.Y(n_6152)
);

INVx2_ASAP7_75t_SL g6153 ( 
.A(n_5650),
.Y(n_6153)
);

AND2x2_ASAP7_75t_L g6154 ( 
.A(n_5637),
.B(n_5227),
.Y(n_6154)
);

HB1xp67_ASAP7_75t_L g6155 ( 
.A(n_5724),
.Y(n_6155)
);

AOI21xp5_ASAP7_75t_L g6156 ( 
.A1(n_5670),
.A2(n_5395),
.B(n_4794),
.Y(n_6156)
);

OAI31xp33_ASAP7_75t_L g6157 ( 
.A1(n_5696),
.A2(n_5407),
.A3(n_5414),
.B(n_5394),
.Y(n_6157)
);

INVx2_ASAP7_75t_L g6158 ( 
.A(n_5748),
.Y(n_6158)
);

AOI22xp33_ASAP7_75t_L g6159 ( 
.A1(n_5701),
.A2(n_4359),
.B1(n_5407),
.B2(n_5394),
.Y(n_6159)
);

AND2x4_ASAP7_75t_L g6160 ( 
.A(n_5777),
.B(n_5572),
.Y(n_6160)
);

NAND4xp25_ASAP7_75t_L g6161 ( 
.A(n_5702),
.B(n_5525),
.C(n_5553),
.D(n_5541),
.Y(n_6161)
);

OAI22xp5_ASAP7_75t_L g6162 ( 
.A1(n_5843),
.A2(n_5529),
.B1(n_4915),
.B2(n_4896),
.Y(n_6162)
);

AOI22xp33_ASAP7_75t_L g6163 ( 
.A1(n_5701),
.A2(n_5427),
.B1(n_5431),
.B2(n_5415),
.Y(n_6163)
);

AND2x2_ASAP7_75t_L g6164 ( 
.A(n_5637),
.B(n_5275),
.Y(n_6164)
);

INVx4_ASAP7_75t_L g6165 ( 
.A(n_5920),
.Y(n_6165)
);

NAND2xp5_ASAP7_75t_L g6166 ( 
.A(n_5630),
.B(n_5348),
.Y(n_6166)
);

INVx1_ASAP7_75t_L g6167 ( 
.A(n_5719),
.Y(n_6167)
);

INVx2_ASAP7_75t_L g6168 ( 
.A(n_5600),
.Y(n_6168)
);

OAI21xp5_ASAP7_75t_L g6169 ( 
.A1(n_5843),
.A2(n_5469),
.B(n_5272),
.Y(n_6169)
);

OAI22xp33_ASAP7_75t_L g6170 ( 
.A1(n_5711),
.A2(n_4909),
.B1(n_5530),
.B2(n_5137),
.Y(n_6170)
);

BUFx3_ASAP7_75t_L g6171 ( 
.A(n_5920),
.Y(n_6171)
);

AOI22xp33_ASAP7_75t_L g6172 ( 
.A1(n_5711),
.A2(n_5427),
.B1(n_5431),
.B2(n_5415),
.Y(n_6172)
);

AOI221xp5_ASAP7_75t_L g6173 ( 
.A1(n_5714),
.A2(n_5431),
.B1(n_5427),
.B2(n_5584),
.C(n_5582),
.Y(n_6173)
);

CKINVDCx16_ASAP7_75t_R g6174 ( 
.A(n_5888),
.Y(n_6174)
);

AND2x2_ASAP7_75t_L g6175 ( 
.A(n_5601),
.B(n_5451),
.Y(n_6175)
);

AND2x2_ASAP7_75t_L g6176 ( 
.A(n_5781),
.B(n_5456),
.Y(n_6176)
);

AOI22xp33_ASAP7_75t_L g6177 ( 
.A1(n_5714),
.A2(n_5649),
.B1(n_5611),
.B2(n_5624),
.Y(n_6177)
);

NAND3xp33_ASAP7_75t_L g6178 ( 
.A(n_5681),
.B(n_5251),
.C(n_5320),
.Y(n_6178)
);

INVx2_ASAP7_75t_L g6179 ( 
.A(n_5600),
.Y(n_6179)
);

NOR2xp33_ASAP7_75t_R g6180 ( 
.A(n_5670),
.B(n_4849),
.Y(n_6180)
);

AND2x2_ASAP7_75t_L g6181 ( 
.A(n_5781),
.B(n_5456),
.Y(n_6181)
);

AOI322xp5_ASAP7_75t_L g6182 ( 
.A1(n_5767),
.A2(n_5565),
.A3(n_5576),
.B1(n_5559),
.B2(n_5588),
.C1(n_5584),
.C2(n_5582),
.Y(n_6182)
);

AND2x2_ASAP7_75t_L g6183 ( 
.A(n_5784),
.B(n_5446),
.Y(n_6183)
);

AND2x4_ASAP7_75t_L g6184 ( 
.A(n_5784),
.B(n_5572),
.Y(n_6184)
);

NAND2xp5_ASAP7_75t_L g6185 ( 
.A(n_5665),
.B(n_5348),
.Y(n_6185)
);

OAI221xp5_ASAP7_75t_L g6186 ( 
.A1(n_5602),
.A2(n_5530),
.B1(n_5320),
.B2(n_5251),
.C(n_4438),
.Y(n_6186)
);

AOI221xp5_ASAP7_75t_L g6187 ( 
.A1(n_5767),
.A2(n_5588),
.B1(n_5596),
.B2(n_5584),
.C(n_5582),
.Y(n_6187)
);

OAI22xp33_ASAP7_75t_L g6188 ( 
.A1(n_5602),
.A2(n_5530),
.B1(n_5137),
.B2(n_5096),
.Y(n_6188)
);

INVx1_ASAP7_75t_L g6189 ( 
.A(n_5722),
.Y(n_6189)
);

AND2x2_ASAP7_75t_L g6190 ( 
.A(n_5790),
.B(n_5446),
.Y(n_6190)
);

BUFx3_ASAP7_75t_L g6191 ( 
.A(n_5920),
.Y(n_6191)
);

OAI31xp33_ASAP7_75t_L g6192 ( 
.A1(n_5678),
.A2(n_5768),
.A3(n_5606),
.B(n_5691),
.Y(n_6192)
);

INVx1_ASAP7_75t_L g6193 ( 
.A(n_5722),
.Y(n_6193)
);

OAI31xp33_ASAP7_75t_L g6194 ( 
.A1(n_5678),
.A2(n_5531),
.A3(n_5538),
.B(n_5527),
.Y(n_6194)
);

INVx1_ASAP7_75t_L g6195 ( 
.A(n_5731),
.Y(n_6195)
);

AND2x4_ASAP7_75t_L g6196 ( 
.A(n_5790),
.B(n_5273),
.Y(n_6196)
);

AOI221xp5_ASAP7_75t_SL g6197 ( 
.A1(n_5684),
.A2(n_4748),
.B1(n_5520),
.B2(n_4944),
.C(n_5270),
.Y(n_6197)
);

AND2x4_ASAP7_75t_L g6198 ( 
.A(n_5674),
.B(n_5273),
.Y(n_6198)
);

AOI21xp5_ASAP7_75t_L g6199 ( 
.A1(n_5831),
.A2(n_5395),
.B(n_5320),
.Y(n_6199)
);

AOI22xp5_ASAP7_75t_L g6200 ( 
.A1(n_5768),
.A2(n_4544),
.B1(n_4903),
.B2(n_4500),
.Y(n_6200)
);

NOR4xp25_ASAP7_75t_SL g6201 ( 
.A(n_5731),
.B(n_4921),
.C(n_4986),
.D(n_4961),
.Y(n_6201)
);

AND2x2_ASAP7_75t_L g6202 ( 
.A(n_5644),
.B(n_5275),
.Y(n_6202)
);

AND2x2_ASAP7_75t_L g6203 ( 
.A(n_5806),
.B(n_5450),
.Y(n_6203)
);

INVx3_ASAP7_75t_L g6204 ( 
.A(n_5704),
.Y(n_6204)
);

INVx1_ASAP7_75t_L g6205 ( 
.A(n_5732),
.Y(n_6205)
);

AOI221xp5_ASAP7_75t_L g6206 ( 
.A1(n_5732),
.A2(n_5597),
.B1(n_5596),
.B2(n_5588),
.C(n_5538),
.Y(n_6206)
);

OAI221xp5_ASAP7_75t_L g6207 ( 
.A1(n_5606),
.A2(n_5320),
.B1(n_5251),
.B2(n_4461),
.C(n_5527),
.Y(n_6207)
);

AOI22xp33_ASAP7_75t_L g6208 ( 
.A1(n_5611),
.A2(n_5545),
.B1(n_5544),
.B2(n_5531),
.Y(n_6208)
);

INVx5_ASAP7_75t_L g6209 ( 
.A(n_5920),
.Y(n_6209)
);

OAI21xp33_ASAP7_75t_L g6210 ( 
.A1(n_5786),
.A2(n_5520),
.B(n_5329),
.Y(n_6210)
);

OR2x2_ASAP7_75t_L g6211 ( 
.A(n_5740),
.B(n_5587),
.Y(n_6211)
);

INVx1_ASAP7_75t_L g6212 ( 
.A(n_5734),
.Y(n_6212)
);

HB1xp67_ASAP7_75t_L g6213 ( 
.A(n_5729),
.Y(n_6213)
);

AOI22xp33_ASAP7_75t_SL g6214 ( 
.A1(n_5691),
.A2(n_4416),
.B1(n_5270),
.B2(n_4500),
.Y(n_6214)
);

OAI31xp33_ASAP7_75t_L g6215 ( 
.A1(n_5691),
.A2(n_5745),
.A3(n_5759),
.B(n_5704),
.Y(n_6215)
);

OAI221xp5_ASAP7_75t_L g6216 ( 
.A1(n_5869),
.A2(n_5547),
.B1(n_5545),
.B2(n_5544),
.C(n_5444),
.Y(n_6216)
);

OAI211xp5_ASAP7_75t_L g6217 ( 
.A1(n_5614),
.A2(n_5618),
.B(n_5688),
.C(n_5650),
.Y(n_6217)
);

AOI22xp33_ASAP7_75t_L g6218 ( 
.A1(n_5624),
.A2(n_5547),
.B1(n_5544),
.B2(n_5437),
.Y(n_6218)
);

NAND4xp25_ASAP7_75t_L g6219 ( 
.A(n_5888),
.B(n_5525),
.C(n_5553),
.D(n_5541),
.Y(n_6219)
);

AO21x2_ASAP7_75t_L g6220 ( 
.A1(n_5887),
.A2(n_5565),
.B(n_5559),
.Y(n_6220)
);

BUFx2_ASAP7_75t_L g6221 ( 
.A(n_5617),
.Y(n_6221)
);

AND2x4_ASAP7_75t_L g6222 ( 
.A(n_5674),
.B(n_5273),
.Y(n_6222)
);

HB1xp67_ASAP7_75t_L g6223 ( 
.A(n_5686),
.Y(n_6223)
);

AOI31xp33_ASAP7_75t_L g6224 ( 
.A1(n_5909),
.A2(n_4758),
.A3(n_4765),
.B(n_4720),
.Y(n_6224)
);

INVx1_ASAP7_75t_L g6225 ( 
.A(n_5734),
.Y(n_6225)
);

OR2x2_ASAP7_75t_L g6226 ( 
.A(n_5741),
.B(n_5496),
.Y(n_6226)
);

AOI22xp33_ASAP7_75t_L g6227 ( 
.A1(n_5638),
.A2(n_5437),
.B1(n_5444),
.B2(n_5436),
.Y(n_6227)
);

INVx2_ASAP7_75t_L g6228 ( 
.A(n_5638),
.Y(n_6228)
);

HB1xp67_ASAP7_75t_L g6229 ( 
.A(n_5695),
.Y(n_6229)
);

INVx2_ASAP7_75t_L g6230 ( 
.A(n_5653),
.Y(n_6230)
);

AOI33xp33_ASAP7_75t_L g6231 ( 
.A1(n_5743),
.A2(n_5396),
.A3(n_5389),
.B1(n_5406),
.B2(n_5405),
.B3(n_5390),
.Y(n_6231)
);

INVx2_ASAP7_75t_L g6232 ( 
.A(n_5653),
.Y(n_6232)
);

INVx1_ASAP7_75t_L g6233 ( 
.A(n_5743),
.Y(n_6233)
);

OAI22xp5_ASAP7_75t_L g6234 ( 
.A1(n_5739),
.A2(n_5838),
.B1(n_5745),
.B2(n_5759),
.Y(n_6234)
);

NAND2xp33_ASAP7_75t_R g6235 ( 
.A(n_5617),
.B(n_5488),
.Y(n_6235)
);

CKINVDCx5p33_ASAP7_75t_R g6236 ( 
.A(n_5888),
.Y(n_6236)
);

INVx1_ASAP7_75t_L g6237 ( 
.A(n_5770),
.Y(n_6237)
);

AOI22xp33_ASAP7_75t_L g6238 ( 
.A1(n_5657),
.A2(n_5437),
.B1(n_5444),
.B2(n_5436),
.Y(n_6238)
);

AOI22xp5_ASAP7_75t_L g6239 ( 
.A1(n_5704),
.A2(n_4903),
.B1(n_4500),
.B2(n_5577),
.Y(n_6239)
);

INVx2_ASAP7_75t_L g6240 ( 
.A(n_5657),
.Y(n_6240)
);

AND2x4_ASAP7_75t_L g6241 ( 
.A(n_5749),
.B(n_5273),
.Y(n_6241)
);

HB1xp67_ASAP7_75t_L g6242 ( 
.A(n_5758),
.Y(n_6242)
);

OR2x2_ASAP7_75t_L g6243 ( 
.A(n_5741),
.B(n_5707),
.Y(n_6243)
);

OAI211xp5_ASAP7_75t_SL g6244 ( 
.A1(n_5749),
.A2(n_5525),
.B(n_5553),
.C(n_5541),
.Y(n_6244)
);

OA21x2_ASAP7_75t_L g6245 ( 
.A1(n_5669),
.A2(n_5576),
.B(n_5565),
.Y(n_6245)
);

OAI22xp5_ASAP7_75t_SL g6246 ( 
.A1(n_5909),
.A2(n_4809),
.B1(n_4987),
.B2(n_4718),
.Y(n_6246)
);

OR2x2_ASAP7_75t_L g6247 ( 
.A(n_5707),
.B(n_5496),
.Y(n_6247)
);

OAI221xp5_ASAP7_75t_L g6248 ( 
.A1(n_5685),
.A2(n_5470),
.B1(n_5476),
.B2(n_5445),
.C(n_5436),
.Y(n_6248)
);

NAND2xp5_ASAP7_75t_L g6249 ( 
.A(n_5685),
.B(n_5452),
.Y(n_6249)
);

OAI31xp33_ASAP7_75t_L g6250 ( 
.A1(n_5745),
.A2(n_5470),
.A3(n_5476),
.B(n_5445),
.Y(n_6250)
);

AOI22xp33_ASAP7_75t_L g6251 ( 
.A1(n_5669),
.A2(n_5470),
.B1(n_5476),
.B2(n_5445),
.Y(n_6251)
);

OAI221xp5_ASAP7_75t_L g6252 ( 
.A1(n_5689),
.A2(n_5597),
.B1(n_5596),
.B2(n_5370),
.C(n_5381),
.Y(n_6252)
);

NAND2xp5_ASAP7_75t_L g6253 ( 
.A(n_5689),
.B(n_5766),
.Y(n_6253)
);

INVxp67_ASAP7_75t_SL g6254 ( 
.A(n_5909),
.Y(n_6254)
);

AOI211xp5_ASAP7_75t_L g6255 ( 
.A1(n_5759),
.A2(n_5577),
.B(n_5281),
.C(n_5371),
.Y(n_6255)
);

OAI22xp33_ASAP7_75t_L g6256 ( 
.A1(n_5797),
.A2(n_5137),
.B1(n_5096),
.B2(n_5058),
.Y(n_6256)
);

NAND3xp33_ASAP7_75t_L g6257 ( 
.A(n_5650),
.B(n_5489),
.C(n_5460),
.Y(n_6257)
);

INVx1_ASAP7_75t_L g6258 ( 
.A(n_5770),
.Y(n_6258)
);

AOI22xp33_ASAP7_75t_L g6259 ( 
.A1(n_5671),
.A2(n_5499),
.B1(n_5500),
.B2(n_5486),
.Y(n_6259)
);

NAND2xp5_ASAP7_75t_L g6260 ( 
.A(n_5766),
.B(n_5725),
.Y(n_6260)
);

INVx2_ASAP7_75t_L g6261 ( 
.A(n_5671),
.Y(n_6261)
);

NAND3xp33_ASAP7_75t_L g6262 ( 
.A(n_5650),
.B(n_5489),
.C(n_5460),
.Y(n_6262)
);

NOR2xp33_ASAP7_75t_R g6263 ( 
.A(n_5688),
.B(n_4730),
.Y(n_6263)
);

AND2x2_ASAP7_75t_L g6264 ( 
.A(n_5644),
.B(n_5655),
.Y(n_6264)
);

AND2x6_ASAP7_75t_SL g6265 ( 
.A(n_5617),
.B(n_4897),
.Y(n_6265)
);

OAI211xp5_ASAP7_75t_L g6266 ( 
.A1(n_5688),
.A2(n_4990),
.B(n_5586),
.C(n_5553),
.Y(n_6266)
);

AOI31xp33_ASAP7_75t_L g6267 ( 
.A1(n_5655),
.A2(n_4739),
.A3(n_4741),
.B(n_5281),
.Y(n_6267)
);

AND2x2_ASAP7_75t_L g6268 ( 
.A(n_5806),
.B(n_5450),
.Y(n_6268)
);

AND2x4_ASAP7_75t_L g6269 ( 
.A(n_5688),
.B(n_5299),
.Y(n_6269)
);

INVxp67_ASAP7_75t_SL g6270 ( 
.A(n_5656),
.Y(n_6270)
);

AO21x2_ASAP7_75t_L g6271 ( 
.A1(n_5900),
.A2(n_5576),
.B(n_5272),
.Y(n_6271)
);

INVx2_ASAP7_75t_SL g6272 ( 
.A(n_5688),
.Y(n_6272)
);

OAI221xp5_ASAP7_75t_L g6273 ( 
.A1(n_5797),
.A2(n_5597),
.B1(n_5352),
.B2(n_5381),
.C(n_5370),
.Y(n_6273)
);

AND2x2_ASAP7_75t_L g6274 ( 
.A(n_5960),
.B(n_5656),
.Y(n_6274)
);

INVx2_ASAP7_75t_SL g6275 ( 
.A(n_5999),
.Y(n_6275)
);

OR2x2_ASAP7_75t_L g6276 ( 
.A(n_5969),
.B(n_5899),
.Y(n_6276)
);

INVx2_ASAP7_75t_L g6277 ( 
.A(n_6055),
.Y(n_6277)
);

INVx1_ASAP7_75t_L g6278 ( 
.A(n_6231),
.Y(n_6278)
);

AND2x2_ASAP7_75t_SL g6279 ( 
.A(n_5986),
.B(n_5619),
.Y(n_6279)
);

INVx1_ASAP7_75t_L g6280 ( 
.A(n_6231),
.Y(n_6280)
);

INVx1_ASAP7_75t_L g6281 ( 
.A(n_5982),
.Y(n_6281)
);

OR2x2_ASAP7_75t_L g6282 ( 
.A(n_6105),
.B(n_5899),
.Y(n_6282)
);

INVx2_ASAP7_75t_L g6283 ( 
.A(n_6055),
.Y(n_6283)
);

NAND2xp5_ASAP7_75t_L g6284 ( 
.A(n_5986),
.B(n_5807),
.Y(n_6284)
);

OR2x2_ASAP7_75t_L g6285 ( 
.A(n_6109),
.B(n_5856),
.Y(n_6285)
);

AND2x4_ASAP7_75t_L g6286 ( 
.A(n_5946),
.B(n_5983),
.Y(n_6286)
);

AND2x2_ASAP7_75t_L g6287 ( 
.A(n_5960),
.B(n_5807),
.Y(n_6287)
);

AND2x4_ASAP7_75t_L g6288 ( 
.A(n_5983),
.B(n_5619),
.Y(n_6288)
);

BUFx2_ASAP7_75t_L g6289 ( 
.A(n_5999),
.Y(n_6289)
);

AND2x4_ASAP7_75t_L g6290 ( 
.A(n_6039),
.B(n_5619),
.Y(n_6290)
);

INVx3_ASAP7_75t_L g6291 ( 
.A(n_6271),
.Y(n_6291)
);

AND2x2_ASAP7_75t_L g6292 ( 
.A(n_5994),
.B(n_5904),
.Y(n_6292)
);

HB1xp67_ASAP7_75t_L g6293 ( 
.A(n_5994),
.Y(n_6293)
);

NOR2xp33_ASAP7_75t_L g6294 ( 
.A(n_6030),
.B(n_5198),
.Y(n_6294)
);

INVx2_ASAP7_75t_L g6295 ( 
.A(n_6271),
.Y(n_6295)
);

AND2x2_ASAP7_75t_L g6296 ( 
.A(n_5992),
.B(n_5904),
.Y(n_6296)
);

AND2x2_ASAP7_75t_L g6297 ( 
.A(n_5992),
.B(n_5947),
.Y(n_6297)
);

AND2x2_ASAP7_75t_L g6298 ( 
.A(n_6068),
.B(n_6095),
.Y(n_6298)
);

INVx1_ASAP7_75t_L g6299 ( 
.A(n_6081),
.Y(n_6299)
);

INVx1_ASAP7_75t_L g6300 ( 
.A(n_5955),
.Y(n_6300)
);

NAND3xp33_ASAP7_75t_L g6301 ( 
.A(n_6032),
.B(n_5664),
.C(n_5627),
.Y(n_6301)
);

AND2x2_ASAP7_75t_L g6302 ( 
.A(n_5943),
.B(n_5808),
.Y(n_6302)
);

INVx1_ASAP7_75t_L g6303 ( 
.A(n_5970),
.Y(n_6303)
);

NAND2xp5_ASAP7_75t_L g6304 ( 
.A(n_5991),
.B(n_5856),
.Y(n_6304)
);

INVx2_ASAP7_75t_L g6305 ( 
.A(n_6013),
.Y(n_6305)
);

NAND2xp5_ASAP7_75t_L g6306 ( 
.A(n_6127),
.B(n_5725),
.Y(n_6306)
);

INVx1_ASAP7_75t_L g6307 ( 
.A(n_5984),
.Y(n_6307)
);

AND2x4_ASAP7_75t_L g6308 ( 
.A(n_6039),
.B(n_5627),
.Y(n_6308)
);

INVx2_ASAP7_75t_L g6309 ( 
.A(n_6013),
.Y(n_6309)
);

INVxp67_ASAP7_75t_SL g6310 ( 
.A(n_5979),
.Y(n_6310)
);

INVx1_ASAP7_75t_L g6311 ( 
.A(n_6150),
.Y(n_6311)
);

AND2x2_ASAP7_75t_L g6312 ( 
.A(n_5943),
.B(n_5808),
.Y(n_6312)
);

INVx1_ASAP7_75t_L g6313 ( 
.A(n_6211),
.Y(n_6313)
);

INVx2_ASAP7_75t_L g6314 ( 
.A(n_6013),
.Y(n_6314)
);

INVx1_ASAP7_75t_L g6315 ( 
.A(n_5942),
.Y(n_6315)
);

AND2x2_ASAP7_75t_L g6316 ( 
.A(n_6084),
.B(n_5822),
.Y(n_6316)
);

INVx2_ASAP7_75t_SL g6317 ( 
.A(n_6013),
.Y(n_6317)
);

INVx1_ASAP7_75t_L g6318 ( 
.A(n_6243),
.Y(n_6318)
);

AND2x2_ASAP7_75t_L g6319 ( 
.A(n_6119),
.B(n_6176),
.Y(n_6319)
);

INVx1_ASAP7_75t_L g6320 ( 
.A(n_6052),
.Y(n_6320)
);

BUFx3_ASAP7_75t_L g6321 ( 
.A(n_6030),
.Y(n_6321)
);

AND2x2_ASAP7_75t_L g6322 ( 
.A(n_6181),
.B(n_5822),
.Y(n_6322)
);

AND2x2_ASAP7_75t_L g6323 ( 
.A(n_6183),
.B(n_5828),
.Y(n_6323)
);

INVx1_ASAP7_75t_L g6324 ( 
.A(n_6052),
.Y(n_6324)
);

AND2x2_ASAP7_75t_L g6325 ( 
.A(n_6190),
.B(n_5828),
.Y(n_6325)
);

INVx2_ASAP7_75t_L g6326 ( 
.A(n_6059),
.Y(n_6326)
);

NOR2x1_ASAP7_75t_L g6327 ( 
.A(n_5951),
.B(n_5627),
.Y(n_6327)
);

AND2x2_ASAP7_75t_L g6328 ( 
.A(n_6038),
.B(n_5830),
.Y(n_6328)
);

NAND2xp5_ASAP7_75t_L g6329 ( 
.A(n_6037),
.B(n_5891),
.Y(n_6329)
);

AND2x2_ASAP7_75t_L g6330 ( 
.A(n_6038),
.B(n_5830),
.Y(n_6330)
);

AND2x2_ASAP7_75t_L g6331 ( 
.A(n_6000),
.B(n_5664),
.Y(n_6331)
);

NAND2xp5_ASAP7_75t_L g6332 ( 
.A(n_6033),
.B(n_5891),
.Y(n_6332)
);

INVx2_ASAP7_75t_L g6333 ( 
.A(n_6059),
.Y(n_6333)
);

INVx1_ASAP7_75t_L g6334 ( 
.A(n_5954),
.Y(n_6334)
);

NAND2xp5_ASAP7_75t_L g6335 ( 
.A(n_5959),
.B(n_5816),
.Y(n_6335)
);

INVx2_ASAP7_75t_L g6336 ( 
.A(n_6059),
.Y(n_6336)
);

INVx2_ASAP7_75t_L g6337 ( 
.A(n_6034),
.Y(n_6337)
);

INVx2_ASAP7_75t_L g6338 ( 
.A(n_6034),
.Y(n_6338)
);

OR2x2_ASAP7_75t_L g6339 ( 
.A(n_6247),
.B(n_5816),
.Y(n_6339)
);

INVx1_ASAP7_75t_L g6340 ( 
.A(n_5956),
.Y(n_6340)
);

OR2x2_ASAP7_75t_L g6341 ( 
.A(n_6226),
.B(n_5852),
.Y(n_6341)
);

NAND2xp5_ASAP7_75t_L g6342 ( 
.A(n_6000),
.B(n_5852),
.Y(n_6342)
);

HB1xp67_ASAP7_75t_L g6343 ( 
.A(n_5958),
.Y(n_6343)
);

AND2x2_ASAP7_75t_L g6344 ( 
.A(n_6000),
.B(n_5664),
.Y(n_6344)
);

AND2x2_ASAP7_75t_L g6345 ( 
.A(n_6065),
.B(n_5747),
.Y(n_6345)
);

AND2x4_ASAP7_75t_L g6346 ( 
.A(n_6204),
.B(n_5882),
.Y(n_6346)
);

INVx1_ASAP7_75t_L g6347 ( 
.A(n_5957),
.Y(n_6347)
);

INVx1_ASAP7_75t_L g6348 ( 
.A(n_5976),
.Y(n_6348)
);

INVx3_ASAP7_75t_L g6349 ( 
.A(n_6053),
.Y(n_6349)
);

INVx2_ASAP7_75t_L g6350 ( 
.A(n_6034),
.Y(n_6350)
);

AND2x2_ASAP7_75t_L g6351 ( 
.A(n_6065),
.B(n_5747),
.Y(n_6351)
);

INVx3_ASAP7_75t_L g6352 ( 
.A(n_6053),
.Y(n_6352)
);

NAND2xp5_ASAP7_75t_L g6353 ( 
.A(n_6021),
.B(n_5884),
.Y(n_6353)
);

AND2x2_ASAP7_75t_L g6354 ( 
.A(n_6196),
.B(n_5751),
.Y(n_6354)
);

AND2x2_ASAP7_75t_L g6355 ( 
.A(n_6196),
.B(n_5751),
.Y(n_6355)
);

AND2x2_ASAP7_75t_L g6356 ( 
.A(n_6196),
.B(n_5738),
.Y(n_6356)
);

AND2x2_ASAP7_75t_L g6357 ( 
.A(n_6011),
.B(n_5738),
.Y(n_6357)
);

INVx2_ASAP7_75t_L g6358 ( 
.A(n_5951),
.Y(n_6358)
);

INVx1_ASAP7_75t_SL g6359 ( 
.A(n_6043),
.Y(n_6359)
);

AND2x2_ASAP7_75t_L g6360 ( 
.A(n_6011),
.B(n_5744),
.Y(n_6360)
);

AND2x2_ASAP7_75t_L g6361 ( 
.A(n_6011),
.B(n_5744),
.Y(n_6361)
);

AND2x2_ASAP7_75t_L g6362 ( 
.A(n_6203),
.B(n_5884),
.Y(n_6362)
);

AND2x2_ASAP7_75t_L g6363 ( 
.A(n_6268),
.B(n_5893),
.Y(n_6363)
);

INVx2_ASAP7_75t_L g6364 ( 
.A(n_5951),
.Y(n_6364)
);

INVx1_ASAP7_75t_SL g6365 ( 
.A(n_6043),
.Y(n_6365)
);

INVx1_ASAP7_75t_L g6366 ( 
.A(n_5980),
.Y(n_6366)
);

AND2x2_ASAP7_75t_L g6367 ( 
.A(n_6145),
.B(n_5893),
.Y(n_6367)
);

NAND2xp5_ASAP7_75t_L g6368 ( 
.A(n_6031),
.B(n_5631),
.Y(n_6368)
);

INVx2_ASAP7_75t_L g6369 ( 
.A(n_6220),
.Y(n_6369)
);

AND2x2_ASAP7_75t_L g6370 ( 
.A(n_5966),
.B(n_5940),
.Y(n_6370)
);

HB1xp67_ASAP7_75t_L g6371 ( 
.A(n_5977),
.Y(n_6371)
);

AND2x4_ASAP7_75t_L g6372 ( 
.A(n_6204),
.B(n_6035),
.Y(n_6372)
);

INVx2_ASAP7_75t_L g6373 ( 
.A(n_6220),
.Y(n_6373)
);

INVx1_ASAP7_75t_L g6374 ( 
.A(n_5998),
.Y(n_6374)
);

AND2x4_ASAP7_75t_L g6375 ( 
.A(n_6204),
.B(n_5882),
.Y(n_6375)
);

NAND2xp5_ASAP7_75t_L g6376 ( 
.A(n_6031),
.B(n_5636),
.Y(n_6376)
);

HB1xp67_ASAP7_75t_L g6377 ( 
.A(n_6041),
.Y(n_6377)
);

INVx2_ASAP7_75t_L g6378 ( 
.A(n_6066),
.Y(n_6378)
);

AND2x2_ASAP7_75t_L g6379 ( 
.A(n_6175),
.B(n_5940),
.Y(n_6379)
);

INVx1_ASAP7_75t_L g6380 ( 
.A(n_6010),
.Y(n_6380)
);

BUFx2_ASAP7_75t_L g6381 ( 
.A(n_6069),
.Y(n_6381)
);

INVx1_ASAP7_75t_L g6382 ( 
.A(n_6018),
.Y(n_6382)
);

NOR2xp67_ASAP7_75t_L g6383 ( 
.A(n_6209),
.B(n_5882),
.Y(n_6383)
);

INVx1_ASAP7_75t_L g6384 ( 
.A(n_6020),
.Y(n_6384)
);

INVx2_ASAP7_75t_L g6385 ( 
.A(n_6066),
.Y(n_6385)
);

AND2x2_ASAP7_75t_L g6386 ( 
.A(n_5961),
.B(n_5897),
.Y(n_6386)
);

INVx1_ASAP7_75t_L g6387 ( 
.A(n_6022),
.Y(n_6387)
);

INVx1_ASAP7_75t_L g6388 ( 
.A(n_6042),
.Y(n_6388)
);

AND2x2_ASAP7_75t_L g6389 ( 
.A(n_5961),
.B(n_5897),
.Y(n_6389)
);

INVx2_ASAP7_75t_L g6390 ( 
.A(n_5942),
.Y(n_6390)
);

INVx2_ASAP7_75t_SL g6391 ( 
.A(n_6269),
.Y(n_6391)
);

AND2x2_ASAP7_75t_L g6392 ( 
.A(n_5961),
.B(n_5623),
.Y(n_6392)
);

INVx1_ASAP7_75t_L g6393 ( 
.A(n_6045),
.Y(n_6393)
);

INVx2_ASAP7_75t_L g6394 ( 
.A(n_5950),
.Y(n_6394)
);

NAND4xp25_ASAP7_75t_L g6395 ( 
.A(n_6129),
.B(n_5623),
.C(n_5632),
.D(n_5628),
.Y(n_6395)
);

AND2x2_ASAP7_75t_L g6396 ( 
.A(n_6054),
.B(n_5632),
.Y(n_6396)
);

INVx3_ASAP7_75t_L g6397 ( 
.A(n_6269),
.Y(n_6397)
);

AND2x2_ASAP7_75t_L g6398 ( 
.A(n_6058),
.B(n_5902),
.Y(n_6398)
);

OR2x2_ASAP7_75t_L g6399 ( 
.A(n_6005),
.B(n_5642),
.Y(n_6399)
);

AND2x2_ASAP7_75t_L g6400 ( 
.A(n_6023),
.B(n_5902),
.Y(n_6400)
);

INVx1_ASAP7_75t_L g6401 ( 
.A(n_6056),
.Y(n_6401)
);

AND2x2_ASAP7_75t_L g6402 ( 
.A(n_6025),
.B(n_5929),
.Y(n_6402)
);

INVx1_ASAP7_75t_L g6403 ( 
.A(n_6060),
.Y(n_6403)
);

INVx1_ASAP7_75t_L g6404 ( 
.A(n_6079),
.Y(n_6404)
);

AND2x2_ASAP7_75t_L g6405 ( 
.A(n_6096),
.B(n_5929),
.Y(n_6405)
);

AND2x2_ASAP7_75t_L g6406 ( 
.A(n_6269),
.B(n_5939),
.Y(n_6406)
);

AND2x2_ASAP7_75t_L g6407 ( 
.A(n_6035),
.B(n_5939),
.Y(n_6407)
);

HB1xp67_ASAP7_75t_L g6408 ( 
.A(n_6041),
.Y(n_6408)
);

NOR2xp67_ASAP7_75t_L g6409 ( 
.A(n_6209),
.B(n_5939),
.Y(n_6409)
);

INVx1_ASAP7_75t_L g6410 ( 
.A(n_6086),
.Y(n_6410)
);

AND2x2_ASAP7_75t_L g6411 ( 
.A(n_6035),
.B(n_5628),
.Y(n_6411)
);

INVx1_ASAP7_75t_L g6412 ( 
.A(n_6092),
.Y(n_6412)
);

NAND2xp5_ASAP7_75t_L g6413 ( 
.A(n_6046),
.B(n_5645),
.Y(n_6413)
);

INVx1_ASAP7_75t_L g6414 ( 
.A(n_6103),
.Y(n_6414)
);

INVx2_ASAP7_75t_L g6415 ( 
.A(n_5950),
.Y(n_6415)
);

NAND2xp5_ASAP7_75t_L g6416 ( 
.A(n_6046),
.B(n_5658),
.Y(n_6416)
);

BUFx3_ASAP7_75t_L g6417 ( 
.A(n_6061),
.Y(n_6417)
);

INVx1_ASAP7_75t_L g6418 ( 
.A(n_6117),
.Y(n_6418)
);

INVx1_ASAP7_75t_SL g6419 ( 
.A(n_6069),
.Y(n_6419)
);

INVx1_ASAP7_75t_L g6420 ( 
.A(n_6118),
.Y(n_6420)
);

NAND2xp5_ASAP7_75t_L g6421 ( 
.A(n_5945),
.B(n_5662),
.Y(n_6421)
);

INVx2_ASAP7_75t_SL g6422 ( 
.A(n_6094),
.Y(n_6422)
);

INVxp67_ASAP7_75t_L g6423 ( 
.A(n_6080),
.Y(n_6423)
);

AND2x2_ASAP7_75t_L g6424 ( 
.A(n_6264),
.B(n_6097),
.Y(n_6424)
);

NOR2xp33_ASAP7_75t_L g6425 ( 
.A(n_6267),
.B(n_5198),
.Y(n_6425)
);

INVx1_ASAP7_75t_L g6426 ( 
.A(n_5965),
.Y(n_6426)
);

INVx2_ASAP7_75t_L g6427 ( 
.A(n_5965),
.Y(n_6427)
);

INVx1_ASAP7_75t_L g6428 ( 
.A(n_6126),
.Y(n_6428)
);

AND2x2_ASAP7_75t_L g6429 ( 
.A(n_6264),
.B(n_5835),
.Y(n_6429)
);

INVx1_ASAP7_75t_L g6430 ( 
.A(n_5972),
.Y(n_6430)
);

NAND2xp5_ASAP7_75t_L g6431 ( 
.A(n_6136),
.B(n_5672),
.Y(n_6431)
);

INVx1_ASAP7_75t_L g6432 ( 
.A(n_5972),
.Y(n_6432)
);

OR2x2_ASAP7_75t_L g6433 ( 
.A(n_6260),
.B(n_5673),
.Y(n_6433)
);

INVxp67_ASAP7_75t_L g6434 ( 
.A(n_6080),
.Y(n_6434)
);

INVx1_ASAP7_75t_L g6435 ( 
.A(n_5974),
.Y(n_6435)
);

INVx1_ASAP7_75t_L g6436 ( 
.A(n_6132),
.Y(n_6436)
);

INVxp67_ASAP7_75t_SL g6437 ( 
.A(n_6016),
.Y(n_6437)
);

AND2x2_ASAP7_75t_L g6438 ( 
.A(n_6097),
.B(n_5835),
.Y(n_6438)
);

INVx2_ASAP7_75t_L g6439 ( 
.A(n_5974),
.Y(n_6439)
);

INVx2_ASAP7_75t_L g6440 ( 
.A(n_5985),
.Y(n_6440)
);

INVx2_ASAP7_75t_SL g6441 ( 
.A(n_6094),
.Y(n_6441)
);

AOI22xp33_ASAP7_75t_L g6442 ( 
.A1(n_5944),
.A2(n_5703),
.B1(n_5705),
.B2(n_5683),
.Y(n_6442)
);

INVx1_ASAP7_75t_L g6443 ( 
.A(n_6138),
.Y(n_6443)
);

INVx1_ASAP7_75t_L g6444 ( 
.A(n_6141),
.Y(n_6444)
);

INVx1_ASAP7_75t_L g6445 ( 
.A(n_6143),
.Y(n_6445)
);

AND2x2_ASAP7_75t_L g6446 ( 
.A(n_6137),
.B(n_5841),
.Y(n_6446)
);

OR2x2_ASAP7_75t_L g6447 ( 
.A(n_6253),
.B(n_5676),
.Y(n_6447)
);

AND2x4_ASAP7_75t_L g6448 ( 
.A(n_6137),
.B(n_6160),
.Y(n_6448)
);

INVx1_ASAP7_75t_L g6449 ( 
.A(n_6149),
.Y(n_6449)
);

BUFx3_ASAP7_75t_L g6450 ( 
.A(n_6112),
.Y(n_6450)
);

NAND2xp5_ASAP7_75t_L g6451 ( 
.A(n_6148),
.B(n_5677),
.Y(n_6451)
);

OR2x2_ASAP7_75t_L g6452 ( 
.A(n_5941),
.B(n_5755),
.Y(n_6452)
);

NAND2xp5_ASAP7_75t_L g6453 ( 
.A(n_6270),
.B(n_5760),
.Y(n_6453)
);

AND2x2_ASAP7_75t_L g6454 ( 
.A(n_6137),
.B(n_5841),
.Y(n_6454)
);

AND2x2_ASAP7_75t_L g6455 ( 
.A(n_6160),
.B(n_5848),
.Y(n_6455)
);

NAND2xp5_ASAP7_75t_L g6456 ( 
.A(n_6122),
.B(n_5761),
.Y(n_6456)
);

INVx1_ASAP7_75t_L g6457 ( 
.A(n_6167),
.Y(n_6457)
);

INVx1_ASAP7_75t_L g6458 ( 
.A(n_6189),
.Y(n_6458)
);

CKINVDCx14_ASAP7_75t_R g6459 ( 
.A(n_6180),
.Y(n_6459)
);

AND2x2_ASAP7_75t_L g6460 ( 
.A(n_6160),
.B(n_5848),
.Y(n_6460)
);

INVxp67_ASAP7_75t_SL g6461 ( 
.A(n_5962),
.Y(n_6461)
);

INVx2_ASAP7_75t_L g6462 ( 
.A(n_5985),
.Y(n_6462)
);

INVx1_ASAP7_75t_L g6463 ( 
.A(n_6193),
.Y(n_6463)
);

INVx1_ASAP7_75t_L g6464 ( 
.A(n_6195),
.Y(n_6464)
);

BUFx2_ASAP7_75t_L g6465 ( 
.A(n_6180),
.Y(n_6465)
);

INVx1_ASAP7_75t_L g6466 ( 
.A(n_6205),
.Y(n_6466)
);

AND2x4_ASAP7_75t_L g6467 ( 
.A(n_6184),
.B(n_5299),
.Y(n_6467)
);

INVx1_ASAP7_75t_L g6468 ( 
.A(n_6212),
.Y(n_6468)
);

OR2x2_ASAP7_75t_L g6469 ( 
.A(n_5948),
.B(n_5762),
.Y(n_6469)
);

OR2x2_ASAP7_75t_L g6470 ( 
.A(n_6099),
.B(n_6249),
.Y(n_6470)
);

AND2x2_ASAP7_75t_L g6471 ( 
.A(n_6184),
.B(n_6221),
.Y(n_6471)
);

AND2x2_ASAP7_75t_L g6472 ( 
.A(n_6184),
.B(n_5860),
.Y(n_6472)
);

AND2x2_ASAP7_75t_L g6473 ( 
.A(n_6133),
.B(n_5860),
.Y(n_6473)
);

INVx2_ASAP7_75t_L g6474 ( 
.A(n_6245),
.Y(n_6474)
);

AND2x4_ASAP7_75t_L g6475 ( 
.A(n_6121),
.B(n_5299),
.Y(n_6475)
);

NAND2xp5_ASAP7_75t_L g6476 ( 
.A(n_6026),
.B(n_6049),
.Y(n_6476)
);

INVx1_ASAP7_75t_L g6477 ( 
.A(n_6225),
.Y(n_6477)
);

AND2x2_ASAP7_75t_L g6478 ( 
.A(n_6133),
.B(n_5861),
.Y(n_6478)
);

AND2x2_ASAP7_75t_L g6479 ( 
.A(n_6154),
.B(n_5861),
.Y(n_6479)
);

BUFx2_ASAP7_75t_SL g6480 ( 
.A(n_6209),
.Y(n_6480)
);

INVx1_ASAP7_75t_L g6481 ( 
.A(n_6233),
.Y(n_6481)
);

BUFx2_ASAP7_75t_L g6482 ( 
.A(n_6263),
.Y(n_6482)
);

OR2x2_ASAP7_75t_SL g6483 ( 
.A(n_6174),
.B(n_5304),
.Y(n_6483)
);

AND2x2_ASAP7_75t_L g6484 ( 
.A(n_6154),
.B(n_5871),
.Y(n_6484)
);

AND2x4_ASAP7_75t_L g6485 ( 
.A(n_6121),
.B(n_5299),
.Y(n_6485)
);

INVx1_ASAP7_75t_SL g6486 ( 
.A(n_6263),
.Y(n_6486)
);

NAND2xp5_ASAP7_75t_L g6487 ( 
.A(n_6026),
.B(n_5764),
.Y(n_6487)
);

OR2x2_ASAP7_75t_L g6488 ( 
.A(n_6085),
.B(n_5771),
.Y(n_6488)
);

AND2x2_ASAP7_75t_L g6489 ( 
.A(n_6164),
.B(n_5871),
.Y(n_6489)
);

OR2x2_ASAP7_75t_L g6490 ( 
.A(n_6124),
.B(n_6128),
.Y(n_6490)
);

HB1xp67_ASAP7_75t_L g6491 ( 
.A(n_6049),
.Y(n_6491)
);

AND2x4_ASAP7_75t_L g6492 ( 
.A(n_6121),
.B(n_5371),
.Y(n_6492)
);

NAND2xp5_ASAP7_75t_L g6493 ( 
.A(n_6050),
.B(n_5776),
.Y(n_6493)
);

OR2x2_ASAP7_75t_L g6494 ( 
.A(n_6185),
.B(n_6166),
.Y(n_6494)
);

BUFx2_ASAP7_75t_L g6495 ( 
.A(n_6088),
.Y(n_6495)
);

INVxp67_ASAP7_75t_L g6496 ( 
.A(n_6142),
.Y(n_6496)
);

AND2x2_ASAP7_75t_L g6497 ( 
.A(n_6164),
.B(n_5875),
.Y(n_6497)
);

INVx2_ASAP7_75t_L g6498 ( 
.A(n_6245),
.Y(n_6498)
);

INVxp67_ASAP7_75t_SL g6499 ( 
.A(n_5962),
.Y(n_6499)
);

AND2x2_ASAP7_75t_L g6500 ( 
.A(n_6202),
.B(n_6198),
.Y(n_6500)
);

AND2x2_ASAP7_75t_L g6501 ( 
.A(n_6202),
.B(n_5875),
.Y(n_6501)
);

INVx2_ASAP7_75t_L g6502 ( 
.A(n_6245),
.Y(n_6502)
);

AND2x2_ASAP7_75t_L g6503 ( 
.A(n_6198),
.B(n_5876),
.Y(n_6503)
);

INVx1_ASAP7_75t_L g6504 ( 
.A(n_6237),
.Y(n_6504)
);

INVx3_ASAP7_75t_L g6505 ( 
.A(n_6198),
.Y(n_6505)
);

AND2x2_ASAP7_75t_L g6506 ( 
.A(n_6222),
.B(n_5876),
.Y(n_6506)
);

INVx3_ASAP7_75t_L g6507 ( 
.A(n_6222),
.Y(n_6507)
);

INVx1_ASAP7_75t_L g6508 ( 
.A(n_6258),
.Y(n_6508)
);

AND2x2_ASAP7_75t_L g6509 ( 
.A(n_6222),
.B(n_6241),
.Y(n_6509)
);

NAND2xp5_ASAP7_75t_L g6510 ( 
.A(n_6050),
.B(n_5780),
.Y(n_6510)
);

INVx1_ASAP7_75t_L g6511 ( 
.A(n_6057),
.Y(n_6511)
);

AND2x2_ASAP7_75t_L g6512 ( 
.A(n_6241),
.B(n_6076),
.Y(n_6512)
);

AOI22xp33_ASAP7_75t_L g6513 ( 
.A1(n_6009),
.A2(n_5703),
.B1(n_5705),
.B2(n_5683),
.Y(n_6513)
);

BUFx2_ASAP7_75t_L g6514 ( 
.A(n_6265),
.Y(n_6514)
);

INVx2_ASAP7_75t_L g6515 ( 
.A(n_6110),
.Y(n_6515)
);

HB1xp67_ASAP7_75t_L g6516 ( 
.A(n_6076),
.Y(n_6516)
);

BUFx2_ASAP7_75t_L g6517 ( 
.A(n_6112),
.Y(n_6517)
);

AND2x2_ASAP7_75t_L g6518 ( 
.A(n_6241),
.B(n_6077),
.Y(n_6518)
);

INVx2_ASAP7_75t_L g6519 ( 
.A(n_6110),
.Y(n_6519)
);

AND2x4_ASAP7_75t_L g6520 ( 
.A(n_6077),
.B(n_5371),
.Y(n_6520)
);

AND2x2_ASAP7_75t_L g6521 ( 
.A(n_6082),
.B(n_5878),
.Y(n_6521)
);

NOR2xp33_ASAP7_75t_L g6522 ( 
.A(n_6165),
.B(n_5198),
.Y(n_6522)
);

AND2x2_ASAP7_75t_L g6523 ( 
.A(n_6082),
.B(n_5878),
.Y(n_6523)
);

AND2x2_ASAP7_75t_L g6524 ( 
.A(n_6108),
.B(n_5491),
.Y(n_6524)
);

AND2x4_ASAP7_75t_SL g6525 ( 
.A(n_6165),
.B(n_6142),
.Y(n_6525)
);

INVx2_ASAP7_75t_L g6526 ( 
.A(n_6110),
.Y(n_6526)
);

NAND2xp5_ASAP7_75t_L g6527 ( 
.A(n_6108),
.B(n_5788),
.Y(n_6527)
);

AND2x2_ASAP7_75t_L g6528 ( 
.A(n_6120),
.B(n_5491),
.Y(n_6528)
);

AND2x2_ASAP7_75t_L g6529 ( 
.A(n_6120),
.B(n_5543),
.Y(n_6529)
);

INVx1_ASAP7_75t_L g6530 ( 
.A(n_6057),
.Y(n_6530)
);

AND2x2_ASAP7_75t_L g6531 ( 
.A(n_6125),
.B(n_5543),
.Y(n_6531)
);

AND2x2_ASAP7_75t_L g6532 ( 
.A(n_6125),
.B(n_5277),
.Y(n_6532)
);

NAND2xp5_ASAP7_75t_L g6533 ( 
.A(n_6070),
.B(n_5792),
.Y(n_6533)
);

INVx2_ASAP7_75t_L g6534 ( 
.A(n_6094),
.Y(n_6534)
);

INVx1_ASAP7_75t_L g6535 ( 
.A(n_6090),
.Y(n_6535)
);

AND2x2_ASAP7_75t_L g6536 ( 
.A(n_6201),
.B(n_5277),
.Y(n_6536)
);

INVx3_ASAP7_75t_L g6537 ( 
.A(n_6152),
.Y(n_6537)
);

INVx1_ASAP7_75t_L g6538 ( 
.A(n_6090),
.Y(n_6538)
);

AND2x4_ASAP7_75t_L g6539 ( 
.A(n_6152),
.B(n_5371),
.Y(n_6539)
);

NAND2xp5_ASAP7_75t_L g6540 ( 
.A(n_6229),
.B(n_6223),
.Y(n_6540)
);

INVx3_ASAP7_75t_L g6541 ( 
.A(n_6153),
.Y(n_6541)
);

OR2x2_ASAP7_75t_L g6542 ( 
.A(n_5988),
.B(n_5796),
.Y(n_6542)
);

BUFx3_ASAP7_75t_L g6543 ( 
.A(n_6209),
.Y(n_6543)
);

AND2x2_ASAP7_75t_L g6544 ( 
.A(n_6051),
.B(n_5546),
.Y(n_6544)
);

AND2x2_ASAP7_75t_SL g6545 ( 
.A(n_6063),
.B(n_4862),
.Y(n_6545)
);

NAND2xp5_ASAP7_75t_L g6546 ( 
.A(n_6213),
.B(n_5799),
.Y(n_6546)
);

AND2x2_ASAP7_75t_L g6547 ( 
.A(n_6171),
.B(n_5546),
.Y(n_6547)
);

INVx2_ASAP7_75t_L g6548 ( 
.A(n_5975),
.Y(n_6548)
);

AND2x4_ASAP7_75t_L g6549 ( 
.A(n_6153),
.B(n_5402),
.Y(n_6549)
);

AND2x2_ASAP7_75t_L g6550 ( 
.A(n_6171),
.B(n_5561),
.Y(n_6550)
);

NAND2xp5_ASAP7_75t_L g6551 ( 
.A(n_6155),
.B(n_5811),
.Y(n_6551)
);

NAND2xp5_ASAP7_75t_L g6552 ( 
.A(n_6242),
.B(n_5812),
.Y(n_6552)
);

INVx1_ASAP7_75t_L g6553 ( 
.A(n_6090),
.Y(n_6553)
);

INVx1_ASAP7_75t_L g6554 ( 
.A(n_5989),
.Y(n_6554)
);

INVxp33_ASAP7_75t_L g6555 ( 
.A(n_6246),
.Y(n_6555)
);

BUFx2_ASAP7_75t_L g6556 ( 
.A(n_6015),
.Y(n_6556)
);

AND2x2_ASAP7_75t_L g6557 ( 
.A(n_6191),
.B(n_5561),
.Y(n_6557)
);

AND2x2_ASAP7_75t_L g6558 ( 
.A(n_6191),
.B(n_5564),
.Y(n_6558)
);

AND2x2_ASAP7_75t_L g6559 ( 
.A(n_6113),
.B(n_5564),
.Y(n_6559)
);

INVx2_ASAP7_75t_L g6560 ( 
.A(n_5975),
.Y(n_6560)
);

NAND2xp5_ASAP7_75t_L g6561 ( 
.A(n_6287),
.B(n_5988),
.Y(n_6561)
);

AND2x2_ASAP7_75t_L g6562 ( 
.A(n_6287),
.B(n_6165),
.Y(n_6562)
);

INVx1_ASAP7_75t_L g6563 ( 
.A(n_6516),
.Y(n_6563)
);

AND2x2_ASAP7_75t_L g6564 ( 
.A(n_6424),
.B(n_6297),
.Y(n_6564)
);

OR2x2_ASAP7_75t_L g6565 ( 
.A(n_6293),
.B(n_6008),
.Y(n_6565)
);

INVx2_ASAP7_75t_L g6566 ( 
.A(n_6326),
.Y(n_6566)
);

NAND2x1_ASAP7_75t_L g6567 ( 
.A(n_6505),
.B(n_6224),
.Y(n_6567)
);

AND2x2_ASAP7_75t_L g6568 ( 
.A(n_6424),
.B(n_6209),
.Y(n_6568)
);

INVx1_ASAP7_75t_L g6569 ( 
.A(n_6474),
.Y(n_6569)
);

NAND2xp5_ASAP7_75t_L g6570 ( 
.A(n_6297),
.B(n_6087),
.Y(n_6570)
);

INVxp67_ASAP7_75t_L g6571 ( 
.A(n_6289),
.Y(n_6571)
);

AND2x2_ASAP7_75t_L g6572 ( 
.A(n_6289),
.B(n_6255),
.Y(n_6572)
);

INVx1_ASAP7_75t_L g6573 ( 
.A(n_6474),
.Y(n_6573)
);

OR2x2_ASAP7_75t_L g6574 ( 
.A(n_6276),
.B(n_6282),
.Y(n_6574)
);

NAND2xp5_ASAP7_75t_L g6575 ( 
.A(n_6367),
.B(n_6098),
.Y(n_6575)
);

INVx1_ASAP7_75t_L g6576 ( 
.A(n_6498),
.Y(n_6576)
);

NAND2xp5_ASAP7_75t_L g6577 ( 
.A(n_6367),
.B(n_5968),
.Y(n_6577)
);

AND2x2_ASAP7_75t_L g6578 ( 
.A(n_6302),
.B(n_6215),
.Y(n_6578)
);

AND2x4_ASAP7_75t_SL g6579 ( 
.A(n_6448),
.B(n_6074),
.Y(n_6579)
);

INVx1_ASAP7_75t_L g6580 ( 
.A(n_6498),
.Y(n_6580)
);

NAND2xp5_ASAP7_75t_L g6581 ( 
.A(n_6302),
.B(n_6017),
.Y(n_6581)
);

INVx1_ASAP7_75t_L g6582 ( 
.A(n_6502),
.Y(n_6582)
);

INVx1_ASAP7_75t_L g6583 ( 
.A(n_6502),
.Y(n_6583)
);

NAND2xp5_ASAP7_75t_L g6584 ( 
.A(n_6312),
.B(n_6177),
.Y(n_6584)
);

INVx2_ASAP7_75t_SL g6585 ( 
.A(n_6509),
.Y(n_6585)
);

INVx2_ASAP7_75t_L g6586 ( 
.A(n_6326),
.Y(n_6586)
);

OAI22xp5_ASAP7_75t_L g6587 ( 
.A1(n_6483),
.A2(n_6001),
.B1(n_5995),
.B2(n_5967),
.Y(n_6587)
);

OR2x2_ASAP7_75t_L g6588 ( 
.A(n_6276),
.B(n_6177),
.Y(n_6588)
);

INVx1_ASAP7_75t_L g6589 ( 
.A(n_6333),
.Y(n_6589)
);

OR2x2_ASAP7_75t_L g6590 ( 
.A(n_6282),
.B(n_6028),
.Y(n_6590)
);

AND2x2_ASAP7_75t_L g6591 ( 
.A(n_6312),
.B(n_6236),
.Y(n_6591)
);

NAND2xp5_ASAP7_75t_L g6592 ( 
.A(n_6328),
.B(n_6330),
.Y(n_6592)
);

INVx1_ASAP7_75t_L g6593 ( 
.A(n_6333),
.Y(n_6593)
);

INVx4_ASAP7_75t_L g6594 ( 
.A(n_6321),
.Y(n_6594)
);

OR2x6_ASAP7_75t_L g6595 ( 
.A(n_6378),
.B(n_6012),
.Y(n_6595)
);

OR3x2_ASAP7_75t_L g6596 ( 
.A(n_6399),
.B(n_6219),
.C(n_6161),
.Y(n_6596)
);

INVx1_ASAP7_75t_L g6597 ( 
.A(n_6336),
.Y(n_6597)
);

INVx1_ASAP7_75t_L g6598 ( 
.A(n_6336),
.Y(n_6598)
);

INVx1_ASAP7_75t_L g6599 ( 
.A(n_6535),
.Y(n_6599)
);

AND2x2_ASAP7_75t_L g6600 ( 
.A(n_6274),
.B(n_6236),
.Y(n_6600)
);

OR2x2_ASAP7_75t_L g6601 ( 
.A(n_6285),
.B(n_6192),
.Y(n_6601)
);

OR2x2_ASAP7_75t_L g6602 ( 
.A(n_6285),
.B(n_6339),
.Y(n_6602)
);

NAND2xp5_ASAP7_75t_L g6603 ( 
.A(n_6328),
.B(n_5964),
.Y(n_6603)
);

OR2x2_ASAP7_75t_L g6604 ( 
.A(n_6339),
.B(n_6083),
.Y(n_6604)
);

HB1xp67_ASAP7_75t_L g6605 ( 
.A(n_6291),
.Y(n_6605)
);

AND2x2_ASAP7_75t_L g6606 ( 
.A(n_6274),
.B(n_6234),
.Y(n_6606)
);

INVx1_ASAP7_75t_SL g6607 ( 
.A(n_6381),
.Y(n_6607)
);

INVx1_ASAP7_75t_L g6608 ( 
.A(n_6535),
.Y(n_6608)
);

NAND2xp5_ASAP7_75t_SL g6609 ( 
.A(n_6291),
.B(n_6007),
.Y(n_6609)
);

NOR2x1_ASAP7_75t_SL g6610 ( 
.A(n_6480),
.B(n_6217),
.Y(n_6610)
);

AND2x2_ASAP7_75t_L g6611 ( 
.A(n_6330),
.B(n_6272),
.Y(n_6611)
);

NAND2xp5_ASAP7_75t_L g6612 ( 
.A(n_6438),
.B(n_6210),
.Y(n_6612)
);

AND2x2_ASAP7_75t_L g6613 ( 
.A(n_6292),
.B(n_6272),
.Y(n_6613)
);

INVx2_ASAP7_75t_L g6614 ( 
.A(n_6291),
.Y(n_6614)
);

INVx1_ASAP7_75t_L g6615 ( 
.A(n_6538),
.Y(n_6615)
);

INVx1_ASAP7_75t_L g6616 ( 
.A(n_6538),
.Y(n_6616)
);

AND2x2_ASAP7_75t_L g6617 ( 
.A(n_6292),
.B(n_6106),
.Y(n_6617)
);

INVx1_ASAP7_75t_L g6618 ( 
.A(n_6553),
.Y(n_6618)
);

OA21x2_ASAP7_75t_L g6619 ( 
.A1(n_6277),
.A2(n_5989),
.B(n_5993),
.Y(n_6619)
);

AND2x2_ASAP7_75t_L g6620 ( 
.A(n_6438),
.B(n_6104),
.Y(n_6620)
);

NAND2xp5_ASAP7_75t_L g6621 ( 
.A(n_6298),
.B(n_5952),
.Y(n_6621)
);

AND2x4_ASAP7_75t_L g6622 ( 
.A(n_6448),
.B(n_6072),
.Y(n_6622)
);

OR2x2_ASAP7_75t_L g6623 ( 
.A(n_6341),
.B(n_6044),
.Y(n_6623)
);

NAND2xp5_ASAP7_75t_L g6624 ( 
.A(n_6298),
.B(n_6006),
.Y(n_6624)
);

AND2x2_ASAP7_75t_L g6625 ( 
.A(n_6429),
.B(n_6197),
.Y(n_6625)
);

OR2x2_ASAP7_75t_L g6626 ( 
.A(n_6341),
.B(n_6067),
.Y(n_6626)
);

INVx2_ASAP7_75t_L g6627 ( 
.A(n_6277),
.Y(n_6627)
);

AND2x2_ASAP7_75t_L g6628 ( 
.A(n_6429),
.B(n_6473),
.Y(n_6628)
);

AND2x2_ASAP7_75t_L g6629 ( 
.A(n_6473),
.B(n_6140),
.Y(n_6629)
);

AND2x2_ASAP7_75t_L g6630 ( 
.A(n_6478),
.B(n_6479),
.Y(n_6630)
);

INVx2_ASAP7_75t_L g6631 ( 
.A(n_6283),
.Y(n_6631)
);

NAND2xp5_ASAP7_75t_L g6632 ( 
.A(n_6316),
.B(n_5963),
.Y(n_6632)
);

NAND2xp5_ASAP7_75t_L g6633 ( 
.A(n_6316),
.B(n_5981),
.Y(n_6633)
);

AND2x2_ASAP7_75t_L g6634 ( 
.A(n_6478),
.B(n_6140),
.Y(n_6634)
);

INVx3_ASAP7_75t_L g6635 ( 
.A(n_6283),
.Y(n_6635)
);

INVx2_ASAP7_75t_L g6636 ( 
.A(n_6553),
.Y(n_6636)
);

OR2x2_ASAP7_75t_L g6637 ( 
.A(n_6281),
.B(n_6151),
.Y(n_6637)
);

AND2x2_ASAP7_75t_L g6638 ( 
.A(n_6479),
.B(n_6147),
.Y(n_6638)
);

INVx1_ASAP7_75t_L g6639 ( 
.A(n_6377),
.Y(n_6639)
);

AND2x2_ASAP7_75t_L g6640 ( 
.A(n_6484),
.B(n_6147),
.Y(n_6640)
);

INVx1_ASAP7_75t_L g6641 ( 
.A(n_6408),
.Y(n_6641)
);

INVx2_ASAP7_75t_L g6642 ( 
.A(n_6505),
.Y(n_6642)
);

OR2x2_ASAP7_75t_L g6643 ( 
.A(n_6281),
.B(n_6318),
.Y(n_6643)
);

INVx2_ASAP7_75t_L g6644 ( 
.A(n_6505),
.Y(n_6644)
);

INVx2_ASAP7_75t_L g6645 ( 
.A(n_6507),
.Y(n_6645)
);

INVx1_ASAP7_75t_L g6646 ( 
.A(n_6491),
.Y(n_6646)
);

INVx1_ASAP7_75t_L g6647 ( 
.A(n_6343),
.Y(n_6647)
);

AND2x2_ASAP7_75t_L g6648 ( 
.A(n_6484),
.B(n_6158),
.Y(n_6648)
);

INVx2_ASAP7_75t_SL g6649 ( 
.A(n_6509),
.Y(n_6649)
);

INVx2_ASAP7_75t_L g6650 ( 
.A(n_6507),
.Y(n_6650)
);

AND2x2_ASAP7_75t_L g6651 ( 
.A(n_6489),
.B(n_5484),
.Y(n_6651)
);

INVx1_ASAP7_75t_L g6652 ( 
.A(n_6371),
.Y(n_6652)
);

INVx2_ASAP7_75t_L g6653 ( 
.A(n_6507),
.Y(n_6653)
);

OR2x2_ASAP7_75t_L g6654 ( 
.A(n_6318),
.B(n_6135),
.Y(n_6654)
);

HB1xp67_ASAP7_75t_L g6655 ( 
.A(n_6495),
.Y(n_6655)
);

AND2x2_ASAP7_75t_L g6656 ( 
.A(n_6489),
.B(n_6497),
.Y(n_6656)
);

AND2x4_ASAP7_75t_L g6657 ( 
.A(n_6448),
.B(n_6078),
.Y(n_6657)
);

AND2x2_ASAP7_75t_L g6658 ( 
.A(n_6497),
.B(n_5484),
.Y(n_6658)
);

AND2x4_ASAP7_75t_L g6659 ( 
.A(n_6500),
.B(n_6158),
.Y(n_6659)
);

NAND2xp33_ASAP7_75t_R g6660 ( 
.A(n_6495),
.B(n_6014),
.Y(n_6660)
);

INVx1_ASAP7_75t_L g6661 ( 
.A(n_6417),
.Y(n_6661)
);

BUFx2_ASAP7_75t_L g6662 ( 
.A(n_6381),
.Y(n_6662)
);

INVx2_ASAP7_75t_L g6663 ( 
.A(n_6295),
.Y(n_6663)
);

INVx1_ASAP7_75t_SL g6664 ( 
.A(n_6370),
.Y(n_6664)
);

INVx2_ASAP7_75t_SL g6665 ( 
.A(n_6500),
.Y(n_6665)
);

AND2x2_ASAP7_75t_L g6666 ( 
.A(n_6501),
.B(n_5517),
.Y(n_6666)
);

AND2x2_ASAP7_75t_L g6667 ( 
.A(n_6501),
.B(n_6319),
.Y(n_6667)
);

INVx1_ASAP7_75t_L g6668 ( 
.A(n_6417),
.Y(n_6668)
);

INVx2_ASAP7_75t_L g6669 ( 
.A(n_6295),
.Y(n_6669)
);

AND2x4_ASAP7_75t_L g6670 ( 
.A(n_6372),
.B(n_5975),
.Y(n_6670)
);

INVx1_ASAP7_75t_L g6671 ( 
.A(n_6390),
.Y(n_6671)
);

INVx1_ASAP7_75t_L g6672 ( 
.A(n_6390),
.Y(n_6672)
);

NAND2xp5_ASAP7_75t_SL g6673 ( 
.A(n_6514),
.B(n_5997),
.Y(n_6673)
);

AND2x2_ASAP7_75t_L g6674 ( 
.A(n_6319),
.B(n_5517),
.Y(n_6674)
);

AND2x2_ASAP7_75t_L g6675 ( 
.A(n_6296),
.B(n_6107),
.Y(n_6675)
);

INVx1_ASAP7_75t_L g6676 ( 
.A(n_6394),
.Y(n_6676)
);

INVx1_ASAP7_75t_L g6677 ( 
.A(n_6394),
.Y(n_6677)
);

AND2x2_ASAP7_75t_L g6678 ( 
.A(n_6296),
.B(n_5566),
.Y(n_6678)
);

AND2x4_ASAP7_75t_L g6679 ( 
.A(n_6372),
.B(n_6254),
.Y(n_6679)
);

INVx1_ASAP7_75t_L g6680 ( 
.A(n_6415),
.Y(n_6680)
);

INVx1_ASAP7_75t_L g6681 ( 
.A(n_6415),
.Y(n_6681)
);

NOR2xp33_ASAP7_75t_L g6682 ( 
.A(n_6459),
.B(n_6004),
.Y(n_6682)
);

NOR2x1_ASAP7_75t_L g6683 ( 
.A(n_6465),
.B(n_6556),
.Y(n_6683)
);

NOR2x1_ASAP7_75t_L g6684 ( 
.A(n_6465),
.B(n_5949),
.Y(n_6684)
);

INVx2_ASAP7_75t_L g6685 ( 
.A(n_6483),
.Y(n_6685)
);

AND2x2_ASAP7_75t_L g6686 ( 
.A(n_6400),
.B(n_5566),
.Y(n_6686)
);

OR2x2_ASAP7_75t_L g6687 ( 
.A(n_6306),
.B(n_6540),
.Y(n_6687)
);

NAND2xp5_ASAP7_75t_L g6688 ( 
.A(n_6322),
.B(n_6027),
.Y(n_6688)
);

INVx1_ASAP7_75t_SL g6689 ( 
.A(n_6370),
.Y(n_6689)
);

INVxp67_ASAP7_75t_L g6690 ( 
.A(n_6517),
.Y(n_6690)
);

AND2x4_ASAP7_75t_SL g6691 ( 
.A(n_6286),
.B(n_5014),
.Y(n_6691)
);

INVx1_ASAP7_75t_L g6692 ( 
.A(n_6427),
.Y(n_6692)
);

AND2x2_ASAP7_75t_L g6693 ( 
.A(n_6400),
.B(n_5594),
.Y(n_6693)
);

INVxp67_ASAP7_75t_L g6694 ( 
.A(n_6517),
.Y(n_6694)
);

AND2x4_ASAP7_75t_L g6695 ( 
.A(n_6372),
.B(n_6257),
.Y(n_6695)
);

INVxp67_ASAP7_75t_SL g6696 ( 
.A(n_6423),
.Y(n_6696)
);

INVx1_ASAP7_75t_L g6697 ( 
.A(n_6427),
.Y(n_6697)
);

AND2x2_ASAP7_75t_L g6698 ( 
.A(n_6398),
.B(n_6131),
.Y(n_6698)
);

OR2x2_ASAP7_75t_L g6699 ( 
.A(n_6335),
.B(n_6329),
.Y(n_6699)
);

HB1xp67_ASAP7_75t_L g6700 ( 
.A(n_6542),
.Y(n_6700)
);

AND2x2_ASAP7_75t_L g6701 ( 
.A(n_6398),
.B(n_6131),
.Y(n_6701)
);

AND2x2_ASAP7_75t_L g6702 ( 
.A(n_6503),
.B(n_6199),
.Y(n_6702)
);

NAND2xp5_ASAP7_75t_L g6703 ( 
.A(n_6322),
.B(n_6071),
.Y(n_6703)
);

HB1xp67_ASAP7_75t_L g6704 ( 
.A(n_6542),
.Y(n_6704)
);

INVx1_ASAP7_75t_L g6705 ( 
.A(n_6439),
.Y(n_6705)
);

OR2x2_ASAP7_75t_L g6706 ( 
.A(n_6284),
.B(n_5971),
.Y(n_6706)
);

INVx2_ASAP7_75t_L g6707 ( 
.A(n_6369),
.Y(n_6707)
);

INVx2_ASAP7_75t_L g6708 ( 
.A(n_6369),
.Y(n_6708)
);

NOR2x1_ASAP7_75t_L g6709 ( 
.A(n_6556),
.B(n_5949),
.Y(n_6709)
);

AND2x2_ASAP7_75t_L g6710 ( 
.A(n_6503),
.B(n_6139),
.Y(n_6710)
);

INVx1_ASAP7_75t_L g6711 ( 
.A(n_6439),
.Y(n_6711)
);

INVx1_ASAP7_75t_L g6712 ( 
.A(n_6440),
.Y(n_6712)
);

INVx2_ASAP7_75t_L g6713 ( 
.A(n_6373),
.Y(n_6713)
);

INVx2_ASAP7_75t_L g6714 ( 
.A(n_6373),
.Y(n_6714)
);

NAND2xp5_ASAP7_75t_L g6715 ( 
.A(n_6323),
.B(n_6071),
.Y(n_6715)
);

INVx1_ASAP7_75t_L g6716 ( 
.A(n_6440),
.Y(n_6716)
);

OR2x2_ASAP7_75t_L g6717 ( 
.A(n_6311),
.B(n_6019),
.Y(n_6717)
);

INVx1_ASAP7_75t_L g6718 ( 
.A(n_6462),
.Y(n_6718)
);

INVx1_ASAP7_75t_SL g6719 ( 
.A(n_6359),
.Y(n_6719)
);

INVx3_ASAP7_75t_L g6720 ( 
.A(n_6346),
.Y(n_6720)
);

AND2x2_ASAP7_75t_L g6721 ( 
.A(n_6506),
.B(n_5594),
.Y(n_6721)
);

NAND2xp5_ASAP7_75t_L g6722 ( 
.A(n_6323),
.B(n_6100),
.Y(n_6722)
);

OAI21xp33_ASAP7_75t_L g6723 ( 
.A1(n_6278),
.A2(n_6139),
.B(n_6073),
.Y(n_6723)
);

AND2x2_ASAP7_75t_L g6724 ( 
.A(n_6506),
.B(n_5586),
.Y(n_6724)
);

NAND2xp5_ASAP7_75t_L g6725 ( 
.A(n_6325),
.B(n_6100),
.Y(n_6725)
);

O2A1O1Ixp33_ASAP7_75t_L g6726 ( 
.A1(n_6278),
.A2(n_6280),
.B(n_6399),
.C(n_6514),
.Y(n_6726)
);

NAND2xp5_ASAP7_75t_L g6727 ( 
.A(n_6325),
.B(n_5953),
.Y(n_6727)
);

AND2x2_ASAP7_75t_L g6728 ( 
.A(n_6407),
.B(n_5586),
.Y(n_6728)
);

INVx1_ASAP7_75t_L g6729 ( 
.A(n_6462),
.Y(n_6729)
);

NOR2xp67_ASAP7_75t_L g6730 ( 
.A(n_6275),
.B(n_6262),
.Y(n_6730)
);

INVx2_ASAP7_75t_L g6731 ( 
.A(n_6349),
.Y(n_6731)
);

NAND2xp5_ASAP7_75t_L g6732 ( 
.A(n_6521),
.B(n_6111),
.Y(n_6732)
);

BUFx2_ASAP7_75t_L g6733 ( 
.A(n_6467),
.Y(n_6733)
);

INVx2_ASAP7_75t_SL g6734 ( 
.A(n_6346),
.Y(n_6734)
);

NAND2xp5_ASAP7_75t_L g6735 ( 
.A(n_6521),
.B(n_6012),
.Y(n_6735)
);

AND2x4_ASAP7_75t_L g6736 ( 
.A(n_6346),
.B(n_6047),
.Y(n_6736)
);

INVx1_ASAP7_75t_L g6737 ( 
.A(n_6300),
.Y(n_6737)
);

INVxp33_ASAP7_75t_L g6738 ( 
.A(n_6286),
.Y(n_6738)
);

INVx1_ASAP7_75t_L g6739 ( 
.A(n_6300),
.Y(n_6739)
);

INVx2_ASAP7_75t_L g6740 ( 
.A(n_6349),
.Y(n_6740)
);

AND2x2_ASAP7_75t_L g6741 ( 
.A(n_6279),
.B(n_6002),
.Y(n_6741)
);

INVx1_ASAP7_75t_L g6742 ( 
.A(n_6303),
.Y(n_6742)
);

INVx1_ASAP7_75t_L g6743 ( 
.A(n_6303),
.Y(n_6743)
);

INVx1_ASAP7_75t_L g6744 ( 
.A(n_6307),
.Y(n_6744)
);

NAND2xp5_ASAP7_75t_L g6745 ( 
.A(n_6523),
.B(n_6102),
.Y(n_6745)
);

INVx1_ASAP7_75t_L g6746 ( 
.A(n_6307),
.Y(n_6746)
);

AND2x2_ASAP7_75t_L g6747 ( 
.A(n_6407),
.B(n_4843),
.Y(n_6747)
);

INVx1_ASAP7_75t_L g6748 ( 
.A(n_6332),
.Y(n_6748)
);

INVx1_ASAP7_75t_L g6749 ( 
.A(n_6523),
.Y(n_6749)
);

INVxp67_ASAP7_75t_L g6750 ( 
.A(n_6450),
.Y(n_6750)
);

INVx2_ASAP7_75t_L g6751 ( 
.A(n_6349),
.Y(n_6751)
);

AND2x4_ASAP7_75t_L g6752 ( 
.A(n_6375),
.B(n_5996),
.Y(n_6752)
);

OR2x2_ASAP7_75t_L g6753 ( 
.A(n_6313),
.B(n_6470),
.Y(n_6753)
);

NAND2xp5_ASAP7_75t_L g6754 ( 
.A(n_6362),
.B(n_6102),
.Y(n_6754)
);

NOR2xp33_ASAP7_75t_L g6755 ( 
.A(n_6365),
.B(n_5198),
.Y(n_6755)
);

NOR2xp67_ASAP7_75t_L g6756 ( 
.A(n_6275),
.B(n_6156),
.Y(n_6756)
);

NAND2xp33_ASAP7_75t_L g6757 ( 
.A(n_6490),
.B(n_6015),
.Y(n_6757)
);

INVx1_ASAP7_75t_L g6758 ( 
.A(n_6512),
.Y(n_6758)
);

OR2x2_ASAP7_75t_L g6759 ( 
.A(n_6470),
.B(n_5329),
.Y(n_6759)
);

INVx2_ASAP7_75t_L g6760 ( 
.A(n_6352),
.Y(n_6760)
);

INVx4_ASAP7_75t_L g6761 ( 
.A(n_6321),
.Y(n_6761)
);

NAND2x1p5_ASAP7_75t_L g6762 ( 
.A(n_6543),
.B(n_4832),
.Y(n_6762)
);

HB1xp67_ASAP7_75t_L g6763 ( 
.A(n_6490),
.Y(n_6763)
);

AND2x2_ASAP7_75t_L g6764 ( 
.A(n_6279),
.B(n_6471),
.Y(n_6764)
);

AND2x2_ASAP7_75t_L g6765 ( 
.A(n_6362),
.B(n_5535),
.Y(n_6765)
);

AND2x2_ASAP7_75t_L g6766 ( 
.A(n_6363),
.B(n_5535),
.Y(n_6766)
);

NAND2xp5_ASAP7_75t_L g6767 ( 
.A(n_6363),
.B(n_5993),
.Y(n_6767)
);

INVxp67_ASAP7_75t_L g6768 ( 
.A(n_6450),
.Y(n_6768)
);

NAND2xp5_ASAP7_75t_L g6769 ( 
.A(n_6544),
.B(n_6178),
.Y(n_6769)
);

AND2x2_ASAP7_75t_L g6770 ( 
.A(n_6402),
.B(n_6405),
.Y(n_6770)
);

AND2x2_ASAP7_75t_L g6771 ( 
.A(n_6402),
.B(n_6405),
.Y(n_6771)
);

INVx1_ASAP7_75t_L g6772 ( 
.A(n_6512),
.Y(n_6772)
);

INVx1_ASAP7_75t_SL g6773 ( 
.A(n_6471),
.Y(n_6773)
);

NAND2xp5_ASAP7_75t_L g6774 ( 
.A(n_6544),
.B(n_6040),
.Y(n_6774)
);

INVx1_ASAP7_75t_SL g6775 ( 
.A(n_6379),
.Y(n_6775)
);

INVxp67_ASAP7_75t_L g6776 ( 
.A(n_6310),
.Y(n_6776)
);

INVx2_ASAP7_75t_L g6777 ( 
.A(n_6352),
.Y(n_6777)
);

AND2x4_ASAP7_75t_L g6778 ( 
.A(n_6375),
.B(n_5402),
.Y(n_6778)
);

NOR2xp33_ASAP7_75t_L g6779 ( 
.A(n_6419),
.B(n_6130),
.Y(n_6779)
);

NOR2x1_ASAP7_75t_SL g6780 ( 
.A(n_6480),
.B(n_6075),
.Y(n_6780)
);

INVx1_ASAP7_75t_L g6781 ( 
.A(n_6518),
.Y(n_6781)
);

AND2x2_ASAP7_75t_L g6782 ( 
.A(n_6446),
.B(n_4802),
.Y(n_6782)
);

NAND2xp5_ASAP7_75t_L g6783 ( 
.A(n_6345),
.B(n_6003),
.Y(n_6783)
);

INVx1_ASAP7_75t_L g6784 ( 
.A(n_6518),
.Y(n_6784)
);

AND2x2_ASAP7_75t_SL g6785 ( 
.A(n_6421),
.B(n_6003),
.Y(n_6785)
);

AND2x2_ASAP7_75t_L g6786 ( 
.A(n_6446),
.B(n_5222),
.Y(n_6786)
);

AND2x2_ASAP7_75t_L g6787 ( 
.A(n_6454),
.B(n_5351),
.Y(n_6787)
);

NOR2xp67_ASAP7_75t_SL g6788 ( 
.A(n_6378),
.B(n_4990),
.Y(n_6788)
);

AND2x4_ASAP7_75t_L g6789 ( 
.A(n_6375),
.B(n_5402),
.Y(n_6789)
);

OR2x2_ASAP7_75t_L g6790 ( 
.A(n_6304),
.B(n_5498),
.Y(n_6790)
);

INVx2_ASAP7_75t_L g6791 ( 
.A(n_6352),
.Y(n_6791)
);

INVx1_ASAP7_75t_SL g6792 ( 
.A(n_6379),
.Y(n_6792)
);

INVx1_ASAP7_75t_L g6793 ( 
.A(n_6511),
.Y(n_6793)
);

AND2x2_ASAP7_75t_L g6794 ( 
.A(n_6454),
.B(n_5222),
.Y(n_6794)
);

INVx2_ASAP7_75t_L g6795 ( 
.A(n_6537),
.Y(n_6795)
);

NAND2xp5_ASAP7_75t_L g6796 ( 
.A(n_6345),
.B(n_6114),
.Y(n_6796)
);

AND2x2_ASAP7_75t_L g6797 ( 
.A(n_6455),
.B(n_5577),
.Y(n_6797)
);

NAND2xp5_ASAP7_75t_L g6798 ( 
.A(n_6351),
.B(n_6157),
.Y(n_6798)
);

AND2x2_ASAP7_75t_L g6799 ( 
.A(n_6455),
.B(n_5577),
.Y(n_6799)
);

NAND2x1_ASAP7_75t_L g6800 ( 
.A(n_6397),
.B(n_6169),
.Y(n_6800)
);

INVx1_ASAP7_75t_L g6801 ( 
.A(n_6511),
.Y(n_6801)
);

INVx1_ASAP7_75t_L g6802 ( 
.A(n_6299),
.Y(n_6802)
);

AND2x2_ASAP7_75t_L g6803 ( 
.A(n_6460),
.B(n_5351),
.Y(n_6803)
);

INVx2_ASAP7_75t_L g6804 ( 
.A(n_6537),
.Y(n_6804)
);

OR2x2_ASAP7_75t_L g6805 ( 
.A(n_6574),
.B(n_6452),
.Y(n_6805)
);

INVx1_ASAP7_75t_L g6806 ( 
.A(n_6602),
.Y(n_6806)
);

NAND2xp5_ASAP7_75t_L g6807 ( 
.A(n_6700),
.B(n_6280),
.Y(n_6807)
);

HB1xp67_ASAP7_75t_L g6808 ( 
.A(n_6564),
.Y(n_6808)
);

INVx1_ASAP7_75t_L g6809 ( 
.A(n_6662),
.Y(n_6809)
);

INVx2_ASAP7_75t_L g6810 ( 
.A(n_6720),
.Y(n_6810)
);

AND2x2_ASAP7_75t_L g6811 ( 
.A(n_6564),
.B(n_6460),
.Y(n_6811)
);

INVx1_ASAP7_75t_L g6812 ( 
.A(n_6630),
.Y(n_6812)
);

XOR2x2_ASAP7_75t_L g6813 ( 
.A(n_6587),
.B(n_6301),
.Y(n_6813)
);

INVx2_ASAP7_75t_L g6814 ( 
.A(n_6720),
.Y(n_6814)
);

INVx1_ASAP7_75t_L g6815 ( 
.A(n_6630),
.Y(n_6815)
);

NAND2xp5_ASAP7_75t_L g6816 ( 
.A(n_6700),
.B(n_6452),
.Y(n_6816)
);

INVx1_ASAP7_75t_L g6817 ( 
.A(n_6655),
.Y(n_6817)
);

INVx2_ASAP7_75t_L g6818 ( 
.A(n_6720),
.Y(n_6818)
);

AND2x2_ASAP7_75t_L g6819 ( 
.A(n_6667),
.B(n_6472),
.Y(n_6819)
);

NAND2x1p5_ASAP7_75t_L g6820 ( 
.A(n_6683),
.B(n_6543),
.Y(n_6820)
);

INVx1_ASAP7_75t_L g6821 ( 
.A(n_6655),
.Y(n_6821)
);

OR2x2_ASAP7_75t_L g6822 ( 
.A(n_6773),
.B(n_6342),
.Y(n_6822)
);

INVx1_ASAP7_75t_L g6823 ( 
.A(n_6628),
.Y(n_6823)
);

INVxp67_ASAP7_75t_L g6824 ( 
.A(n_6704),
.Y(n_6824)
);

OR2x2_ASAP7_75t_L g6825 ( 
.A(n_6607),
.B(n_6353),
.Y(n_6825)
);

NAND2xp5_ASAP7_75t_L g6826 ( 
.A(n_6704),
.B(n_6461),
.Y(n_6826)
);

INVx1_ASAP7_75t_L g6827 ( 
.A(n_6656),
.Y(n_6827)
);

OR2x2_ASAP7_75t_L g6828 ( 
.A(n_6592),
.B(n_6494),
.Y(n_6828)
);

INVx1_ASAP7_75t_L g6829 ( 
.A(n_6770),
.Y(n_6829)
);

AND2x2_ASAP7_75t_L g6830 ( 
.A(n_6771),
.B(n_6472),
.Y(n_6830)
);

NAND2xp5_ASAP7_75t_SL g6831 ( 
.A(n_6664),
.B(n_6064),
.Y(n_6831)
);

INVx1_ASAP7_75t_L g6832 ( 
.A(n_6566),
.Y(n_6832)
);

AND2x4_ASAP7_75t_L g6833 ( 
.A(n_6734),
.B(n_6286),
.Y(n_6833)
);

INVx1_ASAP7_75t_L g6834 ( 
.A(n_6566),
.Y(n_6834)
);

HB1xp67_ASAP7_75t_L g6835 ( 
.A(n_6764),
.Y(n_6835)
);

INVx2_ASAP7_75t_L g6836 ( 
.A(n_6733),
.Y(n_6836)
);

NOR2x1p5_ASAP7_75t_SL g6837 ( 
.A(n_6685),
.B(n_6515),
.Y(n_6837)
);

INVx1_ASAP7_75t_L g6838 ( 
.A(n_6586),
.Y(n_6838)
);

NAND2xp5_ASAP7_75t_L g6839 ( 
.A(n_6763),
.B(n_6499),
.Y(n_6839)
);

INVx3_ASAP7_75t_L g6840 ( 
.A(n_6778),
.Y(n_6840)
);

HB1xp67_ASAP7_75t_L g6841 ( 
.A(n_6764),
.Y(n_6841)
);

INVx1_ASAP7_75t_L g6842 ( 
.A(n_6586),
.Y(n_6842)
);

INVx1_ASAP7_75t_L g6843 ( 
.A(n_6643),
.Y(n_6843)
);

INVx1_ASAP7_75t_L g6844 ( 
.A(n_6731),
.Y(n_6844)
);

AND2x2_ASAP7_75t_L g6845 ( 
.A(n_6674),
.B(n_6351),
.Y(n_6845)
);

NAND2xp5_ASAP7_75t_L g6846 ( 
.A(n_6763),
.B(n_6609),
.Y(n_6846)
);

NAND2xp5_ASAP7_75t_L g6847 ( 
.A(n_6609),
.B(n_6320),
.Y(n_6847)
);

INVx1_ASAP7_75t_L g6848 ( 
.A(n_6731),
.Y(n_6848)
);

INVx2_ASAP7_75t_SL g6849 ( 
.A(n_6613),
.Y(n_6849)
);

NAND2xp5_ASAP7_75t_L g6850 ( 
.A(n_6685),
.B(n_6320),
.Y(n_6850)
);

INVx1_ASAP7_75t_L g6851 ( 
.A(n_6740),
.Y(n_6851)
);

NAND2xp5_ASAP7_75t_L g6852 ( 
.A(n_6589),
.B(n_6324),
.Y(n_6852)
);

INVx3_ASAP7_75t_L g6853 ( 
.A(n_6778),
.Y(n_6853)
);

AOI22xp5_ASAP7_75t_L g6854 ( 
.A1(n_6785),
.A2(n_6545),
.B1(n_6437),
.B2(n_6554),
.Y(n_6854)
);

NAND2xp5_ASAP7_75t_L g6855 ( 
.A(n_6593),
.B(n_6324),
.Y(n_6855)
);

INVx1_ASAP7_75t_L g6856 ( 
.A(n_6740),
.Y(n_6856)
);

AND2x2_ASAP7_75t_L g6857 ( 
.A(n_6678),
.B(n_6406),
.Y(n_6857)
);

AND2x4_ASAP7_75t_SL g6858 ( 
.A(n_6782),
.B(n_6288),
.Y(n_6858)
);

INVxp67_ASAP7_75t_L g6859 ( 
.A(n_6709),
.Y(n_6859)
);

NAND2xp5_ASAP7_75t_L g6860 ( 
.A(n_6597),
.B(n_6598),
.Y(n_6860)
);

INVx1_ASAP7_75t_L g6861 ( 
.A(n_6751),
.Y(n_6861)
);

INVx2_ASAP7_75t_L g6862 ( 
.A(n_6670),
.Y(n_6862)
);

OR2x2_ASAP7_75t_L g6863 ( 
.A(n_6584),
.B(n_6494),
.Y(n_6863)
);

NOR2x1_ASAP7_75t_L g6864 ( 
.A(n_6684),
.B(n_6537),
.Y(n_6864)
);

INVx1_ASAP7_75t_L g6865 ( 
.A(n_6751),
.Y(n_6865)
);

INVx1_ASAP7_75t_L g6866 ( 
.A(n_6760),
.Y(n_6866)
);

INVxp67_ASAP7_75t_L g6867 ( 
.A(n_6600),
.Y(n_6867)
);

NAND2x1_ASAP7_75t_SL g6868 ( 
.A(n_6670),
.B(n_6397),
.Y(n_6868)
);

AND2x2_ASAP7_75t_L g6869 ( 
.A(n_6686),
.B(n_6406),
.Y(n_6869)
);

INVx1_ASAP7_75t_L g6870 ( 
.A(n_6760),
.Y(n_6870)
);

AND2x2_ASAP7_75t_L g6871 ( 
.A(n_6693),
.B(n_6396),
.Y(n_6871)
);

NAND2xp33_ASAP7_75t_L g6872 ( 
.A(n_6719),
.B(n_6331),
.Y(n_6872)
);

INVx1_ASAP7_75t_SL g6873 ( 
.A(n_6689),
.Y(n_6873)
);

HB1xp67_ASAP7_75t_L g6874 ( 
.A(n_6613),
.Y(n_6874)
);

OR2x2_ASAP7_75t_L g6875 ( 
.A(n_6753),
.B(n_6433),
.Y(n_6875)
);

INVx2_ASAP7_75t_SL g6876 ( 
.A(n_6611),
.Y(n_6876)
);

NAND2xp5_ASAP7_75t_L g6877 ( 
.A(n_6785),
.B(n_6299),
.Y(n_6877)
);

OR2x2_ASAP7_75t_L g6878 ( 
.A(n_6590),
.B(n_6433),
.Y(n_6878)
);

INVx1_ASAP7_75t_L g6879 ( 
.A(n_6777),
.Y(n_6879)
);

INVx2_ASAP7_75t_L g6880 ( 
.A(n_6670),
.Y(n_6880)
);

INVx2_ASAP7_75t_L g6881 ( 
.A(n_6734),
.Y(n_6881)
);

NAND3xp33_ASAP7_75t_L g6882 ( 
.A(n_6757),
.B(n_6089),
.C(n_6434),
.Y(n_6882)
);

INVx1_ASAP7_75t_L g6883 ( 
.A(n_6777),
.Y(n_6883)
);

NAND2xp5_ASAP7_75t_L g6884 ( 
.A(n_6698),
.B(n_6337),
.Y(n_6884)
);

AND2x2_ASAP7_75t_L g6885 ( 
.A(n_6765),
.B(n_6396),
.Y(n_6885)
);

INVx1_ASAP7_75t_L g6886 ( 
.A(n_6791),
.Y(n_6886)
);

OAI21xp5_ASAP7_75t_L g6887 ( 
.A1(n_6726),
.A2(n_6545),
.B(n_6554),
.Y(n_6887)
);

INVxp67_ASAP7_75t_L g6888 ( 
.A(n_6595),
.Y(n_6888)
);

AND2x4_ASAP7_75t_L g6889 ( 
.A(n_6585),
.B(n_6288),
.Y(n_6889)
);

AND2x2_ASAP7_75t_L g6890 ( 
.A(n_6766),
.B(n_6357),
.Y(n_6890)
);

INVx2_ASAP7_75t_L g6891 ( 
.A(n_6611),
.Y(n_6891)
);

NAND2xp5_ASAP7_75t_L g6892 ( 
.A(n_6698),
.B(n_6337),
.Y(n_6892)
);

NOR2xp33_ASAP7_75t_L g6893 ( 
.A(n_6594),
.B(n_6288),
.Y(n_6893)
);

OR2x6_ASAP7_75t_L g6894 ( 
.A(n_6776),
.B(n_6385),
.Y(n_6894)
);

AND2x2_ASAP7_75t_L g6895 ( 
.A(n_6702),
.B(n_6357),
.Y(n_6895)
);

NAND2xp5_ASAP7_75t_L g6896 ( 
.A(n_6701),
.B(n_6338),
.Y(n_6896)
);

AND2x4_ASAP7_75t_L g6897 ( 
.A(n_6585),
.B(n_6290),
.Y(n_6897)
);

INVx1_ASAP7_75t_L g6898 ( 
.A(n_6791),
.Y(n_6898)
);

AOI221xp5_ASAP7_75t_L g6899 ( 
.A1(n_6723),
.A2(n_6776),
.B1(n_6673),
.B2(n_6745),
.C(n_6732),
.Y(n_6899)
);

INVx1_ASAP7_75t_L g6900 ( 
.A(n_6642),
.Y(n_6900)
);

INVx2_ASAP7_75t_L g6901 ( 
.A(n_6778),
.Y(n_6901)
);

CKINVDCx16_ASAP7_75t_R g6902 ( 
.A(n_6591),
.Y(n_6902)
);

BUFx3_ASAP7_75t_L g6903 ( 
.A(n_6568),
.Y(n_6903)
);

AND2x2_ASAP7_75t_L g6904 ( 
.A(n_6702),
.B(n_6360),
.Y(n_6904)
);

AND2x2_ASAP7_75t_L g6905 ( 
.A(n_6606),
.B(n_6360),
.Y(n_6905)
);

INVx1_ASAP7_75t_L g6906 ( 
.A(n_6642),
.Y(n_6906)
);

INVx1_ASAP7_75t_SL g6907 ( 
.A(n_6775),
.Y(n_6907)
);

HB1xp67_ASAP7_75t_L g6908 ( 
.A(n_6665),
.Y(n_6908)
);

AND2x2_ASAP7_75t_L g6909 ( 
.A(n_6792),
.B(n_6361),
.Y(n_6909)
);

HB1xp67_ASAP7_75t_L g6910 ( 
.A(n_6665),
.Y(n_6910)
);

OAI32xp33_ASAP7_75t_L g6911 ( 
.A1(n_6660),
.A2(n_6186),
.A3(n_6555),
.B1(n_5987),
.B2(n_6146),
.Y(n_6911)
);

BUFx2_ASAP7_75t_L g6912 ( 
.A(n_6789),
.Y(n_6912)
);

AND2x2_ASAP7_75t_L g6913 ( 
.A(n_6651),
.B(n_6361),
.Y(n_6913)
);

OR2x2_ASAP7_75t_L g6914 ( 
.A(n_6588),
.B(n_6561),
.Y(n_6914)
);

INVx1_ASAP7_75t_L g6915 ( 
.A(n_6644),
.Y(n_6915)
);

OR2x2_ASAP7_75t_L g6916 ( 
.A(n_6722),
.B(n_6447),
.Y(n_6916)
);

NAND2xp5_ASAP7_75t_L g6917 ( 
.A(n_6701),
.B(n_6338),
.Y(n_6917)
);

INVx1_ASAP7_75t_L g6918 ( 
.A(n_6644),
.Y(n_6918)
);

INVx1_ASAP7_75t_L g6919 ( 
.A(n_6645),
.Y(n_6919)
);

NAND2x1p5_ASAP7_75t_L g6920 ( 
.A(n_6594),
.B(n_6761),
.Y(n_6920)
);

INVx1_ASAP7_75t_L g6921 ( 
.A(n_6645),
.Y(n_6921)
);

INVx1_ASAP7_75t_L g6922 ( 
.A(n_6650),
.Y(n_6922)
);

INVxp67_ASAP7_75t_SL g6923 ( 
.A(n_6571),
.Y(n_6923)
);

INVx1_ASAP7_75t_L g6924 ( 
.A(n_6650),
.Y(n_6924)
);

INVx2_ASAP7_75t_SL g6925 ( 
.A(n_6789),
.Y(n_6925)
);

INVx1_ASAP7_75t_SL g6926 ( 
.A(n_6568),
.Y(n_6926)
);

AND2x2_ASAP7_75t_L g6927 ( 
.A(n_6658),
.B(n_6331),
.Y(n_6927)
);

NOR2xp33_ASAP7_75t_SL g6928 ( 
.A(n_6594),
.B(n_6482),
.Y(n_6928)
);

INVx1_ASAP7_75t_L g6929 ( 
.A(n_6653),
.Y(n_6929)
);

INVx1_ASAP7_75t_L g6930 ( 
.A(n_6653),
.Y(n_6930)
);

INVx1_ASAP7_75t_SL g6931 ( 
.A(n_6757),
.Y(n_6931)
);

NAND2xp5_ASAP7_75t_L g6932 ( 
.A(n_6571),
.B(n_6350),
.Y(n_6932)
);

NOR2xp33_ASAP7_75t_L g6933 ( 
.A(n_6761),
.B(n_6738),
.Y(n_6933)
);

NOR2xp33_ASAP7_75t_L g6934 ( 
.A(n_6761),
.B(n_6290),
.Y(n_6934)
);

AND2x2_ASAP7_75t_L g6935 ( 
.A(n_6666),
.B(n_6344),
.Y(n_6935)
);

INVx1_ASAP7_75t_L g6936 ( 
.A(n_6605),
.Y(n_6936)
);

INVx4_ASAP7_75t_L g6937 ( 
.A(n_6679),
.Y(n_6937)
);

INVx2_ASAP7_75t_L g6938 ( 
.A(n_6789),
.Y(n_6938)
);

INVx1_ASAP7_75t_L g6939 ( 
.A(n_6605),
.Y(n_6939)
);

OAI21xp33_ASAP7_75t_L g6940 ( 
.A1(n_6682),
.A2(n_6356),
.B(n_6547),
.Y(n_6940)
);

NAND2xp5_ASAP7_75t_L g6941 ( 
.A(n_6710),
.B(n_6350),
.Y(n_6941)
);

AND2x4_ASAP7_75t_L g6942 ( 
.A(n_6649),
.B(n_6290),
.Y(n_6942)
);

INVx1_ASAP7_75t_L g6943 ( 
.A(n_6749),
.Y(n_6943)
);

NAND2xp5_ASAP7_75t_L g6944 ( 
.A(n_6710),
.B(n_6315),
.Y(n_6944)
);

AND2x2_ASAP7_75t_L g6945 ( 
.A(n_6721),
.B(n_6344),
.Y(n_6945)
);

NAND2xp5_ASAP7_75t_L g6946 ( 
.A(n_6625),
.B(n_6426),
.Y(n_6946)
);

INVx1_ASAP7_75t_L g6947 ( 
.A(n_6758),
.Y(n_6947)
);

INVx2_ASAP7_75t_L g6948 ( 
.A(n_6695),
.Y(n_6948)
);

INVx1_ASAP7_75t_L g6949 ( 
.A(n_6772),
.Y(n_6949)
);

NAND2xp5_ASAP7_75t_L g6950 ( 
.A(n_6690),
.B(n_6430),
.Y(n_6950)
);

OR2x2_ASAP7_75t_L g6951 ( 
.A(n_6725),
.B(n_6447),
.Y(n_6951)
);

AOI22xp5_ASAP7_75t_L g6952 ( 
.A1(n_6673),
.A2(n_6442),
.B1(n_6091),
.B2(n_6513),
.Y(n_6952)
);

AND2x2_ASAP7_75t_L g6953 ( 
.A(n_6620),
.B(n_6411),
.Y(n_6953)
);

INVx1_ASAP7_75t_L g6954 ( 
.A(n_6781),
.Y(n_6954)
);

HB1xp67_ASAP7_75t_L g6955 ( 
.A(n_6629),
.Y(n_6955)
);

INVx2_ASAP7_75t_SL g6956 ( 
.A(n_6695),
.Y(n_6956)
);

NAND2xp5_ASAP7_75t_L g6957 ( 
.A(n_6690),
.B(n_6432),
.Y(n_6957)
);

AND2x2_ASAP7_75t_L g6958 ( 
.A(n_6786),
.B(n_6411),
.Y(n_6958)
);

INVx2_ASAP7_75t_L g6959 ( 
.A(n_6695),
.Y(n_6959)
);

INVx1_ASAP7_75t_L g6960 ( 
.A(n_6784),
.Y(n_6960)
);

NOR2xp33_ASAP7_75t_L g6961 ( 
.A(n_6738),
.B(n_6308),
.Y(n_6961)
);

INVx2_ASAP7_75t_L g6962 ( 
.A(n_6679),
.Y(n_6962)
);

INVxp67_ASAP7_75t_L g6963 ( 
.A(n_6595),
.Y(n_6963)
);

AND2x2_ASAP7_75t_L g6964 ( 
.A(n_6794),
.B(n_6475),
.Y(n_6964)
);

INVx1_ASAP7_75t_L g6965 ( 
.A(n_6629),
.Y(n_6965)
);

AND2x2_ASAP7_75t_L g6966 ( 
.A(n_6797),
.B(n_6475),
.Y(n_6966)
);

INVx2_ASAP7_75t_SL g6967 ( 
.A(n_6679),
.Y(n_6967)
);

INVx1_ASAP7_75t_L g6968 ( 
.A(n_6634),
.Y(n_6968)
);

AND2x4_ASAP7_75t_L g6969 ( 
.A(n_6649),
.B(n_6308),
.Y(n_6969)
);

HB1xp67_ASAP7_75t_L g6970 ( 
.A(n_6634),
.Y(n_6970)
);

AND2x4_ASAP7_75t_L g6971 ( 
.A(n_6562),
.B(n_6308),
.Y(n_6971)
);

INVx1_ASAP7_75t_L g6972 ( 
.A(n_6638),
.Y(n_6972)
);

HB1xp67_ASAP7_75t_L g6973 ( 
.A(n_6638),
.Y(n_6973)
);

INVx2_ASAP7_75t_L g6974 ( 
.A(n_6659),
.Y(n_6974)
);

A2O1A1Ixp33_ASAP7_75t_L g6975 ( 
.A1(n_6800),
.A2(n_6115),
.B(n_6239),
.C(n_6036),
.Y(n_6975)
);

AND2x2_ASAP7_75t_L g6976 ( 
.A(n_6799),
.B(n_6475),
.Y(n_6976)
);

OR2x2_ASAP7_75t_L g6977 ( 
.A(n_6754),
.B(n_6469),
.Y(n_6977)
);

NAND2xp5_ASAP7_75t_L g6978 ( 
.A(n_6694),
.B(n_6435),
.Y(n_6978)
);

INVx1_ASAP7_75t_L g6979 ( 
.A(n_6640),
.Y(n_6979)
);

NOR2xp33_ASAP7_75t_L g6980 ( 
.A(n_6694),
.B(n_6395),
.Y(n_6980)
);

NAND2xp5_ASAP7_75t_L g6981 ( 
.A(n_6640),
.B(n_6340),
.Y(n_6981)
);

INVx1_ASAP7_75t_L g6982 ( 
.A(n_6648),
.Y(n_6982)
);

OA211x2_ASAP7_75t_L g6983 ( 
.A1(n_6567),
.A2(n_6294),
.B(n_6425),
.C(n_6522),
.Y(n_6983)
);

NAND2xp5_ASAP7_75t_L g6984 ( 
.A(n_6648),
.B(n_6340),
.Y(n_6984)
);

AND2x2_ASAP7_75t_L g6985 ( 
.A(n_6578),
.B(n_6485),
.Y(n_6985)
);

INVx1_ASAP7_75t_L g6986 ( 
.A(n_6575),
.Y(n_6986)
);

INVx1_ASAP7_75t_L g6987 ( 
.A(n_6569),
.Y(n_6987)
);

AND2x2_ASAP7_75t_L g6988 ( 
.A(n_6675),
.B(n_6485),
.Y(n_6988)
);

OR2x2_ASAP7_75t_L g6989 ( 
.A(n_6601),
.B(n_6703),
.Y(n_6989)
);

INVx1_ASAP7_75t_L g6990 ( 
.A(n_6573),
.Y(n_6990)
);

INVx3_ASAP7_75t_L g6991 ( 
.A(n_6659),
.Y(n_6991)
);

INVx1_ASAP7_75t_SL g6992 ( 
.A(n_6687),
.Y(n_6992)
);

INVx2_ASAP7_75t_L g6993 ( 
.A(n_6659),
.Y(n_6993)
);

OR2x2_ASAP7_75t_L g6994 ( 
.A(n_6715),
.B(n_6699),
.Y(n_6994)
);

NOR2xp33_ASAP7_75t_L g6995 ( 
.A(n_6750),
.B(n_6482),
.Y(n_6995)
);

INVxp67_ASAP7_75t_L g6996 ( 
.A(n_6595),
.Y(n_6996)
);

NAND2x1p5_ASAP7_75t_L g6997 ( 
.A(n_6661),
.B(n_6486),
.Y(n_6997)
);

NAND2xp5_ASAP7_75t_L g6998 ( 
.A(n_6639),
.B(n_6347),
.Y(n_6998)
);

AND2x2_ASAP7_75t_L g6999 ( 
.A(n_6724),
.B(n_6485),
.Y(n_6999)
);

NOR2xp33_ASAP7_75t_L g7000 ( 
.A(n_6750),
.B(n_6492),
.Y(n_7000)
);

NAND2xp5_ASAP7_75t_L g7001 ( 
.A(n_6641),
.B(n_6646),
.Y(n_7001)
);

INVxp33_ASAP7_75t_L g7002 ( 
.A(n_6779),
.Y(n_7002)
);

OR2x2_ASAP7_75t_L g7003 ( 
.A(n_6767),
.B(n_6469),
.Y(n_7003)
);

INVx2_ASAP7_75t_L g7004 ( 
.A(n_6736),
.Y(n_7004)
);

NOR2xp33_ASAP7_75t_L g7005 ( 
.A(n_6768),
.B(n_6492),
.Y(n_7005)
);

OR2x2_ASAP7_75t_L g7006 ( 
.A(n_6565),
.B(n_6456),
.Y(n_7006)
);

OR2x2_ASAP7_75t_L g7007 ( 
.A(n_6783),
.B(n_6546),
.Y(n_7007)
);

AND2x2_ASAP7_75t_L g7008 ( 
.A(n_6747),
.B(n_6492),
.Y(n_7008)
);

AND2x2_ASAP7_75t_L g7009 ( 
.A(n_6617),
.B(n_6386),
.Y(n_7009)
);

NAND2xp5_ASAP7_75t_L g7010 ( 
.A(n_6696),
.B(n_6347),
.Y(n_7010)
);

OR2x2_ASAP7_75t_L g7011 ( 
.A(n_6769),
.B(n_6551),
.Y(n_7011)
);

INVx1_ASAP7_75t_L g7012 ( 
.A(n_6576),
.Y(n_7012)
);

INVx2_ASAP7_75t_SL g7013 ( 
.A(n_6691),
.Y(n_7013)
);

INVx2_ASAP7_75t_L g7014 ( 
.A(n_6736),
.Y(n_7014)
);

NAND2xp5_ASAP7_75t_L g7015 ( 
.A(n_6696),
.B(n_6348),
.Y(n_7015)
);

OR2x2_ASAP7_75t_L g7016 ( 
.A(n_6604),
.B(n_6431),
.Y(n_7016)
);

AND2x2_ASAP7_75t_L g7017 ( 
.A(n_6617),
.B(n_6386),
.Y(n_7017)
);

INVx1_ASAP7_75t_L g7018 ( 
.A(n_6580),
.Y(n_7018)
);

INVx2_ASAP7_75t_L g7019 ( 
.A(n_6736),
.Y(n_7019)
);

INVx1_ASAP7_75t_L g7020 ( 
.A(n_6582),
.Y(n_7020)
);

OR2x2_ASAP7_75t_L g7021 ( 
.A(n_6623),
.B(n_6451),
.Y(n_7021)
);

INVx1_ASAP7_75t_L g7022 ( 
.A(n_6583),
.Y(n_7022)
);

INVx1_ASAP7_75t_L g7023 ( 
.A(n_6626),
.Y(n_7023)
);

INVx1_ASAP7_75t_L g7024 ( 
.A(n_6636),
.Y(n_7024)
);

OR2x2_ASAP7_75t_L g7025 ( 
.A(n_6805),
.B(n_6581),
.Y(n_7025)
);

AOI32xp33_ASAP7_75t_L g7026 ( 
.A1(n_6846),
.A2(n_6603),
.A3(n_6779),
.B1(n_6741),
.B2(n_6624),
.Y(n_7026)
);

INVx1_ASAP7_75t_SL g7027 ( 
.A(n_6953),
.Y(n_7027)
);

INVx1_ASAP7_75t_L g7028 ( 
.A(n_6808),
.Y(n_7028)
);

AND2x4_ASAP7_75t_L g7029 ( 
.A(n_6889),
.B(n_6385),
.Y(n_7029)
);

INVx1_ASAP7_75t_L g7030 ( 
.A(n_6955),
.Y(n_7030)
);

OR2x2_ASAP7_75t_L g7031 ( 
.A(n_6992),
.B(n_6570),
.Y(n_7031)
);

AND2x4_ASAP7_75t_L g7032 ( 
.A(n_6889),
.B(n_6768),
.Y(n_7032)
);

NAND2xp5_ASAP7_75t_L g7033 ( 
.A(n_6895),
.B(n_6577),
.Y(n_7033)
);

AND2x2_ASAP7_75t_L g7034 ( 
.A(n_6905),
.B(n_6356),
.Y(n_7034)
);

INVx1_ASAP7_75t_L g7035 ( 
.A(n_6970),
.Y(n_7035)
);

AOI22xp5_ASAP7_75t_L g7036 ( 
.A1(n_6899),
.A2(n_6621),
.B1(n_6660),
.B2(n_6727),
.Y(n_7036)
);

XNOR2x1_ASAP7_75t_L g7037 ( 
.A(n_6813),
.B(n_6654),
.Y(n_7037)
);

INVx2_ASAP7_75t_L g7038 ( 
.A(n_6868),
.Y(n_7038)
);

AND2x4_ASAP7_75t_L g7039 ( 
.A(n_6897),
.B(n_6942),
.Y(n_7039)
);

INVxp67_ASAP7_75t_SL g7040 ( 
.A(n_6846),
.Y(n_7040)
);

INVx1_ASAP7_75t_L g7041 ( 
.A(n_6973),
.Y(n_7041)
);

INVx1_ASAP7_75t_L g7042 ( 
.A(n_6874),
.Y(n_7042)
);

NAND2xp5_ASAP7_75t_L g7043 ( 
.A(n_6904),
.B(n_6547),
.Y(n_7043)
);

INVx1_ASAP7_75t_SL g7044 ( 
.A(n_6992),
.Y(n_7044)
);

INVxp67_ASAP7_75t_L g7045 ( 
.A(n_6928),
.Y(n_7045)
);

INVx1_ASAP7_75t_L g7046 ( 
.A(n_6835),
.Y(n_7046)
);

INVx1_ASAP7_75t_L g7047 ( 
.A(n_6841),
.Y(n_7047)
);

AND2x2_ASAP7_75t_L g7048 ( 
.A(n_6811),
.B(n_6550),
.Y(n_7048)
);

OR2x2_ASAP7_75t_L g7049 ( 
.A(n_6875),
.B(n_6706),
.Y(n_7049)
);

INVx1_ASAP7_75t_L g7050 ( 
.A(n_6908),
.Y(n_7050)
);

NOR2xp33_ASAP7_75t_L g7051 ( 
.A(n_6902),
.B(n_6397),
.Y(n_7051)
);

INVx1_ASAP7_75t_L g7052 ( 
.A(n_6910),
.Y(n_7052)
);

NOR2xp67_ASAP7_75t_SL g7053 ( 
.A(n_6809),
.B(n_6668),
.Y(n_7053)
);

INVx1_ASAP7_75t_L g7054 ( 
.A(n_6991),
.Y(n_7054)
);

AND2x2_ASAP7_75t_L g7055 ( 
.A(n_6819),
.B(n_6550),
.Y(n_7055)
);

AND2x2_ASAP7_75t_L g7056 ( 
.A(n_6830),
.B(n_6557),
.Y(n_7056)
);

AOI22xp5_ASAP7_75t_L g7057 ( 
.A1(n_6899),
.A2(n_6798),
.B1(n_6596),
.B2(n_6619),
.Y(n_7057)
);

INVx1_ASAP7_75t_L g7058 ( 
.A(n_6991),
.Y(n_7058)
);

NAND2xp5_ASAP7_75t_L g7059 ( 
.A(n_6931),
.B(n_6557),
.Y(n_7059)
);

INVx1_ASAP7_75t_L g7060 ( 
.A(n_6894),
.Y(n_7060)
);

A2O1A1Ixp33_ASAP7_75t_L g7061 ( 
.A1(n_6837),
.A2(n_6682),
.B(n_6635),
.C(n_6116),
.Y(n_7061)
);

CKINVDCx16_ASAP7_75t_R g7062 ( 
.A(n_7009),
.Y(n_7062)
);

A2O1A1Ixp33_ASAP7_75t_L g7063 ( 
.A1(n_6887),
.A2(n_6635),
.B(n_5973),
.C(n_6688),
.Y(n_7063)
);

INVx2_ASAP7_75t_SL g7064 ( 
.A(n_6858),
.Y(n_7064)
);

OAI22xp5_ASAP7_75t_SL g7065 ( 
.A1(n_6931),
.A2(n_6647),
.B1(n_6652),
.B2(n_6496),
.Y(n_7065)
);

AOI21xp33_ASAP7_75t_SL g7066 ( 
.A1(n_6816),
.A2(n_6755),
.B(n_6717),
.Y(n_7066)
);

HB1xp67_ASAP7_75t_L g7067 ( 
.A(n_6859),
.Y(n_7067)
);

AND2x2_ASAP7_75t_L g7068 ( 
.A(n_6885),
.B(n_6558),
.Y(n_7068)
);

OAI21xp33_ASAP7_75t_L g7069 ( 
.A1(n_6877),
.A2(n_6741),
.B(n_6796),
.Y(n_7069)
);

INVx1_ASAP7_75t_L g7070 ( 
.A(n_6894),
.Y(n_7070)
);

OR2x2_ASAP7_75t_L g7071 ( 
.A(n_6884),
.B(n_6759),
.Y(n_7071)
);

A2O1A1Ixp33_ASAP7_75t_L g7072 ( 
.A1(n_6887),
.A2(n_6635),
.B(n_6774),
.C(n_6636),
.Y(n_7072)
);

NOR2x1_ASAP7_75t_L g7073 ( 
.A(n_6864),
.B(n_6795),
.Y(n_7073)
);

INVx1_ASAP7_75t_L g7074 ( 
.A(n_6894),
.Y(n_7074)
);

INVx2_ASAP7_75t_L g7075 ( 
.A(n_6956),
.Y(n_7075)
);

NAND2xp5_ASAP7_75t_L g7076 ( 
.A(n_6897),
.B(n_6558),
.Y(n_7076)
);

NOR2x1_ASAP7_75t_L g7077 ( 
.A(n_6937),
.B(n_6795),
.Y(n_7077)
);

AND2x2_ASAP7_75t_L g7078 ( 
.A(n_6871),
.B(n_6354),
.Y(n_7078)
);

NAND2xp5_ASAP7_75t_L g7079 ( 
.A(n_6942),
.B(n_6752),
.Y(n_7079)
);

INVx1_ASAP7_75t_L g7080 ( 
.A(n_6965),
.Y(n_7080)
);

OAI22xp33_ASAP7_75t_L g7081 ( 
.A1(n_6816),
.A2(n_6200),
.B1(n_6207),
.B2(n_6101),
.Y(n_7081)
);

INVx2_ASAP7_75t_SL g7082 ( 
.A(n_6969),
.Y(n_7082)
);

NAND2xp5_ASAP7_75t_L g7083 ( 
.A(n_6969),
.B(n_6752),
.Y(n_7083)
);

AOI22xp33_ASAP7_75t_L g7084 ( 
.A1(n_7002),
.A2(n_6619),
.B1(n_6029),
.B2(n_6062),
.Y(n_7084)
);

AOI221xp5_ASAP7_75t_SL g7085 ( 
.A1(n_6859),
.A2(n_6877),
.B1(n_6824),
.B2(n_6807),
.C(n_6839),
.Y(n_7085)
);

NOR2xp33_ASAP7_75t_L g7086 ( 
.A(n_6937),
.B(n_6928),
.Y(n_7086)
);

AND2x2_ASAP7_75t_L g7087 ( 
.A(n_6845),
.B(n_6354),
.Y(n_7087)
);

AND2x2_ASAP7_75t_L g7088 ( 
.A(n_6909),
.B(n_6355),
.Y(n_7088)
);

INVxp67_ASAP7_75t_L g7089 ( 
.A(n_6985),
.Y(n_7089)
);

NOR2xp33_ASAP7_75t_L g7090 ( 
.A(n_6867),
.B(n_6391),
.Y(n_7090)
);

OAI22xp33_ASAP7_75t_L g7091 ( 
.A1(n_6854),
.A2(n_5978),
.B1(n_6735),
.B2(n_5987),
.Y(n_7091)
);

INVx1_ASAP7_75t_L g7092 ( 
.A(n_6968),
.Y(n_7092)
);

INVx1_ASAP7_75t_L g7093 ( 
.A(n_6972),
.Y(n_7093)
);

INVx1_ASAP7_75t_L g7094 ( 
.A(n_6979),
.Y(n_7094)
);

NAND2x1p5_ASAP7_75t_L g7095 ( 
.A(n_6833),
.B(n_6788),
.Y(n_7095)
);

INVx2_ASAP7_75t_L g7096 ( 
.A(n_6840),
.Y(n_7096)
);

INVxp33_ASAP7_75t_L g7097 ( 
.A(n_6997),
.Y(n_7097)
);

AND3x2_ASAP7_75t_L g7098 ( 
.A(n_6824),
.B(n_6755),
.C(n_6804),
.Y(n_7098)
);

INVx3_ASAP7_75t_L g7099 ( 
.A(n_6833),
.Y(n_7099)
);

AND2x2_ASAP7_75t_L g7100 ( 
.A(n_7017),
.B(n_6355),
.Y(n_7100)
);

NAND2xp5_ASAP7_75t_L g7101 ( 
.A(n_6967),
.B(n_6752),
.Y(n_7101)
);

INVx1_ASAP7_75t_L g7102 ( 
.A(n_6982),
.Y(n_7102)
);

AND2x2_ASAP7_75t_L g7103 ( 
.A(n_6890),
.B(n_6389),
.Y(n_7103)
);

NAND4xp75_ASAP7_75t_L g7104 ( 
.A(n_6983),
.B(n_6730),
.C(n_6756),
.D(n_6572),
.Y(n_7104)
);

OAI22xp33_ASAP7_75t_L g7105 ( 
.A1(n_6952),
.A2(n_6672),
.B1(n_6676),
.B2(n_6671),
.Y(n_7105)
);

NAND2x1p5_ASAP7_75t_L g7106 ( 
.A(n_6971),
.B(n_6903),
.Y(n_7106)
);

OAI22xp5_ASAP7_75t_L g7107 ( 
.A1(n_6882),
.A2(n_6596),
.B1(n_6612),
.B2(n_6214),
.Y(n_7107)
);

INVxp67_ASAP7_75t_SL g7108 ( 
.A(n_6872),
.Y(n_7108)
);

INVx2_ASAP7_75t_SL g7109 ( 
.A(n_6869),
.Y(n_7109)
);

INVx1_ASAP7_75t_L g7110 ( 
.A(n_6812),
.Y(n_7110)
);

INVx1_ASAP7_75t_L g7111 ( 
.A(n_6815),
.Y(n_7111)
);

INVx1_ASAP7_75t_L g7112 ( 
.A(n_6878),
.Y(n_7112)
);

HB1xp67_ASAP7_75t_L g7113 ( 
.A(n_7004),
.Y(n_7113)
);

INVx1_ASAP7_75t_L g7114 ( 
.A(n_6912),
.Y(n_7114)
);

INVx1_ASAP7_75t_L g7115 ( 
.A(n_6981),
.Y(n_7115)
);

INVx1_ASAP7_75t_L g7116 ( 
.A(n_6981),
.Y(n_7116)
);

A2O1A1Ixp33_ASAP7_75t_L g7117 ( 
.A1(n_6975),
.A2(n_6716),
.B(n_6697),
.C(n_6680),
.Y(n_7117)
);

AOI22xp33_ASAP7_75t_L g7118 ( 
.A1(n_6989),
.A2(n_6619),
.B1(n_6029),
.B2(n_6062),
.Y(n_7118)
);

INVx1_ASAP7_75t_L g7119 ( 
.A(n_6984),
.Y(n_7119)
);

OAI32xp33_ASAP7_75t_L g7120 ( 
.A1(n_6826),
.A2(n_6637),
.A3(n_6533),
.B1(n_6563),
.B2(n_6536),
.Y(n_7120)
);

NAND4xp25_ASAP7_75t_L g7121 ( 
.A(n_6946),
.B(n_6748),
.C(n_6608),
.D(n_6615),
.Y(n_7121)
);

OR2x2_ASAP7_75t_L g7122 ( 
.A(n_6884),
.B(n_6892),
.Y(n_7122)
);

OAI22xp5_ASAP7_75t_L g7123 ( 
.A1(n_6873),
.A2(n_6907),
.B1(n_6946),
.B2(n_7003),
.Y(n_7123)
);

AND2x2_ASAP7_75t_L g7124 ( 
.A(n_6857),
.B(n_6958),
.Y(n_7124)
);

INVx1_ASAP7_75t_L g7125 ( 
.A(n_6984),
.Y(n_7125)
);

NOR2xp33_ASAP7_75t_L g7126 ( 
.A(n_6867),
.B(n_6391),
.Y(n_7126)
);

INVx1_ASAP7_75t_L g7127 ( 
.A(n_6806),
.Y(n_7127)
);

NOR3x1_ASAP7_75t_L g7128 ( 
.A(n_6849),
.B(n_6633),
.C(n_6632),
.Y(n_7128)
);

INVx1_ASAP7_75t_L g7129 ( 
.A(n_7014),
.Y(n_7129)
);

INVx1_ASAP7_75t_L g7130 ( 
.A(n_7019),
.Y(n_7130)
);

INVx1_ASAP7_75t_L g7131 ( 
.A(n_6923),
.Y(n_7131)
);

INVx1_ASAP7_75t_L g7132 ( 
.A(n_6810),
.Y(n_7132)
);

NAND2x1_ASAP7_75t_L g7133 ( 
.A(n_6840),
.B(n_6539),
.Y(n_7133)
);

NAND2xp5_ASAP7_75t_L g7134 ( 
.A(n_6926),
.B(n_6804),
.Y(n_7134)
);

INVx1_ASAP7_75t_L g7135 ( 
.A(n_6814),
.Y(n_7135)
);

A2O1A1Ixp33_ASAP7_75t_L g7136 ( 
.A1(n_6826),
.A2(n_6712),
.B(n_6677),
.C(n_6692),
.Y(n_7136)
);

AND2x2_ASAP7_75t_L g7137 ( 
.A(n_6945),
.B(n_6389),
.Y(n_7137)
);

NAND2xp5_ASAP7_75t_L g7138 ( 
.A(n_6926),
.B(n_6524),
.Y(n_7138)
);

INVx1_ASAP7_75t_L g7139 ( 
.A(n_6818),
.Y(n_7139)
);

INVx1_ASAP7_75t_L g7140 ( 
.A(n_6892),
.Y(n_7140)
);

NOR2x1p5_ASAP7_75t_SL g7141 ( 
.A(n_6948),
.B(n_6515),
.Y(n_7141)
);

INVx1_ASAP7_75t_L g7142 ( 
.A(n_6896),
.Y(n_7142)
);

NAND2xp5_ASAP7_75t_L g7143 ( 
.A(n_6873),
.B(n_6524),
.Y(n_7143)
);

OR2x2_ASAP7_75t_L g7144 ( 
.A(n_6896),
.B(n_6790),
.Y(n_7144)
);

AOI32xp33_ASAP7_75t_L g7145 ( 
.A1(n_6839),
.A2(n_6170),
.A3(n_6599),
.B1(n_6618),
.B2(n_6616),
.Y(n_7145)
);

OAI22xp33_ASAP7_75t_L g7146 ( 
.A1(n_6914),
.A2(n_6705),
.B1(n_6711),
.B2(n_6681),
.Y(n_7146)
);

AOI22xp5_ASAP7_75t_L g7147 ( 
.A1(n_6807),
.A2(n_6729),
.B1(n_6718),
.B2(n_6530),
.Y(n_7147)
);

INVx1_ASAP7_75t_L g7148 ( 
.A(n_6917),
.Y(n_7148)
);

INVx2_ASAP7_75t_SL g7149 ( 
.A(n_6971),
.Y(n_7149)
);

NAND2xp5_ASAP7_75t_L g7150 ( 
.A(n_6907),
.B(n_6528),
.Y(n_7150)
);

AO221x1_ASAP7_75t_L g7151 ( 
.A1(n_6853),
.A2(n_6024),
.B1(n_6959),
.B2(n_6541),
.C(n_6123),
.Y(n_7151)
);

INVx1_ASAP7_75t_L g7152 ( 
.A(n_6917),
.Y(n_7152)
);

NOR2xp67_ASAP7_75t_L g7153 ( 
.A(n_6853),
.B(n_6876),
.Y(n_7153)
);

NAND3xp33_ASAP7_75t_L g7154 ( 
.A(n_6847),
.B(n_6631),
.C(n_6627),
.Y(n_7154)
);

AND2x2_ASAP7_75t_L g7155 ( 
.A(n_6913),
.B(n_6467),
.Y(n_7155)
);

AOI21xp33_ASAP7_75t_SL g7156 ( 
.A1(n_6997),
.A2(n_6739),
.B(n_6737),
.Y(n_7156)
);

INVx1_ASAP7_75t_L g7157 ( 
.A(n_6974),
.Y(n_7157)
);

OR2x2_ASAP7_75t_L g7158 ( 
.A(n_6941),
.B(n_6488),
.Y(n_7158)
);

AOI32xp33_ASAP7_75t_L g7159 ( 
.A1(n_6831),
.A2(n_6801),
.A3(n_6793),
.B1(n_6622),
.B2(n_6657),
.Y(n_7159)
);

NOR2x1_ASAP7_75t_L g7160 ( 
.A(n_6962),
.B(n_6358),
.Y(n_7160)
);

AND2x2_ASAP7_75t_L g7161 ( 
.A(n_6927),
.B(n_6935),
.Y(n_7161)
);

INVx1_ASAP7_75t_L g7162 ( 
.A(n_6993),
.Y(n_7162)
);

NAND2xp5_ASAP7_75t_L g7163 ( 
.A(n_6925),
.B(n_6528),
.Y(n_7163)
);

INVx1_ASAP7_75t_L g7164 ( 
.A(n_6941),
.Y(n_7164)
);

NOR2xp33_ASAP7_75t_SL g7165 ( 
.A(n_6940),
.B(n_6392),
.Y(n_7165)
);

AND2x2_ASAP7_75t_L g7166 ( 
.A(n_6966),
.B(n_6467),
.Y(n_7166)
);

INVx1_ASAP7_75t_L g7167 ( 
.A(n_6888),
.Y(n_7167)
);

NAND3xp33_ASAP7_75t_L g7168 ( 
.A(n_6847),
.B(n_6631),
.C(n_6627),
.Y(n_7168)
);

INVx1_ASAP7_75t_L g7169 ( 
.A(n_6888),
.Y(n_7169)
);

INVxp33_ASAP7_75t_L g7170 ( 
.A(n_6961),
.Y(n_7170)
);

INVx1_ASAP7_75t_L g7171 ( 
.A(n_6963),
.Y(n_7171)
);

AND2x2_ASAP7_75t_L g7172 ( 
.A(n_6976),
.B(n_6728),
.Y(n_7172)
);

INVxp67_ASAP7_75t_L g7173 ( 
.A(n_6893),
.Y(n_7173)
);

NOR2x1_ASAP7_75t_L g7174 ( 
.A(n_6862),
.B(n_6358),
.Y(n_7174)
);

INVx1_ASAP7_75t_L g7175 ( 
.A(n_6963),
.Y(n_7175)
);

NAND4xp75_ASAP7_75t_SL g7176 ( 
.A(n_7008),
.B(n_6536),
.C(n_6409),
.D(n_6383),
.Y(n_7176)
);

AOI32xp33_ASAP7_75t_L g7177 ( 
.A1(n_6944),
.A2(n_6657),
.A3(n_6622),
.B1(n_6614),
.B2(n_6144),
.Y(n_7177)
);

INVx1_ASAP7_75t_L g7178 ( 
.A(n_6996),
.Y(n_7178)
);

OAI221xp5_ASAP7_75t_L g7179 ( 
.A1(n_6944),
.A2(n_6159),
.B1(n_6144),
.B2(n_6048),
.C(n_6194),
.Y(n_7179)
);

NOR2xp33_ASAP7_75t_L g7180 ( 
.A(n_6934),
.B(n_6525),
.Y(n_7180)
);

NAND2xp5_ASAP7_75t_L g7181 ( 
.A(n_6880),
.B(n_6529),
.Y(n_7181)
);

INVx2_ASAP7_75t_L g7182 ( 
.A(n_6920),
.Y(n_7182)
);

INVx1_ASAP7_75t_L g7183 ( 
.A(n_6996),
.Y(n_7183)
);

AND2x2_ASAP7_75t_L g7184 ( 
.A(n_6988),
.B(n_6525),
.Y(n_7184)
);

OAI32xp33_ASAP7_75t_L g7185 ( 
.A1(n_6977),
.A2(n_6488),
.A3(n_6334),
.B1(n_6552),
.B2(n_6762),
.Y(n_7185)
);

AND2x2_ASAP7_75t_L g7186 ( 
.A(n_6964),
.B(n_6622),
.Y(n_7186)
);

NAND2xp5_ASAP7_75t_L g7187 ( 
.A(n_7023),
.B(n_6529),
.Y(n_7187)
);

NAND2xp5_ASAP7_75t_SL g7188 ( 
.A(n_6863),
.B(n_6657),
.Y(n_7188)
);

OR2x2_ASAP7_75t_L g7189 ( 
.A(n_6828),
.B(n_6453),
.Y(n_7189)
);

INVx1_ASAP7_75t_L g7190 ( 
.A(n_6822),
.Y(n_7190)
);

OAI32xp33_ASAP7_75t_L g7191 ( 
.A1(n_6916),
.A2(n_6334),
.A3(n_6762),
.B1(n_6743),
.B2(n_6744),
.Y(n_7191)
);

AND2x4_ASAP7_75t_L g7192 ( 
.A(n_6999),
.B(n_6579),
.Y(n_7192)
);

OR2x2_ASAP7_75t_L g7193 ( 
.A(n_6825),
.B(n_6476),
.Y(n_7193)
);

OAI22xp33_ASAP7_75t_L g7194 ( 
.A1(n_6994),
.A2(n_6614),
.B1(n_6235),
.B2(n_6188),
.Y(n_7194)
);

OAI22xp5_ASAP7_75t_L g7195 ( 
.A1(n_6951),
.A2(n_6520),
.B1(n_6159),
.B2(n_6539),
.Y(n_7195)
);

AND2x2_ASAP7_75t_L g7196 ( 
.A(n_6891),
.B(n_6787),
.Y(n_7196)
);

NAND2xp33_ASAP7_75t_L g7197 ( 
.A(n_7016),
.B(n_6392),
.Y(n_7197)
);

AOI22xp5_ASAP7_75t_L g7198 ( 
.A1(n_6832),
.A2(n_6669),
.B1(n_6663),
.B2(n_6707),
.Y(n_7198)
);

OR2x2_ASAP7_75t_L g7199 ( 
.A(n_6836),
.B(n_6527),
.Y(n_7199)
);

AND2x4_ASAP7_75t_L g7200 ( 
.A(n_6881),
.B(n_6579),
.Y(n_7200)
);

INVx1_ASAP7_75t_SL g7201 ( 
.A(n_7021),
.Y(n_7201)
);

OAI22xp5_ASAP7_75t_L g7202 ( 
.A1(n_7007),
.A2(n_7006),
.B1(n_7011),
.B2(n_6938),
.Y(n_7202)
);

NAND2xp5_ASAP7_75t_L g7203 ( 
.A(n_6933),
.B(n_6531),
.Y(n_7203)
);

NAND2x1p5_ASAP7_75t_L g7204 ( 
.A(n_7000),
.B(n_6327),
.Y(n_7204)
);

INVx1_ASAP7_75t_L g7205 ( 
.A(n_6829),
.Y(n_7205)
);

AO22x1_ASAP7_75t_L g7206 ( 
.A1(n_6843),
.A2(n_6541),
.B1(n_6746),
.B2(n_6742),
.Y(n_7206)
);

AOI22xp5_ASAP7_75t_L g7207 ( 
.A1(n_6834),
.A2(n_6669),
.B1(n_6663),
.B2(n_6707),
.Y(n_7207)
);

INVx1_ASAP7_75t_L g7208 ( 
.A(n_6823),
.Y(n_7208)
);

AOI32xp33_ASAP7_75t_L g7209 ( 
.A1(n_7024),
.A2(n_6802),
.A3(n_6520),
.B1(n_6348),
.B2(n_6380),
.Y(n_7209)
);

XOR2x2_ASAP7_75t_L g7210 ( 
.A(n_6980),
.B(n_6780),
.Y(n_7210)
);

AND2x2_ASAP7_75t_L g7211 ( 
.A(n_6827),
.B(n_6787),
.Y(n_7211)
);

OR2x2_ASAP7_75t_L g7212 ( 
.A(n_7062),
.B(n_6932),
.Y(n_7212)
);

INVx1_ASAP7_75t_L g7213 ( 
.A(n_7099),
.Y(n_7213)
);

OR2x2_ASAP7_75t_L g7214 ( 
.A(n_7049),
.B(n_7122),
.Y(n_7214)
);

HB1xp67_ASAP7_75t_L g7215 ( 
.A(n_7133),
.Y(n_7215)
);

INVx2_ASAP7_75t_SL g7216 ( 
.A(n_7039),
.Y(n_7216)
);

INVx1_ASAP7_75t_L g7217 ( 
.A(n_7099),
.Y(n_7217)
);

INVx1_ASAP7_75t_L g7218 ( 
.A(n_7138),
.Y(n_7218)
);

NAND3x1_ASAP7_75t_L g7219 ( 
.A(n_7073),
.B(n_7005),
.C(n_6995),
.Y(n_7219)
);

OR2x2_ASAP7_75t_L g7220 ( 
.A(n_7027),
.B(n_6932),
.Y(n_7220)
);

NOR2x1_ASAP7_75t_L g7221 ( 
.A(n_7104),
.B(n_7010),
.Y(n_7221)
);

AND2x2_ASAP7_75t_L g7222 ( 
.A(n_7186),
.B(n_6901),
.Y(n_7222)
);

INVx4_ASAP7_75t_L g7223 ( 
.A(n_7032),
.Y(n_7223)
);

INVx1_ASAP7_75t_SL g7224 ( 
.A(n_7044),
.Y(n_7224)
);

INVxp67_ASAP7_75t_L g7225 ( 
.A(n_7051),
.Y(n_7225)
);

INVx1_ASAP7_75t_L g7226 ( 
.A(n_7059),
.Y(n_7226)
);

OA21x2_ASAP7_75t_L g7227 ( 
.A1(n_7085),
.A2(n_7015),
.B(n_7010),
.Y(n_7227)
);

AOI22xp5_ASAP7_75t_L g7228 ( 
.A1(n_7057),
.A2(n_6842),
.B1(n_6838),
.B2(n_6860),
.Y(n_7228)
);

OAI21x1_ASAP7_75t_L g7229 ( 
.A1(n_7106),
.A2(n_6820),
.B(n_7077),
.Y(n_7229)
);

CKINVDCx16_ASAP7_75t_R g7230 ( 
.A(n_7192),
.Y(n_7230)
);

INVx1_ASAP7_75t_L g7231 ( 
.A(n_7113),
.Y(n_7231)
);

AOI22xp33_ASAP7_75t_L g7232 ( 
.A1(n_7057),
.A2(n_6048),
.B1(n_6713),
.B2(n_6708),
.Y(n_7232)
);

NAND2xp5_ASAP7_75t_L g7233 ( 
.A(n_7085),
.B(n_6817),
.Y(n_7233)
);

INVx1_ASAP7_75t_L g7234 ( 
.A(n_7143),
.Y(n_7234)
);

AND2x2_ASAP7_75t_L g7235 ( 
.A(n_7161),
.B(n_6803),
.Y(n_7235)
);

INVx1_ASAP7_75t_L g7236 ( 
.A(n_7150),
.Y(n_7236)
);

NAND2xp5_ASAP7_75t_L g7237 ( 
.A(n_7036),
.B(n_6821),
.Y(n_7237)
);

HB1xp67_ASAP7_75t_L g7238 ( 
.A(n_7039),
.Y(n_7238)
);

INVx1_ASAP7_75t_L g7239 ( 
.A(n_7144),
.Y(n_7239)
);

NAND2xp5_ASAP7_75t_L g7240 ( 
.A(n_7036),
.B(n_6900),
.Y(n_7240)
);

AND2x2_ASAP7_75t_L g7241 ( 
.A(n_7034),
.B(n_6803),
.Y(n_7241)
);

AND2x4_ASAP7_75t_L g7242 ( 
.A(n_7153),
.B(n_7029),
.Y(n_7242)
);

INVx1_ASAP7_75t_L g7243 ( 
.A(n_7067),
.Y(n_7243)
);

INVx1_ASAP7_75t_L g7244 ( 
.A(n_7193),
.Y(n_7244)
);

OR2x2_ASAP7_75t_L g7245 ( 
.A(n_7158),
.B(n_7001),
.Y(n_7245)
);

INVx6_ASAP7_75t_L g7246 ( 
.A(n_7032),
.Y(n_7246)
);

NAND2xp5_ASAP7_75t_L g7247 ( 
.A(n_7100),
.B(n_6986),
.Y(n_7247)
);

NAND2xp5_ASAP7_75t_L g7248 ( 
.A(n_7124),
.B(n_6920),
.Y(n_7248)
);

NAND2xp5_ASAP7_75t_L g7249 ( 
.A(n_7082),
.B(n_6906),
.Y(n_7249)
);

INVx1_ASAP7_75t_SL g7250 ( 
.A(n_7031),
.Y(n_7250)
);

OR2x2_ASAP7_75t_L g7251 ( 
.A(n_7201),
.B(n_7001),
.Y(n_7251)
);

INVx2_ASAP7_75t_SL g7252 ( 
.A(n_7192),
.Y(n_7252)
);

NOR2xp33_ASAP7_75t_L g7253 ( 
.A(n_7097),
.B(n_7013),
.Y(n_7253)
);

INVx1_ASAP7_75t_L g7254 ( 
.A(n_7141),
.Y(n_7254)
);

AND2x2_ASAP7_75t_L g7255 ( 
.A(n_7048),
.B(n_6532),
.Y(n_7255)
);

INVx1_ASAP7_75t_SL g7256 ( 
.A(n_7025),
.Y(n_7256)
);

INVx2_ASAP7_75t_L g7257 ( 
.A(n_7095),
.Y(n_7257)
);

NAND2xp5_ASAP7_75t_L g7258 ( 
.A(n_7040),
.B(n_7026),
.Y(n_7258)
);

INVx1_ASAP7_75t_L g7259 ( 
.A(n_7188),
.Y(n_7259)
);

INVx1_ASAP7_75t_L g7260 ( 
.A(n_7068),
.Y(n_7260)
);

INVx2_ASAP7_75t_L g7261 ( 
.A(n_7055),
.Y(n_7261)
);

AND2x4_ASAP7_75t_L g7262 ( 
.A(n_7153),
.B(n_6915),
.Y(n_7262)
);

BUFx2_ASAP7_75t_L g7263 ( 
.A(n_7029),
.Y(n_7263)
);

AND2x2_ASAP7_75t_L g7264 ( 
.A(n_7056),
.B(n_7078),
.Y(n_7264)
);

INVx1_ASAP7_75t_L g7265 ( 
.A(n_7079),
.Y(n_7265)
);

INVx1_ASAP7_75t_SL g7266 ( 
.A(n_7083),
.Y(n_7266)
);

INVx2_ASAP7_75t_L g7267 ( 
.A(n_7137),
.Y(n_7267)
);

INVx2_ASAP7_75t_L g7268 ( 
.A(n_7087),
.Y(n_7268)
);

INVx1_ASAP7_75t_L g7269 ( 
.A(n_7134),
.Y(n_7269)
);

AOI222xp33_ASAP7_75t_L g7270 ( 
.A1(n_7154),
.A2(n_6850),
.B1(n_6860),
.B2(n_7012),
.C1(n_6990),
.C2(n_6987),
.Y(n_7270)
);

INVx2_ASAP7_75t_L g7271 ( 
.A(n_7088),
.Y(n_7271)
);

AOI22xp5_ASAP7_75t_L g7272 ( 
.A1(n_7081),
.A2(n_6850),
.B1(n_7020),
.B2(n_7018),
.Y(n_7272)
);

AOI21xp5_ASAP7_75t_L g7273 ( 
.A1(n_7037),
.A2(n_7015),
.B(n_6911),
.Y(n_7273)
);

AND2x4_ASAP7_75t_L g7274 ( 
.A(n_7200),
.B(n_7166),
.Y(n_7274)
);

AND2x2_ASAP7_75t_L g7275 ( 
.A(n_7103),
.B(n_7155),
.Y(n_7275)
);

INVx1_ASAP7_75t_SL g7276 ( 
.A(n_7184),
.Y(n_7276)
);

INVx1_ASAP7_75t_SL g7277 ( 
.A(n_7200),
.Y(n_7277)
);

HB1xp67_ASAP7_75t_L g7278 ( 
.A(n_7089),
.Y(n_7278)
);

HB1xp67_ASAP7_75t_L g7279 ( 
.A(n_7149),
.Y(n_7279)
);

INVx1_ASAP7_75t_SL g7280 ( 
.A(n_7098),
.Y(n_7280)
);

NOR2xp33_ASAP7_75t_SL g7281 ( 
.A(n_7108),
.B(n_6820),
.Y(n_7281)
);

NAND2xp5_ASAP7_75t_L g7282 ( 
.A(n_7072),
.B(n_6918),
.Y(n_7282)
);

NAND2xp5_ASAP7_75t_L g7283 ( 
.A(n_7109),
.B(n_6919),
.Y(n_7283)
);

INVx2_ASAP7_75t_L g7284 ( 
.A(n_7204),
.Y(n_7284)
);

INVx1_ASAP7_75t_L g7285 ( 
.A(n_7101),
.Y(n_7285)
);

INVx1_ASAP7_75t_L g7286 ( 
.A(n_7076),
.Y(n_7286)
);

INVx1_ASAP7_75t_L g7287 ( 
.A(n_7043),
.Y(n_7287)
);

INVx1_ASAP7_75t_L g7288 ( 
.A(n_7071),
.Y(n_7288)
);

AND2x2_ASAP7_75t_L g7289 ( 
.A(n_7172),
.B(n_6532),
.Y(n_7289)
);

OAI221xp5_ASAP7_75t_L g7290 ( 
.A1(n_7063),
.A2(n_6855),
.B1(n_6852),
.B2(n_6844),
.C(n_6851),
.Y(n_7290)
);

NOR2xp33_ASAP7_75t_L g7291 ( 
.A(n_7170),
.B(n_6691),
.Y(n_7291)
);

AND2x2_ASAP7_75t_L g7292 ( 
.A(n_7064),
.B(n_6559),
.Y(n_7292)
);

INVx1_ASAP7_75t_SL g7293 ( 
.A(n_7189),
.Y(n_7293)
);

AOI22xp5_ASAP7_75t_L g7294 ( 
.A1(n_7107),
.A2(n_7022),
.B1(n_6856),
.B2(n_6861),
.Y(n_7294)
);

INVx1_ASAP7_75t_SL g7295 ( 
.A(n_7210),
.Y(n_7295)
);

AND2x2_ASAP7_75t_L g7296 ( 
.A(n_7196),
.B(n_6559),
.Y(n_7296)
);

NAND2xp5_ASAP7_75t_L g7297 ( 
.A(n_7177),
.B(n_6921),
.Y(n_7297)
);

INVx2_ASAP7_75t_L g7298 ( 
.A(n_7038),
.Y(n_7298)
);

INVx1_ASAP7_75t_L g7299 ( 
.A(n_7187),
.Y(n_7299)
);

OR2x2_ASAP7_75t_L g7300 ( 
.A(n_7123),
.B(n_6950),
.Y(n_7300)
);

INVx1_ASAP7_75t_L g7301 ( 
.A(n_7112),
.Y(n_7301)
);

OR2x2_ASAP7_75t_L g7302 ( 
.A(n_7033),
.B(n_6950),
.Y(n_7302)
);

INVx1_ASAP7_75t_L g7303 ( 
.A(n_7065),
.Y(n_7303)
);

INVx1_ASAP7_75t_L g7304 ( 
.A(n_7065),
.Y(n_7304)
);

INVx1_ASAP7_75t_L g7305 ( 
.A(n_7181),
.Y(n_7305)
);

AND2x2_ASAP7_75t_L g7306 ( 
.A(n_7211),
.B(n_7075),
.Y(n_7306)
);

NOR2xp33_ASAP7_75t_L g7307 ( 
.A(n_7045),
.B(n_6539),
.Y(n_7307)
);

AND2x2_ASAP7_75t_L g7308 ( 
.A(n_7190),
.B(n_6520),
.Y(n_7308)
);

INVx1_ASAP7_75t_L g7309 ( 
.A(n_7046),
.Y(n_7309)
);

AO22x1_ASAP7_75t_L g7310 ( 
.A1(n_7128),
.A2(n_6924),
.B1(n_6929),
.B2(n_6922),
.Y(n_7310)
);

OAI21x1_ASAP7_75t_L g7311 ( 
.A1(n_7174),
.A2(n_6541),
.B(n_6852),
.Y(n_7311)
);

AND2x2_ASAP7_75t_L g7312 ( 
.A(n_7114),
.B(n_6549),
.Y(n_7312)
);

CKINVDCx16_ASAP7_75t_R g7313 ( 
.A(n_7165),
.Y(n_7313)
);

OAI21xp33_ASAP7_75t_L g7314 ( 
.A1(n_7159),
.A2(n_6531),
.B(n_6549),
.Y(n_7314)
);

INVx3_ASAP7_75t_L g7315 ( 
.A(n_7096),
.Y(n_7315)
);

AND2x2_ASAP7_75t_L g7316 ( 
.A(n_7090),
.B(n_6549),
.Y(n_7316)
);

INVx1_ASAP7_75t_L g7317 ( 
.A(n_7047),
.Y(n_7317)
);

NAND2xp5_ASAP7_75t_SL g7318 ( 
.A(n_7066),
.B(n_6317),
.Y(n_7318)
);

BUFx3_ASAP7_75t_L g7319 ( 
.A(n_7163),
.Y(n_7319)
);

OR2x2_ASAP7_75t_L g7320 ( 
.A(n_7140),
.B(n_6957),
.Y(n_7320)
);

INVx2_ASAP7_75t_SL g7321 ( 
.A(n_7160),
.Y(n_7321)
);

INVx1_ASAP7_75t_SL g7322 ( 
.A(n_7197),
.Y(n_7322)
);

AOI22xp33_ASAP7_75t_L g7323 ( 
.A1(n_7151),
.A2(n_7179),
.B1(n_7154),
.B2(n_7168),
.Y(n_7323)
);

INVx1_ASAP7_75t_SL g7324 ( 
.A(n_7199),
.Y(n_7324)
);

OAI22xp5_ASAP7_75t_L g7325 ( 
.A1(n_7069),
.A2(n_6855),
.B1(n_6978),
.B2(n_6957),
.Y(n_7325)
);

INVx1_ASAP7_75t_L g7326 ( 
.A(n_7202),
.Y(n_7326)
);

AND2x2_ASAP7_75t_L g7327 ( 
.A(n_7126),
.B(n_6610),
.Y(n_7327)
);

INVx1_ASAP7_75t_L g7328 ( 
.A(n_7028),
.Y(n_7328)
);

AND2x2_ASAP7_75t_L g7329 ( 
.A(n_7180),
.B(n_6947),
.Y(n_7329)
);

INVx2_ASAP7_75t_L g7330 ( 
.A(n_7042),
.Y(n_7330)
);

NOR2xp67_ASAP7_75t_L g7331 ( 
.A(n_7156),
.B(n_6317),
.Y(n_7331)
);

NAND2xp5_ASAP7_75t_L g7332 ( 
.A(n_7142),
.B(n_6930),
.Y(n_7332)
);

INVx1_ASAP7_75t_L g7333 ( 
.A(n_7206),
.Y(n_7333)
);

AND2x2_ASAP7_75t_L g7334 ( 
.A(n_7066),
.B(n_6949),
.Y(n_7334)
);

NOR3xp33_ASAP7_75t_L g7335 ( 
.A(n_7069),
.B(n_6978),
.C(n_6939),
.Y(n_7335)
);

AND2x2_ASAP7_75t_L g7336 ( 
.A(n_7148),
.B(n_6954),
.Y(n_7336)
);

NAND3xp33_ASAP7_75t_L g7337 ( 
.A(n_7168),
.B(n_6936),
.C(n_6865),
.Y(n_7337)
);

INVx1_ASAP7_75t_L g7338 ( 
.A(n_7198),
.Y(n_7338)
);

INVx1_ASAP7_75t_SL g7339 ( 
.A(n_7203),
.Y(n_7339)
);

INVx2_ASAP7_75t_SL g7340 ( 
.A(n_7050),
.Y(n_7340)
);

INVx2_ASAP7_75t_L g7341 ( 
.A(n_7030),
.Y(n_7341)
);

NAND2xp5_ASAP7_75t_L g7342 ( 
.A(n_7152),
.B(n_6848),
.Y(n_7342)
);

NOR2xp33_ASAP7_75t_L g7343 ( 
.A(n_7120),
.B(n_6364),
.Y(n_7343)
);

OR2x2_ASAP7_75t_L g7344 ( 
.A(n_7164),
.B(n_6960),
.Y(n_7344)
);

AND2x2_ASAP7_75t_L g7345 ( 
.A(n_7086),
.B(n_6943),
.Y(n_7345)
);

INVx1_ASAP7_75t_L g7346 ( 
.A(n_7198),
.Y(n_7346)
);

NOR2x1_ASAP7_75t_L g7347 ( 
.A(n_7176),
.B(n_6866),
.Y(n_7347)
);

INVx2_ASAP7_75t_SL g7348 ( 
.A(n_7052),
.Y(n_7348)
);

NOR2x1_ASAP7_75t_L g7349 ( 
.A(n_7121),
.B(n_6870),
.Y(n_7349)
);

INVxp67_ASAP7_75t_L g7350 ( 
.A(n_7053),
.Y(n_7350)
);

NAND2xp5_ASAP7_75t_L g7351 ( 
.A(n_7156),
.B(n_6879),
.Y(n_7351)
);

NOR2xp33_ASAP7_75t_L g7352 ( 
.A(n_7131),
.B(n_6364),
.Y(n_7352)
);

INVx1_ASAP7_75t_L g7353 ( 
.A(n_7207),
.Y(n_7353)
);

NOR2x1_ASAP7_75t_L g7354 ( 
.A(n_7121),
.B(n_6883),
.Y(n_7354)
);

INVx1_ASAP7_75t_L g7355 ( 
.A(n_7207),
.Y(n_7355)
);

INVx4_ASAP7_75t_L g7356 ( 
.A(n_7182),
.Y(n_7356)
);

INVx2_ASAP7_75t_SL g7357 ( 
.A(n_7060),
.Y(n_7357)
);

AND2x2_ASAP7_75t_L g7358 ( 
.A(n_7173),
.B(n_6886),
.Y(n_7358)
);

INVx1_ASAP7_75t_L g7359 ( 
.A(n_7129),
.Y(n_7359)
);

INVx3_ASAP7_75t_L g7360 ( 
.A(n_7070),
.Y(n_7360)
);

INVxp67_ASAP7_75t_L g7361 ( 
.A(n_7074),
.Y(n_7361)
);

OR2x2_ASAP7_75t_L g7362 ( 
.A(n_7035),
.B(n_6998),
.Y(n_7362)
);

INVx1_ASAP7_75t_L g7363 ( 
.A(n_7130),
.Y(n_7363)
);

AO22x1_ASAP7_75t_L g7364 ( 
.A1(n_7041),
.A2(n_6898),
.B1(n_6309),
.B2(n_6314),
.Y(n_7364)
);

INVx1_ASAP7_75t_L g7365 ( 
.A(n_7147),
.Y(n_7365)
);

INVx2_ASAP7_75t_L g7366 ( 
.A(n_7054),
.Y(n_7366)
);

NAND3xp33_ASAP7_75t_L g7367 ( 
.A(n_7061),
.B(n_6713),
.C(n_6708),
.Y(n_7367)
);

HB1xp67_ASAP7_75t_L g7368 ( 
.A(n_7058),
.Y(n_7368)
);

CKINVDCx16_ASAP7_75t_R g7369 ( 
.A(n_7147),
.Y(n_7369)
);

CKINVDCx16_ASAP7_75t_R g7370 ( 
.A(n_7127),
.Y(n_7370)
);

INVx1_ASAP7_75t_SL g7371 ( 
.A(n_7132),
.Y(n_7371)
);

OR2x2_ASAP7_75t_L g7372 ( 
.A(n_7135),
.B(n_6998),
.Y(n_7372)
);

INVx1_ASAP7_75t_L g7373 ( 
.A(n_7139),
.Y(n_7373)
);

AND2x2_ASAP7_75t_L g7374 ( 
.A(n_7205),
.B(n_6305),
.Y(n_7374)
);

NAND2xp5_ASAP7_75t_L g7375 ( 
.A(n_7146),
.B(n_6366),
.Y(n_7375)
);

INVx2_ASAP7_75t_L g7376 ( 
.A(n_7157),
.Y(n_7376)
);

INVx4_ASAP7_75t_L g7377 ( 
.A(n_7167),
.Y(n_7377)
);

NOR2xp33_ASAP7_75t_L g7378 ( 
.A(n_7185),
.B(n_6305),
.Y(n_7378)
);

INVx1_ASAP7_75t_SL g7379 ( 
.A(n_7162),
.Y(n_7379)
);

INVx1_ASAP7_75t_L g7380 ( 
.A(n_7169),
.Y(n_7380)
);

INVx1_ASAP7_75t_L g7381 ( 
.A(n_7171),
.Y(n_7381)
);

OR2x2_ASAP7_75t_L g7382 ( 
.A(n_7110),
.B(n_6368),
.Y(n_7382)
);

AND2x2_ASAP7_75t_L g7383 ( 
.A(n_7208),
.B(n_6309),
.Y(n_7383)
);

INVx2_ASAP7_75t_L g7384 ( 
.A(n_7111),
.Y(n_7384)
);

OA21x2_ASAP7_75t_L g7385 ( 
.A1(n_7117),
.A2(n_6714),
.B(n_6314),
.Y(n_7385)
);

AOI22xp5_ASAP7_75t_L g7386 ( 
.A1(n_7323),
.A2(n_7369),
.B1(n_7254),
.B2(n_7266),
.Y(n_7386)
);

INVx1_ASAP7_75t_SL g7387 ( 
.A(n_7214),
.Y(n_7387)
);

INVx1_ASAP7_75t_L g7388 ( 
.A(n_7263),
.Y(n_7388)
);

AOI221x1_ASAP7_75t_L g7389 ( 
.A1(n_7273),
.A2(n_7178),
.B1(n_7183),
.B2(n_7175),
.C(n_7136),
.Y(n_7389)
);

NAND3xp33_ASAP7_75t_L g7390 ( 
.A(n_7227),
.B(n_7118),
.C(n_7084),
.Y(n_7390)
);

INVx2_ASAP7_75t_L g7391 ( 
.A(n_7246),
.Y(n_7391)
);

NOR2xp33_ASAP7_75t_L g7392 ( 
.A(n_7246),
.B(n_7191),
.Y(n_7392)
);

NOR2xp67_ASAP7_75t_L g7393 ( 
.A(n_7223),
.B(n_7238),
.Y(n_7393)
);

INVx1_ASAP7_75t_L g7394 ( 
.A(n_7296),
.Y(n_7394)
);

AOI322xp5_ASAP7_75t_L g7395 ( 
.A1(n_7232),
.A2(n_7105),
.A3(n_7091),
.B1(n_6714),
.B2(n_7194),
.C1(n_7119),
.C2(n_7116),
.Y(n_7395)
);

OAI222xp33_ASAP7_75t_L g7396 ( 
.A1(n_7349),
.A2(n_7145),
.B1(n_7195),
.B2(n_7209),
.C1(n_6560),
.C2(n_6548),
.Y(n_7396)
);

OAI22xp5_ASAP7_75t_L g7397 ( 
.A1(n_7250),
.A2(n_7125),
.B1(n_7115),
.B2(n_7092),
.Y(n_7397)
);

INVx1_ASAP7_75t_SL g7398 ( 
.A(n_7256),
.Y(n_7398)
);

INVx2_ASAP7_75t_L g7399 ( 
.A(n_7223),
.Y(n_7399)
);

OAI31xp33_ASAP7_75t_L g7400 ( 
.A1(n_7365),
.A2(n_7367),
.A3(n_7337),
.B(n_7240),
.Y(n_7400)
);

OR2x2_ASAP7_75t_L g7401 ( 
.A(n_7277),
.B(n_7080),
.Y(n_7401)
);

OAI22xp5_ASAP7_75t_L g7402 ( 
.A1(n_7250),
.A2(n_7094),
.B1(n_7102),
.B2(n_7093),
.Y(n_7402)
);

AOI32xp33_ASAP7_75t_L g7403 ( 
.A1(n_7354),
.A2(n_6366),
.A3(n_6382),
.B1(n_6380),
.B2(n_6374),
.Y(n_7403)
);

INVx1_ASAP7_75t_SL g7404 ( 
.A(n_7256),
.Y(n_7404)
);

NAND2xp33_ASAP7_75t_L g7405 ( 
.A(n_7219),
.B(n_6422),
.Y(n_7405)
);

NAND2xp5_ASAP7_75t_L g7406 ( 
.A(n_7230),
.B(n_6548),
.Y(n_7406)
);

OR2x2_ASAP7_75t_L g7407 ( 
.A(n_7277),
.B(n_6376),
.Y(n_7407)
);

AOI22xp33_ASAP7_75t_L g7408 ( 
.A1(n_7367),
.A2(n_6560),
.B1(n_6187),
.B2(n_6173),
.Y(n_7408)
);

INVx1_ASAP7_75t_L g7409 ( 
.A(n_7212),
.Y(n_7409)
);

INVx1_ASAP7_75t_L g7410 ( 
.A(n_7255),
.Y(n_7410)
);

INVxp67_ASAP7_75t_SL g7411 ( 
.A(n_7215),
.Y(n_7411)
);

AND2x2_ASAP7_75t_L g7412 ( 
.A(n_7275),
.B(n_6422),
.Y(n_7412)
);

NOR2xp33_ASAP7_75t_L g7413 ( 
.A(n_7281),
.B(n_6413),
.Y(n_7413)
);

NAND2xp5_ASAP7_75t_L g7414 ( 
.A(n_7242),
.B(n_6416),
.Y(n_7414)
);

NAND2xp5_ASAP7_75t_L g7415 ( 
.A(n_7242),
.B(n_6493),
.Y(n_7415)
);

AND2x2_ASAP7_75t_L g7416 ( 
.A(n_7289),
.B(n_6441),
.Y(n_7416)
);

INVx1_ASAP7_75t_L g7417 ( 
.A(n_7279),
.Y(n_7417)
);

INVx1_ASAP7_75t_SL g7418 ( 
.A(n_7385),
.Y(n_7418)
);

OAI221xp5_ASAP7_75t_L g7419 ( 
.A1(n_7237),
.A2(n_6510),
.B1(n_6487),
.B2(n_6526),
.C(n_6519),
.Y(n_7419)
);

NAND2xp5_ASAP7_75t_L g7420 ( 
.A(n_7252),
.B(n_7216),
.Y(n_7420)
);

AND2x2_ASAP7_75t_L g7421 ( 
.A(n_7274),
.B(n_6441),
.Y(n_7421)
);

NAND2xp5_ASAP7_75t_L g7422 ( 
.A(n_7274),
.B(n_6504),
.Y(n_7422)
);

INVx1_ASAP7_75t_L g7423 ( 
.A(n_7264),
.Y(n_7423)
);

AND2x2_ASAP7_75t_L g7424 ( 
.A(n_7222),
.B(n_6519),
.Y(n_7424)
);

AOI21xp5_ASAP7_75t_L g7425 ( 
.A1(n_7237),
.A2(n_6526),
.B(n_6534),
.Y(n_7425)
);

OAI32xp33_ASAP7_75t_L g7426 ( 
.A1(n_7240),
.A2(n_6384),
.A3(n_6387),
.B1(n_6382),
.B2(n_6374),
.Y(n_7426)
);

OA21x2_ASAP7_75t_L g7427 ( 
.A1(n_7233),
.A2(n_6534),
.B(n_6387),
.Y(n_7427)
);

INVxp67_ASAP7_75t_L g7428 ( 
.A(n_7281),
.Y(n_7428)
);

AOI22xp5_ASAP7_75t_L g7429 ( 
.A1(n_7266),
.A2(n_5990),
.B1(n_6235),
.B2(n_6384),
.Y(n_7429)
);

NAND2xp5_ASAP7_75t_L g7430 ( 
.A(n_7276),
.B(n_6388),
.Y(n_7430)
);

AOI21xp33_ASAP7_75t_SL g7431 ( 
.A1(n_7313),
.A2(n_6093),
.B(n_6388),
.Y(n_7431)
);

OAI21xp33_ASAP7_75t_L g7432 ( 
.A1(n_7314),
.A2(n_7276),
.B(n_7224),
.Y(n_7432)
);

NAND2xp5_ASAP7_75t_L g7433 ( 
.A(n_7324),
.B(n_6393),
.Y(n_7433)
);

AOI22xp5_ASAP7_75t_L g7434 ( 
.A1(n_7370),
.A2(n_6401),
.B1(n_6403),
.B2(n_6393),
.Y(n_7434)
);

NAND2xp5_ASAP7_75t_L g7435 ( 
.A(n_7324),
.B(n_7293),
.Y(n_7435)
);

NOR2xp67_ASAP7_75t_L g7436 ( 
.A(n_7321),
.B(n_6401),
.Y(n_7436)
);

INVx1_ASAP7_75t_L g7437 ( 
.A(n_7306),
.Y(n_7437)
);

AOI221xp5_ASAP7_75t_L g7438 ( 
.A1(n_7325),
.A2(n_6410),
.B1(n_6412),
.B2(n_6404),
.C(n_6403),
.Y(n_7438)
);

INVx1_ASAP7_75t_L g7439 ( 
.A(n_7220),
.Y(n_7439)
);

OAI22xp33_ASAP7_75t_L g7440 ( 
.A1(n_7228),
.A2(n_6410),
.B1(n_6412),
.B2(n_6404),
.Y(n_7440)
);

INVx1_ASAP7_75t_L g7441 ( 
.A(n_7251),
.Y(n_7441)
);

AOI221xp5_ASAP7_75t_L g7442 ( 
.A1(n_7325),
.A2(n_7282),
.B1(n_7233),
.B2(n_7297),
.C(n_7338),
.Y(n_7442)
);

AND2x2_ASAP7_75t_L g7443 ( 
.A(n_7235),
.B(n_6414),
.Y(n_7443)
);

NAND2xp5_ASAP7_75t_L g7444 ( 
.A(n_7293),
.B(n_6414),
.Y(n_7444)
);

INVx1_ASAP7_75t_SL g7445 ( 
.A(n_7385),
.Y(n_7445)
);

INVx1_ASAP7_75t_L g7446 ( 
.A(n_7245),
.Y(n_7446)
);

AOI22xp33_ASAP7_75t_L g7447 ( 
.A1(n_7346),
.A2(n_6163),
.B1(n_6172),
.B2(n_6168),
.Y(n_7447)
);

INVx1_ASAP7_75t_L g7448 ( 
.A(n_7292),
.Y(n_7448)
);

NOR2xp33_ASAP7_75t_L g7449 ( 
.A(n_7224),
.B(n_6418),
.Y(n_7449)
);

INVx1_ASAP7_75t_L g7450 ( 
.A(n_7308),
.Y(n_7450)
);

INVx1_ASAP7_75t_L g7451 ( 
.A(n_7315),
.Y(n_7451)
);

AOI21xp5_ASAP7_75t_L g7452 ( 
.A1(n_7282),
.A2(n_6420),
.B(n_6418),
.Y(n_7452)
);

AND2x2_ASAP7_75t_L g7453 ( 
.A(n_7241),
.B(n_6420),
.Y(n_7453)
);

INVx1_ASAP7_75t_L g7454 ( 
.A(n_7315),
.Y(n_7454)
);

AND2x2_ASAP7_75t_L g7455 ( 
.A(n_7316),
.B(n_6428),
.Y(n_7455)
);

HB1xp67_ASAP7_75t_L g7456 ( 
.A(n_7227),
.Y(n_7456)
);

INVx1_ASAP7_75t_L g7457 ( 
.A(n_7262),
.Y(n_7457)
);

O2A1O1Ixp5_ASAP7_75t_L g7458 ( 
.A1(n_7310),
.A2(n_6428),
.B(n_6443),
.C(n_6436),
.Y(n_7458)
);

NAND2xp5_ASAP7_75t_L g7459 ( 
.A(n_7322),
.B(n_7280),
.Y(n_7459)
);

OAI221xp5_ASAP7_75t_L g7460 ( 
.A1(n_7297),
.A2(n_6468),
.B1(n_6477),
.B2(n_6466),
.C(n_6464),
.Y(n_7460)
);

INVx1_ASAP7_75t_L g7461 ( 
.A(n_7262),
.Y(n_7461)
);

NAND2xp5_ASAP7_75t_L g7462 ( 
.A(n_7322),
.B(n_6436),
.Y(n_7462)
);

NAND2x1_ASAP7_75t_L g7463 ( 
.A(n_7312),
.B(n_6443),
.Y(n_7463)
);

INVx3_ASAP7_75t_L g7464 ( 
.A(n_7229),
.Y(n_7464)
);

OR2x2_ASAP7_75t_L g7465 ( 
.A(n_7379),
.B(n_6444),
.Y(n_7465)
);

OAI22xp5_ASAP7_75t_L g7466 ( 
.A1(n_7339),
.A2(n_6445),
.B1(n_6449),
.B2(n_6444),
.Y(n_7466)
);

NAND2xp5_ASAP7_75t_L g7467 ( 
.A(n_7280),
.B(n_6445),
.Y(n_7467)
);

INVx1_ASAP7_75t_L g7468 ( 
.A(n_7267),
.Y(n_7468)
);

NOR2xp67_ASAP7_75t_L g7469 ( 
.A(n_7350),
.B(n_6449),
.Y(n_7469)
);

INVx2_ASAP7_75t_L g7470 ( 
.A(n_7311),
.Y(n_7470)
);

INVx2_ASAP7_75t_L g7471 ( 
.A(n_7372),
.Y(n_7471)
);

NAND2xp5_ASAP7_75t_L g7472 ( 
.A(n_7379),
.B(n_6457),
.Y(n_7472)
);

AOI22xp33_ASAP7_75t_L g7473 ( 
.A1(n_7353),
.A2(n_6163),
.B1(n_6172),
.B2(n_6168),
.Y(n_7473)
);

INVx1_ASAP7_75t_L g7474 ( 
.A(n_7334),
.Y(n_7474)
);

O2A1O1Ixp33_ASAP7_75t_L g7475 ( 
.A1(n_7258),
.A2(n_6464),
.B(n_6457),
.C(n_6463),
.Y(n_7475)
);

INVx2_ASAP7_75t_SL g7476 ( 
.A(n_7261),
.Y(n_7476)
);

INVx1_ASAP7_75t_L g7477 ( 
.A(n_7278),
.Y(n_7477)
);

NAND2xp5_ASAP7_75t_L g7478 ( 
.A(n_7339),
.B(n_6458),
.Y(n_7478)
);

OR2x2_ASAP7_75t_L g7479 ( 
.A(n_7302),
.B(n_6458),
.Y(n_7479)
);

OAI221xp5_ASAP7_75t_L g7480 ( 
.A1(n_7337),
.A2(n_6466),
.B1(n_6477),
.B2(n_6468),
.C(n_6463),
.Y(n_7480)
);

OAI32xp33_ASAP7_75t_L g7481 ( 
.A1(n_7258),
.A2(n_6481),
.A3(n_6508),
.B1(n_6244),
.B2(n_6162),
.Y(n_7481)
);

OAI21xp5_ASAP7_75t_L g7482 ( 
.A1(n_7221),
.A2(n_7347),
.B(n_7307),
.Y(n_7482)
);

NAND3xp33_ASAP7_75t_L g7483 ( 
.A(n_7355),
.B(n_6508),
.C(n_6481),
.Y(n_7483)
);

AOI21xp33_ASAP7_75t_L g7484 ( 
.A1(n_7270),
.A2(n_6228),
.B(n_6179),
.Y(n_7484)
);

OAI21xp5_ASAP7_75t_SL g7485 ( 
.A1(n_7270),
.A2(n_6266),
.B(n_6256),
.Y(n_7485)
);

OAI22xp5_ASAP7_75t_L g7486 ( 
.A1(n_7239),
.A2(n_5819),
.B1(n_5829),
.B2(n_5785),
.Y(n_7486)
);

NAND2xp5_ASAP7_75t_L g7487 ( 
.A(n_7364),
.B(n_5814),
.Y(n_7487)
);

O2A1O1Ixp5_ASAP7_75t_L g7488 ( 
.A1(n_7318),
.A2(n_6228),
.B(n_6230),
.C(n_6179),
.Y(n_7488)
);

OR2x2_ASAP7_75t_L g7489 ( 
.A(n_7300),
.B(n_5815),
.Y(n_7489)
);

INVx1_ASAP7_75t_L g7490 ( 
.A(n_7249),
.Y(n_7490)
);

NOR2xp33_ASAP7_75t_L g7491 ( 
.A(n_7377),
.B(n_4840),
.Y(n_7491)
);

INVx1_ASAP7_75t_L g7492 ( 
.A(n_7249),
.Y(n_7492)
);

AOI22xp5_ASAP7_75t_L g7493 ( 
.A1(n_7295),
.A2(n_6230),
.B1(n_6240),
.B2(n_6232),
.Y(n_7493)
);

NOR2xp33_ASAP7_75t_L g7494 ( 
.A(n_7377),
.B(n_5877),
.Y(n_7494)
);

AOI21xp33_ASAP7_75t_L g7495 ( 
.A1(n_7351),
.A2(n_6240),
.B(n_6232),
.Y(n_7495)
);

INVx1_ASAP7_75t_L g7496 ( 
.A(n_7351),
.Y(n_7496)
);

NAND2xp5_ASAP7_75t_L g7497 ( 
.A(n_7271),
.B(n_5892),
.Y(n_7497)
);

INVx2_ASAP7_75t_L g7498 ( 
.A(n_7319),
.Y(n_7498)
);

INVx2_ASAP7_75t_L g7499 ( 
.A(n_7268),
.Y(n_7499)
);

INVx1_ASAP7_75t_SL g7500 ( 
.A(n_7295),
.Y(n_7500)
);

NOR2xp67_ASAP7_75t_SL g7501 ( 
.A(n_7231),
.B(n_5014),
.Y(n_7501)
);

OAI221xp5_ASAP7_75t_SL g7502 ( 
.A1(n_7272),
.A2(n_6182),
.B1(n_6250),
.B2(n_6206),
.C(n_6261),
.Y(n_7502)
);

AOI22xp33_ASAP7_75t_SL g7503 ( 
.A1(n_7360),
.A2(n_6261),
.B1(n_6273),
.B2(n_6252),
.Y(n_7503)
);

AND2x2_ASAP7_75t_L g7504 ( 
.A(n_7327),
.B(n_5916),
.Y(n_7504)
);

NOR3xp33_ASAP7_75t_SL g7505 ( 
.A(n_7290),
.B(n_6216),
.C(n_6248),
.Y(n_7505)
);

OAI22xp5_ASAP7_75t_L g7506 ( 
.A1(n_7288),
.A2(n_7257),
.B1(n_7294),
.B2(n_7371),
.Y(n_7506)
);

INVx1_ASAP7_75t_L g7507 ( 
.A(n_7368),
.Y(n_7507)
);

OAI322xp33_ASAP7_75t_L g7508 ( 
.A1(n_7303),
.A2(n_5901),
.A3(n_5933),
.B1(n_5905),
.B2(n_5906),
.C1(n_5823),
.C2(n_5885),
.Y(n_7508)
);

NAND2x1p5_ASAP7_75t_L g7509 ( 
.A(n_7371),
.B(n_4832),
.Y(n_7509)
);

AOI22xp5_ASAP7_75t_L g7510 ( 
.A1(n_7357),
.A2(n_6134),
.B1(n_5716),
.B2(n_5742),
.Y(n_7510)
);

AND2x2_ASAP7_75t_L g7511 ( 
.A(n_7260),
.B(n_5918),
.Y(n_7511)
);

AOI22xp5_ASAP7_75t_L g7512 ( 
.A1(n_7361),
.A2(n_7360),
.B1(n_7265),
.B2(n_7376),
.Y(n_7512)
);

OAI32xp33_ASAP7_75t_L g7513 ( 
.A1(n_7335),
.A2(n_5829),
.A3(n_5832),
.B1(n_5819),
.B2(n_5785),
.Y(n_7513)
);

INVx1_ASAP7_75t_L g7514 ( 
.A(n_7247),
.Y(n_7514)
);

NOR2xp33_ASAP7_75t_L g7515 ( 
.A(n_7356),
.B(n_5923),
.Y(n_7515)
);

OR2x2_ASAP7_75t_L g7516 ( 
.A(n_7259),
.B(n_5928),
.Y(n_7516)
);

INVx1_ASAP7_75t_L g7517 ( 
.A(n_7283),
.Y(n_7517)
);

INVx1_ASAP7_75t_L g7518 ( 
.A(n_7320),
.Y(n_7518)
);

NAND2xp5_ASAP7_75t_L g7519 ( 
.A(n_7244),
.B(n_5930),
.Y(n_7519)
);

NAND2xp5_ASAP7_75t_L g7520 ( 
.A(n_7331),
.B(n_5832),
.Y(n_7520)
);

OAI221xp5_ASAP7_75t_L g7521 ( 
.A1(n_7380),
.A2(n_6227),
.B1(n_6238),
.B2(n_6218),
.C(n_6208),
.Y(n_7521)
);

INVx1_ASAP7_75t_L g7522 ( 
.A(n_7213),
.Y(n_7522)
);

OR2x2_ASAP7_75t_L g7523 ( 
.A(n_7217),
.B(n_5837),
.Y(n_7523)
);

INVx1_ASAP7_75t_L g7524 ( 
.A(n_7358),
.Y(n_7524)
);

AND2x2_ASAP7_75t_L g7525 ( 
.A(n_7329),
.B(n_5402),
.Y(n_7525)
);

BUFx2_ASAP7_75t_L g7526 ( 
.A(n_7356),
.Y(n_7526)
);

NOR2xp33_ASAP7_75t_L g7527 ( 
.A(n_7284),
.B(n_5837),
.Y(n_7527)
);

AOI221xp5_ASAP7_75t_L g7528 ( 
.A1(n_7375),
.A2(n_6227),
.B1(n_6238),
.B2(n_6218),
.C(n_6208),
.Y(n_7528)
);

NAND3xp33_ASAP7_75t_L g7529 ( 
.A(n_7304),
.B(n_6259),
.C(n_6251),
.Y(n_7529)
);

XNOR2xp5_ASAP7_75t_L g7530 ( 
.A(n_7387),
.B(n_7326),
.Y(n_7530)
);

NOR2x1p5_ASAP7_75t_L g7531 ( 
.A(n_7406),
.B(n_7435),
.Y(n_7531)
);

OAI22xp5_ASAP7_75t_L g7532 ( 
.A1(n_7387),
.A2(n_7298),
.B1(n_7269),
.B2(n_7243),
.Y(n_7532)
);

OAI222xp33_ASAP7_75t_L g7533 ( 
.A1(n_7418),
.A2(n_7333),
.B1(n_7375),
.B2(n_7225),
.C1(n_7362),
.C2(n_7226),
.Y(n_7533)
);

AOI221x1_ASAP7_75t_L g7534 ( 
.A1(n_7390),
.A2(n_7381),
.B1(n_7359),
.B2(n_7363),
.C(n_7301),
.Y(n_7534)
);

AOI221xp5_ASAP7_75t_L g7535 ( 
.A1(n_7390),
.A2(n_7378),
.B1(n_7343),
.B2(n_7342),
.C(n_7373),
.Y(n_7535)
);

NAND2xp33_ASAP7_75t_L g7536 ( 
.A(n_7404),
.B(n_7248),
.Y(n_7536)
);

NAND2xp5_ASAP7_75t_SL g7537 ( 
.A(n_7400),
.B(n_7340),
.Y(n_7537)
);

INVx1_ASAP7_75t_L g7538 ( 
.A(n_7393),
.Y(n_7538)
);

NAND2xp5_ASAP7_75t_L g7539 ( 
.A(n_7404),
.B(n_7336),
.Y(n_7539)
);

AOI21xp33_ASAP7_75t_SL g7540 ( 
.A1(n_7400),
.A2(n_7291),
.B(n_7344),
.Y(n_7540)
);

NAND3xp33_ASAP7_75t_L g7541 ( 
.A(n_7456),
.B(n_7253),
.C(n_7352),
.Y(n_7541)
);

INVx1_ASAP7_75t_L g7542 ( 
.A(n_7418),
.Y(n_7542)
);

OR2x2_ASAP7_75t_L g7543 ( 
.A(n_7500),
.B(n_7382),
.Y(n_7543)
);

OR2x2_ASAP7_75t_L g7544 ( 
.A(n_7398),
.B(n_7332),
.Y(n_7544)
);

AOI22xp5_ASAP7_75t_L g7545 ( 
.A1(n_7445),
.A2(n_7285),
.B1(n_7234),
.B2(n_7236),
.Y(n_7545)
);

AOI21xp5_ASAP7_75t_L g7546 ( 
.A1(n_7445),
.A2(n_7342),
.B(n_7348),
.Y(n_7546)
);

AOI21xp5_ASAP7_75t_L g7547 ( 
.A1(n_7405),
.A2(n_7383),
.B(n_7374),
.Y(n_7547)
);

INVxp67_ASAP7_75t_L g7548 ( 
.A(n_7424),
.Y(n_7548)
);

INVx2_ASAP7_75t_L g7549 ( 
.A(n_7509),
.Y(n_7549)
);

INVx2_ASAP7_75t_L g7550 ( 
.A(n_7509),
.Y(n_7550)
);

OAI22xp33_ASAP7_75t_L g7551 ( 
.A1(n_7386),
.A2(n_7384),
.B1(n_7366),
.B2(n_7218),
.Y(n_7551)
);

INVxp67_ASAP7_75t_L g7552 ( 
.A(n_7526),
.Y(n_7552)
);

INVx1_ASAP7_75t_L g7553 ( 
.A(n_7411),
.Y(n_7553)
);

NOR2xp33_ASAP7_75t_L g7554 ( 
.A(n_7391),
.B(n_7441),
.Y(n_7554)
);

AOI221xp5_ASAP7_75t_L g7555 ( 
.A1(n_7484),
.A2(n_7305),
.B1(n_7317),
.B2(n_7328),
.C(n_7309),
.Y(n_7555)
);

INVx2_ASAP7_75t_L g7556 ( 
.A(n_7443),
.Y(n_7556)
);

OAI22xp5_ASAP7_75t_L g7557 ( 
.A1(n_7429),
.A2(n_7330),
.B1(n_7341),
.B2(n_7286),
.Y(n_7557)
);

AND2x2_ASAP7_75t_L g7558 ( 
.A(n_7525),
.B(n_7345),
.Y(n_7558)
);

AND2x2_ASAP7_75t_L g7559 ( 
.A(n_7412),
.B(n_7287),
.Y(n_7559)
);

INVx1_ASAP7_75t_L g7560 ( 
.A(n_7453),
.Y(n_7560)
);

OAI21xp5_ASAP7_75t_L g7561 ( 
.A1(n_7482),
.A2(n_7299),
.B(n_5842),
.Y(n_7561)
);

NOR2xp33_ASAP7_75t_SL g7562 ( 
.A(n_7432),
.B(n_4832),
.Y(n_7562)
);

INVx2_ASAP7_75t_SL g7563 ( 
.A(n_7401),
.Y(n_7563)
);

AOI211xp5_ASAP7_75t_L g7564 ( 
.A1(n_7396),
.A2(n_5839),
.B(n_5844),
.C(n_5842),
.Y(n_7564)
);

OAI21xp5_ASAP7_75t_L g7565 ( 
.A1(n_7413),
.A2(n_5844),
.B(n_5839),
.Y(n_7565)
);

OAI211xp5_ASAP7_75t_SL g7566 ( 
.A1(n_7442),
.A2(n_6259),
.B(n_6251),
.C(n_5847),
.Y(n_7566)
);

OR2x2_ASAP7_75t_L g7567 ( 
.A(n_7407),
.B(n_5845),
.Y(n_7567)
);

AOI21xp5_ASAP7_75t_L g7568 ( 
.A1(n_7452),
.A2(n_5847),
.B(n_5845),
.Y(n_7568)
);

NAND2xp5_ASAP7_75t_L g7569 ( 
.A(n_7423),
.B(n_5849),
.Y(n_7569)
);

OAI221xp5_ASAP7_75t_SL g7570 ( 
.A1(n_7395),
.A2(n_5716),
.B1(n_5750),
.B2(n_5742),
.C(n_5710),
.Y(n_7570)
);

INVx1_ASAP7_75t_L g7571 ( 
.A(n_7420),
.Y(n_7571)
);

AOI22xp33_ASAP7_75t_SL g7572 ( 
.A1(n_7529),
.A2(n_5750),
.B1(n_5757),
.B2(n_5710),
.Y(n_7572)
);

NOR2xp33_ASAP7_75t_L g7573 ( 
.A(n_7446),
.B(n_5849),
.Y(n_7573)
);

INVx1_ASAP7_75t_L g7574 ( 
.A(n_7430),
.Y(n_7574)
);

AND2x2_ASAP7_75t_L g7575 ( 
.A(n_7421),
.B(n_5850),
.Y(n_7575)
);

INVxp67_ASAP7_75t_L g7576 ( 
.A(n_7449),
.Y(n_7576)
);

INVx1_ASAP7_75t_SL g7577 ( 
.A(n_7455),
.Y(n_7577)
);

NAND2xp5_ASAP7_75t_L g7578 ( 
.A(n_7471),
.B(n_7476),
.Y(n_7578)
);

OAI21xp33_ASAP7_75t_SL g7579 ( 
.A1(n_7403),
.A2(n_5855),
.B(n_5850),
.Y(n_7579)
);

OAI21xp5_ASAP7_75t_L g7580 ( 
.A1(n_7428),
.A2(n_5858),
.B(n_5855),
.Y(n_7580)
);

AND2x2_ASAP7_75t_L g7581 ( 
.A(n_7416),
.B(n_5858),
.Y(n_7581)
);

INVx2_ASAP7_75t_L g7582 ( 
.A(n_7479),
.Y(n_7582)
);

NOR2xp33_ASAP7_75t_L g7583 ( 
.A(n_7451),
.B(n_7454),
.Y(n_7583)
);

OAI22xp5_ASAP7_75t_L g7584 ( 
.A1(n_7439),
.A2(n_5915),
.B1(n_5934),
.B2(n_5913),
.Y(n_7584)
);

AOI22x1_ASAP7_75t_L g7585 ( 
.A1(n_7399),
.A2(n_5915),
.B1(n_5934),
.B2(n_5913),
.Y(n_7585)
);

INVx2_ASAP7_75t_L g7586 ( 
.A(n_7465),
.Y(n_7586)
);

AOI22xp33_ASAP7_75t_L g7587 ( 
.A1(n_7528),
.A2(n_5769),
.B1(n_5795),
.B2(n_5757),
.Y(n_7587)
);

NAND2xp5_ASAP7_75t_L g7588 ( 
.A(n_7437),
.B(n_5866),
.Y(n_7588)
);

OAI21xp33_ASAP7_75t_SL g7589 ( 
.A1(n_7434),
.A2(n_5867),
.B(n_5866),
.Y(n_7589)
);

AND2x2_ASAP7_75t_L g7590 ( 
.A(n_7394),
.B(n_5867),
.Y(n_7590)
);

INVxp33_ASAP7_75t_L g7591 ( 
.A(n_7491),
.Y(n_7591)
);

NAND2xp5_ASAP7_75t_L g7592 ( 
.A(n_7388),
.B(n_5870),
.Y(n_7592)
);

AND2x2_ASAP7_75t_L g7593 ( 
.A(n_7450),
.B(n_5870),
.Y(n_7593)
);

NAND4xp25_ASAP7_75t_L g7594 ( 
.A(n_7389),
.B(n_5114),
.C(n_4729),
.D(n_5873),
.Y(n_7594)
);

INVx2_ASAP7_75t_SL g7595 ( 
.A(n_7463),
.Y(n_7595)
);

INVx1_ASAP7_75t_L g7596 ( 
.A(n_7444),
.Y(n_7596)
);

NAND2xp5_ASAP7_75t_L g7597 ( 
.A(n_7518),
.B(n_5873),
.Y(n_7597)
);

OR2x2_ASAP7_75t_L g7598 ( 
.A(n_7459),
.B(n_5874),
.Y(n_7598)
);

INVxp67_ASAP7_75t_L g7599 ( 
.A(n_7392),
.Y(n_7599)
);

INVx3_ASAP7_75t_L g7600 ( 
.A(n_7499),
.Y(n_7600)
);

AOI22xp5_ASAP7_75t_L g7601 ( 
.A1(n_7496),
.A2(n_5834),
.B1(n_5795),
.B2(n_5813),
.Y(n_7601)
);

OR2x2_ASAP7_75t_L g7602 ( 
.A(n_7422),
.B(n_5874),
.Y(n_7602)
);

CKINVDCx16_ASAP7_75t_R g7603 ( 
.A(n_7506),
.Y(n_7603)
);

AOI32xp33_ASAP7_75t_L g7604 ( 
.A1(n_7474),
.A2(n_5938),
.A3(n_5937),
.B1(n_5896),
.B2(n_5813),
.Y(n_7604)
);

AND2x4_ASAP7_75t_L g7605 ( 
.A(n_7498),
.B(n_7457),
.Y(n_7605)
);

OR2x2_ASAP7_75t_L g7606 ( 
.A(n_7414),
.B(n_5896),
.Y(n_7606)
);

OAI221xp5_ASAP7_75t_L g7607 ( 
.A1(n_7512),
.A2(n_5938),
.B1(n_5937),
.B2(n_5769),
.C(n_5834),
.Y(n_7607)
);

INVx1_ASAP7_75t_SL g7608 ( 
.A(n_7415),
.Y(n_7608)
);

OAI22xp5_ASAP7_75t_L g7609 ( 
.A1(n_7468),
.A2(n_5396),
.B1(n_5405),
.B2(n_5390),
.Y(n_7609)
);

NAND2xp33_ASAP7_75t_SL g7610 ( 
.A(n_7501),
.B(n_4931),
.Y(n_7610)
);

A2O1A1Ixp33_ASAP7_75t_L g7611 ( 
.A1(n_7529),
.A2(n_5823),
.B(n_5840),
.C(n_5825),
.Y(n_7611)
);

INVx1_ASAP7_75t_L g7612 ( 
.A(n_7433),
.Y(n_7612)
);

NAND2xp5_ASAP7_75t_L g7613 ( 
.A(n_7461),
.B(n_7410),
.Y(n_7613)
);

AOI22xp33_ASAP7_75t_L g7614 ( 
.A1(n_7521),
.A2(n_5936),
.B1(n_5840),
.B2(n_5853),
.Y(n_7614)
);

OAI21xp33_ASAP7_75t_L g7615 ( 
.A1(n_7485),
.A2(n_5853),
.B(n_5825),
.Y(n_7615)
);

OAI321xp33_ASAP7_75t_L g7616 ( 
.A1(n_7502),
.A2(n_5885),
.A3(n_5872),
.B1(n_5907),
.B2(n_5894),
.C(n_5863),
.Y(n_7616)
);

AOI211xp5_ASAP7_75t_L g7617 ( 
.A1(n_7481),
.A2(n_5014),
.B(n_5936),
.C(n_5872),
.Y(n_7617)
);

NAND2x1p5_ASAP7_75t_L g7618 ( 
.A(n_7417),
.B(n_4832),
.Y(n_7618)
);

NAND3xp33_ASAP7_75t_L g7619 ( 
.A(n_7425),
.B(n_5894),
.C(n_5863),
.Y(n_7619)
);

OAI221xp5_ASAP7_75t_L g7620 ( 
.A1(n_7467),
.A2(n_5907),
.B1(n_5924),
.B2(n_5912),
.C(n_5911),
.Y(n_7620)
);

OR2x2_ASAP7_75t_L g7621 ( 
.A(n_7462),
.B(n_5373),
.Y(n_7621)
);

OAI22xp5_ASAP7_75t_L g7622 ( 
.A1(n_7477),
.A2(n_7507),
.B1(n_7409),
.B2(n_7524),
.Y(n_7622)
);

AOI22xp5_ASAP7_75t_L g7623 ( 
.A1(n_7427),
.A2(n_5912),
.B1(n_5924),
.B2(n_5911),
.Y(n_7623)
);

NAND2xp5_ASAP7_75t_L g7624 ( 
.A(n_7436),
.B(n_7493),
.Y(n_7624)
);

AOI22xp5_ASAP7_75t_SL g7625 ( 
.A1(n_7448),
.A2(n_5014),
.B1(n_5453),
.B2(n_5425),
.Y(n_7625)
);

INVx2_ASAP7_75t_L g7626 ( 
.A(n_7489),
.Y(n_7626)
);

INVx1_ASAP7_75t_L g7627 ( 
.A(n_7478),
.Y(n_7627)
);

INVx1_ASAP7_75t_L g7628 ( 
.A(n_7472),
.Y(n_7628)
);

O2A1O1Ixp5_ASAP7_75t_L g7629 ( 
.A1(n_7458),
.A2(n_5931),
.B(n_5935),
.C(n_5365),
.Y(n_7629)
);

NOR2xp33_ASAP7_75t_L g7630 ( 
.A(n_7490),
.B(n_5931),
.Y(n_7630)
);

INVx2_ASAP7_75t_L g7631 ( 
.A(n_7464),
.Y(n_7631)
);

AND2x2_ASAP7_75t_SL g7632 ( 
.A(n_7514),
.B(n_5014),
.Y(n_7632)
);

NAND2xp5_ASAP7_75t_L g7633 ( 
.A(n_7492),
.B(n_7469),
.Y(n_7633)
);

AOI21xp33_ASAP7_75t_L g7634 ( 
.A1(n_7470),
.A2(n_5935),
.B(n_5499),
.Y(n_7634)
);

OAI32xp33_ASAP7_75t_L g7635 ( 
.A1(n_7516),
.A2(n_5424),
.A3(n_5373),
.B1(n_5474),
.B2(n_5452),
.Y(n_7635)
);

INVx1_ASAP7_75t_L g7636 ( 
.A(n_7427),
.Y(n_7636)
);

INVx1_ASAP7_75t_L g7637 ( 
.A(n_7487),
.Y(n_7637)
);

NAND2xp5_ASAP7_75t_L g7638 ( 
.A(n_7464),
.B(n_5406),
.Y(n_7638)
);

OAI211xp5_ASAP7_75t_L g7639 ( 
.A1(n_7485),
.A2(n_4969),
.B(n_4982),
.C(n_5005),
.Y(n_7639)
);

OAI21xp33_ASAP7_75t_L g7640 ( 
.A1(n_7517),
.A2(n_5024),
.B(n_5365),
.Y(n_7640)
);

INVx1_ASAP7_75t_L g7641 ( 
.A(n_7483),
.Y(n_7641)
);

INVx1_ASAP7_75t_L g7642 ( 
.A(n_7483),
.Y(n_7642)
);

OR2x2_ASAP7_75t_L g7643 ( 
.A(n_7402),
.B(n_5424),
.Y(n_7643)
);

OR2x2_ASAP7_75t_L g7644 ( 
.A(n_7397),
.B(n_5474),
.Y(n_7644)
);

OAI22xp5_ASAP7_75t_L g7645 ( 
.A1(n_7419),
.A2(n_5409),
.B1(n_5417),
.B2(n_5411),
.Y(n_7645)
);

INVx1_ASAP7_75t_L g7646 ( 
.A(n_7488),
.Y(n_7646)
);

AOI22xp5_ASAP7_75t_L g7647 ( 
.A1(n_7408),
.A2(n_5499),
.B1(n_5500),
.B2(n_5486),
.Y(n_7647)
);

INVx1_ASAP7_75t_L g7648 ( 
.A(n_7520),
.Y(n_7648)
);

OR2x2_ASAP7_75t_L g7649 ( 
.A(n_7522),
.B(n_5590),
.Y(n_7649)
);

INVx1_ASAP7_75t_L g7650 ( 
.A(n_7466),
.Y(n_7650)
);

OAI22xp33_ASAP7_75t_SL g7651 ( 
.A1(n_7460),
.A2(n_5500),
.B1(n_5505),
.B2(n_5486),
.Y(n_7651)
);

NAND2xp5_ASAP7_75t_L g7652 ( 
.A(n_7504),
.B(n_7431),
.Y(n_7652)
);

NAND2xp5_ASAP7_75t_SL g7653 ( 
.A(n_7440),
.B(n_5425),
.Y(n_7653)
);

OAI32xp33_ASAP7_75t_L g7654 ( 
.A1(n_7519),
.A2(n_5127),
.A3(n_5002),
.B1(n_4906),
.B2(n_4930),
.Y(n_7654)
);

INVx1_ASAP7_75t_L g7655 ( 
.A(n_7515),
.Y(n_7655)
);

AOI221xp5_ASAP7_75t_L g7656 ( 
.A1(n_7495),
.A2(n_7426),
.B1(n_7508),
.B2(n_7480),
.C(n_7447),
.Y(n_7656)
);

NOR2xp33_ASAP7_75t_L g7657 ( 
.A(n_7508),
.B(n_7497),
.Y(n_7657)
);

NAND2xp5_ASAP7_75t_L g7658 ( 
.A(n_7511),
.B(n_5409),
.Y(n_7658)
);

NAND2xp5_ASAP7_75t_L g7659 ( 
.A(n_7527),
.B(n_5411),
.Y(n_7659)
);

AND2x2_ASAP7_75t_L g7660 ( 
.A(n_7603),
.B(n_7494),
.Y(n_7660)
);

NOR2xp33_ASAP7_75t_L g7661 ( 
.A(n_7548),
.B(n_7523),
.Y(n_7661)
);

INVx1_ASAP7_75t_L g7662 ( 
.A(n_7636),
.Y(n_7662)
);

AOI22xp33_ASAP7_75t_L g7663 ( 
.A1(n_7542),
.A2(n_7473),
.B1(n_7503),
.B2(n_7510),
.Y(n_7663)
);

NAND2xp5_ASAP7_75t_L g7664 ( 
.A(n_7600),
.B(n_7577),
.Y(n_7664)
);

NAND2xp5_ASAP7_75t_L g7665 ( 
.A(n_7600),
.B(n_7505),
.Y(n_7665)
);

OR2x2_ASAP7_75t_L g7666 ( 
.A(n_7543),
.B(n_7486),
.Y(n_7666)
);

AND2x4_ASAP7_75t_L g7667 ( 
.A(n_7563),
.B(n_7475),
.Y(n_7667)
);

HB1xp67_ASAP7_75t_L g7668 ( 
.A(n_7530),
.Y(n_7668)
);

AND2x2_ASAP7_75t_L g7669 ( 
.A(n_7558),
.B(n_7559),
.Y(n_7669)
);

AND2x2_ASAP7_75t_L g7670 ( 
.A(n_7556),
.B(n_7438),
.Y(n_7670)
);

INVx1_ASAP7_75t_SL g7671 ( 
.A(n_7544),
.Y(n_7671)
);

AOI22xp33_ASAP7_75t_L g7672 ( 
.A1(n_7566),
.A2(n_5514),
.B1(n_5521),
.B2(n_5505),
.Y(n_7672)
);

BUFx2_ASAP7_75t_L g7673 ( 
.A(n_7605),
.Y(n_7673)
);

NAND2x1_ASAP7_75t_SL g7674 ( 
.A(n_7605),
.B(n_7582),
.Y(n_7674)
);

OR2x2_ASAP7_75t_L g7675 ( 
.A(n_7539),
.B(n_7537),
.Y(n_7675)
);

INVx1_ASAP7_75t_L g7676 ( 
.A(n_7536),
.Y(n_7676)
);

INVx1_ASAP7_75t_L g7677 ( 
.A(n_7578),
.Y(n_7677)
);

INVx1_ASAP7_75t_L g7678 ( 
.A(n_7652),
.Y(n_7678)
);

INVx1_ASAP7_75t_SL g7679 ( 
.A(n_7608),
.Y(n_7679)
);

AND2x4_ASAP7_75t_L g7680 ( 
.A(n_7595),
.B(n_5425),
.Y(n_7680)
);

INVx1_ASAP7_75t_L g7681 ( 
.A(n_7531),
.Y(n_7681)
);

INVx1_ASAP7_75t_L g7682 ( 
.A(n_7560),
.Y(n_7682)
);

NAND2xp5_ASAP7_75t_L g7683 ( 
.A(n_7546),
.B(n_7513),
.Y(n_7683)
);

NOR2xp33_ASAP7_75t_L g7684 ( 
.A(n_7533),
.B(n_5425),
.Y(n_7684)
);

AND2x2_ASAP7_75t_L g7685 ( 
.A(n_7586),
.B(n_5453),
.Y(n_7685)
);

AND2x2_ASAP7_75t_L g7686 ( 
.A(n_7554),
.B(n_5453),
.Y(n_7686)
);

NOR2xp33_ASAP7_75t_L g7687 ( 
.A(n_7540),
.B(n_5453),
.Y(n_7687)
);

AND2x4_ASAP7_75t_L g7688 ( 
.A(n_7626),
.B(n_5471),
.Y(n_7688)
);

NOR2xp33_ASAP7_75t_L g7689 ( 
.A(n_7553),
.B(n_5471),
.Y(n_7689)
);

NAND2xp5_ASAP7_75t_L g7690 ( 
.A(n_7547),
.B(n_5417),
.Y(n_7690)
);

INVx1_ASAP7_75t_SL g7691 ( 
.A(n_7624),
.Y(n_7691)
);

NOR2xp33_ASAP7_75t_L g7692 ( 
.A(n_7541),
.B(n_5471),
.Y(n_7692)
);

INVx2_ASAP7_75t_L g7693 ( 
.A(n_7618),
.Y(n_7693)
);

OR2x2_ASAP7_75t_L g7694 ( 
.A(n_7613),
.B(n_5590),
.Y(n_7694)
);

INVx1_ASAP7_75t_L g7695 ( 
.A(n_7641),
.Y(n_7695)
);

INVx1_ASAP7_75t_L g7696 ( 
.A(n_7642),
.Y(n_7696)
);

OAI21xp5_ASAP7_75t_SL g7697 ( 
.A1(n_7535),
.A2(n_5511),
.B(n_5471),
.Y(n_7697)
);

AND2x2_ASAP7_75t_L g7698 ( 
.A(n_7571),
.B(n_5511),
.Y(n_7698)
);

OAI22xp5_ASAP7_75t_L g7699 ( 
.A1(n_7545),
.A2(n_5599),
.B1(n_5422),
.B2(n_5426),
.Y(n_7699)
);

NOR2x1_ASAP7_75t_L g7700 ( 
.A(n_7551),
.B(n_5419),
.Y(n_7700)
);

AND2x2_ASAP7_75t_L g7701 ( 
.A(n_7625),
.B(n_5511),
.Y(n_7701)
);

NOR2xp33_ASAP7_75t_L g7702 ( 
.A(n_7599),
.B(n_5511),
.Y(n_7702)
);

NOR2xp33_ASAP7_75t_L g7703 ( 
.A(n_7538),
.B(n_5419),
.Y(n_7703)
);

INVx2_ASAP7_75t_L g7704 ( 
.A(n_7567),
.Y(n_7704)
);

INVx1_ASAP7_75t_L g7705 ( 
.A(n_7581),
.Y(n_7705)
);

OR2x2_ASAP7_75t_L g7706 ( 
.A(n_7532),
.B(n_5498),
.Y(n_7706)
);

NAND2xp5_ASAP7_75t_L g7707 ( 
.A(n_7632),
.B(n_5422),
.Y(n_7707)
);

INVx1_ASAP7_75t_L g7708 ( 
.A(n_7545),
.Y(n_7708)
);

NOR2xp33_ASAP7_75t_L g7709 ( 
.A(n_7576),
.B(n_5426),
.Y(n_7709)
);

NAND2xp5_ASAP7_75t_L g7710 ( 
.A(n_7575),
.B(n_5428),
.Y(n_7710)
);

NAND2xp5_ASAP7_75t_L g7711 ( 
.A(n_7646),
.B(n_7593),
.Y(n_7711)
);

NOR2xp33_ASAP7_75t_L g7712 ( 
.A(n_7615),
.B(n_5428),
.Y(n_7712)
);

INVx1_ASAP7_75t_L g7713 ( 
.A(n_7631),
.Y(n_7713)
);

AOI221x1_ASAP7_75t_SL g7714 ( 
.A1(n_7557),
.A2(n_5599),
.B1(n_5434),
.B2(n_5435),
.C(n_5432),
.Y(n_7714)
);

INVxp67_ASAP7_75t_SL g7715 ( 
.A(n_7633),
.Y(n_7715)
);

AOI21xp5_ASAP7_75t_L g7716 ( 
.A1(n_7653),
.A2(n_5432),
.B(n_5429),
.Y(n_7716)
);

AND2x2_ASAP7_75t_L g7717 ( 
.A(n_7552),
.B(n_7596),
.Y(n_7717)
);

NAND2xp5_ASAP7_75t_L g7718 ( 
.A(n_7534),
.B(n_5429),
.Y(n_7718)
);

OR2x2_ASAP7_75t_L g7719 ( 
.A(n_7644),
.B(n_5434),
.Y(n_7719)
);

OR2x2_ASAP7_75t_L g7720 ( 
.A(n_7643),
.B(n_5435),
.Y(n_7720)
);

INVx1_ASAP7_75t_L g7721 ( 
.A(n_7598),
.Y(n_7721)
);

OR2x2_ASAP7_75t_L g7722 ( 
.A(n_7621),
.B(n_5443),
.Y(n_7722)
);

NAND2xp5_ASAP7_75t_L g7723 ( 
.A(n_7590),
.B(n_5443),
.Y(n_7723)
);

INVx1_ASAP7_75t_L g7724 ( 
.A(n_7619),
.Y(n_7724)
);

INVxp67_ASAP7_75t_L g7725 ( 
.A(n_7562),
.Y(n_7725)
);

AND2x2_ASAP7_75t_L g7726 ( 
.A(n_7612),
.B(n_5117),
.Y(n_7726)
);

OR2x2_ASAP7_75t_L g7727 ( 
.A(n_7649),
.B(n_5457),
.Y(n_7727)
);

NAND2xp5_ASAP7_75t_L g7728 ( 
.A(n_7564),
.B(n_7574),
.Y(n_7728)
);

NAND2xp5_ASAP7_75t_L g7729 ( 
.A(n_7628),
.B(n_5457),
.Y(n_7729)
);

NAND2xp5_ASAP7_75t_L g7730 ( 
.A(n_7630),
.B(n_5462),
.Y(n_7730)
);

NAND2xp5_ASAP7_75t_L g7731 ( 
.A(n_7627),
.B(n_5462),
.Y(n_7731)
);

NAND2xp5_ASAP7_75t_L g7732 ( 
.A(n_7573),
.B(n_5466),
.Y(n_7732)
);

NAND2xp5_ASAP7_75t_L g7733 ( 
.A(n_7617),
.B(n_5466),
.Y(n_7733)
);

AND2x4_ASAP7_75t_L g7734 ( 
.A(n_7549),
.B(n_4832),
.Y(n_7734)
);

INVx2_ASAP7_75t_L g7735 ( 
.A(n_7606),
.Y(n_7735)
);

INVx1_ASAP7_75t_L g7736 ( 
.A(n_7615),
.Y(n_7736)
);

NOR2xp33_ASAP7_75t_L g7737 ( 
.A(n_7570),
.B(n_5468),
.Y(n_7737)
);

BUFx2_ASAP7_75t_L g7738 ( 
.A(n_7610),
.Y(n_7738)
);

INVx2_ASAP7_75t_L g7739 ( 
.A(n_7602),
.Y(n_7739)
);

AND2x4_ASAP7_75t_L g7740 ( 
.A(n_7550),
.B(n_5468),
.Y(n_7740)
);

AOI222xp33_ASAP7_75t_L g7741 ( 
.A1(n_7616),
.A2(n_5514),
.B1(n_5521),
.B2(n_5505),
.C1(n_5381),
.C2(n_5352),
.Y(n_7741)
);

NAND2xp5_ASAP7_75t_L g7742 ( 
.A(n_7648),
.B(n_5477),
.Y(n_7742)
);

INVxp67_ASAP7_75t_SL g7743 ( 
.A(n_7657),
.Y(n_7743)
);

INVx1_ASAP7_75t_L g7744 ( 
.A(n_7658),
.Y(n_7744)
);

NAND2xp5_ASAP7_75t_L g7745 ( 
.A(n_7655),
.B(n_7637),
.Y(n_7745)
);

AND2x2_ASAP7_75t_L g7746 ( 
.A(n_7583),
.B(n_5117),
.Y(n_7746)
);

INVxp67_ASAP7_75t_SL g7747 ( 
.A(n_7597),
.Y(n_7747)
);

NOR2xp33_ASAP7_75t_L g7748 ( 
.A(n_7622),
.B(n_5477),
.Y(n_7748)
);

INVx1_ASAP7_75t_L g7749 ( 
.A(n_7638),
.Y(n_7749)
);

NAND2xp5_ASAP7_75t_L g7750 ( 
.A(n_7568),
.B(n_5482),
.Y(n_7750)
);

NAND2xp5_ASAP7_75t_L g7751 ( 
.A(n_7656),
.B(n_5482),
.Y(n_7751)
);

INVx1_ASAP7_75t_L g7752 ( 
.A(n_7569),
.Y(n_7752)
);

INVx2_ASAP7_75t_L g7753 ( 
.A(n_7585),
.Y(n_7753)
);

INVx2_ASAP7_75t_L g7754 ( 
.A(n_7629),
.Y(n_7754)
);

NAND2x1_ASAP7_75t_SL g7755 ( 
.A(n_7650),
.B(n_5304),
.Y(n_7755)
);

INVx1_ASAP7_75t_L g7756 ( 
.A(n_7659),
.Y(n_7756)
);

INVx2_ASAP7_75t_L g7757 ( 
.A(n_7588),
.Y(n_7757)
);

NAND2x1p5_ASAP7_75t_L g7758 ( 
.A(n_7592),
.B(n_4906),
.Y(n_7758)
);

INVx1_ASAP7_75t_L g7759 ( 
.A(n_7623),
.Y(n_7759)
);

AND2x2_ASAP7_75t_L g7760 ( 
.A(n_7591),
.B(n_5304),
.Y(n_7760)
);

NOR2xp67_ASAP7_75t_L g7761 ( 
.A(n_7639),
.B(n_7594),
.Y(n_7761)
);

NAND2xp5_ASAP7_75t_L g7762 ( 
.A(n_7555),
.B(n_7561),
.Y(n_7762)
);

NOR2xp33_ASAP7_75t_L g7763 ( 
.A(n_7607),
.B(n_7579),
.Y(n_7763)
);

NAND2xp5_ASAP7_75t_L g7764 ( 
.A(n_7604),
.B(n_5492),
.Y(n_7764)
);

AND2x2_ASAP7_75t_L g7765 ( 
.A(n_7580),
.B(n_5304),
.Y(n_7765)
);

OR2x2_ASAP7_75t_L g7766 ( 
.A(n_7565),
.B(n_7645),
.Y(n_7766)
);

NAND2xp5_ASAP7_75t_L g7767 ( 
.A(n_7640),
.B(n_5492),
.Y(n_7767)
);

INVxp67_ASAP7_75t_L g7768 ( 
.A(n_7601),
.Y(n_7768)
);

INVx1_ASAP7_75t_L g7769 ( 
.A(n_7623),
.Y(n_7769)
);

NAND2xp5_ASAP7_75t_L g7770 ( 
.A(n_7614),
.B(n_5493),
.Y(n_7770)
);

AOI21xp5_ASAP7_75t_L g7771 ( 
.A1(n_7664),
.A2(n_7579),
.B(n_7589),
.Y(n_7771)
);

NAND3xp33_ASAP7_75t_L g7772 ( 
.A(n_7673),
.B(n_7572),
.C(n_7587),
.Y(n_7772)
);

NAND3xp33_ASAP7_75t_L g7773 ( 
.A(n_7708),
.B(n_7611),
.C(n_7601),
.Y(n_7773)
);

NOR3xp33_ASAP7_75t_L g7774 ( 
.A(n_7660),
.B(n_7634),
.C(n_7589),
.Y(n_7774)
);

AOI21xp5_ASAP7_75t_L g7775 ( 
.A1(n_7671),
.A2(n_7584),
.B(n_7609),
.Y(n_7775)
);

INVx1_ASAP7_75t_L g7776 ( 
.A(n_7674),
.Y(n_7776)
);

AOI211xp5_ASAP7_75t_L g7777 ( 
.A1(n_7671),
.A2(n_7651),
.B(n_7635),
.C(n_7620),
.Y(n_7777)
);

NOR4xp25_ASAP7_75t_SL g7778 ( 
.A(n_7738),
.B(n_7654),
.C(n_7647),
.D(n_4950),
.Y(n_7778)
);

NAND2xp5_ASAP7_75t_L g7779 ( 
.A(n_7669),
.B(n_7688),
.Y(n_7779)
);

NOR3xp33_ASAP7_75t_L g7780 ( 
.A(n_7668),
.B(n_7647),
.C(n_5521),
.Y(n_7780)
);

NOR3x1_ASAP7_75t_L g7781 ( 
.A(n_7675),
.B(n_5469),
.C(n_4792),
.Y(n_7781)
);

NOR2xp67_ASAP7_75t_L g7782 ( 
.A(n_7676),
.B(n_5493),
.Y(n_7782)
);

NAND2xp33_ASAP7_75t_L g7783 ( 
.A(n_7679),
.B(n_5494),
.Y(n_7783)
);

NAND2xp5_ASAP7_75t_L g7784 ( 
.A(n_7688),
.B(n_5494),
.Y(n_7784)
);

AOI21xp5_ASAP7_75t_L g7785 ( 
.A1(n_7684),
.A2(n_5504),
.B(n_5501),
.Y(n_7785)
);

AOI211xp5_ASAP7_75t_L g7786 ( 
.A1(n_7679),
.A2(n_5469),
.B(n_5052),
.C(n_5501),
.Y(n_7786)
);

NAND4xp25_ASAP7_75t_L g7787 ( 
.A(n_7687),
.B(n_5161),
.C(n_4466),
.D(n_5127),
.Y(n_7787)
);

NOR2x1_ASAP7_75t_SL g7788 ( 
.A(n_7666),
.B(n_5504),
.Y(n_7788)
);

AOI22xp5_ASAP7_75t_L g7789 ( 
.A1(n_7743),
.A2(n_7691),
.B1(n_7754),
.B2(n_7663),
.Y(n_7789)
);

NOR2xp33_ASAP7_75t_L g7790 ( 
.A(n_7691),
.B(n_5539),
.Y(n_7790)
);

NAND3xp33_ASAP7_75t_SL g7791 ( 
.A(n_7665),
.B(n_5514),
.C(n_5352),
.Y(n_7791)
);

INVx1_ASAP7_75t_L g7792 ( 
.A(n_7667),
.Y(n_7792)
);

NOR2xp33_ASAP7_75t_L g7793 ( 
.A(n_7695),
.B(n_5539),
.Y(n_7793)
);

NOR3xp33_ASAP7_75t_L g7794 ( 
.A(n_7711),
.B(n_5370),
.C(n_5330),
.Y(n_7794)
);

AOI22xp5_ASAP7_75t_L g7795 ( 
.A1(n_7760),
.A2(n_5542),
.B1(n_5539),
.B2(n_5383),
.Y(n_7795)
);

INVx2_ASAP7_75t_L g7796 ( 
.A(n_7686),
.Y(n_7796)
);

BUFx3_ASAP7_75t_L g7797 ( 
.A(n_7713),
.Y(n_7797)
);

NAND2xp5_ASAP7_75t_L g7798 ( 
.A(n_7667),
.B(n_5508),
.Y(n_7798)
);

NAND4xp25_ASAP7_75t_SL g7799 ( 
.A(n_7762),
.B(n_5508),
.C(n_5515),
.D(n_5510),
.Y(n_7799)
);

INVxp33_ASAP7_75t_L g7800 ( 
.A(n_7702),
.Y(n_7800)
);

OAI21xp5_ASAP7_75t_SL g7801 ( 
.A1(n_7697),
.A2(n_5127),
.B(n_5002),
.Y(n_7801)
);

AOI221xp5_ASAP7_75t_L g7802 ( 
.A1(n_7736),
.A2(n_5384),
.B1(n_5383),
.B2(n_5330),
.C(n_5510),
.Y(n_7802)
);

AOI322xp5_ASAP7_75t_L g7803 ( 
.A1(n_7759),
.A2(n_5383),
.A3(n_5384),
.B1(n_5330),
.B2(n_5393),
.C1(n_5518),
.C2(n_5515),
.Y(n_7803)
);

INVxp33_ASAP7_75t_L g7804 ( 
.A(n_7692),
.Y(n_7804)
);

OAI21xp5_ASAP7_75t_L g7805 ( 
.A1(n_7718),
.A2(n_7696),
.B(n_7661),
.Y(n_7805)
);

NAND2xp5_ASAP7_75t_SL g7806 ( 
.A(n_7680),
.B(n_5518),
.Y(n_7806)
);

INVxp67_ASAP7_75t_L g7807 ( 
.A(n_7689),
.Y(n_7807)
);

AO22x2_ASAP7_75t_L g7808 ( 
.A1(n_7769),
.A2(n_7662),
.B1(n_7768),
.B2(n_7678),
.Y(n_7808)
);

NAND2xp5_ASAP7_75t_SL g7809 ( 
.A(n_7680),
.B(n_5519),
.Y(n_7809)
);

INVx1_ASAP7_75t_L g7810 ( 
.A(n_7706),
.Y(n_7810)
);

OAI21xp5_ASAP7_75t_SL g7811 ( 
.A1(n_7697),
.A2(n_5127),
.B(n_5002),
.Y(n_7811)
);

INVxp67_ASAP7_75t_SL g7812 ( 
.A(n_7683),
.Y(n_7812)
);

OAI211xp5_ASAP7_75t_L g7813 ( 
.A1(n_7715),
.A2(n_5025),
.B(n_5449),
.C(n_5416),
.Y(n_7813)
);

NAND2xp5_ASAP7_75t_L g7814 ( 
.A(n_7685),
.B(n_5519),
.Y(n_7814)
);

NAND4xp25_ASAP7_75t_L g7815 ( 
.A(n_7761),
.B(n_5161),
.C(n_4466),
.D(n_5002),
.Y(n_7815)
);

AND2x2_ASAP7_75t_L g7816 ( 
.A(n_7698),
.B(n_5072),
.Y(n_7816)
);

NAND3xp33_ASAP7_75t_SL g7817 ( 
.A(n_7681),
.B(n_5384),
.C(n_5185),
.Y(n_7817)
);

OAI31xp33_ASAP7_75t_L g7818 ( 
.A1(n_7724),
.A2(n_7763),
.A3(n_7765),
.B(n_7749),
.Y(n_7818)
);

NAND4xp25_ASAP7_75t_L g7819 ( 
.A(n_7677),
.B(n_5047),
.C(n_5046),
.D(n_4547),
.Y(n_7819)
);

AOI21xp33_ASAP7_75t_SL g7820 ( 
.A1(n_7728),
.A2(n_5449),
.B(n_5416),
.Y(n_7820)
);

NAND2xp5_ASAP7_75t_SL g7821 ( 
.A(n_7734),
.B(n_5524),
.Y(n_7821)
);

NAND2xp5_ASAP7_75t_L g7822 ( 
.A(n_7746),
.B(n_5524),
.Y(n_7822)
);

NAND2xp5_ASAP7_75t_L g7823 ( 
.A(n_7747),
.B(n_5528),
.Y(n_7823)
);

NAND2xp5_ASAP7_75t_L g7824 ( 
.A(n_7704),
.B(n_5528),
.Y(n_7824)
);

XNOR2x2_ASAP7_75t_L g7825 ( 
.A(n_7745),
.B(n_7670),
.Y(n_7825)
);

NAND5xp2_ASAP7_75t_L g7826 ( 
.A(n_7717),
.B(n_5120),
.C(n_4728),
.D(n_4598),
.E(n_4585),
.Y(n_7826)
);

NOR4xp25_ASAP7_75t_SL g7827 ( 
.A(n_7705),
.B(n_5550),
.C(n_5554),
.D(n_5549),
.Y(n_7827)
);

AOI22xp5_ASAP7_75t_L g7828 ( 
.A1(n_7682),
.A2(n_5542),
.B1(n_5539),
.B2(n_5416),
.Y(n_7828)
);

O2A1O1Ixp33_ASAP7_75t_L g7829 ( 
.A1(n_7753),
.A2(n_5550),
.B(n_5554),
.C(n_5549),
.Y(n_7829)
);

NAND4xp75_ASAP7_75t_L g7830 ( 
.A(n_7721),
.B(n_5416),
.C(n_5449),
.D(n_5106),
.Y(n_7830)
);

OAI221xp5_ASAP7_75t_L g7831 ( 
.A1(n_7755),
.A2(n_5449),
.B1(n_5558),
.B2(n_5569),
.C(n_5562),
.Y(n_7831)
);

AND4x1_ASAP7_75t_L g7832 ( 
.A(n_7744),
.B(n_5073),
.C(n_4547),
.D(n_4947),
.Y(n_7832)
);

NOR2xp33_ASAP7_75t_L g7833 ( 
.A(n_7735),
.B(n_5542),
.Y(n_7833)
);

NOR2xp33_ASAP7_75t_L g7834 ( 
.A(n_7739),
.B(n_5542),
.Y(n_7834)
);

AOI22xp5_ASAP7_75t_L g7835 ( 
.A1(n_7757),
.A2(n_5562),
.B1(n_5569),
.B2(n_5558),
.Y(n_7835)
);

HB1xp67_ASAP7_75t_L g7836 ( 
.A(n_7700),
.Y(n_7836)
);

INVx1_ASAP7_75t_L g7837 ( 
.A(n_7726),
.Y(n_7837)
);

HB1xp67_ASAP7_75t_L g7838 ( 
.A(n_7734),
.Y(n_7838)
);

INVx1_ASAP7_75t_L g7839 ( 
.A(n_7694),
.Y(n_7839)
);

INVx1_ASAP7_75t_L g7840 ( 
.A(n_7750),
.Y(n_7840)
);

O2A1O1Ixp33_ASAP7_75t_L g7841 ( 
.A1(n_7693),
.A2(n_5571),
.B(n_5580),
.C(n_5570),
.Y(n_7841)
);

INVx1_ASAP7_75t_SL g7842 ( 
.A(n_7766),
.Y(n_7842)
);

NAND2xp5_ASAP7_75t_SL g7843 ( 
.A(n_7701),
.B(n_5570),
.Y(n_7843)
);

NOR3xp33_ASAP7_75t_L g7844 ( 
.A(n_7752),
.B(n_5580),
.C(n_5571),
.Y(n_7844)
);

OR2x2_ASAP7_75t_L g7845 ( 
.A(n_7690),
.B(n_7758),
.Y(n_7845)
);

XNOR2x1_ASAP7_75t_L g7846 ( 
.A(n_7751),
.B(n_7756),
.Y(n_7846)
);

AOI22xp5_ASAP7_75t_L g7847 ( 
.A1(n_7751),
.A2(n_5532),
.B1(n_5534),
.B2(n_5509),
.Y(n_7847)
);

BUFx2_ASAP7_75t_L g7848 ( 
.A(n_7758),
.Y(n_7848)
);

AOI211x1_ASAP7_75t_SL g7849 ( 
.A1(n_7699),
.A2(n_4943),
.B(n_5091),
.C(n_5084),
.Y(n_7849)
);

NOR2x1_ASAP7_75t_L g7850 ( 
.A(n_7748),
.B(n_7729),
.Y(n_7850)
);

NOR2xp33_ASAP7_75t_L g7851 ( 
.A(n_7719),
.B(n_5073),
.Y(n_7851)
);

NAND4xp25_ASAP7_75t_L g7852 ( 
.A(n_7714),
.B(n_5065),
.C(n_4588),
.D(n_4402),
.Y(n_7852)
);

AOI211xp5_ASAP7_75t_L g7853 ( 
.A1(n_7737),
.A2(n_5091),
.B(n_5129),
.C(n_5084),
.Y(n_7853)
);

NAND2xp5_ASAP7_75t_L g7854 ( 
.A(n_7714),
.B(n_5509),
.Y(n_7854)
);

NOR3x1_ASAP7_75t_L g7855 ( 
.A(n_7731),
.B(n_5109),
.C(n_5006),
.Y(n_7855)
);

INVx2_ASAP7_75t_L g7856 ( 
.A(n_7727),
.Y(n_7856)
);

INVx1_ASAP7_75t_L g7857 ( 
.A(n_7750),
.Y(n_7857)
);

NAND4xp25_ASAP7_75t_L g7858 ( 
.A(n_7725),
.B(n_7709),
.C(n_7703),
.D(n_7742),
.Y(n_7858)
);

NAND4xp25_ASAP7_75t_L g7859 ( 
.A(n_7712),
.B(n_4588),
.C(n_4573),
.D(n_4678),
.Y(n_7859)
);

NOR2xp33_ASAP7_75t_L g7860 ( 
.A(n_7720),
.B(n_5551),
.Y(n_7860)
);

INVx2_ASAP7_75t_L g7861 ( 
.A(n_7722),
.Y(n_7861)
);

NAND2xp5_ASAP7_75t_L g7862 ( 
.A(n_7808),
.B(n_7740),
.Y(n_7862)
);

NAND2xp5_ASAP7_75t_L g7863 ( 
.A(n_7808),
.B(n_7740),
.Y(n_7863)
);

NAND3xp33_ASAP7_75t_L g7864 ( 
.A(n_7789),
.B(n_7733),
.C(n_7699),
.Y(n_7864)
);

NOR2x1p5_ASAP7_75t_SL g7865 ( 
.A(n_7776),
.B(n_7764),
.Y(n_7865)
);

INVx1_ASAP7_75t_L g7866 ( 
.A(n_7825),
.Y(n_7866)
);

NAND4xp25_ASAP7_75t_L g7867 ( 
.A(n_7842),
.B(n_7767),
.C(n_7770),
.D(n_7730),
.Y(n_7867)
);

NOR3xp33_ASAP7_75t_L g7868 ( 
.A(n_7779),
.B(n_7707),
.C(n_7710),
.Y(n_7868)
);

INVx1_ASAP7_75t_L g7869 ( 
.A(n_7792),
.Y(n_7869)
);

A2O1A1Ixp33_ASAP7_75t_L g7870 ( 
.A1(n_7790),
.A2(n_7732),
.B(n_7723),
.C(n_7716),
.Y(n_7870)
);

NAND2x1_ASAP7_75t_L g7871 ( 
.A(n_7848),
.B(n_7672),
.Y(n_7871)
);

NAND2xp5_ASAP7_75t_L g7872 ( 
.A(n_7842),
.B(n_7741),
.Y(n_7872)
);

INVx1_ASAP7_75t_L g7873 ( 
.A(n_7797),
.Y(n_7873)
);

NAND2xp67_ASAP7_75t_SL g7874 ( 
.A(n_7816),
.B(n_7741),
.Y(n_7874)
);

NAND2xp5_ASAP7_75t_L g7875 ( 
.A(n_7838),
.B(n_7836),
.Y(n_7875)
);

NOR2xp33_ASAP7_75t_L g7876 ( 
.A(n_7804),
.B(n_5551),
.Y(n_7876)
);

NAND2x1p5_ASAP7_75t_L g7877 ( 
.A(n_7839),
.B(n_5006),
.Y(n_7877)
);

NAND2xp5_ASAP7_75t_L g7878 ( 
.A(n_7788),
.B(n_5393),
.Y(n_7878)
);

NOR2x1_ASAP7_75t_L g7879 ( 
.A(n_7858),
.B(n_5458),
.Y(n_7879)
);

HB1xp67_ASAP7_75t_L g7880 ( 
.A(n_7782),
.Y(n_7880)
);

AOI22xp5_ASAP7_75t_L g7881 ( 
.A1(n_7812),
.A2(n_5509),
.B1(n_5534),
.B2(n_5532),
.Y(n_7881)
);

NAND2xp5_ASAP7_75t_L g7882 ( 
.A(n_7810),
.B(n_5393),
.Y(n_7882)
);

NOR2xp33_ASAP7_75t_L g7883 ( 
.A(n_7773),
.B(n_5551),
.Y(n_7883)
);

AND2x2_ASAP7_75t_L g7884 ( 
.A(n_7796),
.B(n_7855),
.Y(n_7884)
);

AND2x2_ASAP7_75t_L g7885 ( 
.A(n_7837),
.B(n_5393),
.Y(n_7885)
);

NOR3xp33_ASAP7_75t_L g7886 ( 
.A(n_7805),
.B(n_5130),
.C(n_4638),
.Y(n_7886)
);

OAI211xp5_ASAP7_75t_SL g7887 ( 
.A1(n_7818),
.A2(n_4678),
.B(n_5149),
.C(n_5109),
.Y(n_7887)
);

NAND2xp5_ASAP7_75t_L g7888 ( 
.A(n_7771),
.B(n_5393),
.Y(n_7888)
);

AOI322xp5_ASAP7_75t_L g7889 ( 
.A1(n_7793),
.A2(n_5393),
.A3(n_4853),
.B1(n_4891),
.B2(n_4856),
.C1(n_4894),
.C2(n_4865),
.Y(n_7889)
);

OAI21x1_ASAP7_75t_L g7890 ( 
.A1(n_7775),
.A2(n_5458),
.B(n_5551),
.Y(n_7890)
);

NAND4xp25_ASAP7_75t_L g7891 ( 
.A(n_7772),
.B(n_4573),
.C(n_4546),
.D(n_4638),
.Y(n_7891)
);

NAND4xp25_ASAP7_75t_L g7892 ( 
.A(n_7777),
.B(n_4412),
.C(n_4642),
.D(n_4628),
.Y(n_7892)
);

AND4x1_ASAP7_75t_L g7893 ( 
.A(n_7805),
.B(n_4973),
.C(n_4978),
.D(n_4968),
.Y(n_7893)
);

INVx1_ASAP7_75t_L g7894 ( 
.A(n_7850),
.Y(n_7894)
);

AOI211xp5_ASAP7_75t_L g7895 ( 
.A1(n_7774),
.A2(n_5091),
.B(n_5129),
.C(n_5084),
.Y(n_7895)
);

OAI21xp33_ASAP7_75t_L g7896 ( 
.A1(n_7800),
.A2(n_5186),
.B(n_5149),
.Y(n_7896)
);

NOR2xp67_ASAP7_75t_L g7897 ( 
.A(n_7807),
.B(n_5186),
.Y(n_7897)
);

NAND3xp33_ASAP7_75t_SL g7898 ( 
.A(n_7845),
.B(n_5132),
.C(n_5090),
.Y(n_7898)
);

NAND2xp5_ASAP7_75t_L g7899 ( 
.A(n_7833),
.B(n_5458),
.Y(n_7899)
);

AOI21xp5_ASAP7_75t_L g7900 ( 
.A1(n_7783),
.A2(n_5458),
.B(n_5509),
.Y(n_7900)
);

INVx2_ASAP7_75t_SL g7901 ( 
.A(n_7861),
.Y(n_7901)
);

NOR4xp25_ASAP7_75t_L g7902 ( 
.A(n_7840),
.B(n_5177),
.C(n_5179),
.D(n_5176),
.Y(n_7902)
);

AOI21xp5_ASAP7_75t_L g7903 ( 
.A1(n_7798),
.A2(n_5534),
.B(n_5532),
.Y(n_7903)
);

INVx1_ASAP7_75t_L g7904 ( 
.A(n_7846),
.Y(n_7904)
);

NAND2xp5_ASAP7_75t_SL g7905 ( 
.A(n_7856),
.B(n_5084),
.Y(n_7905)
);

INVx1_ASAP7_75t_L g7906 ( 
.A(n_7857),
.Y(n_7906)
);

NOR2xp33_ASAP7_75t_L g7907 ( 
.A(n_7834),
.B(n_5563),
.Y(n_7907)
);

NAND2xp5_ASAP7_75t_SL g7908 ( 
.A(n_7853),
.B(n_5084),
.Y(n_7908)
);

NOR3xp33_ASAP7_75t_L g7909 ( 
.A(n_7780),
.B(n_4853),
.C(n_4845),
.Y(n_7909)
);

INVxp33_ASAP7_75t_L g7910 ( 
.A(n_7823),
.Y(n_7910)
);

NOR3xp33_ASAP7_75t_L g7911 ( 
.A(n_7791),
.B(n_4853),
.C(n_4845),
.Y(n_7911)
);

NAND4xp25_ASAP7_75t_L g7912 ( 
.A(n_7851),
.B(n_4973),
.C(n_4978),
.D(n_4968),
.Y(n_7912)
);

NAND2xp5_ASAP7_75t_L g7913 ( 
.A(n_7785),
.B(n_5532),
.Y(n_7913)
);

NOR2xp33_ASAP7_75t_L g7914 ( 
.A(n_7814),
.B(n_5563),
.Y(n_7914)
);

NOR4xp75_ASAP7_75t_SL g7915 ( 
.A(n_7824),
.B(n_5095),
.C(n_4996),
.D(n_4578),
.Y(n_7915)
);

AOI221x1_ASAP7_75t_L g7916 ( 
.A1(n_7844),
.A2(n_5129),
.B1(n_5165),
.B2(n_5091),
.C(n_5176),
.Y(n_7916)
);

AOI211xp5_ASAP7_75t_L g7917 ( 
.A1(n_7831),
.A2(n_5129),
.B(n_5165),
.C(n_5091),
.Y(n_7917)
);

AOI21xp5_ASAP7_75t_L g7918 ( 
.A1(n_7843),
.A2(n_5552),
.B(n_5534),
.Y(n_7918)
);

INVx2_ASAP7_75t_L g7919 ( 
.A(n_7784),
.Y(n_7919)
);

AND2x2_ASAP7_75t_L g7920 ( 
.A(n_7778),
.B(n_5072),
.Y(n_7920)
);

INVx3_ASAP7_75t_L g7921 ( 
.A(n_7822),
.Y(n_7921)
);

AOI22xp5_ASAP7_75t_L g7922 ( 
.A1(n_7860),
.A2(n_5585),
.B1(n_5552),
.B2(n_5563),
.Y(n_7922)
);

NAND4xp75_ASAP7_75t_L g7923 ( 
.A(n_7781),
.B(n_5106),
.C(n_5595),
.D(n_5563),
.Y(n_7923)
);

OAI21xp33_ASAP7_75t_L g7924 ( 
.A1(n_7801),
.A2(n_4996),
.B(n_5036),
.Y(n_7924)
);

NAND3xp33_ASAP7_75t_L g7925 ( 
.A(n_7794),
.B(n_5595),
.C(n_5165),
.Y(n_7925)
);

OR2x2_ASAP7_75t_L g7926 ( 
.A(n_7852),
.B(n_5552),
.Y(n_7926)
);

INVx1_ASAP7_75t_L g7927 ( 
.A(n_7854),
.Y(n_7927)
);

AOI22xp5_ASAP7_75t_L g7928 ( 
.A1(n_7854),
.A2(n_5585),
.B1(n_5552),
.B2(n_5595),
.Y(n_7928)
);

NAND2xp5_ASAP7_75t_SL g7929 ( 
.A(n_7829),
.B(n_5129),
.Y(n_7929)
);

NAND2xp5_ASAP7_75t_L g7930 ( 
.A(n_7827),
.B(n_5585),
.Y(n_7930)
);

NAND2xp5_ASAP7_75t_L g7931 ( 
.A(n_7806),
.B(n_5585),
.Y(n_7931)
);

INVx1_ASAP7_75t_L g7932 ( 
.A(n_7809),
.Y(n_7932)
);

NAND2xp5_ASAP7_75t_SL g7933 ( 
.A(n_7847),
.B(n_5165),
.Y(n_7933)
);

NAND3xp33_ASAP7_75t_L g7934 ( 
.A(n_7803),
.B(n_5595),
.C(n_5165),
.Y(n_7934)
);

NAND3xp33_ASAP7_75t_L g7935 ( 
.A(n_7821),
.B(n_4856),
.C(n_4845),
.Y(n_7935)
);

NOR2xp33_ASAP7_75t_L g7936 ( 
.A(n_7817),
.B(n_4856),
.Y(n_7936)
);

INVxp33_ASAP7_75t_SL g7937 ( 
.A(n_7835),
.Y(n_7937)
);

INVx1_ASAP7_75t_L g7938 ( 
.A(n_7841),
.Y(n_7938)
);

OAI211xp5_ASAP7_75t_SL g7939 ( 
.A1(n_7849),
.A2(n_4522),
.B(n_5179),
.C(n_5177),
.Y(n_7939)
);

NAND4xp25_ASAP7_75t_L g7940 ( 
.A(n_7786),
.B(n_7787),
.C(n_7815),
.D(n_7811),
.Y(n_7940)
);

AOI221xp5_ASAP7_75t_L g7941 ( 
.A1(n_7862),
.A2(n_7799),
.B1(n_7820),
.B2(n_7802),
.C(n_7795),
.Y(n_7941)
);

NOR3xp33_ASAP7_75t_L g7942 ( 
.A(n_7866),
.B(n_7813),
.C(n_7859),
.Y(n_7942)
);

NAND3xp33_ASAP7_75t_L g7943 ( 
.A(n_7863),
.B(n_7828),
.C(n_7832),
.Y(n_7943)
);

OAI221xp5_ASAP7_75t_L g7944 ( 
.A1(n_7875),
.A2(n_7819),
.B1(n_7826),
.B2(n_7830),
.C(n_5120),
.Y(n_7944)
);

NAND3xp33_ASAP7_75t_SL g7945 ( 
.A(n_7904),
.B(n_7872),
.C(n_7894),
.Y(n_7945)
);

NAND4xp25_ASAP7_75t_L g7946 ( 
.A(n_7864),
.B(n_7826),
.C(n_4412),
.D(n_4368),
.Y(n_7946)
);

OR2x2_ASAP7_75t_L g7947 ( 
.A(n_7877),
.B(n_4865),
.Y(n_7947)
);

NOR3xp33_ASAP7_75t_L g7948 ( 
.A(n_7873),
.B(n_4891),
.C(n_4865),
.Y(n_7948)
);

NOR3xp33_ASAP7_75t_L g7949 ( 
.A(n_7901),
.B(n_4894),
.C(n_4891),
.Y(n_7949)
);

INVx1_ASAP7_75t_L g7950 ( 
.A(n_7877),
.Y(n_7950)
);

NAND2xp5_ASAP7_75t_L g7951 ( 
.A(n_7880),
.B(n_4894),
.Y(n_7951)
);

NOR2xp33_ASAP7_75t_L g7952 ( 
.A(n_7878),
.B(n_4935),
.Y(n_7952)
);

NOR3xp33_ASAP7_75t_L g7953 ( 
.A(n_7869),
.B(n_7906),
.C(n_7921),
.Y(n_7953)
);

AOI21xp5_ASAP7_75t_L g7954 ( 
.A1(n_7905),
.A2(n_5183),
.B(n_5181),
.Y(n_7954)
);

NOR4xp25_ASAP7_75t_L g7955 ( 
.A(n_7867),
.B(n_5183),
.C(n_5191),
.D(n_5181),
.Y(n_7955)
);

NAND3xp33_ASAP7_75t_L g7956 ( 
.A(n_7868),
.B(n_4936),
.C(n_4935),
.Y(n_7956)
);

AOI32xp33_ASAP7_75t_L g7957 ( 
.A1(n_7884),
.A2(n_4910),
.A3(n_4927),
.B1(n_4918),
.B2(n_4895),
.Y(n_7957)
);

AOI211xp5_ASAP7_75t_L g7958 ( 
.A1(n_7910),
.A2(n_4910),
.B(n_4918),
.C(n_4895),
.Y(n_7958)
);

NAND4xp25_ASAP7_75t_L g7959 ( 
.A(n_7897),
.B(n_4615),
.C(n_4945),
.D(n_4927),
.Y(n_7959)
);

AOI221x1_ASAP7_75t_L g7960 ( 
.A1(n_7932),
.A2(n_5191),
.B1(n_5158),
.B2(n_5104),
.C(n_5034),
.Y(n_7960)
);

NAND5xp2_ASAP7_75t_L g7961 ( 
.A(n_7895),
.B(n_7883),
.C(n_7920),
.D(n_7888),
.E(n_7876),
.Y(n_7961)
);

NAND4xp25_ASAP7_75t_L g7962 ( 
.A(n_7882),
.B(n_4615),
.C(n_4948),
.D(n_4945),
.Y(n_7962)
);

NOR3xp33_ASAP7_75t_L g7963 ( 
.A(n_7921),
.B(n_4936),
.C(n_4935),
.Y(n_7963)
);

NAND3xp33_ASAP7_75t_L g7964 ( 
.A(n_7871),
.B(n_4942),
.C(n_4936),
.Y(n_7964)
);

NOR2x1p5_ASAP7_75t_L g7965 ( 
.A(n_7898),
.B(n_4979),
.Y(n_7965)
);

NOR3xp33_ASAP7_75t_L g7966 ( 
.A(n_7919),
.B(n_7927),
.C(n_7938),
.Y(n_7966)
);

NOR2xp33_ASAP7_75t_L g7967 ( 
.A(n_7923),
.B(n_4942),
.Y(n_7967)
);

OAI21xp5_ASAP7_75t_L g7968 ( 
.A1(n_7870),
.A2(n_4970),
.B(n_4942),
.Y(n_7968)
);

NOR3xp33_ASAP7_75t_L g7969 ( 
.A(n_7879),
.B(n_4983),
.C(n_4970),
.Y(n_7969)
);

AOI21xp5_ASAP7_75t_L g7970 ( 
.A1(n_7937),
.A2(n_4417),
.B(n_4970),
.Y(n_7970)
);

NOR2x1_ASAP7_75t_L g7971 ( 
.A(n_7874),
.B(n_4948),
.Y(n_7971)
);

NOR2xp33_ASAP7_75t_SL g7972 ( 
.A(n_7940),
.B(n_4996),
.Y(n_7972)
);

NAND4xp25_ASAP7_75t_L g7973 ( 
.A(n_7940),
.B(n_4180),
.C(n_4420),
.D(n_4694),
.Y(n_7973)
);

AOI211x1_ASAP7_75t_L g7974 ( 
.A1(n_7896),
.A2(n_4858),
.B(n_4800),
.C(n_4801),
.Y(n_7974)
);

AOI221x1_ASAP7_75t_L g7975 ( 
.A1(n_7887),
.A2(n_5158),
.B1(n_5104),
.B2(n_5034),
.C(n_5048),
.Y(n_7975)
);

O2A1O1Ixp33_ASAP7_75t_SL g7976 ( 
.A1(n_7929),
.A2(n_4565),
.B(n_4400),
.C(n_4499),
.Y(n_7976)
);

NAND4xp75_ASAP7_75t_L g7977 ( 
.A(n_7865),
.B(n_5106),
.C(n_4417),
.D(n_4858),
.Y(n_7977)
);

NAND3xp33_ASAP7_75t_L g7978 ( 
.A(n_7917),
.B(n_4984),
.C(n_4983),
.Y(n_7978)
);

AOI211xp5_ASAP7_75t_L g7979 ( 
.A1(n_7934),
.A2(n_5103),
.B(n_5138),
.C(n_5028),
.Y(n_7979)
);

NOR3xp33_ASAP7_75t_SL g7980 ( 
.A(n_7908),
.B(n_7930),
.C(n_7933),
.Y(n_7980)
);

NAND3xp33_ASAP7_75t_L g7981 ( 
.A(n_7936),
.B(n_4984),
.C(n_4983),
.Y(n_7981)
);

NAND4xp75_ASAP7_75t_L g7982 ( 
.A(n_7885),
.B(n_4417),
.C(n_4702),
.D(n_4697),
.Y(n_7982)
);

NAND3xp33_ASAP7_75t_L g7983 ( 
.A(n_7926),
.B(n_4991),
.C(n_4984),
.Y(n_7983)
);

AOI221x1_ASAP7_75t_SL g7984 ( 
.A1(n_7913),
.A2(n_4994),
.B1(n_5007),
.B2(n_4998),
.C(n_4991),
.Y(n_7984)
);

NAND2xp5_ASAP7_75t_L g7985 ( 
.A(n_7914),
.B(n_4991),
.Y(n_7985)
);

INVx1_ASAP7_75t_SL g7986 ( 
.A(n_7931),
.Y(n_7986)
);

AND3x1_ASAP7_75t_L g7987 ( 
.A(n_7924),
.B(n_4887),
.C(n_4878),
.Y(n_7987)
);

NOR3xp33_ASAP7_75t_L g7988 ( 
.A(n_7899),
.B(n_4998),
.C(n_4994),
.Y(n_7988)
);

O2A1O1Ixp33_ASAP7_75t_L g7989 ( 
.A1(n_7907),
.A2(n_5120),
.B(n_4728),
.C(n_5096),
.Y(n_7989)
);

NOR2xp33_ASAP7_75t_L g7990 ( 
.A(n_7925),
.B(n_4994),
.Y(n_7990)
);

OAI22xp5_ASAP7_75t_L g7991 ( 
.A1(n_7935),
.A2(n_4998),
.B1(n_5015),
.B2(n_5007),
.Y(n_7991)
);

OAI211xp5_ASAP7_75t_SL g7992 ( 
.A1(n_7918),
.A2(n_4468),
.B(n_4454),
.C(n_4481),
.Y(n_7992)
);

NAND2xp5_ASAP7_75t_L g7993 ( 
.A(n_7886),
.B(n_5007),
.Y(n_7993)
);

NOR2xp67_ASAP7_75t_L g7994 ( 
.A(n_7912),
.B(n_5104),
.Y(n_7994)
);

NAND2xp5_ASAP7_75t_L g7995 ( 
.A(n_7916),
.B(n_5015),
.Y(n_7995)
);

AOI21xp33_ASAP7_75t_L g7996 ( 
.A1(n_7928),
.A2(n_5059),
.B(n_5015),
.Y(n_7996)
);

INVx1_ASAP7_75t_L g7997 ( 
.A(n_7890),
.Y(n_7997)
);

NAND3xp33_ASAP7_75t_L g7998 ( 
.A(n_7903),
.B(n_5068),
.C(n_5059),
.Y(n_7998)
);

NOR4xp75_ASAP7_75t_L g7999 ( 
.A(n_7915),
.B(n_4468),
.C(n_4887),
.D(n_4878),
.Y(n_7999)
);

NOR3xp33_ASAP7_75t_L g8000 ( 
.A(n_7939),
.B(n_5068),
.C(n_5059),
.Y(n_8000)
);

NAND2xp5_ASAP7_75t_L g8001 ( 
.A(n_7902),
.B(n_5068),
.Y(n_8001)
);

NOR3xp33_ASAP7_75t_L g8002 ( 
.A(n_7892),
.B(n_5094),
.C(n_5076),
.Y(n_8002)
);

NOR2xp33_ASAP7_75t_L g8003 ( 
.A(n_7893),
.B(n_5076),
.Y(n_8003)
);

AOI21xp5_ASAP7_75t_L g8004 ( 
.A1(n_7900),
.A2(n_5094),
.B(n_5076),
.Y(n_8004)
);

NAND4xp25_ASAP7_75t_L g8005 ( 
.A(n_7889),
.B(n_4180),
.C(n_4420),
.D(n_4694),
.Y(n_8005)
);

NAND2xp5_ASAP7_75t_L g8006 ( 
.A(n_7911),
.B(n_5094),
.Y(n_8006)
);

NAND3xp33_ASAP7_75t_L g8007 ( 
.A(n_7909),
.B(n_5147),
.C(n_5118),
.Y(n_8007)
);

NAND4xp75_ASAP7_75t_L g8008 ( 
.A(n_7922),
.B(n_4702),
.C(n_4703),
.D(n_4697),
.Y(n_8008)
);

NAND2xp5_ASAP7_75t_L g8009 ( 
.A(n_7881),
.B(n_5118),
.Y(n_8009)
);

NAND4xp25_ASAP7_75t_L g8010 ( 
.A(n_7912),
.B(n_4180),
.C(n_4694),
.D(n_4452),
.Y(n_8010)
);

AOI21xp5_ASAP7_75t_L g8011 ( 
.A1(n_7891),
.A2(n_5147),
.B(n_5118),
.Y(n_8011)
);

NAND2xp5_ASAP7_75t_L g8012 ( 
.A(n_7866),
.B(n_5147),
.Y(n_8012)
);

AOI21xp5_ASAP7_75t_L g8013 ( 
.A1(n_7866),
.A2(n_5172),
.B(n_5152),
.Y(n_8013)
);

NOR4xp25_ASAP7_75t_SL g8014 ( 
.A(n_7866),
.B(n_5018),
.C(n_4868),
.D(n_4698),
.Y(n_8014)
);

NAND4xp75_ASAP7_75t_L g8015 ( 
.A(n_7865),
.B(n_4703),
.C(n_4274),
.D(n_4416),
.Y(n_8015)
);

NAND2x1p5_ASAP7_75t_L g8016 ( 
.A(n_7894),
.B(n_4399),
.Y(n_8016)
);

NAND3xp33_ASAP7_75t_L g8017 ( 
.A(n_7866),
.B(n_5172),
.C(n_5152),
.Y(n_8017)
);

NAND4xp25_ASAP7_75t_L g8018 ( 
.A(n_7866),
.B(n_4180),
.C(n_5034),
.D(n_4979),
.Y(n_8018)
);

INVx1_ASAP7_75t_L g8019 ( 
.A(n_7971),
.Y(n_8019)
);

NAND2xp5_ASAP7_75t_L g8020 ( 
.A(n_7950),
.B(n_8014),
.Y(n_8020)
);

AOI211xp5_ASAP7_75t_L g8021 ( 
.A1(n_7961),
.A2(n_4633),
.B(n_5034),
.C(n_4979),
.Y(n_8021)
);

NAND4xp25_ASAP7_75t_L g8022 ( 
.A(n_7953),
.B(n_7972),
.C(n_7945),
.D(n_7942),
.Y(n_8022)
);

INVx2_ASAP7_75t_L g8023 ( 
.A(n_8016),
.Y(n_8023)
);

NAND2xp5_ASAP7_75t_L g8024 ( 
.A(n_7966),
.B(n_5152),
.Y(n_8024)
);

NOR3xp33_ASAP7_75t_SL g8025 ( 
.A(n_7943),
.B(n_5018),
.C(n_4470),
.Y(n_8025)
);

NOR3x1_ASAP7_75t_L g8026 ( 
.A(n_8012),
.B(n_4454),
.C(n_4481),
.Y(n_8026)
);

AOI221xp5_ASAP7_75t_L g8027 ( 
.A1(n_7944),
.A2(n_5172),
.B1(n_4904),
.B2(n_4907),
.C(n_4899),
.Y(n_8027)
);

INVx1_ASAP7_75t_L g8028 ( 
.A(n_7947),
.Y(n_8028)
);

AOI221x1_ASAP7_75t_L g8029 ( 
.A1(n_7997),
.A2(n_5104),
.B1(n_5158),
.B2(n_5048),
.C(n_4979),
.Y(n_8029)
);

NOR3xp33_ASAP7_75t_L g8030 ( 
.A(n_7986),
.B(n_4899),
.C(n_4815),
.Y(n_8030)
);

NAND3xp33_ASAP7_75t_SL g8031 ( 
.A(n_7941),
.B(n_4904),
.C(n_4815),
.Y(n_8031)
);

OAI21xp5_ASAP7_75t_L g8032 ( 
.A1(n_7951),
.A2(n_5032),
.B(n_4907),
.Y(n_8032)
);

AOI211xp5_ASAP7_75t_L g8033 ( 
.A1(n_8017),
.A2(n_5048),
.B(n_4800),
.C(n_4801),
.Y(n_8033)
);

NOR2xp33_ASAP7_75t_L g8034 ( 
.A(n_8016),
.B(n_5032),
.Y(n_8034)
);

AOI221xp5_ASAP7_75t_L g8035 ( 
.A1(n_8013),
.A2(n_5033),
.B1(n_5110),
.B2(n_5101),
.C(n_5048),
.Y(n_8035)
);

INVx1_ASAP7_75t_L g8036 ( 
.A(n_8001),
.Y(n_8036)
);

OAI211xp5_ASAP7_75t_SL g8037 ( 
.A1(n_7980),
.A2(n_4482),
.B(n_4492),
.C(n_4526),
.Y(n_8037)
);

NAND4xp25_ASAP7_75t_SL g8038 ( 
.A(n_7975),
.B(n_4793),
.C(n_4813),
.D(n_4806),
.Y(n_8038)
);

NAND4xp25_ASAP7_75t_L g8039 ( 
.A(n_7984),
.B(n_4407),
.C(n_4648),
.D(n_4647),
.Y(n_8039)
);

OAI211xp5_ASAP7_75t_L g8040 ( 
.A1(n_7995),
.A2(n_4806),
.B(n_4813),
.C(n_4793),
.Y(n_8040)
);

INVx1_ASAP7_75t_L g8041 ( 
.A(n_8003),
.Y(n_8041)
);

NOR3xp33_ASAP7_75t_L g8042 ( 
.A(n_7952),
.B(n_5101),
.C(n_5033),
.Y(n_8042)
);

NOR3xp33_ASAP7_75t_SL g8043 ( 
.A(n_7977),
.B(n_5018),
.C(n_4470),
.Y(n_8043)
);

NAND3xp33_ASAP7_75t_L g8044 ( 
.A(n_7967),
.B(n_5110),
.C(n_4574),
.Y(n_8044)
);

OAI211xp5_ASAP7_75t_L g8045 ( 
.A1(n_8018),
.A2(n_4831),
.B(n_4846),
.C(n_4814),
.Y(n_8045)
);

NOR4xp25_ASAP7_75t_L g8046 ( 
.A(n_7993),
.B(n_5030),
.C(n_5038),
.D(n_4995),
.Y(n_8046)
);

OAI211xp5_ASAP7_75t_SL g8047 ( 
.A1(n_7985),
.A2(n_4482),
.B(n_4492),
.C(n_4526),
.Y(n_8047)
);

AOI21xp5_ASAP7_75t_L g8048 ( 
.A1(n_7990),
.A2(n_4416),
.B(n_4995),
.Y(n_8048)
);

AOI221xp5_ASAP7_75t_L g8049 ( 
.A1(n_7984),
.A2(n_5041),
.B1(n_5044),
.B2(n_5038),
.C(n_5030),
.Y(n_8049)
);

AND4x1_ASAP7_75t_L g8050 ( 
.A(n_7979),
.B(n_4831),
.C(n_4846),
.D(n_4814),
.Y(n_8050)
);

NAND2xp5_ASAP7_75t_SL g8051 ( 
.A(n_7994),
.B(n_4868),
.Y(n_8051)
);

NAND5xp2_ASAP7_75t_L g8052 ( 
.A(n_7949),
.B(n_4728),
.C(n_4630),
.D(n_4875),
.E(n_5096),
.Y(n_8052)
);

INVx1_ASAP7_75t_L g8053 ( 
.A(n_7999),
.Y(n_8053)
);

NAND4xp25_ASAP7_75t_L g8054 ( 
.A(n_7946),
.B(n_4407),
.C(n_4648),
.D(n_4647),
.Y(n_8054)
);

NAND2xp5_ASAP7_75t_L g8055 ( 
.A(n_7955),
.B(n_5190),
.Y(n_8055)
);

NOR4xp25_ASAP7_75t_L g8056 ( 
.A(n_7992),
.B(n_5044),
.C(n_5041),
.D(n_4875),
.Y(n_8056)
);

O2A1O1Ixp33_ASAP7_75t_L g8057 ( 
.A1(n_8009),
.A2(n_5137),
.B(n_5058),
.C(n_5004),
.Y(n_8057)
);

NAND4xp25_ASAP7_75t_L g8058 ( 
.A(n_7964),
.B(n_4407),
.C(n_5158),
.D(n_4439),
.Y(n_8058)
);

NAND3xp33_ASAP7_75t_SL g8059 ( 
.A(n_7969),
.B(n_4559),
.C(n_4506),
.Y(n_8059)
);

NOR3xp33_ASAP7_75t_L g8060 ( 
.A(n_8006),
.B(n_4407),
.C(n_4506),
.Y(n_8060)
);

NAND2xp5_ASAP7_75t_L g8061 ( 
.A(n_7948),
.B(n_4416),
.Y(n_8061)
);

AOI21xp5_ASAP7_75t_L g8062 ( 
.A1(n_7970),
.A2(n_4274),
.B(n_5075),
.Y(n_8062)
);

INVx1_ASAP7_75t_L g8063 ( 
.A(n_7965),
.Y(n_8063)
);

NOR3xp33_ASAP7_75t_L g8064 ( 
.A(n_7983),
.B(n_4564),
.C(n_4559),
.Y(n_8064)
);

AND4x1_ASAP7_75t_L g8065 ( 
.A(n_7958),
.B(n_5151),
.C(n_5171),
.D(n_5143),
.Y(n_8065)
);

NAND4xp25_ASAP7_75t_L g8066 ( 
.A(n_7962),
.B(n_4408),
.C(n_4439),
.D(n_5143),
.Y(n_8066)
);

INVx1_ASAP7_75t_L g8067 ( 
.A(n_7956),
.Y(n_8067)
);

NAND2xp5_ASAP7_75t_SL g8068 ( 
.A(n_7968),
.B(n_4868),
.Y(n_8068)
);

O2A1O1Ixp5_ASAP7_75t_SL g8069 ( 
.A1(n_7996),
.A2(n_4455),
.B(n_4527),
.C(n_4499),
.Y(n_8069)
);

NOR3xp33_ASAP7_75t_L g8070 ( 
.A(n_8008),
.B(n_7982),
.C(n_7981),
.Y(n_8070)
);

INVx1_ASAP7_75t_L g8071 ( 
.A(n_7963),
.Y(n_8071)
);

NAND3xp33_ASAP7_75t_SL g8072 ( 
.A(n_8002),
.B(n_4564),
.C(n_4384),
.Y(n_8072)
);

NAND4xp75_ASAP7_75t_L g8073 ( 
.A(n_7960),
.B(n_4273),
.C(n_4274),
.D(n_4270),
.Y(n_8073)
);

AND2x2_ASAP7_75t_L g8074 ( 
.A(n_7987),
.B(n_5075),
.Y(n_8074)
);

OAI221xp5_ASAP7_75t_L g8075 ( 
.A1(n_7978),
.A2(n_5137),
.B1(n_5004),
.B2(n_5058),
.C(n_4837),
.Y(n_8075)
);

AOI211xp5_ASAP7_75t_SL g8076 ( 
.A1(n_7954),
.A2(n_4499),
.B(n_4527),
.C(n_4455),
.Y(n_8076)
);

NAND3xp33_ASAP7_75t_L g8077 ( 
.A(n_8000),
.B(n_4574),
.C(n_4563),
.Y(n_8077)
);

NOR2x1_ASAP7_75t_L g8078 ( 
.A(n_7959),
.B(n_5004),
.Y(n_8078)
);

AOI221xp5_ASAP7_75t_L g8079 ( 
.A1(n_8011),
.A2(n_4684),
.B1(n_4698),
.B2(n_4700),
.C(n_4550),
.Y(n_8079)
);

NAND5xp2_ASAP7_75t_L g8080 ( 
.A(n_7988),
.B(n_4630),
.C(n_5169),
.D(n_5164),
.E(n_5018),
.Y(n_8080)
);

AOI222xp33_ASAP7_75t_L g8081 ( 
.A1(n_7998),
.A2(n_4666),
.B1(n_4700),
.B2(n_4684),
.C1(n_4643),
.C2(n_4655),
.Y(n_8081)
);

AOI22xp5_ASAP7_75t_L g8082 ( 
.A1(n_8019),
.A2(n_8070),
.B1(n_8063),
.B2(n_8022),
.Y(n_8082)
);

OAI21xp33_ASAP7_75t_L g8083 ( 
.A1(n_8053),
.A2(n_7973),
.B(n_7957),
.Y(n_8083)
);

NAND2xp5_ASAP7_75t_L g8084 ( 
.A(n_8036),
.B(n_8004),
.Y(n_8084)
);

AOI22xp33_ASAP7_75t_L g8085 ( 
.A1(n_8028),
.A2(n_8007),
.B1(n_7991),
.B2(n_8005),
.Y(n_8085)
);

AOI22xp5_ASAP7_75t_L g8086 ( 
.A1(n_8041),
.A2(n_8015),
.B1(n_8010),
.B2(n_7976),
.Y(n_8086)
);

INVx1_ASAP7_75t_L g8087 ( 
.A(n_8024),
.Y(n_8087)
);

AOI221xp5_ASAP7_75t_L g8088 ( 
.A1(n_8020),
.A2(n_7989),
.B1(n_7974),
.B2(n_4430),
.C(n_4596),
.Y(n_8088)
);

AO22x2_ASAP7_75t_L g8089 ( 
.A1(n_8023),
.A2(n_4384),
.B1(n_5139),
.B2(n_5107),
.Y(n_8089)
);

OAI21xp33_ASAP7_75t_L g8090 ( 
.A1(n_8078),
.A2(n_5151),
.B(n_5171),
.Y(n_8090)
);

NAND3xp33_ASAP7_75t_L g8091 ( 
.A(n_8067),
.B(n_4574),
.C(n_4563),
.Y(n_8091)
);

NOR2x1_ASAP7_75t_SL g8092 ( 
.A(n_8071),
.B(n_5004),
.Y(n_8092)
);

INVx1_ASAP7_75t_L g8093 ( 
.A(n_8055),
.Y(n_8093)
);

OAI22xp5_ASAP7_75t_L g8094 ( 
.A1(n_8043),
.A2(n_4385),
.B1(n_4274),
.B2(n_5107),
.Y(n_8094)
);

NOR2x1_ASAP7_75t_L g8095 ( 
.A(n_8031),
.B(n_5004),
.Y(n_8095)
);

NAND2xp5_ASAP7_75t_L g8096 ( 
.A(n_8025),
.B(n_4563),
.Y(n_8096)
);

OAI211xp5_ASAP7_75t_L g8097 ( 
.A1(n_8051),
.A2(n_4399),
.B(n_5139),
.C(n_5099),
.Y(n_8097)
);

XNOR2xp5_ASAP7_75t_L g8098 ( 
.A(n_8065),
.B(n_4830),
.Y(n_8098)
);

XNOR2xp5_ASAP7_75t_L g8099 ( 
.A(n_8074),
.B(n_4830),
.Y(n_8099)
);

INVxp67_ASAP7_75t_SL g8100 ( 
.A(n_8034),
.Y(n_8100)
);

INVx1_ASAP7_75t_L g8101 ( 
.A(n_8068),
.Y(n_8101)
);

NOR2xp33_ASAP7_75t_R g8102 ( 
.A(n_8038),
.B(n_4652),
.Y(n_8102)
);

AOI22xp5_ASAP7_75t_L g8103 ( 
.A1(n_8061),
.A2(n_4868),
.B1(n_5099),
.B2(n_5093),
.Y(n_8103)
);

INVx2_ASAP7_75t_L g8104 ( 
.A(n_8026),
.Y(n_8104)
);

O2A1O1Ixp33_ASAP7_75t_L g8105 ( 
.A1(n_8062),
.A2(n_5058),
.B(n_4837),
.C(n_4830),
.Y(n_8105)
);

INVx1_ASAP7_75t_L g8106 ( 
.A(n_8030),
.Y(n_8106)
);

NOR2xp33_ASAP7_75t_R g8107 ( 
.A(n_8072),
.B(n_4652),
.Y(n_8107)
);

INVx1_ASAP7_75t_L g8108 ( 
.A(n_8044),
.Y(n_8108)
);

INVx1_ASAP7_75t_SL g8109 ( 
.A(n_8032),
.Y(n_8109)
);

INVx1_ASAP7_75t_L g8110 ( 
.A(n_8066),
.Y(n_8110)
);

AOI22xp33_ASAP7_75t_L g8111 ( 
.A1(n_8042),
.A2(n_4868),
.B1(n_4188),
.B2(n_4574),
.Y(n_8111)
);

AOI222xp33_ASAP7_75t_L g8112 ( 
.A1(n_8079),
.A2(n_4399),
.B1(n_5093),
.B2(n_4578),
.C1(n_4643),
.C2(n_4655),
.Y(n_8112)
);

AOI22xp5_ASAP7_75t_L g8113 ( 
.A1(n_8037),
.A2(n_4868),
.B1(n_5058),
.B2(n_4270),
.Y(n_8113)
);

AOI211xp5_ASAP7_75t_SL g8114 ( 
.A1(n_8021),
.A2(n_4455),
.B(n_4527),
.C(n_4499),
.Y(n_8114)
);

AND2x2_ASAP7_75t_L g8115 ( 
.A(n_8056),
.B(n_4868),
.Y(n_8115)
);

INVx1_ASAP7_75t_L g8116 ( 
.A(n_8050),
.Y(n_8116)
);

INVx1_ASAP7_75t_L g8117 ( 
.A(n_8029),
.Y(n_8117)
);

INVx1_ASAP7_75t_L g8118 ( 
.A(n_8058),
.Y(n_8118)
);

INVx1_ASAP7_75t_L g8119 ( 
.A(n_8048),
.Y(n_8119)
);

NAND2xp5_ASAP7_75t_L g8120 ( 
.A(n_8060),
.B(n_4563),
.Y(n_8120)
);

AOI22xp33_ASAP7_75t_SL g8121 ( 
.A1(n_8040),
.A2(n_4868),
.B1(n_4430),
.B2(n_4550),
.Y(n_8121)
);

OAI21xp5_ASAP7_75t_L g8122 ( 
.A1(n_8077),
.A2(n_4273),
.B(n_4270),
.Y(n_8122)
);

NOR2xp33_ASAP7_75t_R g8123 ( 
.A(n_8059),
.B(n_4652),
.Y(n_8123)
);

AND2x4_ASAP7_75t_L g8124 ( 
.A(n_8064),
.B(n_4442),
.Y(n_8124)
);

HB1xp67_ASAP7_75t_L g8125 ( 
.A(n_8046),
.Y(n_8125)
);

NAND2xp33_ASAP7_75t_L g8126 ( 
.A(n_8049),
.B(n_4868),
.Y(n_8126)
);

NAND2xp5_ASAP7_75t_L g8127 ( 
.A(n_8027),
.B(n_4273),
.Y(n_8127)
);

AOI22xp5_ASAP7_75t_L g8128 ( 
.A1(n_8047),
.A2(n_4270),
.B1(n_4837),
.B2(n_4830),
.Y(n_8128)
);

AOI221xp5_ASAP7_75t_SL g8129 ( 
.A1(n_8117),
.A2(n_8083),
.B1(n_8116),
.B2(n_8085),
.C(n_8118),
.Y(n_8129)
);

INVx2_ASAP7_75t_L g8130 ( 
.A(n_8104),
.Y(n_8130)
);

INVx1_ASAP7_75t_L g8131 ( 
.A(n_8125),
.Y(n_8131)
);

INVx1_ASAP7_75t_L g8132 ( 
.A(n_8100),
.Y(n_8132)
);

INVx1_ASAP7_75t_L g8133 ( 
.A(n_8084),
.Y(n_8133)
);

NAND2x1p5_ASAP7_75t_SL g8134 ( 
.A(n_8095),
.B(n_8080),
.Y(n_8134)
);

INVx1_ASAP7_75t_L g8135 ( 
.A(n_8119),
.Y(n_8135)
);

AND2x2_ASAP7_75t_L g8136 ( 
.A(n_8092),
.B(n_8033),
.Y(n_8136)
);

NOR2x1_ASAP7_75t_L g8137 ( 
.A(n_8093),
.B(n_8052),
.Y(n_8137)
);

INVx2_ASAP7_75t_L g8138 ( 
.A(n_8124),
.Y(n_8138)
);

INVxp67_ASAP7_75t_L g8139 ( 
.A(n_8082),
.Y(n_8139)
);

OR2x2_ASAP7_75t_L g8140 ( 
.A(n_8096),
.B(n_8045),
.Y(n_8140)
);

INVx1_ASAP7_75t_L g8141 ( 
.A(n_8109),
.Y(n_8141)
);

INVx1_ASAP7_75t_L g8142 ( 
.A(n_8099),
.Y(n_8142)
);

NAND4xp75_ASAP7_75t_L g8143 ( 
.A(n_8087),
.B(n_8106),
.C(n_8110),
.D(n_8108),
.Y(n_8143)
);

INVx1_ASAP7_75t_L g8144 ( 
.A(n_8086),
.Y(n_8144)
);

INVx1_ASAP7_75t_L g8145 ( 
.A(n_8126),
.Y(n_8145)
);

AND2x2_ASAP7_75t_L g8146 ( 
.A(n_8115),
.B(n_8076),
.Y(n_8146)
);

INVx1_ASAP7_75t_L g8147 ( 
.A(n_8101),
.Y(n_8147)
);

NAND2xp5_ASAP7_75t_L g8148 ( 
.A(n_8088),
.B(n_8069),
.Y(n_8148)
);

NOR3xp33_ASAP7_75t_L g8149 ( 
.A(n_8094),
.B(n_8075),
.C(n_8057),
.Y(n_8149)
);

INVxp33_ASAP7_75t_L g8150 ( 
.A(n_8102),
.Y(n_8150)
);

INVx3_ASAP7_75t_L g8151 ( 
.A(n_8124),
.Y(n_8151)
);

INVx2_ASAP7_75t_L g8152 ( 
.A(n_8098),
.Y(n_8152)
);

INVxp67_ASAP7_75t_SL g8153 ( 
.A(n_8120),
.Y(n_8153)
);

AOI22xp5_ASAP7_75t_L g8154 ( 
.A1(n_8103),
.A2(n_8081),
.B1(n_8073),
.B2(n_8035),
.Y(n_8154)
);

XOR2x1_ASAP7_75t_L g8155 ( 
.A(n_8107),
.B(n_8076),
.Y(n_8155)
);

INVx2_ASAP7_75t_L g8156 ( 
.A(n_8127),
.Y(n_8156)
);

INVx1_ASAP7_75t_L g8157 ( 
.A(n_8123),
.Y(n_8157)
);

NOR2x1_ASAP7_75t_L g8158 ( 
.A(n_8097),
.B(n_8090),
.Y(n_8158)
);

NAND2x1p5_ASAP7_75t_SL g8159 ( 
.A(n_8114),
.B(n_8081),
.Y(n_8159)
);

NAND4xp75_ASAP7_75t_L g8160 ( 
.A(n_8113),
.B(n_8039),
.C(n_8054),
.D(n_4273),
.Y(n_8160)
);

INVx1_ASAP7_75t_SL g8161 ( 
.A(n_8121),
.Y(n_8161)
);

AND2x2_ASAP7_75t_L g8162 ( 
.A(n_8089),
.B(n_5160),
.Y(n_8162)
);

AND2x4_ASAP7_75t_L g8163 ( 
.A(n_8128),
.B(n_4442),
.Y(n_8163)
);

INVx3_ASAP7_75t_L g8164 ( 
.A(n_8089),
.Y(n_8164)
);

AND2x4_ASAP7_75t_L g8165 ( 
.A(n_8122),
.B(n_4442),
.Y(n_8165)
);

AOI211xp5_ASAP7_75t_SL g8166 ( 
.A1(n_8131),
.A2(n_8105),
.B(n_8112),
.C(n_8091),
.Y(n_8166)
);

NOR3xp33_ASAP7_75t_L g8167 ( 
.A(n_8132),
.B(n_8111),
.C(n_4527),
.Y(n_8167)
);

NOR5xp2_ASAP7_75t_L g8168 ( 
.A(n_8139),
.B(n_4182),
.C(n_4184),
.D(n_4124),
.E(n_4052),
.Y(n_8168)
);

AND2x2_ASAP7_75t_L g8169 ( 
.A(n_8131),
.B(n_5160),
.Y(n_8169)
);

HB1xp67_ASAP7_75t_L g8170 ( 
.A(n_8164),
.Y(n_8170)
);

AND3x1_ASAP7_75t_L g8171 ( 
.A(n_8132),
.B(n_4512),
.C(n_4511),
.Y(n_8171)
);

A2O1A1Ixp33_ASAP7_75t_L g8172 ( 
.A1(n_8164),
.A2(n_4581),
.B(n_4534),
.C(n_4566),
.Y(n_8172)
);

NAND4xp75_ASAP7_75t_L g8173 ( 
.A(n_8129),
.B(n_4333),
.C(n_4332),
.D(n_4188),
.Y(n_8173)
);

NAND3xp33_ASAP7_75t_L g8174 ( 
.A(n_8141),
.B(n_4837),
.C(n_4830),
.Y(n_8174)
);

NAND4xp75_ASAP7_75t_L g8175 ( 
.A(n_8137),
.B(n_4333),
.C(n_4332),
.D(n_4188),
.Y(n_8175)
);

AOI22xp33_ASAP7_75t_L g8176 ( 
.A1(n_8141),
.A2(n_4188),
.B1(n_4283),
.B2(n_4296),
.Y(n_8176)
);

NOR3xp33_ASAP7_75t_L g8177 ( 
.A(n_8133),
.B(n_4577),
.C(n_4602),
.Y(n_8177)
);

NOR2x1p5_ASAP7_75t_L g8178 ( 
.A(n_8143),
.B(n_4442),
.Y(n_8178)
);

NAND4xp25_ASAP7_75t_L g8179 ( 
.A(n_8147),
.B(n_8144),
.C(n_8136),
.D(n_8130),
.Y(n_8179)
);

OAI322xp33_ASAP7_75t_L g8180 ( 
.A1(n_8147),
.A2(n_4566),
.A3(n_4534),
.B1(n_4385),
.B2(n_4315),
.C1(n_4363),
.C2(n_4355),
.Y(n_8180)
);

NAND3xp33_ASAP7_75t_L g8181 ( 
.A(n_8135),
.B(n_4837),
.C(n_4550),
.Y(n_8181)
);

NAND4xp25_ASAP7_75t_L g8182 ( 
.A(n_8158),
.B(n_4560),
.C(n_4569),
.D(n_4555),
.Y(n_8182)
);

NOR3xp33_ASAP7_75t_L g8183 ( 
.A(n_8142),
.B(n_4577),
.C(n_4602),
.Y(n_8183)
);

NAND5xp2_ASAP7_75t_L g8184 ( 
.A(n_8149),
.B(n_4630),
.C(n_5164),
.D(n_5169),
.E(n_5160),
.Y(n_8184)
);

AND3x4_ASAP7_75t_L g8185 ( 
.A(n_8152),
.B(n_4674),
.C(n_4439),
.Y(n_8185)
);

NOR2x1_ASAP7_75t_L g8186 ( 
.A(n_8151),
.B(n_4355),
.Y(n_8186)
);

NAND4xp75_ASAP7_75t_L g8187 ( 
.A(n_8157),
.B(n_4333),
.C(n_4332),
.D(n_4283),
.Y(n_8187)
);

NAND4xp25_ASAP7_75t_L g8188 ( 
.A(n_8140),
.B(n_4560),
.C(n_4569),
.D(n_4555),
.Y(n_8188)
);

INVx1_ASAP7_75t_L g8189 ( 
.A(n_8134),
.Y(n_8189)
);

NOR3xp33_ASAP7_75t_L g8190 ( 
.A(n_8153),
.B(n_4618),
.C(n_4609),
.Y(n_8190)
);

NAND4xp75_ASAP7_75t_L g8191 ( 
.A(n_8138),
.B(n_8156),
.C(n_8145),
.D(n_8146),
.Y(n_8191)
);

NOR3xp33_ASAP7_75t_L g8192 ( 
.A(n_8151),
.B(n_4618),
.C(n_4609),
.Y(n_8192)
);

NAND3xp33_ASAP7_75t_L g8193 ( 
.A(n_8150),
.B(n_4550),
.C(n_4442),
.Y(n_8193)
);

NOR3xp33_ASAP7_75t_L g8194 ( 
.A(n_8161),
.B(n_4629),
.C(n_4621),
.Y(n_8194)
);

NOR2xp33_ASAP7_75t_L g8195 ( 
.A(n_8155),
.B(n_4442),
.Y(n_8195)
);

OAI21xp5_ASAP7_75t_L g8196 ( 
.A1(n_8148),
.A2(n_4283),
.B(n_4582),
.Y(n_8196)
);

INVx1_ASAP7_75t_L g8197 ( 
.A(n_8159),
.Y(n_8197)
);

AND2x2_ASAP7_75t_L g8198 ( 
.A(n_8162),
.B(n_5160),
.Y(n_8198)
);

INVx1_ASAP7_75t_L g8199 ( 
.A(n_8154),
.Y(n_8199)
);

AND2x4_ASAP7_75t_L g8200 ( 
.A(n_8163),
.B(n_4550),
.Y(n_8200)
);

OAI22xp33_ASAP7_75t_L g8201 ( 
.A1(n_8189),
.A2(n_8197),
.B1(n_8166),
.B2(n_8179),
.Y(n_8201)
);

INVx1_ASAP7_75t_L g8202 ( 
.A(n_8170),
.Y(n_8202)
);

INVx1_ASAP7_75t_L g8203 ( 
.A(n_8178),
.Y(n_8203)
);

INVxp67_ASAP7_75t_SL g8204 ( 
.A(n_8199),
.Y(n_8204)
);

NAND2xp5_ASAP7_75t_L g8205 ( 
.A(n_8191),
.B(n_8163),
.Y(n_8205)
);

INVx1_ASAP7_75t_SL g8206 ( 
.A(n_8195),
.Y(n_8206)
);

XNOR2xp5_ASAP7_75t_L g8207 ( 
.A(n_8171),
.B(n_8160),
.Y(n_8207)
);

INVx1_ASAP7_75t_L g8208 ( 
.A(n_8169),
.Y(n_8208)
);

INVx1_ASAP7_75t_L g8209 ( 
.A(n_8186),
.Y(n_8209)
);

CKINVDCx20_ASAP7_75t_R g8210 ( 
.A(n_8193),
.Y(n_8210)
);

INVx1_ASAP7_75t_L g8211 ( 
.A(n_8167),
.Y(n_8211)
);

AND2x4_ASAP7_75t_L g8212 ( 
.A(n_8200),
.B(n_8165),
.Y(n_8212)
);

AOI221xp5_ASAP7_75t_L g8213 ( 
.A1(n_8200),
.A2(n_8165),
.B1(n_4550),
.B2(n_4558),
.C(n_4661),
.Y(n_8213)
);

NAND2xp5_ASAP7_75t_L g8214 ( 
.A(n_8183),
.B(n_4283),
.Y(n_8214)
);

HB1xp67_ASAP7_75t_L g8215 ( 
.A(n_8185),
.Y(n_8215)
);

BUFx6f_ASAP7_75t_L g8216 ( 
.A(n_8174),
.Y(n_8216)
);

INVx1_ASAP7_75t_L g8217 ( 
.A(n_8177),
.Y(n_8217)
);

OAI22xp5_ASAP7_75t_L g8218 ( 
.A1(n_8173),
.A2(n_4596),
.B1(n_4646),
.B2(n_4558),
.Y(n_8218)
);

BUFx2_ASAP7_75t_L g8219 ( 
.A(n_8196),
.Y(n_8219)
);

INVxp67_ASAP7_75t_L g8220 ( 
.A(n_8190),
.Y(n_8220)
);

HB1xp67_ASAP7_75t_L g8221 ( 
.A(n_8194),
.Y(n_8221)
);

NOR3xp33_ASAP7_75t_L g8222 ( 
.A(n_8181),
.B(n_3910),
.C(n_3895),
.Y(n_8222)
);

AO221x1_ASAP7_75t_L g8223 ( 
.A1(n_8184),
.A2(n_4661),
.B1(n_4646),
.B2(n_4596),
.C(n_4558),
.Y(n_8223)
);

NOR2xp33_ASAP7_75t_L g8224 ( 
.A(n_8198),
.B(n_4558),
.Y(n_8224)
);

AOI322xp5_ASAP7_75t_L g8225 ( 
.A1(n_8204),
.A2(n_8192),
.A3(n_8176),
.B1(n_8172),
.B2(n_8168),
.C1(n_8188),
.C2(n_8182),
.Y(n_8225)
);

AOI322xp5_ASAP7_75t_L g8226 ( 
.A1(n_8202),
.A2(n_8175),
.A3(n_8187),
.B1(n_8180),
.B2(n_4570),
.C1(n_4545),
.C2(n_4512),
.Y(n_8226)
);

INVx2_ASAP7_75t_L g8227 ( 
.A(n_8212),
.Y(n_8227)
);

AOI322xp5_ASAP7_75t_L g8228 ( 
.A1(n_8201),
.A2(n_4570),
.A3(n_4545),
.B1(n_4511),
.B2(n_4629),
.C1(n_4635),
.C2(n_4621),
.Y(n_8228)
);

OAI322xp33_ASAP7_75t_L g8229 ( 
.A1(n_8209),
.A2(n_4315),
.A3(n_4363),
.B1(n_4581),
.B2(n_4558),
.C1(n_4646),
.C2(n_4596),
.Y(n_8229)
);

AOI22xp5_ASAP7_75t_L g8230 ( 
.A1(n_8205),
.A2(n_4558),
.B1(n_4661),
.B2(n_4596),
.Y(n_8230)
);

OA22x2_ASAP7_75t_L g8231 ( 
.A1(n_8207),
.A2(n_4671),
.B1(n_4631),
.B2(n_4635),
.Y(n_8231)
);

OAI322xp33_ASAP7_75t_SL g8232 ( 
.A1(n_8208),
.A2(n_5160),
.A3(n_4701),
.B1(n_4586),
.B2(n_4696),
.C1(n_4582),
.C2(n_4590),
.Y(n_8232)
);

AOI22xp5_ASAP7_75t_L g8233 ( 
.A1(n_8210),
.A2(n_4596),
.B1(n_4646),
.B2(n_4661),
.Y(n_8233)
);

AND2x2_ASAP7_75t_L g8234 ( 
.A(n_8223),
.B(n_5160),
.Y(n_8234)
);

INVx2_ASAP7_75t_L g8235 ( 
.A(n_8212),
.Y(n_8235)
);

NAND4xp25_ASAP7_75t_L g8236 ( 
.A(n_8206),
.B(n_4631),
.C(n_4594),
.D(n_4592),
.Y(n_8236)
);

HB1xp67_ASAP7_75t_L g8237 ( 
.A(n_8215),
.Y(n_8237)
);

HB1xp67_ASAP7_75t_L g8238 ( 
.A(n_8203),
.Y(n_8238)
);

NOR2x1_ASAP7_75t_L g8239 ( 
.A(n_8211),
.B(n_4674),
.Y(n_8239)
);

OAI221xp5_ASAP7_75t_L g8240 ( 
.A1(n_8219),
.A2(n_4646),
.B1(n_4661),
.B2(n_4333),
.C(n_4332),
.Y(n_8240)
);

A2O1A1Ixp33_ASAP7_75t_L g8241 ( 
.A1(n_8221),
.A2(n_4671),
.B(n_4646),
.C(n_4661),
.Y(n_8241)
);

AOI22xp5_ASAP7_75t_L g8242 ( 
.A1(n_8237),
.A2(n_8216),
.B1(n_8217),
.B2(n_8220),
.Y(n_8242)
);

AOI22xp5_ASAP7_75t_L g8243 ( 
.A1(n_8227),
.A2(n_8216),
.B1(n_8224),
.B2(n_8222),
.Y(n_8243)
);

INVx1_ASAP7_75t_L g8244 ( 
.A(n_8235),
.Y(n_8244)
);

AOI22xp5_ASAP7_75t_L g8245 ( 
.A1(n_8238),
.A2(n_8216),
.B1(n_8214),
.B2(n_8213),
.Y(n_8245)
);

AND4x1_ASAP7_75t_L g8246 ( 
.A(n_8239),
.B(n_8218),
.C(n_4600),
.D(n_4592),
.Y(n_8246)
);

OAI22x1_ASAP7_75t_L g8247 ( 
.A1(n_8234),
.A2(n_4530),
.B1(n_4532),
.B2(n_4552),
.Y(n_8247)
);

INVx2_ASAP7_75t_L g8248 ( 
.A(n_8230),
.Y(n_8248)
);

INVx2_ASAP7_75t_L g8249 ( 
.A(n_8231),
.Y(n_8249)
);

AOI22xp33_ASAP7_75t_L g8250 ( 
.A1(n_8233),
.A2(n_4296),
.B1(n_4651),
.B2(n_4653),
.Y(n_8250)
);

INVx2_ASAP7_75t_L g8251 ( 
.A(n_8225),
.Y(n_8251)
);

INVx2_ASAP7_75t_L g8252 ( 
.A(n_8226),
.Y(n_8252)
);

BUFx2_ASAP7_75t_L g8253 ( 
.A(n_8241),
.Y(n_8253)
);

INVxp67_ASAP7_75t_SL g8254 ( 
.A(n_8236),
.Y(n_8254)
);

NOR3xp33_ASAP7_75t_L g8255 ( 
.A(n_8244),
.B(n_8229),
.C(n_8240),
.Y(n_8255)
);

OR2x6_ASAP7_75t_L g8256 ( 
.A(n_8251),
.B(n_8249),
.Y(n_8256)
);

OAI21xp33_ASAP7_75t_SL g8257 ( 
.A1(n_8242),
.A2(n_8228),
.B(n_8232),
.Y(n_8257)
);

AND2x2_ASAP7_75t_SL g8258 ( 
.A(n_8252),
.B(n_4671),
.Y(n_8258)
);

INVx1_ASAP7_75t_L g8259 ( 
.A(n_8245),
.Y(n_8259)
);

AOI221x1_ASAP7_75t_L g8260 ( 
.A1(n_8248),
.A2(n_4594),
.B1(n_4600),
.B2(n_4168),
.C(n_4650),
.Y(n_8260)
);

OR5x1_ASAP7_75t_L g8261 ( 
.A(n_8243),
.B(n_4591),
.C(n_4597),
.D(n_4370),
.E(n_4390),
.Y(n_8261)
);

OAI221xp5_ASAP7_75t_L g8262 ( 
.A1(n_8254),
.A2(n_4147),
.B1(n_4108),
.B2(n_4107),
.C(n_4696),
.Y(n_8262)
);

NAND3xp33_ASAP7_75t_L g8263 ( 
.A(n_8253),
.B(n_8246),
.C(n_8250),
.Y(n_8263)
);

OR3x1_ASAP7_75t_L g8264 ( 
.A(n_8247),
.B(n_3935),
.C(n_3925),
.Y(n_8264)
);

NAND4xp25_ASAP7_75t_SL g8265 ( 
.A(n_8242),
.B(n_4653),
.C(n_4649),
.D(n_4645),
.Y(n_8265)
);

NAND3xp33_ASAP7_75t_SL g8266 ( 
.A(n_8242),
.B(n_4645),
.C(n_4637),
.Y(n_8266)
);

OAI22xp5_ASAP7_75t_L g8267 ( 
.A1(n_8256),
.A2(n_4674),
.B1(n_4637),
.B2(n_4649),
.Y(n_8267)
);

NAND2xp5_ASAP7_75t_L g8268 ( 
.A(n_8256),
.B(n_4650),
.Y(n_8268)
);

OAI22xp5_ASAP7_75t_SL g8269 ( 
.A1(n_8259),
.A2(n_4176),
.B1(n_4158),
.B2(n_4024),
.Y(n_8269)
);

INVx1_ASAP7_75t_L g8270 ( 
.A(n_8263),
.Y(n_8270)
);

CKINVDCx20_ASAP7_75t_R g8271 ( 
.A(n_8257),
.Y(n_8271)
);

OAI21xp5_ASAP7_75t_L g8272 ( 
.A1(n_8255),
.A2(n_4651),
.B(n_4528),
.Y(n_8272)
);

OAI21xp33_ASAP7_75t_L g8273 ( 
.A1(n_8258),
.A2(n_4682),
.B(n_4681),
.Y(n_8273)
);

OAI22xp5_ASAP7_75t_L g8274 ( 
.A1(n_8264),
.A2(n_4674),
.B1(n_3955),
.B2(n_4024),
.Y(n_8274)
);

NAND2xp5_ASAP7_75t_L g8275 ( 
.A(n_8266),
.B(n_8260),
.Y(n_8275)
);

AOI22xp33_ASAP7_75t_SL g8276 ( 
.A1(n_8271),
.A2(n_8262),
.B1(n_8265),
.B2(n_8261),
.Y(n_8276)
);

AOI22x1_ASAP7_75t_L g8277 ( 
.A1(n_8270),
.A2(n_3955),
.B1(n_4122),
.B2(n_3966),
.Y(n_8277)
);

OAI22xp5_ASAP7_75t_SL g8278 ( 
.A1(n_8275),
.A2(n_4176),
.B1(n_4158),
.B2(n_3966),
.Y(n_8278)
);

NAND2xp5_ASAP7_75t_L g8279 ( 
.A(n_8268),
.B(n_4296),
.Y(n_8279)
);

OAI22xp5_ASAP7_75t_L g8280 ( 
.A1(n_8272),
.A2(n_4699),
.B1(n_4007),
.B2(n_4024),
.Y(n_8280)
);

OAI22x1_ASAP7_75t_L g8281 ( 
.A1(n_8269),
.A2(n_4530),
.B1(n_4552),
.B2(n_4540),
.Y(n_8281)
);

OAI22xp33_ASAP7_75t_L g8282 ( 
.A1(n_8279),
.A2(n_8274),
.B1(n_8267),
.B2(n_8273),
.Y(n_8282)
);

INVx1_ASAP7_75t_L g8283 ( 
.A(n_8276),
.Y(n_8283)
);

AOI21xp5_ASAP7_75t_L g8284 ( 
.A1(n_8283),
.A2(n_8278),
.B(n_8280),
.Y(n_8284)
);

NOR2xp33_ASAP7_75t_L g8285 ( 
.A(n_8282),
.B(n_8277),
.Y(n_8285)
);

AOI22xp5_ASAP7_75t_L g8286 ( 
.A1(n_8285),
.A2(n_8281),
.B1(n_3966),
.B2(n_4007),
.Y(n_8286)
);

AO22x2_ASAP7_75t_L g8287 ( 
.A1(n_8284),
.A2(n_4528),
.B1(n_4518),
.B2(n_4530),
.Y(n_8287)
);

OAI21xp5_ASAP7_75t_L g8288 ( 
.A1(n_8286),
.A2(n_4528),
.B(n_4518),
.Y(n_8288)
);

INVx1_ASAP7_75t_L g8289 ( 
.A(n_8288),
.Y(n_8289)
);

AOI221xp5_ASAP7_75t_L g8290 ( 
.A1(n_8289),
.A2(n_8287),
.B1(n_4532),
.B2(n_4530),
.C(n_4552),
.Y(n_8290)
);

AOI22xp33_ASAP7_75t_L g8291 ( 
.A1(n_8290),
.A2(n_4620),
.B1(n_4532),
.B2(n_4540),
.Y(n_8291)
);

AOI211xp5_ASAP7_75t_L g8292 ( 
.A1(n_8291),
.A2(n_3884),
.B(n_4013),
.C(n_4041),
.Y(n_8292)
);


endmodule