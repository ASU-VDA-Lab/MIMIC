module fake_jpeg_29851_n_187 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_187);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_11),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx8_ASAP7_75t_SL g69 ( 
.A(n_0),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_24),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_0),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_69),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_79),
.Y(n_86)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_1),
.Y(n_79)
);

INVx6_ASAP7_75t_SL g80 ( 
.A(n_54),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_80),
.B(n_56),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

BUFx16f_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_26),
.C(n_49),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_72),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

AND2x4_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_56),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_88),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_80),
.A2(n_85),
.B1(n_76),
.B2(n_82),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_89),
.A2(n_58),
.B1(n_75),
.B2(n_27),
.Y(n_110)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

OR2x2_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_70),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_94),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_84),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_66),
.B1(n_54),
.B2(n_70),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_96),
.A2(n_66),
.B1(n_73),
.B2(n_61),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_99),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_62),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_102),
.A2(n_108),
.B1(n_109),
.B2(n_10),
.Y(n_133)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

BUFx12_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_9),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_60),
.B(n_57),
.C(n_55),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_107),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_100),
.A2(n_68),
.B1(n_67),
.B2(n_65),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_68),
.B1(n_63),
.B2(n_59),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_115),
.B1(n_117),
.B2(n_9),
.Y(n_132)
);

AO22x1_ASAP7_75t_SL g112 ( 
.A1(n_92),
.A2(n_75),
.B1(n_23),
.B2(n_29),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_87),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_75),
.B1(n_3),
.B2(n_5),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_74),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_118),
.B(n_8),
.Y(n_127)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_119),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_120),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_133),
.B1(n_40),
.B2(n_37),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_2),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_122),
.B(n_123),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_7),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_30),
.B(n_48),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_124),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_22),
.C(n_44),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_16),
.C(n_21),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_131),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_114),
.B(n_8),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_130),
.B(n_135),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_132),
.A2(n_41),
.B1(n_17),
.B2(n_19),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_107),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_136),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_11),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_104),
.B(n_52),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_106),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_139),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_103),
.B(n_12),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_14),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_141),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_15),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_143),
.A2(n_150),
.B1(n_125),
.B2(n_38),
.Y(n_165)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_146),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_142),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_142),
.Y(n_148)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_133),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_160),
.Y(n_170)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_158),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_124),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_159),
.A2(n_152),
.B(n_161),
.Y(n_167)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_129),
.C(n_128),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_150),
.C(n_144),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_169),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_35),
.B1(n_39),
.B2(n_143),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_152),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_148),
.B(n_156),
.Y(n_169)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_175),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_172),
.B(n_153),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_179),
.B(n_177),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_180),
.A2(n_172),
.B(n_170),
.Y(n_181)
);

OAI21xp33_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_174),
.B(n_178),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_164),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_173),
.C(n_170),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_173),
.B1(n_162),
.B2(n_171),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_163),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_168),
.Y(n_187)
);


endmodule