module fake_jpeg_8383_n_140 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_140);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_15),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_28),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_0),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_45),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_71),
.Y(n_72)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_1),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_49),
.B(n_40),
.C(n_4),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_73),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_46),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_41),
.B1(n_46),
.B2(n_47),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_42),
.B1(n_50),
.B2(n_53),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_71),
.B(n_47),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_86),
.Y(n_110)
);

NAND3xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_1),
.C(n_2),
.Y(n_86)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_91),
.Y(n_117)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_68),
.A2(n_57),
.B1(n_54),
.B2(n_44),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_59),
.B1(n_55),
.B2(n_48),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_57),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_93),
.A2(n_2),
.B(n_3),
.Y(n_102)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_98),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_116),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_105),
.A2(n_113),
.B1(n_118),
.B2(n_80),
.Y(n_119)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_115),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_76),
.A2(n_43),
.B1(n_38),
.B2(n_5),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_87),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_119),
.A2(n_117),
.B1(n_99),
.B2(n_104),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_123),
.A2(n_124),
.B(n_120),
.Y(n_125)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_110),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_121),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_127),
.B(n_6),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_106),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_130),
.A2(n_112),
.B(n_100),
.Y(n_131)
);

OAI21x1_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_6),
.B(n_7),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_7),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_112),
.B(n_100),
.Y(n_134)
);

NOR3xp33_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_101),
.C(n_111),
.Y(n_135)
);

AOI321xp33_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_121),
.A3(n_81),
.B1(n_114),
.B2(n_85),
.C(n_103),
.Y(n_136)
);

AO21x1_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_74),
.B(n_10),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_8),
.B(n_11),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_14),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_36),
.B(n_17),
.Y(n_140)
);


endmodule