module fake_ariane_1044_n_828 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_828);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_828;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_760;
wire n_591;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_584;
wire n_528;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_756;
wire n_466;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_151;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_158;
wire n_259;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_271;
wire n_507;
wire n_465;
wire n_486;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_365;
wire n_238;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_780;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_705;
wire n_630;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_747;
wire n_741;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_742;
wire n_716;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_804;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_793;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_317;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_10),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_131),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_128),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_146),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_90),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_74),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_121),
.Y(n_158)
);

NOR2xp67_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_81),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_63),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_69),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_11),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_92),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_50),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_107),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_38),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_58),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_95),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_18),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_122),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_83),
.Y(n_172)
);

BUFx10_ASAP7_75t_L g173 ( 
.A(n_61),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_133),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_32),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_94),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_4),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_144),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_101),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_100),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_98),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_106),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_7),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_33),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_72),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_123),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_34),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_149),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_64),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_97),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_86),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_134),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_37),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_87),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_3),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_116),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_26),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_143),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_40),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_43),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_77),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_52),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_112),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_1),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_137),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_108),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_28),
.B(n_119),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_65),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_12),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_68),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_80),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g214 ( 
.A(n_117),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_141),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_154),
.Y(n_216)
);

OAI22x1_ASAP7_75t_SL g217 ( 
.A1(n_151),
.A2(n_184),
.B1(n_178),
.B2(n_162),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_160),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_160),
.Y(n_220)
);

OA21x2_ASAP7_75t_L g221 ( 
.A1(n_156),
.A2(n_0),
.B(n_1),
.Y(n_221)
);

AND2x4_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_0),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_160),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_173),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_153),
.B(n_17),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_183),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_186),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_206),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_173),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_161),
.Y(n_230)
);

AND2x4_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_2),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_192),
.B(n_2),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_214),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_174),
.B(n_3),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_160),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_195),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_160),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_165),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_166),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_160),
.Y(n_241)
);

OAI21x1_ASAP7_75t_L g242 ( 
.A1(n_168),
.A2(n_82),
.B(n_148),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_169),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_171),
.Y(n_244)
);

OAI22x1_ASAP7_75t_SL g245 ( 
.A1(n_213),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_245)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

BUFx8_ASAP7_75t_SL g247 ( 
.A(n_152),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_177),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_194),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_185),
.B(n_5),
.Y(n_250)
);

OAI22x1_ASAP7_75t_SL g251 ( 
.A1(n_189),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_191),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_193),
.Y(n_253)
);

AND2x4_ASAP7_75t_L g254 ( 
.A(n_201),
.B(n_8),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_212),
.B(n_9),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_203),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_210),
.Y(n_257)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_194),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_155),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_194),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_194),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_157),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_158),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_247),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_247),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_229),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_229),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_230),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_R g269 ( 
.A(n_233),
.B(n_163),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_233),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_224),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_226),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_237),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_216),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_237),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_230),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_263),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_259),
.Y(n_278)
);

NAND2xp33_ASAP7_75t_R g279 ( 
.A(n_234),
.B(n_164),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_259),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_200),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_262),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_226),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_R g284 ( 
.A(n_262),
.B(n_167),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_262),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_217),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_224),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_230),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_257),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_243),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_R g291 ( 
.A(n_225),
.B(n_170),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_243),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_246),
.B(n_172),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_248),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_216),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_R g296 ( 
.A(n_260),
.B(n_175),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_230),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_254),
.B(n_176),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_248),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_252),
.Y(n_300)
);

AND2x6_ASAP7_75t_L g301 ( 
.A(n_254),
.B(n_194),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_230),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_226),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_R g304 ( 
.A(n_260),
.B(n_179),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_252),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_228),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_216),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_216),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_256),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_216),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_218),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_222),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_240),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_226),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_268),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_301),
.B(n_232),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_276),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_288),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_290),
.B(n_254),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_297),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_292),
.B(n_235),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_294),
.B(n_235),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_278),
.B(n_246),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_302),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_295),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_299),
.B(n_246),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_274),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_274),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_280),
.B(n_246),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_282),
.B(n_246),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_285),
.B(n_250),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_271),
.B(n_244),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_281),
.B(n_239),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_307),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_312),
.B(n_269),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_291),
.B(n_222),
.Y(n_336)
);

A2O1A1Ixp33_ASAP7_75t_L g337 ( 
.A1(n_305),
.A2(n_255),
.B(n_250),
.C(n_231),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_313),
.B(n_222),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_300),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_272),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_279),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_287),
.B(n_231),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_309),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_283),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_301),
.B(n_255),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_303),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_314),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_277),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_308),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_266),
.B(n_231),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_310),
.Y(n_351)
);

INVxp33_ASAP7_75t_L g352 ( 
.A(n_306),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_311),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_301),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_298),
.B(n_239),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_275),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_301),
.B(n_253),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_301),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_296),
.B(n_304),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_267),
.B(n_253),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_296),
.B(n_218),
.Y(n_361)
);

INVxp33_ASAP7_75t_L g362 ( 
.A(n_284),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_304),
.B(n_218),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_284),
.B(n_218),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_289),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_293),
.B(n_261),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_270),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_273),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_279),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_264),
.B(n_218),
.Y(n_370)
);

OR2x6_ASAP7_75t_L g371 ( 
.A(n_265),
.B(n_245),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_286),
.B(n_256),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_301),
.B(n_261),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_313),
.B(n_256),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_290),
.B(n_256),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_290),
.B(n_256),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_295),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_290),
.B(n_226),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_313),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_290),
.B(n_227),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_301),
.B(n_219),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_271),
.B(n_242),
.Y(n_382)
);

NOR2x1p5_ASAP7_75t_L g383 ( 
.A(n_264),
.B(n_251),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_301),
.B(n_219),
.Y(n_384)
);

NAND3xp33_ASAP7_75t_L g385 ( 
.A(n_279),
.B(n_227),
.C(n_221),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_356),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_242),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_333),
.B(n_220),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_315),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_369),
.B(n_220),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_341),
.B(n_223),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_317),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_358),
.B(n_223),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_354),
.B(n_236),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_331),
.B(n_227),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_355),
.B(n_227),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_337),
.B(n_227),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_376),
.B(n_180),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_328),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_339),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_362),
.B(n_181),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_318),
.Y(n_402)
);

NOR3xp33_ASAP7_75t_SL g403 ( 
.A(n_367),
.B(n_207),
.C(n_187),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_359),
.B(n_188),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_336),
.B(n_332),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_340),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_316),
.A2(n_205),
.B1(n_190),
.B2(n_196),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_325),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_323),
.B(n_198),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_366),
.A2(n_221),
.B(n_249),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_366),
.A2(n_221),
.B(n_249),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_329),
.B(n_199),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_L g413 ( 
.A1(n_316),
.A2(n_345),
.B1(n_385),
.B2(n_357),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_344),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_379),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_349),
.B(n_202),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_327),
.Y(n_417)
);

BUFx4f_ASAP7_75t_L g418 ( 
.A(n_349),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_320),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_368),
.B(n_204),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_328),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_338),
.B(n_208),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_353),
.B(n_221),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_356),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_348),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_365),
.Y(n_426)
);

NOR2x2_ASAP7_75t_L g427 ( 
.A(n_371),
.B(n_9),
.Y(n_427)
);

AND2x2_ASAP7_75t_SL g428 ( 
.A(n_372),
.B(n_209),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_L g429 ( 
.A1(n_382),
.A2(n_241),
.B1(n_238),
.B2(n_236),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_324),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_360),
.B(n_238),
.Y(n_431)
);

NAND3xp33_ASAP7_75t_SL g432 ( 
.A(n_335),
.B(n_241),
.C(n_11),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_346),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_343),
.Y(n_434)
);

BUFx12f_ASAP7_75t_L g435 ( 
.A(n_371),
.Y(n_435)
);

AND2x2_ASAP7_75t_SL g436 ( 
.A(n_349),
.B(n_10),
.Y(n_436)
);

AO22x2_ASAP7_75t_L g437 ( 
.A1(n_350),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_347),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_328),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_325),
.Y(n_440)
);

NAND2xp33_ASAP7_75t_L g441 ( 
.A(n_330),
.B(n_194),
.Y(n_441)
);

O2A1O1Ixp33_ASAP7_75t_L g442 ( 
.A1(n_342),
.A2(n_159),
.B(n_14),
.C(n_15),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_321),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_373),
.B(n_258),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_322),
.B(n_352),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_334),
.B(n_258),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_319),
.A2(n_258),
.B1(n_15),
.B2(n_16),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_351),
.B(n_258),
.Y(n_448)
);

INVx2_ASAP7_75t_SL g449 ( 
.A(n_370),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_325),
.Y(n_450)
);

INVx5_ASAP7_75t_L g451 ( 
.A(n_377),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_377),
.Y(n_452)
);

BUFx12f_ASAP7_75t_SL g453 ( 
.A(n_371),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_378),
.B(n_258),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g455 ( 
.A(n_380),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_377),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_364),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_361),
.B(n_13),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_373),
.B(n_16),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_428),
.A2(n_363),
.B1(n_375),
.B2(n_381),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_406),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_415),
.B(n_326),
.Y(n_462)
);

O2A1O1Ixp33_ASAP7_75t_L g463 ( 
.A1(n_426),
.A2(n_384),
.B(n_381),
.C(n_382),
.Y(n_463)
);

O2A1O1Ixp33_ASAP7_75t_L g464 ( 
.A1(n_422),
.A2(n_384),
.B(n_383),
.C(n_21),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_405),
.B(n_449),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_388),
.B(n_19),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_386),
.B(n_20),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_388),
.B(n_22),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_386),
.B(n_23),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_444),
.A2(n_24),
.B(n_25),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_418),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_444),
.A2(n_27),
.B(n_29),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_391),
.B(n_30),
.Y(n_473)
);

O2A1O1Ixp33_ASAP7_75t_L g474 ( 
.A1(n_442),
.A2(n_443),
.B(n_402),
.C(n_389),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_424),
.B(n_31),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_414),
.Y(n_476)
);

O2A1O1Ixp33_ASAP7_75t_L g477 ( 
.A1(n_392),
.A2(n_35),
.B(n_36),
.C(n_39),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_433),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_410),
.A2(n_41),
.B(n_42),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_419),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_407),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_481)
);

A2O1A1Ixp33_ASAP7_75t_SL g482 ( 
.A1(n_420),
.A2(n_150),
.B(n_48),
.C(n_49),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_424),
.B(n_47),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_425),
.B(n_147),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_408),
.Y(n_485)
);

NAND2xp33_ASAP7_75t_L g486 ( 
.A(n_459),
.B(n_51),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_408),
.Y(n_487)
);

A2O1A1Ixp33_ASAP7_75t_SL g488 ( 
.A1(n_401),
.A2(n_145),
.B(n_54),
.C(n_55),
.Y(n_488)
);

BUFx12f_ASAP7_75t_L g489 ( 
.A(n_435),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_417),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_430),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_391),
.B(n_431),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_400),
.B(n_445),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_418),
.B(n_53),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_434),
.Y(n_495)
);

CKINVDCx8_ASAP7_75t_R g496 ( 
.A(n_451),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_438),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_408),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_413),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_499)
);

AOI21x1_ASAP7_75t_L g500 ( 
.A1(n_423),
.A2(n_60),
.B(n_62),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_397),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_394),
.A2(n_66),
.B(n_67),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_416),
.B(n_70),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_455),
.B(n_457),
.Y(n_504)
);

OR2x6_ASAP7_75t_L g505 ( 
.A(n_437),
.B(n_71),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_436),
.B(n_451),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_453),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_390),
.B(n_73),
.Y(n_508)
);

BUFx4f_ASAP7_75t_L g509 ( 
.A(n_450),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_399),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_451),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_399),
.Y(n_512)
);

O2A1O1Ixp33_ASAP7_75t_L g513 ( 
.A1(n_459),
.A2(n_75),
.B(n_76),
.C(n_78),
.Y(n_513)
);

CKINVDCx6p67_ASAP7_75t_R g514 ( 
.A(n_404),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_421),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_437),
.B(n_79),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_390),
.B(n_84),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_403),
.B(n_85),
.Y(n_518)
);

INVx1_ASAP7_75t_SL g519 ( 
.A(n_507),
.Y(n_519)
);

AOI21x1_ASAP7_75t_L g520 ( 
.A1(n_466),
.A2(n_411),
.B(n_395),
.Y(n_520)
);

OAI21x1_ASAP7_75t_L g521 ( 
.A1(n_479),
.A2(n_394),
.B(n_454),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_480),
.Y(n_522)
);

AOI22x1_ASAP7_75t_L g523 ( 
.A1(n_502),
.A2(n_421),
.B1(n_439),
.B2(n_452),
.Y(n_523)
);

INVx5_ASAP7_75t_L g524 ( 
.A(n_511),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_496),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_478),
.Y(n_526)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_500),
.A2(n_517),
.B(n_508),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_485),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_463),
.A2(n_429),
.B(n_393),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_511),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_485),
.Y(n_531)
);

AOI22x1_ASAP7_75t_L g532 ( 
.A1(n_510),
.A2(n_440),
.B1(n_456),
.B2(n_387),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_491),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g534 ( 
.A1(n_468),
.A2(n_393),
.B(n_458),
.Y(n_534)
);

OAI21x1_ASAP7_75t_L g535 ( 
.A1(n_473),
.A2(n_396),
.B(n_448),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_461),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g537 ( 
.A(n_493),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_485),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_465),
.B(n_412),
.Y(n_539)
);

NAND2x1p5_ASAP7_75t_L g540 ( 
.A(n_509),
.B(n_387),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_487),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_492),
.B(n_409),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_474),
.A2(n_398),
.B(n_441),
.Y(n_543)
);

OA21x2_ASAP7_75t_L g544 ( 
.A1(n_501),
.A2(n_470),
.B(n_472),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_506),
.B(n_432),
.Y(n_545)
);

AO21x2_ASAP7_75t_L g546 ( 
.A1(n_460),
.A2(n_447),
.B(n_446),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_511),
.Y(n_547)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_499),
.A2(n_88),
.B(n_89),
.Y(n_548)
);

BUFx2_ASAP7_75t_R g549 ( 
.A(n_504),
.Y(n_549)
);

AO21x2_ASAP7_75t_L g550 ( 
.A1(n_488),
.A2(n_91),
.B(n_93),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_462),
.B(n_96),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_509),
.Y(n_552)
);

BUFx12f_ASAP7_75t_L g553 ( 
.A(n_489),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_487),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_495),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_487),
.Y(n_556)
);

AO21x2_ASAP7_75t_L g557 ( 
.A1(n_482),
.A2(n_99),
.B(n_102),
.Y(n_557)
);

INVx4_ASAP7_75t_L g558 ( 
.A(n_498),
.Y(n_558)
);

AO21x2_ASAP7_75t_L g559 ( 
.A1(n_486),
.A2(n_103),
.B(n_104),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_514),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_498),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_497),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_498),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_471),
.Y(n_564)
);

OA21x2_ASAP7_75t_L g565 ( 
.A1(n_476),
.A2(n_105),
.B(n_109),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_510),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_537),
.B(n_467),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_522),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_526),
.Y(n_569)
);

AOI21x1_ASAP7_75t_L g570 ( 
.A1(n_520),
.A2(n_481),
.B(n_518),
.Y(n_570)
);

BUFx2_ASAP7_75t_SL g571 ( 
.A(n_525),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_526),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_533),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_536),
.A2(n_505),
.B1(n_516),
.B2(n_490),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_552),
.B(n_512),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_536),
.Y(n_576)
);

AO21x1_ASAP7_75t_L g577 ( 
.A1(n_548),
.A2(n_543),
.B(n_529),
.Y(n_577)
);

AOI21x1_ASAP7_75t_L g578 ( 
.A1(n_520),
.A2(n_515),
.B(n_503),
.Y(n_578)
);

HB1xp67_ASAP7_75t_SL g579 ( 
.A(n_549),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_553),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_555),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_541),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_562),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_530),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_530),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_547),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_540),
.Y(n_587)
);

INVx6_ASAP7_75t_L g588 ( 
.A(n_524),
.Y(n_588)
);

OAI22xp33_ASAP7_75t_L g589 ( 
.A1(n_539),
.A2(n_505),
.B1(n_484),
.B2(n_483),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_541),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_565),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_547),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_565),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_540),
.Y(n_594)
);

AOI21x1_ASAP7_75t_L g595 ( 
.A1(n_527),
.A2(n_513),
.B(n_477),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_542),
.A2(n_512),
.B1(n_475),
.B2(n_469),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_540),
.B(n_494),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_565),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_519),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_554),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_525),
.Y(n_601)
);

AO21x1_ASAP7_75t_L g602 ( 
.A1(n_548),
.A2(n_464),
.B(n_111),
.Y(n_602)
);

OAI21x1_ASAP7_75t_L g603 ( 
.A1(n_535),
.A2(n_110),
.B(n_113),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_541),
.Y(n_604)
);

NAND2x1p5_ASAP7_75t_L g605 ( 
.A(n_524),
.B(n_114),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_544),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_544),
.Y(n_607)
);

OR2x6_ASAP7_75t_L g608 ( 
.A(n_597),
.B(n_552),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_580),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_604),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_580),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_601),
.B(n_567),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_589),
.A2(n_545),
.B1(n_551),
.B2(n_566),
.Y(n_613)
);

INVx4_ASAP7_75t_R g614 ( 
.A(n_579),
.Y(n_614)
);

CKINVDCx16_ASAP7_75t_R g615 ( 
.A(n_601),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_571),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_581),
.B(n_564),
.Y(n_617)
);

CKINVDCx16_ASAP7_75t_R g618 ( 
.A(n_599),
.Y(n_618)
);

OR2x2_ASAP7_75t_L g619 ( 
.A(n_581),
.B(n_554),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_604),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_584),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_R g622 ( 
.A(n_588),
.B(n_560),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_583),
.Y(n_623)
);

CKINVDCx16_ASAP7_75t_R g624 ( 
.A(n_597),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_583),
.B(n_568),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g626 ( 
.A1(n_574),
.A2(n_566),
.B1(n_560),
.B2(n_532),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_573),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_596),
.A2(n_569),
.B1(n_576),
.B2(n_572),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_582),
.Y(n_629)
);

INVx6_ASAP7_75t_SL g630 ( 
.A(n_575),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_R g631 ( 
.A(n_588),
.B(n_553),
.Y(n_631)
);

NAND3xp33_ASAP7_75t_SL g632 ( 
.A(n_602),
.B(n_577),
.C(n_605),
.Y(n_632)
);

BUFx2_ASAP7_75t_L g633 ( 
.A(n_582),
.Y(n_633)
);

BUFx4f_ASAP7_75t_L g634 ( 
.A(n_588),
.Y(n_634)
);

INVx11_ASAP7_75t_L g635 ( 
.A(n_588),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_585),
.Y(n_636)
);

NAND2xp33_ASAP7_75t_SL g637 ( 
.A(n_582),
.B(n_566),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_569),
.B(n_556),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_572),
.A2(n_576),
.B1(n_546),
.B2(n_577),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_586),
.B(n_564),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_602),
.A2(n_546),
.B1(n_559),
.B2(n_561),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_587),
.A2(n_524),
.B1(n_561),
.B2(n_538),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_606),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_592),
.B(n_524),
.Y(n_644)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_600),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_575),
.A2(n_546),
.B1(n_559),
.B2(n_561),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_575),
.B(n_524),
.Y(n_647)
);

XNOR2xp5_ASAP7_75t_L g648 ( 
.A(n_605),
.B(n_427),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_578),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_582),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_587),
.B(n_528),
.Y(n_651)
);

OAI21xp33_ASAP7_75t_L g652 ( 
.A1(n_570),
.A2(n_538),
.B(n_531),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_R g653 ( 
.A(n_587),
.B(n_556),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_582),
.Y(n_654)
);

CKINVDCx16_ASAP7_75t_R g655 ( 
.A(n_590),
.Y(n_655)
);

BUFx12f_ASAP7_75t_L g656 ( 
.A(n_590),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_590),
.Y(n_657)
);

BUFx10_ASAP7_75t_L g658 ( 
.A(n_590),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_590),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_625),
.B(n_627),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_624),
.B(n_643),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_613),
.A2(n_594),
.B1(n_559),
.B2(n_538),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_611),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_643),
.Y(n_664)
);

BUFx2_ASAP7_75t_L g665 ( 
.A(n_622),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_623),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_638),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_610),
.B(n_607),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_617),
.B(n_594),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_638),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_620),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_610),
.B(n_607),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_650),
.B(n_606),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_636),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_619),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_657),
.B(n_578),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_612),
.B(n_594),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_618),
.B(n_531),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_628),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_640),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_649),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_629),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_633),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_639),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_608),
.B(n_598),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_608),
.Y(n_686)
);

INVx8_ASAP7_75t_L g687 ( 
.A(n_608),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_615),
.B(n_531),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_659),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_659),
.B(n_541),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_655),
.B(n_528),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_621),
.B(n_613),
.Y(n_692)
);

BUFx2_ASAP7_75t_SL g693 ( 
.A(n_609),
.Y(n_693)
);

OR2x6_ASAP7_75t_L g694 ( 
.A(n_626),
.B(n_605),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_659),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_645),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_644),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_651),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_654),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_647),
.B(n_541),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_661),
.B(n_616),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_661),
.B(n_648),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_660),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_660),
.B(n_626),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_667),
.Y(n_705)
);

NOR2x1p5_ASAP7_75t_L g706 ( 
.A(n_692),
.B(n_614),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_670),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_668),
.B(n_641),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_681),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_675),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_685),
.B(n_686),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_685),
.B(n_646),
.Y(n_712)
);

AND2x6_ASAP7_75t_L g713 ( 
.A(n_662),
.B(n_593),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_680),
.B(n_658),
.Y(n_714)
);

HB1xp67_ASAP7_75t_L g715 ( 
.A(n_668),
.Y(n_715)
);

OAI221xp5_ASAP7_75t_L g716 ( 
.A1(n_674),
.A2(n_632),
.B1(n_652),
.B2(n_642),
.C(n_634),
.Y(n_716)
);

NAND2x1p5_ASAP7_75t_L g717 ( 
.A(n_665),
.B(n_634),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_681),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_677),
.B(n_698),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_671),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_690),
.B(n_637),
.Y(n_721)
);

OR2x2_ASAP7_75t_L g722 ( 
.A(n_698),
.B(n_632),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_697),
.B(n_642),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_682),
.B(n_656),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_678),
.B(n_658),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_666),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_696),
.B(n_631),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_683),
.B(n_598),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_664),
.Y(n_729)
);

NAND2x1_ASAP7_75t_L g730 ( 
.A(n_705),
.B(n_694),
.Y(n_730)
);

OAI21xp5_ASAP7_75t_L g731 ( 
.A1(n_713),
.A2(n_694),
.B(n_684),
.Y(n_731)
);

NOR2x1_ASAP7_75t_L g732 ( 
.A(n_706),
.B(n_699),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_707),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_719),
.B(n_693),
.Y(n_734)
);

OAI33xp33_ASAP7_75t_L g735 ( 
.A1(n_710),
.A2(n_679),
.A3(n_669),
.B1(n_688),
.B2(n_663),
.B3(n_664),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_703),
.B(n_715),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_715),
.B(n_672),
.Y(n_737)
);

NOR2x1_ASAP7_75t_L g738 ( 
.A(n_727),
.B(n_689),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_704),
.B(n_672),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_720),
.B(n_673),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_711),
.B(n_694),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_711),
.B(n_673),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_701),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_702),
.B(n_663),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_711),
.B(n_695),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_726),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_729),
.B(n_676),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_746),
.Y(n_748)
);

NAND2xp33_ASAP7_75t_L g749 ( 
.A(n_732),
.B(n_717),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_744),
.B(n_717),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_742),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_733),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_731),
.A2(n_721),
.B1(n_716),
.B2(n_723),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_740),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_731),
.A2(n_721),
.B1(n_724),
.B2(n_725),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_737),
.B(n_708),
.Y(n_756)
);

AOI211xp5_ASAP7_75t_L g757 ( 
.A1(n_735),
.A2(n_734),
.B(n_725),
.C(n_722),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_738),
.B(n_714),
.Y(n_758)
);

OAI21xp33_ASAP7_75t_L g759 ( 
.A1(n_757),
.A2(n_740),
.B(n_747),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_753),
.A2(n_735),
.B1(n_757),
.B2(n_713),
.Y(n_760)
);

OAI21xp33_ASAP7_75t_SL g761 ( 
.A1(n_754),
.A2(n_743),
.B(n_736),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_752),
.Y(n_762)
);

O2A1O1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_755),
.A2(n_747),
.B(n_684),
.C(n_739),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_756),
.B(n_745),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_749),
.A2(n_713),
.B1(n_708),
.B2(n_712),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_760),
.B(n_758),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_762),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_764),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_759),
.B(n_751),
.Y(n_769)
);

AOI31xp33_ASAP7_75t_L g770 ( 
.A1(n_761),
.A2(n_750),
.A3(n_758),
.B(n_741),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_763),
.B(n_748),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_768),
.B(n_769),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_766),
.B(n_765),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_770),
.B(n_730),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_767),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_772),
.B(n_771),
.Y(n_776)
);

NOR3xp33_ASAP7_75t_L g777 ( 
.A(n_773),
.B(n_689),
.C(n_695),
.Y(n_777)
);

AOI221xp5_ASAP7_75t_L g778 ( 
.A1(n_776),
.A2(n_775),
.B1(n_774),
.B2(n_712),
.C(n_726),
.Y(n_778)
);

A2O1A1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_777),
.A2(n_774),
.B(n_712),
.C(n_741),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_776),
.A2(n_687),
.B(n_691),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_780),
.B(n_778),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_779),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_778),
.Y(n_783)
);

NOR4xp25_ASAP7_75t_L g784 ( 
.A(n_778),
.B(n_556),
.C(n_528),
.D(n_676),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_780),
.Y(n_785)
);

NOR2x1_ASAP7_75t_L g786 ( 
.A(n_780),
.B(n_558),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_785),
.B(n_713),
.Y(n_787)
);

AND3x4_ASAP7_75t_L g788 ( 
.A(n_783),
.B(n_700),
.C(n_690),
.Y(n_788)
);

AOI21xp33_ASAP7_75t_SL g789 ( 
.A1(n_782),
.A2(n_687),
.B(n_603),
.Y(n_789)
);

NOR3xp33_ASAP7_75t_L g790 ( 
.A(n_781),
.B(n_558),
.C(n_603),
.Y(n_790)
);

OAI211xp5_ASAP7_75t_SL g791 ( 
.A1(n_786),
.A2(n_728),
.B(n_713),
.C(n_595),
.Y(n_791)
);

OR2x2_ASAP7_75t_L g792 ( 
.A(n_784),
.B(n_700),
.Y(n_792)
);

NOR2xp67_ASAP7_75t_L g793 ( 
.A(n_787),
.B(n_784),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_792),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_790),
.Y(n_795)
);

OAI221xp5_ASAP7_75t_L g796 ( 
.A1(n_789),
.A2(n_595),
.B1(n_523),
.B2(n_718),
.C(n_709),
.Y(n_796)
);

INVxp33_ASAP7_75t_SL g797 ( 
.A(n_788),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_791),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_794),
.Y(n_799)
);

XNOR2x1_ASAP7_75t_L g800 ( 
.A(n_793),
.B(n_700),
.Y(n_800)
);

NAND3xp33_ASAP7_75t_SL g801 ( 
.A(n_798),
.B(n_653),
.C(n_558),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_795),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_796),
.Y(n_803)
);

XOR2xp5_ASAP7_75t_L g804 ( 
.A(n_797),
.B(n_563),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_794),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_794),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_794),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_794),
.B(n_690),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_799),
.B(n_557),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_805),
.B(n_635),
.Y(n_810)
);

OAI31xp33_ASAP7_75t_L g811 ( 
.A1(n_802),
.A2(n_718),
.A3(n_709),
.B(n_593),
.Y(n_811)
);

AO22x2_ASAP7_75t_L g812 ( 
.A1(n_806),
.A2(n_557),
.B1(n_550),
.B2(n_591),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_807),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_803),
.A2(n_630),
.B1(n_687),
.B2(n_557),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_804),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_800),
.A2(n_630),
.B1(n_687),
.B2(n_550),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_808),
.B(n_563),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_813),
.A2(n_801),
.B1(n_550),
.B2(n_544),
.Y(n_818)
);

AOI22x1_ASAP7_75t_L g819 ( 
.A1(n_809),
.A2(n_563),
.B1(n_118),
.B2(n_120),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_SL g820 ( 
.A1(n_810),
.A2(n_563),
.B1(n_591),
.B2(n_125),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_815),
.B(n_115),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_816),
.A2(n_527),
.B1(n_563),
.B2(n_535),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_SL g823 ( 
.A1(n_821),
.A2(n_814),
.B1(n_817),
.B2(n_811),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_SL g824 ( 
.A1(n_820),
.A2(n_812),
.B1(n_126),
.B2(n_127),
.Y(n_824)
);

OAI21xp5_ASAP7_75t_L g825 ( 
.A1(n_824),
.A2(n_819),
.B(n_818),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_825),
.A2(n_823),
.B1(n_822),
.B2(n_812),
.Y(n_826)
);

AOI221xp5_ASAP7_75t_L g827 ( 
.A1(n_826),
.A2(n_124),
.B1(n_129),
.B2(n_130),
.C(n_132),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_827),
.A2(n_534),
.B1(n_521),
.B2(n_135),
.Y(n_828)
);


endmodule