module fake_jpeg_14642_n_91 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_91);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_91;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_5),
.B(n_9),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_2),
.B(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_7),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_14),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_24),
.A2(n_31),
.B(n_22),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_18),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_33),
.Y(n_37)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_27),
.A2(n_29),
.B1(n_12),
.B2(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_L g29 ( 
.A1(n_16),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx24_ASAP7_75t_SL g48 ( 
.A(n_30),
.Y(n_48)
);

NAND2xp33_ASAP7_75t_SL g31 ( 
.A(n_18),
.B(n_4),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_21),
.C(n_20),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_21),
.C(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_5),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_39),
.Y(n_63)
);

A2O1A1O1Ixp25_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_22),
.B(n_21),
.C(n_19),
.D(n_17),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_20),
.C(n_9),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_25),
.A2(n_16),
.B1(n_15),
.B2(n_12),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_8),
.B1(n_10),
.B2(n_44),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_26),
.A2(n_21),
.B1(n_19),
.B2(n_13),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_52),
.B1(n_23),
.B2(n_20),
.Y(n_54)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_50),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_17),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_30),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_51),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_23),
.A2(n_24),
.B1(n_13),
.B2(n_8),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_59),
.B1(n_60),
.B2(n_37),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_6),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_56),
.B(n_57),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_7),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_46),
.C(n_56),
.Y(n_70)
);

OAI22x1_ASAP7_75t_SL g60 ( 
.A1(n_38),
.A2(n_10),
.B1(n_39),
.B2(n_42),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_37),
.A2(n_51),
.B(n_41),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_64),
.B(n_58),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_66),
.A2(n_67),
.B1(n_74),
.B2(n_55),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_41),
.B1(n_34),
.B2(n_52),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_48),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_70),
.C(n_73),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_62),
.A2(n_46),
.B1(n_54),
.B2(n_63),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_65),
.B(n_70),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_SL g71 ( 
.A(n_57),
.B(n_61),
.C(n_62),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_73),
.Y(n_80)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_72),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_53),
.B1(n_62),
.B2(n_64),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_55),
.B1(n_65),
.B2(n_67),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_77),
.B(n_78),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_79),
.A2(n_80),
.B(n_77),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_80),
.C(n_79),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_82),
.B(n_76),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_84),
.B(n_87),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_86),
.C(n_83),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_81),
.Y(n_87)
);

BUFx24_ASAP7_75t_SL g90 ( 
.A(n_89),
.Y(n_90)
);

NAND2x1_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_88),
.Y(n_91)
);


endmodule