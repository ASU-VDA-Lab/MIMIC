module fake_jpeg_24077_n_167 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_167);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_10),
.B(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_0),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_36),
.A2(n_40),
.B(n_20),
.C(n_29),
.Y(n_65)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_38),
.B(n_48),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_2),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_14),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_25),
.B1(n_31),
.B2(n_19),
.Y(n_58)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_49),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_46),
.Y(n_75)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_16),
.B1(n_28),
.B2(n_29),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_51),
.A2(n_74),
.B1(n_78),
.B2(n_32),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_2),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_56),
.A2(n_46),
.B(n_33),
.C(n_32),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_15),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_57),
.B(n_26),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_58),
.A2(n_17),
.B(n_32),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_61),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_25),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_65),
.B(n_3),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_20),
.Y(n_66)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_70),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_28),
.C(n_31),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_17),
.C(n_15),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_18),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_21),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_21),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_24),
.Y(n_73)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_37),
.A2(n_24),
.B1(n_22),
.B2(n_19),
.Y(n_74)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_35),
.A2(n_22),
.B1(n_21),
.B2(n_32),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_85),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_86),
.A2(n_60),
.B1(n_52),
.B2(n_62),
.Y(n_102)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_97),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_62),
.A2(n_67),
.B(n_54),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_76),
.C(n_78),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_64),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_93),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_91),
.B(n_92),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_96),
.B(n_56),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_54),
.B(n_46),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_99),
.Y(n_115)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_100),
.A2(n_65),
.B1(n_68),
.B2(n_78),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_85),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_84),
.B(n_72),
.Y(n_129)
);

XOR2x2_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_54),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_104),
.B(n_91),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_93),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_106),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_89),
.A2(n_88),
.B1(n_92),
.B2(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_117),
.Y(n_120)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_78),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_116),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_114),
.C(n_98),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_56),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_55),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_94),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_76),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_80),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_124),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_121),
.A2(n_129),
.B1(n_112),
.B2(n_60),
.Y(n_142)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_122),
.B(n_125),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_81),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_126),
.A2(n_108),
.B(n_107),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_84),
.C(n_53),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_132),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_81),
.Y(n_131)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_52),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_120),
.A2(n_111),
.B(n_126),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_119),
.C(n_127),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_141),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_128),
.A2(n_103),
.B(n_109),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_142),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_127),
.A2(n_101),
.B1(n_114),
.B2(n_116),
.Y(n_143)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_124),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_145),
.B(n_149),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_136),
.C(n_139),
.Y(n_157)
);

NAND4xp25_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_123),
.C(n_121),
.D(n_59),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_148),
.A2(n_150),
.B1(n_141),
.B2(n_75),
.Y(n_153)
);

AO221x1_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_75),
.B1(n_4),
.B2(n_3),
.C(n_130),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_153),
.A2(n_154),
.B(n_151),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_151),
.A2(n_139),
.B1(n_140),
.B2(n_144),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_146),
.B(n_137),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_155),
.B(n_147),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_157),
.B(n_158),
.C(n_145),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_137),
.C(n_83),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_159),
.B(n_162),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_160),
.A2(n_161),
.B(n_156),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_152),
.C(n_83),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_163),
.A2(n_79),
.B(n_6),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_13),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_164),
.Y(n_167)
);


endmodule