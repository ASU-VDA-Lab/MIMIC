module real_aes_7696_n_286 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_286);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_286;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_800;
wire n_778;
wire n_618;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_503;
wire n_635;
wire n_287;
wire n_357;
wire n_386;
wire n_673;
wire n_905;
wire n_518;
wire n_792;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_852;
wire n_766;
wire n_919;
wire n_857;
wire n_461;
wire n_908;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_886;
wire n_856;
wire n_594;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_626;
wire n_292;
wire n_400;
wire n_539;
wire n_625;
wire n_289;
wire n_462;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_726;
wire n_369;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_316;
wire n_656;
wire n_532;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_298;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_898;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_649;
wire n_749;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_915;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_498;
wire n_691;
wire n_765;
wire n_481;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_653;
wire n_365;
wire n_526;
wire n_637;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_922;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_314;
wire n_753;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_639;
wire n_587;
wire n_546;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_0), .A2(n_77), .B1(n_424), .B2(n_631), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_1), .A2(n_43), .B1(n_433), .B2(n_434), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_2), .Y(n_403) );
AOI22xp33_ASAP7_75t_SL g428 ( .A1(n_3), .A2(n_276), .B1(n_429), .B2(n_431), .Y(n_428) );
AOI22xp33_ASAP7_75t_SL g629 ( .A1(n_4), .A2(n_102), .B1(n_344), .B2(n_610), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_5), .A2(n_170), .B1(n_507), .B2(n_919), .Y(n_918) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_6), .A2(n_126), .B1(n_426), .B2(n_433), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g790 ( .A1(n_7), .A2(n_791), .B1(n_815), .B2(n_816), .Y(n_790) );
INVx1_ASAP7_75t_L g815 ( .A(n_7), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_8), .A2(n_221), .B1(n_689), .B2(n_691), .Y(n_688) );
CKINVDCx20_ASAP7_75t_R g379 ( .A(n_9), .Y(n_379) );
INVx1_ASAP7_75t_L g390 ( .A(n_10), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_11), .A2(n_96), .B1(n_349), .B2(n_353), .Y(n_348) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_12), .Y(n_525) );
AOI22xp33_ASAP7_75t_SL g594 ( .A1(n_13), .A2(n_128), .B1(n_448), .B2(n_595), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_14), .A2(n_284), .B1(n_326), .B2(n_610), .Y(n_609) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_15), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_16), .Y(n_405) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_17), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g652 ( .A(n_18), .Y(n_652) );
CKINVDCx20_ASAP7_75t_R g657 ( .A(n_19), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_20), .A2(n_134), .B1(n_411), .B2(n_578), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_21), .A2(n_34), .B1(n_434), .B2(n_503), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_22), .A2(n_150), .B1(n_486), .B2(n_839), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_23), .A2(n_217), .B1(n_422), .B2(n_446), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_24), .A2(n_127), .B1(n_495), .B2(n_542), .Y(n_541) );
AOI22x1_ASAP7_75t_L g736 ( .A1(n_25), .A2(n_737), .B1(n_767), .B2(n_768), .Y(n_736) );
INVx1_ASAP7_75t_L g767 ( .A(n_25), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_26), .A2(n_280), .B1(n_531), .B2(n_626), .Y(n_783) );
AO22x2_ASAP7_75t_L g321 ( .A1(n_27), .A2(n_91), .B1(n_313), .B2(n_318), .Y(n_321) );
INVx1_ASAP7_75t_L g864 ( .A(n_27), .Y(n_864) );
CKINVDCx20_ASAP7_75t_R g789 ( .A(n_28), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_29), .A2(n_249), .B1(n_433), .B2(n_434), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_30), .A2(n_181), .B1(n_307), .B2(n_324), .Y(n_306) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_31), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g590 ( .A(n_32), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_33), .A2(n_268), .B1(n_344), .B2(n_566), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_35), .A2(n_136), .B1(n_324), .B2(n_472), .Y(n_471) );
AOI22xp33_ASAP7_75t_SL g633 ( .A1(n_36), .A2(n_46), .B1(n_341), .B2(n_498), .Y(n_633) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_37), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_38), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_39), .B(n_381), .Y(n_380) );
CKINVDCx20_ASAP7_75t_R g588 ( .A(n_40), .Y(n_588) );
INVx1_ASAP7_75t_L g359 ( .A(n_41), .Y(n_359) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_42), .Y(n_386) );
AO22x2_ASAP7_75t_L g323 ( .A1(n_44), .A2(n_93), .B1(n_313), .B2(n_314), .Y(n_323) );
INVx1_ASAP7_75t_L g865 ( .A(n_44), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_45), .A2(n_101), .B1(n_544), .B2(n_607), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_47), .A2(n_162), .B1(n_326), .B2(n_635), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_48), .A2(n_208), .B1(n_549), .B2(n_745), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_49), .Y(n_837) );
AOI22xp33_ASAP7_75t_SL g914 ( .A1(n_50), .A2(n_107), .B1(n_497), .B2(n_691), .Y(n_914) );
AOI211xp5_ASAP7_75t_L g286 ( .A1(n_51), .A2(n_287), .B(n_295), .C(n_866), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_52), .Y(n_570) );
AOI22xp33_ASAP7_75t_SL g882 ( .A1(n_53), .A2(n_204), .B1(n_422), .B2(n_424), .Y(n_882) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_54), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_55), .B(n_451), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_56), .A2(n_197), .B1(n_694), .B2(n_917), .Y(n_916) );
CKINVDCx20_ASAP7_75t_R g363 ( .A(n_57), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_58), .A2(n_216), .B1(n_350), .B2(n_472), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_59), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_60), .A2(n_90), .B1(n_331), .B2(n_422), .Y(n_421) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_61), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_62), .A2(n_109), .B1(n_308), .B2(n_468), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_63), .A2(n_235), .B1(n_382), .B2(n_448), .Y(n_447) );
AOI22xp33_ASAP7_75t_SL g470 ( .A1(n_64), .A2(n_241), .B1(n_429), .B2(n_431), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_65), .A2(n_173), .B1(n_340), .B2(n_343), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_66), .A2(n_174), .B1(n_587), .B2(n_626), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_67), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_68), .A2(n_132), .B1(n_464), .B2(n_745), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_69), .B(n_381), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_70), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_71), .A2(n_88), .B1(n_382), .B2(n_679), .Y(n_678) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_72), .Y(n_711) );
CKINVDCx20_ASAP7_75t_R g873 ( .A(n_73), .Y(n_873) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_74), .A2(n_137), .B1(n_417), .B2(n_578), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g592 ( .A(n_75), .Y(n_592) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_76), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g831 ( .A(n_78), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_79), .A2(n_227), .B1(n_597), .B2(n_599), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_80), .A2(n_129), .B1(n_307), .B2(n_331), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_81), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_82), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_83), .A2(n_193), .B1(n_329), .B2(n_334), .Y(n_328) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_84), .Y(n_722) );
AOI222xp33_ASAP7_75t_L g787 ( .A1(n_85), .A2(n_159), .B1(n_168), .B2(n_368), .C1(n_448), .C2(n_788), .Y(n_787) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_86), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_87), .A2(n_194), .B1(n_424), .B2(n_426), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_89), .A2(n_153), .B1(n_459), .B2(n_572), .Y(n_571) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_92), .Y(n_682) );
AOI22xp33_ASAP7_75t_SL g913 ( .A1(n_94), .A2(n_190), .B1(n_604), .B2(n_687), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_95), .A2(n_171), .B1(n_502), .B2(n_503), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_97), .Y(n_799) );
AND2x2_ASAP7_75t_L g293 ( .A(n_98), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g803 ( .A(n_99), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_100), .A2(n_200), .B1(n_497), .B2(n_827), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_103), .A2(n_198), .B1(n_353), .B2(n_750), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g905 ( .A(n_104), .Y(n_905) );
INVx1_ASAP7_75t_L g290 ( .A(n_105), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_106), .A2(n_175), .B1(n_422), .B2(n_726), .Y(n_785) );
INVx1_ASAP7_75t_L g802 ( .A(n_108), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_110), .A2(n_154), .B1(n_341), .B2(n_343), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_111), .A2(n_135), .B1(n_383), .B2(n_654), .Y(n_653) );
CKINVDCx20_ASAP7_75t_R g833 ( .A(n_112), .Y(n_833) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_113), .A2(n_272), .B1(n_383), .B2(n_411), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_114), .A2(n_244), .B1(n_542), .B2(n_562), .Y(n_561) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_115), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_116), .A2(n_195), .B1(n_824), .B2(n_825), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_117), .A2(n_251), .B1(n_624), .B2(n_848), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_118), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g906 ( .A(n_119), .Y(n_906) );
AOI22xp33_ASAP7_75t_SL g879 ( .A1(n_120), .A2(n_123), .B1(n_411), .B2(n_626), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_121), .A2(n_231), .B1(n_505), .B2(n_508), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_122), .B(n_455), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_124), .A2(n_226), .B1(n_334), .B2(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_125), .B(n_598), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_130), .A2(n_133), .B1(n_544), .B2(n_778), .Y(n_777) );
OA22x2_ASAP7_75t_L g643 ( .A1(n_131), .A2(n_644), .B1(n_645), .B2(n_665), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_131), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_138), .A2(n_140), .B1(n_811), .B2(n_812), .Y(n_810) );
INVxp67_ASAP7_75t_L g895 ( .A(n_139), .Y(n_895) );
XOR2x2_ASAP7_75t_L g897 ( .A(n_139), .B(n_898), .Y(n_897) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_141), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_142), .B(n_622), .Y(n_621) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_143), .Y(n_760) );
XNOR2x2_ASAP7_75t_L g819 ( .A(n_144), .B(n_820), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g372 ( .A(n_145), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_146), .A2(n_242), .B1(n_426), .B2(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g294 ( .A(n_147), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_148), .B(n_486), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_149), .Y(n_834) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_151), .A2(n_303), .B1(n_397), .B2(n_398), .Y(n_302) );
INVx1_ASAP7_75t_L g397 ( .A(n_151), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_152), .B(n_877), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_155), .A2(n_218), .B1(n_497), .B2(n_499), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_156), .Y(n_740) );
AND2x6_ASAP7_75t_L g289 ( .A(n_157), .B(n_290), .Y(n_289) );
HB1xp67_ASAP7_75t_L g858 ( .A(n_157), .Y(n_858) );
AO22x2_ASAP7_75t_L g312 ( .A1(n_158), .A2(n_230), .B1(n_313), .B2(n_314), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_160), .A2(n_191), .B1(n_549), .B2(n_694), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g903 ( .A(n_161), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_163), .A2(n_184), .B1(n_340), .B2(n_343), .Y(n_339) );
AOI22xp33_ASAP7_75t_SL g842 ( .A1(n_164), .A2(n_248), .B1(n_843), .B2(n_845), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_165), .B(n_624), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_166), .A2(n_261), .B1(n_350), .B2(n_424), .Y(n_663) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_167), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_169), .A2(n_215), .B1(n_374), .B2(n_566), .Y(n_661) );
INVx1_ASAP7_75t_L g696 ( .A(n_172), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_176), .A2(n_189), .B1(n_458), .B2(n_459), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g672 ( .A(n_177), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_178), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_179), .Y(n_829) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_180), .A2(n_211), .B1(n_341), .B2(n_717), .Y(n_716) );
AOI22xp33_ASAP7_75t_SL g885 ( .A1(n_182), .A2(n_256), .B1(n_542), .B2(n_811), .Y(n_885) );
AOI22xp33_ASAP7_75t_SL g886 ( .A1(n_183), .A2(n_265), .B1(n_326), .B2(n_426), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_185), .A2(n_285), .B1(n_464), .B2(n_466), .Y(n_463) );
INVx1_ASAP7_75t_L g481 ( .A(n_186), .Y(n_481) );
AO22x2_ASAP7_75t_L g317 ( .A1(n_187), .A2(n_253), .B1(n_313), .B2(n_318), .Y(n_317) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_188), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_192), .A2(n_277), .B1(n_549), .B2(n_552), .Y(n_548) );
AOI22xp5_ASAP7_75t_SL g474 ( .A1(n_196), .A2(n_475), .B1(n_510), .B2(n_511), .Y(n_474) );
INVx1_ASAP7_75t_L g511 ( .A(n_196), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_199), .Y(n_798) );
AOI22xp5_ASAP7_75t_L g520 ( .A1(n_201), .A2(n_521), .B1(n_554), .B2(n_555), .Y(n_520) );
INVx1_ASAP7_75t_L g554 ( .A(n_201), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g910 ( .A(n_202), .Y(n_910) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_203), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_205), .Y(n_656) );
AOI22xp33_ASAP7_75t_SL g883 ( .A1(n_206), .A2(n_233), .B1(n_498), .B2(n_635), .Y(n_883) );
AOI22xp33_ASAP7_75t_SL g874 ( .A1(n_207), .A2(n_255), .B1(n_458), .B2(n_578), .Y(n_874) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_209), .A2(n_228), .B1(n_411), .B2(n_578), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_210), .Y(n_795) );
INVx1_ASAP7_75t_L g484 ( .A(n_212), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_213), .Y(n_748) );
XOR2xp5_ASAP7_75t_SL g867 ( .A(n_214), .B(n_868), .Y(n_867) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_219), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_220), .A2(n_243), .B1(n_499), .B2(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_222), .B(n_451), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_223), .A2(n_260), .B1(n_686), .B2(n_687), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_224), .Y(n_727) );
INVx1_ASAP7_75t_L g478 ( .A(n_225), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g648 ( .A(n_229), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g862 ( .A(n_230), .B(n_863), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_232), .A2(n_238), .B1(n_334), .B2(n_424), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g901 ( .A(n_234), .Y(n_901) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_236), .Y(n_762) );
INVx1_ASAP7_75t_L g558 ( .A(n_237), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_239), .A2(n_281), .B1(n_353), .B2(n_544), .Y(n_808) );
INVx1_ASAP7_75t_L g435 ( .A(n_240), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_245), .Y(n_473) );
OA22x2_ASAP7_75t_L g581 ( .A1(n_246), .A2(n_582), .B1(n_583), .B2(n_612), .Y(n_581) );
CKINVDCx20_ASAP7_75t_R g582 ( .A(n_246), .Y(n_582) );
INVx1_ASAP7_75t_L g483 ( .A(n_247), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_250), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_252), .B(n_382), .Y(n_800) );
INVx1_ASAP7_75t_L g861 ( .A(n_253), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_254), .A2(n_270), .B1(n_422), .B2(n_566), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_257), .A2(n_262), .B1(n_334), .B2(n_433), .Y(n_664) );
CKINVDCx20_ASAP7_75t_R g909 ( .A(n_258), .Y(n_909) );
INVx1_ASAP7_75t_L g489 ( .A(n_259), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_263), .B(n_587), .Y(n_907) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_264), .Y(n_720) );
INVx1_ASAP7_75t_L g313 ( .A(n_266), .Y(n_313) );
INVx1_ASAP7_75t_L g315 ( .A(n_266), .Y(n_315) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_267), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_269), .Y(n_535) );
INVx1_ASAP7_75t_L g490 ( .A(n_271), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g618 ( .A(n_273), .Y(n_618) );
CKINVDCx20_ASAP7_75t_R g674 ( .A(n_274), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_275), .Y(n_676) );
OA22x2_ASAP7_75t_L g699 ( .A1(n_278), .A2(n_700), .B1(n_701), .B2(n_702), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_278), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_279), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g414 ( .A(n_282), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_283), .Y(n_766) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
HB1xp67_ASAP7_75t_L g857 ( .A(n_290), .Y(n_857) );
OAI21xp5_ASAP7_75t_L g893 ( .A1(n_291), .A2(n_856), .B(n_894), .Y(n_893) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_292), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_734), .B1(n_851), .B2(n_852), .C(n_853), .Y(n_295) );
INVx1_ASAP7_75t_L g851 ( .A(n_296), .Y(n_851) );
XNOR2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_513), .Y(n_296) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B1(n_437), .B2(n_512), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_302), .B1(n_399), .B2(n_436), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g398 ( .A(n_303), .Y(n_398) );
AND2x2_ASAP7_75t_SL g303 ( .A(n_304), .B(n_357), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_305), .B(n_338), .Y(n_304) );
NAND2xp33_ASAP7_75t_SL g305 ( .A(n_306), .B(n_328), .Y(n_305) );
BUFx3_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx3_ASAP7_75t_L g495 ( .A(n_308), .Y(n_495) );
INVx3_ASAP7_75t_L g605 ( .A(n_308), .Y(n_605) );
BUFx6f_ASAP7_75t_L g824 ( .A(n_308), .Y(n_824) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g425 ( .A(n_309), .Y(n_425) );
BUFx2_ASAP7_75t_SL g686 ( .A(n_309), .Y(n_686) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_319), .Y(n_309) );
AND2x6_ASAP7_75t_L g331 ( .A(n_310), .B(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g341 ( .A(n_310), .B(n_342), .Y(n_341) );
AND2x6_ASAP7_75t_L g370 ( .A(n_310), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_316), .Y(n_310) );
AND2x2_ASAP7_75t_L g327 ( .A(n_311), .B(n_317), .Y(n_327) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_312), .B(n_317), .Y(n_337) );
AND2x2_ASAP7_75t_L g346 ( .A(n_312), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g378 ( .A(n_312), .B(n_321), .Y(n_378) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g318 ( .A(n_315), .Y(n_318) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g347 ( .A(n_317), .Y(n_347) );
INVx1_ASAP7_75t_L g377 ( .A(n_317), .Y(n_377) );
AND2x4_ASAP7_75t_L g326 ( .A(n_319), .B(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g335 ( .A(n_319), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g345 ( .A(n_319), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_319), .B(n_346), .Y(n_731) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
OR2x2_ASAP7_75t_L g333 ( .A(n_320), .B(n_323), .Y(n_333) );
AND2x2_ASAP7_75t_L g342 ( .A(n_320), .B(n_323), .Y(n_342) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g371 ( .A(n_321), .B(n_323), .Y(n_371) );
AND2x2_ASAP7_75t_L g376 ( .A(n_322), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g389 ( .A(n_322), .Y(n_389) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g356 ( .A(n_323), .Y(n_356) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx3_ASAP7_75t_L g433 ( .A(n_326), .Y(n_433) );
BUFx3_ASAP7_75t_L g503 ( .A(n_326), .Y(n_503) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_326), .Y(n_551) );
INVx1_ASAP7_75t_L g362 ( .A(n_327), .Y(n_362) );
NAND2x1p5_ASAP7_75t_L g365 ( .A(n_327), .B(n_342), .Y(n_365) );
AND2x4_ASAP7_75t_L g453 ( .A(n_327), .B(n_332), .Y(n_453) );
AND2x6_ASAP7_75t_L g456 ( .A(n_327), .B(n_342), .Y(n_456) );
INVx4_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx4_ASAP7_75t_L g542 ( .A(n_330), .Y(n_542) );
OAI21xp33_ASAP7_75t_SL g651 ( .A1(n_330), .A2(n_652), .B(n_653), .Y(n_651) );
INVx2_ASAP7_75t_SL g694 ( .A(n_330), .Y(n_694) );
INVx11_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx11_ASAP7_75t_L g465 ( .A(n_331), .Y(n_465) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g361 ( .A(n_333), .B(n_362), .Y(n_361) );
BUFx3_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx2_ASAP7_75t_L g426 ( .A(n_335), .Y(n_426) );
BUFx3_ASAP7_75t_L g468 ( .A(n_335), .Y(n_468) );
BUFx3_ASAP7_75t_L g631 ( .A(n_335), .Y(n_631) );
BUFx2_ASAP7_75t_SL g687 ( .A(n_335), .Y(n_687) );
BUFx2_ASAP7_75t_SL g825 ( .A(n_335), .Y(n_825) );
AND2x2_ASAP7_75t_L g472 ( .A(n_336), .B(n_389), .Y(n_472) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OR2x6_ASAP7_75t_L g355 ( .A(n_337), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_348), .Y(n_338) );
BUFx3_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx6_ASAP7_75t_L g430 ( .A(n_341), .Y(n_430) );
BUFx3_ASAP7_75t_L g507 ( .A(n_341), .Y(n_507) );
BUFx3_ASAP7_75t_L g566 ( .A(n_341), .Y(n_566) );
AND2x2_ASAP7_75t_L g352 ( .A(n_342), .B(n_346), .Y(n_352) );
BUFx3_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx3_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx3_ASAP7_75t_L g422 ( .A(n_345), .Y(n_422) );
BUFx3_ASAP7_75t_L g466 ( .A(n_345), .Y(n_466) );
BUFx3_ASAP7_75t_L g920 ( .A(n_345), .Y(n_920) );
INVx1_ASAP7_75t_L g396 ( .A(n_347), .Y(n_396) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx2_ASAP7_75t_L g750 ( .A(n_350), .Y(n_750) );
INVx5_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx3_ASAP7_75t_L g431 ( .A(n_351), .Y(n_431) );
INVx4_ASAP7_75t_L g498 ( .A(n_351), .Y(n_498) );
BUFx3_ASAP7_75t_L g545 ( .A(n_351), .Y(n_545) );
INVx1_ASAP7_75t_L g717 ( .A(n_351), .Y(n_717) );
INVx8_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx4f_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
BUFx2_ASAP7_75t_L g434 ( .A(n_354), .Y(n_434) );
BUFx2_ASAP7_75t_L g499 ( .A(n_354), .Y(n_499) );
BUFx2_ASAP7_75t_L g827 ( .A(n_354), .Y(n_827) );
INVx6_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_SL g607 ( .A(n_355), .Y(n_607) );
INVx1_ASAP7_75t_SL g635 ( .A(n_355), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_355), .A2(n_393), .B1(n_656), .B2(n_657), .Y(n_655) );
INVx1_ASAP7_75t_L g691 ( .A(n_355), .Y(n_691) );
INVx1_ASAP7_75t_L g460 ( .A(n_356), .Y(n_460) );
NOR3xp33_ASAP7_75t_L g357 ( .A(n_358), .B(n_366), .C(n_385), .Y(n_357) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_360), .B1(n_363), .B2(n_364), .Y(n_358) );
INVx1_ASAP7_75t_L g755 ( .A(n_360), .Y(n_755) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx3_ASAP7_75t_L g404 ( .A(n_361), .Y(n_404) );
INVx2_ASAP7_75t_L g480 ( .A(n_361), .Y(n_480) );
OAI221xp5_ASAP7_75t_L g568 ( .A1(n_361), .A2(n_364), .B1(n_569), .B2(n_570), .C(n_571), .Y(n_568) );
INVx2_ASAP7_75t_L g527 ( .A(n_364), .Y(n_527) );
BUFx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g407 ( .A(n_365), .Y(n_407) );
OAI221xp5_ASAP7_75t_SL g366 ( .A1(n_367), .A2(n_372), .B1(n_373), .B2(n_379), .C(n_380), .Y(n_366) );
OAI221xp5_ASAP7_75t_SL g482 ( .A1(n_367), .A2(n_373), .B1(n_483), .B2(n_484), .C(n_485), .Y(n_482) );
OAI221xp5_ASAP7_75t_SL g528 ( .A1(n_367), .A2(n_529), .B1(n_530), .B2(n_532), .C(n_533), .Y(n_528) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx4_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OAI21xp5_ASAP7_75t_SL g408 ( .A1(n_369), .A2(n_409), .B(n_410), .Y(n_408) );
BUFx2_ASAP7_75t_L g677 ( .A(n_369), .Y(n_677) );
INVx4_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_370), .Y(n_446) );
BUFx3_ASAP7_75t_L g575 ( .A(n_370), .Y(n_575) );
INVx2_ASAP7_75t_L g617 ( .A(n_370), .Y(n_617) );
INVx2_ASAP7_75t_L g797 ( .A(n_370), .Y(n_797) );
INVx1_ASAP7_75t_L g394 ( .A(n_371), .Y(n_394) );
AND2x4_ASAP7_75t_L g412 ( .A(n_371), .B(n_396), .Y(n_412) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
BUFx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_375), .Y(n_417) );
BUFx4f_ASAP7_75t_SL g458 ( .A(n_375), .Y(n_458) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_375), .Y(n_531) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_375), .Y(n_587) );
AND2x4_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
INVx1_ASAP7_75t_L g384 ( .A(n_377), .Y(n_384) );
AND2x4_ASAP7_75t_L g383 ( .A(n_378), .B(n_384), .Y(n_383) );
NAND2x1p5_ASAP7_75t_L g388 ( .A(n_378), .B(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g459 ( .A(n_378), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g761 ( .A(n_381), .Y(n_761) );
BUFx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_383), .Y(n_487) );
BUFx12f_ASAP7_75t_L g578 ( .A(n_383), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B1(n_390), .B2(n_391), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_387), .A2(n_491), .B1(n_909), .B2(n_910), .Y(n_908) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_388), .A2(n_414), .B1(n_415), .B2(n_418), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_388), .A2(n_489), .B1(n_490), .B2(n_491), .Y(n_488) );
INVx4_ASAP7_75t_L g537 ( .A(n_388), .Y(n_537) );
BUFx3_ASAP7_75t_L g713 ( .A(n_388), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_391), .A2(n_535), .B1(n_536), .B2(n_538), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g763 ( .A1(n_391), .A2(n_764), .B1(n_765), .B2(n_766), .Y(n_763) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g491 ( .A(n_392), .Y(n_491) );
CKINVDCx16_ASAP7_75t_R g392 ( .A(n_393), .Y(n_392) );
BUFx2_ASAP7_75t_L g804 ( .A(n_393), .Y(n_804) );
OR2x6_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g436 ( .A(n_399), .Y(n_436) );
XOR2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_435), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_419), .Y(n_400) );
NOR3xp33_ASAP7_75t_L g401 ( .A(n_402), .B(n_408), .C(n_413), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_404), .B1(n_405), .B2(n_406), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_404), .A2(n_648), .B1(n_649), .B2(n_650), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_404), .A2(n_526), .B1(n_794), .B2(n_795), .Y(n_793) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_406), .A2(n_478), .B1(n_479), .B2(n_481), .Y(n_477) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g650 ( .A(n_407), .Y(n_650) );
BUFx2_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
BUFx2_ASAP7_75t_SL g448 ( .A(n_412), .Y(n_448) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_412), .Y(n_572) );
OAI221xp5_ASAP7_75t_L g796 ( .A1(n_415), .A2(n_797), .B1(n_798), .B2(n_799), .C(n_800), .Y(n_796) );
INVx2_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_SL g758 ( .A(n_416), .Y(n_758) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_420), .B(n_427), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_423), .Y(n_420) );
INVx1_ASAP7_75t_L g813 ( .A(n_422), .Y(n_813) );
INVx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx3_ASAP7_75t_L g562 ( .A(n_425), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_432), .Y(n_427) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g778 ( .A(n_430), .Y(n_778) );
INVx3_ASAP7_75t_L g811 ( .A(n_430), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g832 ( .A1(n_430), .A2(n_729), .B1(n_833), .B2(n_834), .Y(n_832) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_433), .Y(n_742) );
INVx4_ASAP7_75t_L g512 ( .A(n_437), .Y(n_512) );
XOR2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_474), .Y(n_437) );
INVx2_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
INVx3_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
XOR2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_473), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_442), .B(n_461), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_443), .B(n_449), .Y(n_442) );
OAI21xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_445), .B(n_447), .Y(n_443) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_SL g589 ( .A(n_446), .Y(n_589) );
NAND3xp33_ASAP7_75t_L g449 ( .A(n_450), .B(n_454), .C(n_457), .Y(n_449) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx5_ASAP7_75t_L g598 ( .A(n_452), .Y(n_598) );
INVx2_ASAP7_75t_L g622 ( .A(n_452), .Y(n_622) );
INVx2_ASAP7_75t_L g848 ( .A(n_452), .Y(n_848) );
INVx4_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx4f_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_SL g600 ( .A(n_456), .Y(n_600) );
BUFx2_ASAP7_75t_L g624 ( .A(n_456), .Y(n_624) );
BUFx2_ASAP7_75t_L g595 ( .A(n_459), .Y(n_595) );
BUFx3_ASAP7_75t_L g626 ( .A(n_459), .Y(n_626) );
BUFx2_ASAP7_75t_L g654 ( .A(n_459), .Y(n_654) );
INVx1_ASAP7_75t_L g844 ( .A(n_459), .Y(n_844) );
NOR2x1_ASAP7_75t_L g461 ( .A(n_462), .B(n_469), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_467), .Y(n_462) );
INVx4_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g502 ( .A(n_465), .Y(n_502) );
INVx5_ASAP7_75t_SL g610 ( .A(n_465), .Y(n_610) );
INVx1_ASAP7_75t_L g726 ( .A(n_465), .Y(n_726) );
INVx1_ASAP7_75t_L g509 ( .A(n_466), .Y(n_509) );
INVx2_ASAP7_75t_L g553 ( .A(n_468), .Y(n_553) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_468), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVx1_ASAP7_75t_SL g510 ( .A(n_475), .Y(n_510) );
AND2x2_ASAP7_75t_SL g475 ( .A(n_476), .B(n_492), .Y(n_475) );
NOR3xp33_ASAP7_75t_L g476 ( .A(n_477), .B(n_482), .C(n_488), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_479), .A2(n_524), .B1(n_525), .B2(n_526), .Y(n_523) );
OAI22xp5_ASAP7_75t_SL g704 ( .A1(n_479), .A2(n_526), .B1(n_705), .B2(n_706), .Y(n_704) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_SL g673 ( .A(n_480), .Y(n_673) );
INVx2_ASAP7_75t_L g902 ( .A(n_480), .Y(n_902) );
INVx1_ASAP7_75t_L g591 ( .A(n_486), .Y(n_591) );
BUFx4f_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_491), .A2(n_536), .B1(n_681), .B2(n_682), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_500), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_496), .Y(n_493) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g690 ( .A(n_498), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_504), .Y(n_500) );
BUFx2_ASAP7_75t_L g917 ( .A(n_503), .Y(n_917) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OAI221xp5_ASAP7_75t_SL g746 ( .A1(n_506), .A2(n_729), .B1(n_747), .B2(n_748), .C(n_749), .Y(n_746) );
INVx3_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B1(n_639), .B2(n_733), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OAI22xp5_ASAP7_75t_SL g515 ( .A1(n_516), .A2(n_517), .B1(n_579), .B2(n_580), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
OAI22xp5_ASAP7_75t_SL g518 ( .A1(n_519), .A2(n_520), .B1(n_556), .B2(n_557), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g555 ( .A(n_521), .Y(n_555) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_539), .Y(n_521) );
NOR3xp33_ASAP7_75t_L g522 ( .A(n_523), .B(n_528), .C(n_534), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_526), .A2(n_672), .B1(n_673), .B2(n_674), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_526), .A2(n_753), .B1(n_754), .B2(n_756), .Y(n_752) );
OAI22xp5_ASAP7_75t_L g900 ( .A1(n_526), .A2(n_901), .B1(n_902), .B2(n_903), .Y(n_900) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
OAI22xp33_ASAP7_75t_L g710 ( .A1(n_530), .A2(n_711), .B1(n_712), .B2(n_713), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_531), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_536), .A2(n_802), .B1(n_803), .B2(n_804), .Y(n_801) );
INVx3_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g765 ( .A(n_537), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_540), .B(n_546), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
INVx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
INVx4_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g828 ( .A1(n_550), .A2(n_829), .B1(n_830), .B2(n_831), .Y(n_828) );
INVx4_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
XNOR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
NOR4xp75_ASAP7_75t_L g559 ( .A(n_560), .B(n_564), .C(n_568), .D(n_573), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_561), .B(n_563), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_565), .B(n_567), .Y(n_564) );
INVx1_ASAP7_75t_SL g846 ( .A(n_572), .Y(n_846) );
OAI21xp5_ASAP7_75t_SL g573 ( .A1(n_574), .A2(n_576), .B(n_577), .Y(n_573) );
OAI21xp33_ASAP7_75t_L g707 ( .A1(n_574), .A2(n_708), .B(n_709), .Y(n_707) );
OAI21xp5_ASAP7_75t_SL g872 ( .A1(n_574), .A2(n_873), .B(n_874), .Y(n_872) );
INVx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
BUFx4f_ASAP7_75t_SL g788 ( .A(n_578), .Y(n_788) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_613), .B1(n_637), .B2(n_638), .Y(n_580) );
INVx1_ASAP7_75t_L g637 ( .A(n_581), .Y(n_637) );
INVx1_ASAP7_75t_SL g612 ( .A(n_583), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_601), .Y(n_583) );
NOR2x1_ASAP7_75t_L g584 ( .A(n_585), .B(n_593), .Y(n_584) );
OAI222xp33_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_588), .B1(n_589), .B2(n_590), .C1(n_591), .C2(n_592), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
BUFx2_ASAP7_75t_L g679 ( .A(n_587), .Y(n_679) );
INVx4_ASAP7_75t_L g840 ( .A(n_587), .Y(n_840) );
OAI222xp33_ASAP7_75t_L g757 ( .A1(n_589), .A2(n_758), .B1(n_759), .B2(n_760), .C1(n_761), .C2(n_762), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_SL g877 ( .A(n_600), .Y(n_877) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_602), .B(n_608), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_606), .Y(n_602) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OAI221xp5_ASAP7_75t_SL g739 ( .A1(n_605), .A2(n_740), .B1(n_741), .B2(n_743), .C(n_744), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .Y(n_608) );
INVx1_ASAP7_75t_L g830 ( .A(n_610), .Y(n_830) );
INVx3_ASAP7_75t_L g638 ( .A(n_613), .Y(n_638) );
XOR2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_636), .Y(n_613) );
NAND2x1_ASAP7_75t_SL g614 ( .A(n_615), .B(n_627), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_616), .B(n_620), .Y(n_615) );
OAI21xp5_ASAP7_75t_SL g616 ( .A1(n_617), .A2(n_618), .B(n_619), .Y(n_616) );
OAI21xp5_ASAP7_75t_SL g836 ( .A1(n_617), .A2(n_837), .B(n_838), .Y(n_836) );
NAND3xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .C(n_625), .Y(n_620) );
NOR2x1_ASAP7_75t_L g627 ( .A(n_628), .B(n_632), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g733 ( .A(n_639), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_641), .B1(n_666), .B2(n_732), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g665 ( .A(n_645), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_658), .Y(n_645) );
NOR3xp33_ASAP7_75t_L g646 ( .A(n_647), .B(n_651), .C(n_655), .Y(n_646) );
OA211x2_ASAP7_75t_L g780 ( .A1(n_650), .A2(n_781), .B(n_782), .C(n_783), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_659), .B(n_662), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx1_ASAP7_75t_L g732 ( .A(n_666), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .B1(n_697), .B2(n_698), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
XOR2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_696), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_683), .Y(n_669) );
NOR3xp33_ASAP7_75t_L g670 ( .A(n_671), .B(n_675), .C(n_680), .Y(n_670) );
OAI21xp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_677), .B(n_678), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_692), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_688), .Y(n_684) );
INVx1_ASAP7_75t_L g721 ( .A(n_686), .Y(n_721) );
INVx1_ASAP7_75t_SL g723 ( .A(n_687), .Y(n_723) );
INVx3_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_693), .B(n_695), .Y(n_692) );
INVx1_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_714), .Y(n_702) );
NOR3xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_707), .C(n_710), .Y(n_703) );
NOR3xp33_ASAP7_75t_L g714 ( .A(n_715), .B(n_719), .C(n_724), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_718), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_721), .B1(n_722), .B2(n_723), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_727), .B1(n_728), .B2(n_729), .Y(n_724) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g852 ( .A(n_734), .Y(n_852) );
AOI22xp5_ASAP7_75t_SL g734 ( .A1(n_735), .A2(n_819), .B1(n_849), .B2(n_850), .Y(n_734) );
INVx1_ASAP7_75t_L g849 ( .A(n_735), .Y(n_849) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_769), .B1(n_770), .B2(n_818), .Y(n_735) );
INVx2_ASAP7_75t_L g818 ( .A(n_736), .Y(n_818) );
INVx1_ASAP7_75t_SL g768 ( .A(n_737), .Y(n_768) );
AND2x2_ASAP7_75t_SL g737 ( .A(n_738), .B(n_751), .Y(n_737) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_746), .Y(n_738) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NOR3xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_757), .C(n_763), .Y(n_751) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
OAI221xp5_ASAP7_75t_L g904 ( .A1(n_761), .A2(n_797), .B1(n_905), .B2(n_906), .C(n_907), .Y(n_904) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
OAI22xp5_ASAP7_75t_SL g770 ( .A1(n_771), .A2(n_772), .B1(n_790), .B2(n_817), .Y(n_770) );
INVx1_ASAP7_75t_SL g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
XOR2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_789), .Y(n_774) );
NAND4xp75_ASAP7_75t_L g775 ( .A(n_776), .B(n_780), .C(n_784), .D(n_787), .Y(n_775) );
AND2x2_ASAP7_75t_L g776 ( .A(n_777), .B(n_779), .Y(n_776) );
AND2x2_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .Y(n_784) );
INVx1_ASAP7_75t_L g817 ( .A(n_790), .Y(n_817) );
INVx2_ASAP7_75t_L g816 ( .A(n_791), .Y(n_816) );
AND2x2_ASAP7_75t_SL g791 ( .A(n_792), .B(n_805), .Y(n_791) );
NOR3xp33_ASAP7_75t_L g792 ( .A(n_793), .B(n_796), .C(n_801), .Y(n_792) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_806), .B(n_809), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_810), .B(n_814), .Y(n_809) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx2_ASAP7_75t_L g850 ( .A(n_819), .Y(n_850) );
NAND2xp5_ASAP7_75t_SL g820 ( .A(n_821), .B(n_835), .Y(n_820) );
NOR3xp33_ASAP7_75t_L g821 ( .A(n_822), .B(n_828), .C(n_832), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_823), .B(n_826), .Y(n_822) );
NOR2xp33_ASAP7_75t_L g835 ( .A(n_836), .B(n_841), .Y(n_835) );
INVx3_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_842), .B(n_847), .Y(n_841) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_SL g853 ( .A(n_854), .Y(n_853) );
NOR2x1_ASAP7_75t_L g854 ( .A(n_855), .B(n_859), .Y(n_854) );
OR2x2_ASAP7_75t_SL g923 ( .A(n_855), .B(n_860), .Y(n_923) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_856), .B(n_858), .Y(n_855) );
CKINVDCx20_ASAP7_75t_R g889 ( .A(n_856), .Y(n_889) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_857), .B(n_891), .Y(n_894) );
CKINVDCx16_ASAP7_75t_R g891 ( .A(n_858), .Y(n_891) );
CKINVDCx20_ASAP7_75t_R g859 ( .A(n_860), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_861), .B(n_862), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_864), .B(n_865), .Y(n_863) );
OAI322xp33_ASAP7_75t_L g866 ( .A1(n_867), .A2(n_887), .A3(n_890), .B1(n_892), .B2(n_895), .C1(n_896), .C2(n_921), .Y(n_866) );
HB1xp67_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_871), .B(n_880), .Y(n_870) );
NOR2xp67_ASAP7_75t_L g871 ( .A(n_872), .B(n_875), .Y(n_871) );
NAND3xp33_ASAP7_75t_L g875 ( .A(n_876), .B(n_878), .C(n_879), .Y(n_875) );
NOR2x1_ASAP7_75t_L g880 ( .A(n_881), .B(n_884), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_882), .B(n_883), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_885), .B(n_886), .Y(n_884) );
HB1xp67_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
HB1xp67_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
CKINVDCx20_ASAP7_75t_R g892 ( .A(n_893), .Y(n_892) );
INVx2_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_899), .B(n_911), .Y(n_898) );
NOR3xp33_ASAP7_75t_L g899 ( .A(n_900), .B(n_904), .C(n_908), .Y(n_899) );
NOR2xp33_ASAP7_75t_L g911 ( .A(n_912), .B(n_915), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_913), .B(n_914), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_916), .B(n_918), .Y(n_915) );
BUFx4f_ASAP7_75t_SL g919 ( .A(n_920), .Y(n_919) );
CKINVDCx20_ASAP7_75t_R g921 ( .A(n_922), .Y(n_921) );
CKINVDCx20_ASAP7_75t_R g922 ( .A(n_923), .Y(n_922) );
endmodule