module fake_netlist_5_390_n_772 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_772);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_772;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_146;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_452;
wire n_525;
wire n_493;
wire n_397;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_155;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_443;
wire n_372;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_433;
wire n_604;
wire n_368;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_147;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_150;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_579;
wire n_250;
wire n_394;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_428;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_185;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_169;
wire n_550;
wire n_522;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_344;
wire n_287;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_145;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_432;
wire n_164;
wire n_553;
wire n_395;
wire n_727;
wire n_311;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_144;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_517;
wire n_482;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_571;
wire n_461;
wire n_333;
wire n_477;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_151;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_730;
wire n_729;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_647;
wire n_480;
wire n_607;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_707;
wire n_710;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_453;
wire n_403;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_148;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_766;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_162;
wire n_759;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_64),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_139),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_89),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_26),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_86),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_22),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_75),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_115),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_36),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_76),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_88),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_16),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_17),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_90),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_35),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_126),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_43),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_104),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_74),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_98),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_72),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_124),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_11),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_133),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_13),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_11),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_21),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_62),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_130),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_0),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_23),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_4),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_15),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_138),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_23),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_83),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_3),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_100),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_109),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_131),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_97),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_46),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_95),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_65),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_116),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_27),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_154),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_0),
.Y(n_199)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_160),
.Y(n_201)
);

AND2x4_ASAP7_75t_L g202 ( 
.A(n_154),
.B(n_25),
.Y(n_202)
);

AND2x4_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_28),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_191),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_145),
.Y(n_206)
);

AND2x4_ASAP7_75t_L g207 ( 
.A(n_148),
.B(n_29),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_149),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_183),
.B(n_1),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_150),
.Y(n_210)
);

AND2x4_ASAP7_75t_L g211 ( 
.A(n_153),
.B(n_30),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_155),
.Y(n_213)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_170),
.B(n_1),
.Y(n_215)
);

AND2x4_ASAP7_75t_L g216 ( 
.A(n_171),
.B(n_31),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_159),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g219 ( 
.A(n_152),
.Y(n_219)
);

AND2x6_ASAP7_75t_L g220 ( 
.A(n_178),
.B(n_180),
.Y(n_220)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_157),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_172),
.B(n_2),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_2),
.Y(n_223)
);

AND2x4_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_32),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_175),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_158),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_164),
.B(n_3),
.Y(n_230)
);

BUFx8_ASAP7_75t_SL g231 ( 
.A(n_152),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_144),
.B(n_4),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_182),
.B(n_5),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_161),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g235 ( 
.A(n_182),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_144),
.B(n_5),
.Y(n_236)
);

AND2x2_ASAP7_75t_SL g237 ( 
.A(n_209),
.B(n_166),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_162),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_198),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_146),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_198),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_198),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_204),
.B(n_146),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_147),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_230),
.A2(n_196),
.B1(n_193),
.B2(n_179),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_199),
.A2(n_174),
.B1(n_176),
.B2(n_181),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_198),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_222),
.A2(n_185),
.B1(n_187),
.B2(n_189),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_217),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_201),
.B(n_147),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_219),
.A2(n_185),
.B1(n_187),
.B2(n_189),
.Y(n_252)
);

NAND3x1_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_6),
.C(n_7),
.Y(n_253)
);

AND2x2_ASAP7_75t_SL g254 ( 
.A(n_203),
.B(n_151),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_197),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_151),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_231),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_184),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_219),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_202),
.A2(n_195),
.B1(n_184),
.B2(n_173),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_235),
.A2(n_195),
.B1(n_169),
.B2(n_168),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_L g262 ( 
.A1(n_215),
.A2(n_163),
.B1(n_7),
.B2(n_8),
.Y(n_262)
);

BUFx6f_ASAP7_75t_SL g263 ( 
.A(n_202),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_33),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_232),
.Y(n_265)
);

AND2x4_ASAP7_75t_L g266 ( 
.A(n_202),
.B(n_34),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_235),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_223),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_198),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_233),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_270)
);

AO22x2_ASAP7_75t_L g271 ( 
.A1(n_203),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_236),
.A2(n_14),
.B1(n_17),
.B2(n_18),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_203),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_205),
.Y(n_274)
);

AO22x2_ASAP7_75t_L g275 ( 
.A1(n_207),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_207),
.A2(n_22),
.B1(n_24),
.B2(n_37),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_L g277 ( 
.A1(n_208),
.A2(n_24),
.B1(n_38),
.B2(n_39),
.Y(n_277)
);

OAI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_207),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_L g279 ( 
.A1(n_218),
.A2(n_227),
.B1(n_210),
.B2(n_200),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_234),
.B(n_44),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_L g281 ( 
.A1(n_218),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_281)
);

AO22x2_ASAP7_75t_L g282 ( 
.A1(n_211),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_211),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_239),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_242),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_247),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_238),
.B(n_234),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_243),
.B(n_234),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_241),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_241),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_245),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_241),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_274),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_256),
.B(n_234),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_274),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_251),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_240),
.B(n_254),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_266),
.B(n_211),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_258),
.B(n_200),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_257),
.B(n_216),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_251),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_255),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_252),
.Y(n_304)
);

XOR2x2_ASAP7_75t_L g305 ( 
.A(n_253),
.B(n_231),
.Y(n_305)
);

NAND2x1p5_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_216),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_255),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_266),
.Y(n_308)
);

AND2x4_ASAP7_75t_L g309 ( 
.A(n_283),
.B(n_216),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_250),
.B(n_244),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_249),
.B(n_200),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_264),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_279),
.A2(n_224),
.B(n_200),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_263),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_261),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_265),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_263),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_276),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_280),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_265),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_282),
.Y(n_321)
);

AND2x2_ASAP7_75t_SL g322 ( 
.A(n_237),
.B(n_224),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_260),
.B(n_200),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_282),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_278),
.B(n_224),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_271),
.Y(n_326)
);

INVxp33_ASAP7_75t_L g327 ( 
.A(n_271),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_275),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_275),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_281),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_273),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_277),
.Y(n_332)
);

INVxp33_ASAP7_75t_L g333 ( 
.A(n_270),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_259),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_246),
.B(n_213),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_267),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_270),
.B(n_218),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_268),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_248),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_272),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_262),
.B(n_213),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_272),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_239),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_239),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_238),
.B(n_213),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_239),
.Y(n_346)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_319),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_294),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_308),
.B(n_310),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_289),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_299),
.B(n_220),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_284),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_295),
.B(n_227),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_298),
.B(n_227),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_316),
.Y(n_355)
);

AND2x2_ASAP7_75t_SL g356 ( 
.A(n_322),
.B(n_206),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_299),
.B(n_220),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_309),
.A2(n_220),
.B1(n_210),
.B2(n_206),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_296),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_325),
.A2(n_337),
.B(n_309),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_297),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_298),
.B(n_205),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_306),
.Y(n_363)
);

AND2x4_ASAP7_75t_L g364 ( 
.A(n_309),
.B(n_55),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_302),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_322),
.B(n_205),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_285),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_286),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_341),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_301),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_306),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_319),
.B(n_220),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_303),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_312),
.B(n_210),
.Y(n_374)
);

INVx2_ASAP7_75t_SL g375 ( 
.A(n_329),
.Y(n_375)
);

BUFx4f_ASAP7_75t_L g376 ( 
.A(n_319),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_288),
.Y(n_377)
);

AND2x4_ASAP7_75t_L g378 ( 
.A(n_331),
.B(n_56),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_319),
.B(n_220),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_339),
.Y(n_380)
);

AND2x2_ASAP7_75t_SL g381 ( 
.A(n_330),
.B(n_206),
.Y(n_381)
);

OAI21x1_ASAP7_75t_L g382 ( 
.A1(n_313),
.A2(n_220),
.B(n_226),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_338),
.B(n_210),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_307),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_318),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_316),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_343),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_325),
.A2(n_221),
.B(n_214),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_344),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_329),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_346),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_335),
.B(n_57),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_328),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_290),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_291),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_293),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_287),
.B(n_206),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_287),
.B(n_206),
.Y(n_398)
);

AND2x2_ASAP7_75t_SL g399 ( 
.A(n_321),
.B(n_212),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_300),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_314),
.Y(n_401)
);

BUFx12f_ASAP7_75t_SL g402 ( 
.A(n_311),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_328),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_326),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_332),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_342),
.B(n_212),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_334),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_324),
.B(n_58),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_324),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_336),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_317),
.B(n_59),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_327),
.B(n_212),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_345),
.B(n_323),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_345),
.B(n_212),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_410),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_355),
.B(n_320),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_363),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_364),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_362),
.B(n_323),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_363),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_362),
.B(n_327),
.Y(n_421)
);

INVx5_ASAP7_75t_L g422 ( 
.A(n_347),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_390),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_408),
.Y(n_424)
);

AND2x6_ASAP7_75t_L g425 ( 
.A(n_364),
.B(n_333),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_350),
.B(n_333),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_349),
.B(n_334),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_354),
.B(n_213),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_356),
.B(n_292),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_403),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_385),
.B(n_369),
.Y(n_431)
);

INVx6_ASAP7_75t_L g432 ( 
.A(n_364),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_363),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_361),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_361),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_361),
.Y(n_436)
);

INVxp67_ASAP7_75t_SL g437 ( 
.A(n_371),
.Y(n_437)
);

NAND2x1_ASAP7_75t_L g438 ( 
.A(n_347),
.B(n_212),
.Y(n_438)
);

INVx4_ASAP7_75t_L g439 ( 
.A(n_371),
.Y(n_439)
);

AND2x6_ASAP7_75t_L g440 ( 
.A(n_364),
.B(n_226),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_403),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_403),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_354),
.B(n_353),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_371),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_411),
.B(n_349),
.Y(n_445)
);

OR2x6_ASAP7_75t_L g446 ( 
.A(n_408),
.B(n_305),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_376),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_353),
.B(n_347),
.Y(n_448)
);

CKINVDCx6p67_ASAP7_75t_R g449 ( 
.A(n_407),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_412),
.B(n_292),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_347),
.B(n_213),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_401),
.Y(n_452)
);

AND2x6_ASAP7_75t_L g453 ( 
.A(n_378),
.B(n_226),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_412),
.B(n_340),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_365),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_380),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_365),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_408),
.B(n_315),
.Y(n_458)
);

OR2x6_ASAP7_75t_L g459 ( 
.A(n_408),
.B(n_305),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_411),
.B(n_315),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_365),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_348),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_389),
.Y(n_463)
);

OR2x6_ASAP7_75t_L g464 ( 
.A(n_360),
.B(n_340),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_389),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_406),
.B(n_214),
.Y(n_466)
);

AND2x4_ASAP7_75t_SL g467 ( 
.A(n_378),
.B(n_304),
.Y(n_467)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_409),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_406),
.B(n_214),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_389),
.Y(n_470)
);

NAND2x1p5_ASAP7_75t_L g471 ( 
.A(n_422),
.B(n_376),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_424),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_L g473 ( 
.A1(n_464),
.A2(n_356),
.B1(n_405),
.B2(n_381),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_449),
.Y(n_474)
);

INVx6_ASAP7_75t_L g475 ( 
.A(n_417),
.Y(n_475)
);

BUFx4f_ASAP7_75t_SL g476 ( 
.A(n_415),
.Y(n_476)
);

NAND2x1p5_ASAP7_75t_L g477 ( 
.A(n_422),
.B(n_376),
.Y(n_477)
);

INVx4_ASAP7_75t_L g478 ( 
.A(n_422),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_434),
.Y(n_479)
);

CKINVDCx11_ASAP7_75t_R g480 ( 
.A(n_446),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_452),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_417),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_430),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_454),
.Y(n_484)
);

BUFx12f_ASAP7_75t_L g485 ( 
.A(n_460),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_441),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_425),
.A2(n_356),
.B1(n_366),
.B2(n_413),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_468),
.Y(n_488)
);

INVx2_ASAP7_75t_SL g489 ( 
.A(n_417),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_467),
.Y(n_490)
);

INVx4_ASAP7_75t_L g491 ( 
.A(n_422),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_468),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_417),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_434),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_420),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_435),
.Y(n_496)
);

BUFx12f_ASAP7_75t_L g497 ( 
.A(n_460),
.Y(n_497)
);

NAND2x1p5_ASAP7_75t_L g498 ( 
.A(n_418),
.B(n_376),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_426),
.B(n_407),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_467),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_420),
.Y(n_501)
);

BUFx2_ASAP7_75t_SL g502 ( 
.A(n_452),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g503 ( 
.A(n_450),
.Y(n_503)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_427),
.Y(n_504)
);

INVx5_ASAP7_75t_L g505 ( 
.A(n_425),
.Y(n_505)
);

BUFx5_ASAP7_75t_L g506 ( 
.A(n_425),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_420),
.Y(n_507)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_420),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_458),
.Y(n_509)
);

BUFx4_ASAP7_75t_SL g510 ( 
.A(n_446),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_442),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_433),
.Y(n_512)
);

NAND2x1_ASAP7_75t_L g513 ( 
.A(n_432),
.B(n_352),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_435),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_425),
.A2(n_366),
.B1(n_413),
.B2(n_369),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_433),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_433),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_458),
.Y(n_518)
);

OR2x2_ASAP7_75t_L g519 ( 
.A(n_421),
.B(n_370),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_484),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_476),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_479),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_478),
.A2(n_443),
.B(n_448),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_499),
.A2(n_464),
.B1(n_429),
.B2(n_460),
.Y(n_524)
);

CKINVDCx6p67_ASAP7_75t_R g525 ( 
.A(n_485),
.Y(n_525)
);

OAI22xp33_ASAP7_75t_L g526 ( 
.A1(n_503),
.A2(n_464),
.B1(n_416),
.B2(n_446),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_476),
.Y(n_527)
);

OAI22xp33_ASAP7_75t_L g528 ( 
.A1(n_504),
.A2(n_459),
.B1(n_456),
.B2(n_304),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_481),
.Y(n_529)
);

INVx8_ASAP7_75t_L g530 ( 
.A(n_493),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_479),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_519),
.A2(n_429),
.B1(n_425),
.B2(n_445),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_493),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_509),
.A2(n_445),
.B1(n_458),
.B2(n_392),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_494),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_473),
.A2(n_437),
.B1(n_432),
.B2(n_418),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_518),
.A2(n_386),
.B(n_431),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_473),
.B(n_360),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_SL g539 ( 
.A1(n_485),
.A2(n_459),
.B1(n_431),
.B2(n_378),
.Y(n_539)
);

INVx1_ASAP7_75t_SL g540 ( 
.A(n_474),
.Y(n_540)
);

INVx6_ASAP7_75t_L g541 ( 
.A(n_508),
.Y(n_541)
);

BUFx2_ASAP7_75t_SL g542 ( 
.A(n_481),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_494),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_517),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_496),
.Y(n_545)
);

BUFx8_ASAP7_75t_L g546 ( 
.A(n_497),
.Y(n_546)
);

INVx6_ASAP7_75t_L g547 ( 
.A(n_508),
.Y(n_547)
);

NAND2x1p5_ASAP7_75t_L g548 ( 
.A(n_478),
.B(n_439),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_483),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_515),
.A2(n_432),
.B1(n_419),
.B2(n_497),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_472),
.A2(n_392),
.B1(n_459),
.B2(n_405),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_486),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_487),
.B(n_405),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_472),
.A2(n_392),
.B1(n_378),
.B2(n_456),
.Y(n_554)
);

BUFx2_ASAP7_75t_SL g555 ( 
.A(n_507),
.Y(n_555)
);

OAI22xp33_ASAP7_75t_L g556 ( 
.A1(n_490),
.A2(n_462),
.B1(n_437),
.B2(n_401),
.Y(n_556)
);

BUFx12f_ASAP7_75t_L g557 ( 
.A(n_480),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_517),
.Y(n_558)
);

BUFx12f_ASAP7_75t_L g559 ( 
.A(n_480),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_493),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_SL g561 ( 
.A1(n_490),
.A2(n_381),
.B1(n_392),
.B2(n_453),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_502),
.A2(n_411),
.B1(n_400),
.B2(n_402),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_511),
.B(n_455),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_538),
.A2(n_381),
.B1(n_383),
.B2(n_384),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_538),
.A2(n_383),
.B1(n_384),
.B2(n_373),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_526),
.A2(n_500),
.B1(n_411),
.B2(n_401),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_520),
.Y(n_567)
);

OAI21xp33_ASAP7_75t_L g568 ( 
.A1(n_537),
.A2(n_373),
.B(n_359),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_539),
.A2(n_348),
.B1(n_359),
.B2(n_453),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_549),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_524),
.B(n_423),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_520),
.B(n_393),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_552),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_557),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_557),
.Y(n_575)
);

OR2x2_ASAP7_75t_SL g576 ( 
.A(n_559),
.B(n_510),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_SL g577 ( 
.A1(n_559),
.A2(n_453),
.B1(n_505),
.B2(n_500),
.Y(n_577)
);

OAI22xp33_ASAP7_75t_L g578 ( 
.A1(n_550),
.A2(n_505),
.B1(n_439),
.B2(n_457),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_553),
.A2(n_528),
.B1(n_551),
.B2(n_532),
.Y(n_579)
);

BUFx6f_ASAP7_75t_SL g580 ( 
.A(n_521),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_563),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_553),
.B(n_393),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_554),
.A2(n_400),
.B1(n_453),
.B2(n_374),
.Y(n_583)
);

AO22x1_ASAP7_75t_L g584 ( 
.A1(n_546),
.A2(n_453),
.B1(n_507),
.B2(n_505),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_534),
.A2(n_400),
.B1(n_374),
.B2(n_440),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_529),
.B(n_404),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_SL g587 ( 
.A1(n_561),
.A2(n_388),
.B(n_358),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_563),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_SL g589 ( 
.A1(n_546),
.A2(n_505),
.B1(n_506),
.B2(n_440),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_L g590 ( 
.A1(n_523),
.A2(n_428),
.B(n_466),
.Y(n_590)
);

AOI222xp33_ASAP7_75t_L g591 ( 
.A1(n_546),
.A2(n_404),
.B1(n_399),
.B2(n_388),
.C1(n_440),
.C2(n_391),
.Y(n_591)
);

OAI222xp33_ASAP7_75t_L g592 ( 
.A1(n_562),
.A2(n_498),
.B1(n_358),
.B2(n_513),
.C1(n_447),
.C2(n_436),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_525),
.A2(n_440),
.B1(n_399),
.B2(n_391),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_536),
.A2(n_447),
.B1(n_444),
.B2(n_433),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_530),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_529),
.B(n_399),
.Y(n_596)
);

OAI22xp33_ASAP7_75t_L g597 ( 
.A1(n_525),
.A2(n_444),
.B1(n_436),
.B2(n_461),
.Y(n_597)
);

INVx1_ASAP7_75t_SL g598 ( 
.A(n_540),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_542),
.B(n_501),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_556),
.A2(n_444),
.B1(n_498),
.B2(n_409),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_522),
.Y(n_601)
);

OAI21xp5_ASAP7_75t_SL g602 ( 
.A1(n_527),
.A2(n_409),
.B(n_469),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_SL g603 ( 
.A1(n_527),
.A2(n_506),
.B1(n_440),
.B2(n_444),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_530),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_522),
.A2(n_461),
.B1(n_470),
.B2(n_463),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_SL g606 ( 
.A1(n_548),
.A2(n_409),
.B(n_471),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_530),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_L g608 ( 
.A1(n_521),
.A2(n_475),
.B1(n_488),
.B2(n_492),
.Y(n_608)
);

OAI22xp33_ASAP7_75t_L g609 ( 
.A1(n_531),
.A2(n_470),
.B1(n_463),
.B2(n_465),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_555),
.B(n_501),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_531),
.A2(n_465),
.B1(n_514),
.B2(n_496),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_541),
.A2(n_506),
.B1(n_395),
.B2(n_402),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_598),
.B(n_402),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_566),
.A2(n_506),
.B1(n_541),
.B2(n_547),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_579),
.A2(n_569),
.B1(n_593),
.B2(n_565),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_568),
.A2(n_506),
.B1(n_395),
.B2(n_547),
.Y(n_616)
);

NOR3xp33_ASAP7_75t_L g617 ( 
.A(n_602),
.B(n_508),
.C(n_397),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_571),
.A2(n_506),
.B1(n_547),
.B2(n_541),
.Y(n_618)
);

AND2x2_ASAP7_75t_SL g619 ( 
.A(n_569),
.B(n_493),
.Y(n_619)
);

AOI221x1_ASAP7_75t_L g620 ( 
.A1(n_594),
.A2(n_414),
.B1(n_398),
.B2(n_397),
.C(n_533),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_SL g621 ( 
.A1(n_580),
.A2(n_541),
.B1(n_547),
.B2(n_548),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_SL g622 ( 
.A1(n_580),
.A2(n_471),
.B1(n_477),
.B2(n_530),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_581),
.B(n_535),
.Y(n_623)
);

OAI222xp33_ASAP7_75t_L g624 ( 
.A1(n_582),
.A2(n_545),
.B1(n_543),
.B2(n_535),
.C1(n_560),
.C2(n_533),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_591),
.A2(n_475),
.B1(n_394),
.B2(n_396),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_578),
.A2(n_475),
.B1(n_394),
.B2(n_396),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_572),
.B(n_543),
.Y(n_627)
);

OAI22xp33_ASAP7_75t_L g628 ( 
.A1(n_587),
.A2(n_545),
.B1(n_477),
.B2(n_492),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_SL g629 ( 
.A1(n_596),
.A2(n_488),
.B1(n_495),
.B2(n_517),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_SL g630 ( 
.A1(n_600),
.A2(n_516),
.B1(n_495),
.B2(n_517),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_578),
.A2(n_396),
.B1(n_394),
.B2(n_367),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_SL g632 ( 
.A1(n_567),
.A2(n_495),
.B1(n_516),
.B2(n_489),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_574),
.A2(n_482),
.B1(n_489),
.B2(n_512),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_585),
.A2(n_387),
.B1(n_352),
.B2(n_367),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g635 ( 
.A1(n_565),
.A2(n_482),
.B1(n_512),
.B2(n_491),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_564),
.A2(n_514),
.B1(n_228),
.B2(n_226),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_588),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_SL g638 ( 
.A1(n_588),
.A2(n_495),
.B1(n_516),
.B2(n_560),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_SL g639 ( 
.A1(n_570),
.A2(n_516),
.B1(n_533),
.B2(n_560),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_564),
.A2(n_226),
.B1(n_228),
.B2(n_398),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_SL g641 ( 
.A1(n_573),
.A2(n_558),
.B1(n_544),
.B2(n_491),
.Y(n_641)
);

NAND3xp33_ASAP7_75t_SL g642 ( 
.A(n_575),
.B(n_414),
.C(n_438),
.Y(n_642)
);

OA211x2_ASAP7_75t_L g643 ( 
.A1(n_590),
.A2(n_451),
.B(n_379),
.C(n_372),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g644 ( 
.A1(n_612),
.A2(n_583),
.B1(n_577),
.B2(n_576),
.Y(n_644)
);

NAND3xp33_ASAP7_75t_L g645 ( 
.A(n_586),
.B(n_608),
.C(n_603),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_601),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_599),
.B(n_544),
.Y(n_647)
);

OAI211xp5_ASAP7_75t_L g648 ( 
.A1(n_606),
.A2(n_375),
.B(n_228),
.C(n_351),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_637),
.Y(n_649)
);

NAND3xp33_ASAP7_75t_L g650 ( 
.A(n_615),
.B(n_610),
.C(n_589),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_L g651 ( 
.A1(n_642),
.A2(n_597),
.B(n_592),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_627),
.B(n_611),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_623),
.B(n_611),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_619),
.B(n_597),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_646),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_647),
.B(n_618),
.Y(n_656)
);

OAI221xp5_ASAP7_75t_SL g657 ( 
.A1(n_616),
.A2(n_605),
.B1(n_609),
.B2(n_351),
.C(n_357),
.Y(n_657)
);

AOI221xp5_ASAP7_75t_L g658 ( 
.A1(n_644),
.A2(n_228),
.B1(n_584),
.B2(n_609),
.C(n_387),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_624),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_619),
.B(n_605),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_628),
.B(n_614),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_613),
.B(n_544),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_628),
.B(n_544),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_L g664 ( 
.A1(n_645),
.A2(n_633),
.B1(n_640),
.B2(n_625),
.Y(n_664)
);

OAI21xp33_ASAP7_75t_L g665 ( 
.A1(n_640),
.A2(n_228),
.B(n_595),
.Y(n_665)
);

NAND4xp25_ASAP7_75t_L g666 ( 
.A(n_643),
.B(n_607),
.C(n_377),
.D(n_352),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_R g667 ( 
.A(n_636),
.B(n_595),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_621),
.B(n_607),
.Y(n_668)
);

NAND3xp33_ASAP7_75t_L g669 ( 
.A(n_617),
.B(n_604),
.C(n_595),
.Y(n_669)
);

NAND3xp33_ASAP7_75t_L g670 ( 
.A(n_620),
.B(n_639),
.C(n_638),
.Y(n_670)
);

NAND3xp33_ASAP7_75t_L g671 ( 
.A(n_641),
.B(n_604),
.C(n_595),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_629),
.B(n_558),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_636),
.B(n_632),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_648),
.B(n_622),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_630),
.B(n_558),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_631),
.B(n_558),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_649),
.B(n_635),
.Y(n_677)
);

NAND3xp33_ASAP7_75t_L g678 ( 
.A(n_650),
.B(n_626),
.C(n_634),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_655),
.B(n_656),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_659),
.Y(n_680)
);

NAND4xp75_ASAP7_75t_L g681 ( 
.A(n_674),
.B(n_604),
.C(n_379),
.D(n_372),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_661),
.B(n_604),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_662),
.B(n_60),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_672),
.B(n_61),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_668),
.B(n_63),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_668),
.B(n_66),
.Y(n_686)
);

OAI211xp5_ASAP7_75t_SL g687 ( 
.A1(n_651),
.A2(n_387),
.B(n_377),
.C(n_368),
.Y(n_687)
);

NAND3xp33_ASAP7_75t_L g688 ( 
.A(n_669),
.B(n_368),
.C(n_352),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_664),
.A2(n_387),
.B1(n_367),
.B2(n_377),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_652),
.B(n_367),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_653),
.B(n_654),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_663),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_660),
.B(n_368),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_679),
.B(n_672),
.Y(n_694)
);

NAND3xp33_ASAP7_75t_L g695 ( 
.A(n_691),
.B(n_674),
.C(n_670),
.Y(n_695)
);

OAI22xp33_ASAP7_75t_L g696 ( 
.A1(n_689),
.A2(n_654),
.B1(n_673),
.B2(n_671),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_692),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_680),
.Y(n_698)
);

NOR4xp25_ASAP7_75t_L g699 ( 
.A(n_678),
.B(n_665),
.C(n_658),
.D(n_657),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_677),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_690),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_682),
.B(n_666),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_684),
.B(n_675),
.Y(n_703)
);

XOR2x2_ASAP7_75t_L g704 ( 
.A(n_685),
.B(n_676),
.Y(n_704)
);

XOR2x2_ASAP7_75t_L g705 ( 
.A(n_704),
.B(n_695),
.Y(n_705)
);

XOR2x2_ASAP7_75t_L g706 ( 
.A(n_704),
.B(n_686),
.Y(n_706)
);

XNOR2x1_ASAP7_75t_L g707 ( 
.A(n_698),
.B(n_683),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_696),
.B(n_693),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_700),
.B(n_689),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_709),
.Y(n_710)
);

XOR2x2_ASAP7_75t_L g711 ( 
.A(n_705),
.B(n_702),
.Y(n_711)
);

OA22x2_ASAP7_75t_L g712 ( 
.A1(n_708),
.A2(n_706),
.B1(n_703),
.B2(n_701),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_707),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_710),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_710),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_712),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_713),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_716),
.A2(n_696),
.B1(n_702),
.B2(n_711),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_714),
.Y(n_719)
);

AO22x2_ASAP7_75t_L g720 ( 
.A1(n_717),
.A2(n_715),
.B1(n_714),
.B2(n_697),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_719),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_720),
.Y(n_722)
);

HB1xp67_ASAP7_75t_L g723 ( 
.A(n_718),
.Y(n_723)
);

OAI22xp33_ASAP7_75t_L g724 ( 
.A1(n_718),
.A2(n_688),
.B1(n_699),
.B2(n_694),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_723),
.A2(n_681),
.B1(n_687),
.B2(n_676),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_724),
.B(n_667),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_721),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_722),
.A2(n_667),
.B1(n_491),
.B2(n_478),
.Y(n_728)
);

NOR2xp67_ASAP7_75t_L g729 ( 
.A(n_722),
.B(n_67),
.Y(n_729)
);

AO22x2_ASAP7_75t_L g730 ( 
.A1(n_722),
.A2(n_375),
.B1(n_377),
.B2(n_368),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_723),
.A2(n_382),
.B1(n_221),
.B2(n_214),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_726),
.A2(n_382),
.B1(n_221),
.B2(n_214),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_729),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_727),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_730),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_725),
.A2(n_221),
.B1(n_69),
.B2(n_71),
.Y(n_736)
);

HB1xp67_ASAP7_75t_L g737 ( 
.A(n_728),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_731),
.Y(n_738)
);

AO22x2_ASAP7_75t_L g739 ( 
.A1(n_734),
.A2(n_68),
.B1(n_73),
.B2(n_77),
.Y(n_739)
);

AO22x2_ASAP7_75t_L g740 ( 
.A1(n_735),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_740)
);

AND4x1_ASAP7_75t_L g741 ( 
.A(n_736),
.B(n_81),
.C(n_82),
.D(n_84),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_733),
.A2(n_221),
.B1(n_87),
.B2(n_91),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_737),
.B(n_85),
.Y(n_743)
);

AND5x1_ASAP7_75t_L g744 ( 
.A(n_732),
.B(n_143),
.C(n_93),
.D(n_94),
.E(n_96),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_738),
.B(n_142),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_733),
.B(n_92),
.Y(n_746)
);

AO22x2_ASAP7_75t_L g747 ( 
.A1(n_734),
.A2(n_99),
.B1(n_102),
.B2(n_103),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_743),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_745),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_746),
.B(n_105),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_740),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_739),
.A2(n_106),
.B1(n_107),
.B2(n_111),
.Y(n_752)
);

INVx5_ASAP7_75t_L g753 ( 
.A(n_747),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_741),
.B(n_112),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_742),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_751),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_753),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_753),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_754),
.A2(n_744),
.B1(n_114),
.B2(n_117),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_752),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_755),
.A2(n_113),
.B1(n_118),
.B2(n_119),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_757),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_758),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_756),
.B(n_748),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_SL g765 ( 
.A1(n_762),
.A2(n_760),
.B1(n_749),
.B2(n_750),
.Y(n_765)
);

AOI31xp33_ASAP7_75t_L g766 ( 
.A1(n_763),
.A2(n_759),
.A3(n_761),
.B(n_123),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_764),
.A2(n_120),
.B1(n_121),
.B2(n_125),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_765),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_768),
.A2(n_767),
.B1(n_766),
.B2(n_129),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_769),
.Y(n_770)
);

AOI221x1_ASAP7_75t_L g771 ( 
.A1(n_770),
.A2(n_127),
.B1(n_128),
.B2(n_132),
.C(n_134),
.Y(n_771)
);

AOI211xp5_ASAP7_75t_L g772 ( 
.A1(n_771),
.A2(n_135),
.B(n_136),
.C(n_137),
.Y(n_772)
);


endmodule