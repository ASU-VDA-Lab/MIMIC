module real_jpeg_10318_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_301, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_301;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_249;
wire n_78;
wire n_166;
wire n_176;
wire n_286;
wire n_292;
wire n_221;
wire n_215;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_297;
wire n_240;
wire n_55;
wire n_125;
wire n_180;
wire n_58;
wire n_52;
wire n_209;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_295;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_1),
.A2(n_47),
.B(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_1),
.B(n_47),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_1),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_1),
.A2(n_74),
.B1(n_77),
.B2(n_151),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_1),
.A2(n_33),
.B(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_1),
.B(n_33),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_1),
.B(n_197),
.Y(n_196)
);

AOI21xp33_ASAP7_75t_L g216 ( 
.A1(n_1),
.A2(n_30),
.B(n_34),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_1),
.A2(n_27),
.B1(n_36),
.B2(n_153),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_2),
.A2(n_47),
.B1(n_48),
.B2(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_2),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_2),
.A2(n_59),
.B1(n_60),
.B2(n_142),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_142),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_2),
.A2(n_27),
.B1(n_36),
.B2(n_142),
.Y(n_238)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_4),
.A2(n_47),
.B1(n_48),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_4),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_4),
.A2(n_59),
.B1(n_60),
.B2(n_63),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_63),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_5),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_5),
.A2(n_27),
.B1(n_36),
.B2(n_51),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_5),
.A2(n_51),
.B1(n_59),
.B2(n_60),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_7),
.A2(n_27),
.B1(n_36),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_39),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_7),
.A2(n_39),
.B1(n_47),
.B2(n_48),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_7),
.A2(n_39),
.B1(n_59),
.B2(n_60),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_SL g56 ( 
.A1(n_8),
.A2(n_47),
.B(n_57),
.C(n_58),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_8),
.B(n_47),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_8),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_58)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

BUFx6f_ASAP7_75t_SL g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_53),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_11),
.A2(n_53),
.B1(n_59),
.B2(n_60),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_13),
.A2(n_59),
.B1(n_60),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_13),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_13),
.A2(n_47),
.B1(n_48),
.B2(n_133),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_133),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_13),
.A2(n_27),
.B1(n_36),
.B2(n_133),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_14),
.A2(n_27),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_14),
.A2(n_37),
.B1(n_59),
.B2(n_60),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_14),
.A2(n_37),
.B1(n_47),
.B2(n_48),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_16),
.A2(n_27),
.B1(n_36),
.B2(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_16),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_16),
.A2(n_59),
.B1(n_60),
.B2(n_117),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_16),
.A2(n_47),
.B1(n_48),
.B2(n_117),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_16),
.A2(n_33),
.B1(n_34),
.B2(n_117),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_17),
.A2(n_27),
.B1(n_36),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_17),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_17),
.A2(n_59),
.B1(n_60),
.B2(n_84),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_17),
.A2(n_47),
.B1(n_48),
.B2(n_84),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_17),
.A2(n_33),
.B1(n_34),
.B2(n_84),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_99),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_98),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_85),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_22),
.B(n_85),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_65),
.C(n_70),
.Y(n_22)
);

FAx1_ASAP7_75t_SL g121 ( 
.A(n_23),
.B(n_65),
.CI(n_70),
.CON(n_121),
.SN(n_121)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_40),
.B2(n_41),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_24),
.A2(n_25),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_25),
.B(n_54),
.C(n_64),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_32),
.B1(n_35),
.B2(n_38),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_26),
.A2(n_32),
.B1(n_35),
.B2(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_26),
.A2(n_32),
.B1(n_38),
.B2(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_26),
.A2(n_32),
.B1(n_83),
.B2(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_26),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_26),
.A2(n_32),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_26),
.A2(n_32),
.B1(n_116),
.B2(n_250),
.Y(n_267)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B(n_31),
.C(n_32),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_29),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_27),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g215 ( 
.A1(n_27),
.A2(n_29),
.B(n_153),
.C(n_216),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_29),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_32),
.Y(n_197)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_44),
.Y(n_45)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_54),
.B1(n_55),
.B2(n_64),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_46),
.B1(n_50),
.B2(n_52),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_46),
.B1(n_50),
.B2(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_43),
.A2(n_46),
.B1(n_52),
.B2(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_43),
.A2(n_46),
.B1(n_67),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_43),
.A2(n_46),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_43),
.A2(n_46),
.B1(n_177),
.B2(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_43),
.A2(n_46),
.B1(n_193),
.B2(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_43),
.A2(n_46),
.B1(n_234),
.B2(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_43),
.A2(n_46),
.B1(n_120),
.B2(n_246),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_44),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_44),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_45),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_46),
.B(n_153),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_47),
.B(n_49),
.Y(n_181)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_48),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_54),
.A2(n_55),
.B1(n_93),
.B2(n_95),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_58),
.B(n_62),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_58),
.B1(n_62),
.B2(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_58),
.B1(n_69),
.B2(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_56),
.A2(n_58),
.B1(n_80),
.B2(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_56),
.A2(n_58),
.B1(n_139),
.B2(n_141),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_56),
.A2(n_58),
.B1(n_141),
.B2(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_56),
.A2(n_58),
.B1(n_166),
.B2(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_56),
.A2(n_58),
.B1(n_173),
.B2(n_205),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_56),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_56),
.A2(n_58),
.B1(n_113),
.B2(n_256),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_57),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_58),
.B(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_58),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_59),
.B(n_61),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_59),
.B(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_60),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_65),
.A2(n_66),
.B(n_68),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_81),
.B(n_82),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_71),
.A2(n_72),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_79),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_73),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_73),
.A2(n_81),
.B1(n_82),
.B2(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_73),
.A2(n_79),
.B1(n_81),
.B2(n_281),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_77),
.B(n_78),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_74),
.A2(n_77),
.B1(n_78),
.B2(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_74),
.A2(n_77),
.B1(n_132),
.B2(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_74),
.A2(n_77),
.B1(n_135),
.B2(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_74),
.A2(n_77),
.B1(n_168),
.B2(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_74),
.A2(n_77),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_74),
.A2(n_77),
.B1(n_111),
.B2(n_220),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_75),
.A2(n_76),
.B1(n_131),
.B2(n_134),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_75),
.A2(n_76),
.B1(n_185),
.B2(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_77),
.B(n_153),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_79),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_82),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_97),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_91),
.B1(n_92),
.B2(n_96),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_89),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_93),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_122),
.B(n_298),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_121),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_101),
.B(n_121),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_106),
.C(n_107),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_102),
.B(n_106),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_107),
.A2(n_108),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_114),
.C(n_118),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_109),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_110),
.B(n_112),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_114),
.A2(n_115),
.B1(n_118),
.B2(n_119),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_121),
.Y(n_300)
);

AOI321xp33_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_275),
.A3(n_286),
.B1(n_292),
.B2(n_297),
.C(n_301),
.Y(n_122)
);

NOR3xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_240),
.C(n_271),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_209),
.B(n_239),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_187),
.B(n_208),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_170),
.B(n_186),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_160),
.B(n_169),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_148),
.B(n_159),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_136),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_130),
.B(n_136),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_143),
.B2(n_147),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_137),
.B(n_147),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_140),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_143),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_154),
.B(n_158),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_152),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_161),
.B(n_162),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_163),
.B(n_171),
.Y(n_186)
);

FAx1_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_165),
.CI(n_167),
.CON(n_163),
.SN(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_171),
.Y(n_188)
);

FAx1_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_174),
.CI(n_178),
.CON(n_171),
.SN(n_171)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_176),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_183),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_188),
.B(n_189),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_201),
.B2(n_202),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_204),
.C(n_206),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_194),
.B1(n_195),
.B2(n_200),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_192),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_198),
.C(n_200),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_197),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_199),
.Y(n_219)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_206),
.B2(n_207),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_203),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_204),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_205),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_210),
.B(n_211),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_224),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_213),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_213),
.B(n_223),
.C(n_224),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_217),
.B2(n_218),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_214),
.B(n_218),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_221),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_235),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_232),
.B2(n_233),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_232),
.C(n_235),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_230),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_238),
.Y(n_249)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

AOI21xp33_ASAP7_75t_L g293 ( 
.A1(n_241),
.A2(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_258),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_242),
.B(n_258),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_253),
.C(n_257),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_252),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_247),
.B1(n_248),
.B2(n_251),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_245),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_SL g269 ( 
.A(n_247),
.B(n_251),
.C(n_252),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_257),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_255),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_269),
.B2(n_270),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_262),
.C(n_270),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_266),
.C(n_268),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_265),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_269),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_273),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_283),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_276),
.B(n_283),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_280),
.C(n_282),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_277),
.A2(n_278),
.B1(n_280),
.B2(n_291),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_280),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_287),
.A2(n_293),
.B(n_296),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_288),
.B(n_289),
.Y(n_296)
);


endmodule