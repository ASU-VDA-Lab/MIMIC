module fake_jpeg_24163_n_233 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_233);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_233;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_17),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_7),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_40),
.Y(n_57)
);

OR2x2_ASAP7_75t_SL g40 ( 
.A(n_20),
.B(n_0),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx5_ASAP7_75t_SL g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_28),
.A2(n_7),
.B(n_1),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_34),
.C(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_8),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_45),
.B(n_24),
.Y(n_64)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_30),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_18),
.B1(n_27),
.B2(n_25),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_50),
.A2(n_51),
.B1(n_60),
.B2(n_63),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_47),
.A2(n_30),
.B1(n_28),
.B2(n_19),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_23),
.B(n_26),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_59),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_42),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_19),
.B1(n_36),
.B2(n_34),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_52),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_26),
.B1(n_33),
.B2(n_16),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_66),
.Y(n_81)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_18),
.B1(n_21),
.B2(n_22),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_68),
.A2(n_76),
.B1(n_4),
.B2(n_5),
.Y(n_106)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_77),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_40),
.A2(n_19),
.B1(n_32),
.B2(n_31),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_72),
.A2(n_33),
.B(n_2),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_45),
.B(n_31),
.Y(n_73)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_38),
.B(n_24),
.Y(n_74)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_25),
.Y(n_75)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_27),
.B1(n_23),
.B2(n_22),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_39),
.B(n_21),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_39),
.B(n_16),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_79),
.Y(n_89)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_87),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_33),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_93),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_90),
.B(n_80),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_91),
.B(n_99),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_33),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_9),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_109),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_97),
.B(n_53),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_57),
.A2(n_0),
.B(n_3),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_106),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_57),
.B(n_4),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_64),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_100),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_55),
.B(n_4),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_88),
.A2(n_76),
.B1(n_70),
.B2(n_67),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_119),
.B1(n_131),
.B2(n_136),
.Y(n_140)
);

AO22x1_ASAP7_75t_SL g115 ( 
.A1(n_86),
.A2(n_63),
.B1(n_51),
.B2(n_60),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_115),
.A2(n_92),
.B1(n_101),
.B2(n_96),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_116),
.B(n_109),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_53),
.B1(n_48),
.B2(n_70),
.Y(n_119)
);

OA21x2_ASAP7_75t_L g120 ( 
.A1(n_90),
.A2(n_97),
.B(n_99),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_120),
.A2(n_134),
.B(n_81),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_129),
.C(n_92),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_53),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_94),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_85),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_130),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_97),
.A2(n_66),
.B1(n_69),
.B2(n_49),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_98),
.Y(n_132)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_5),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_101),
.A2(n_69),
.B1(n_49),
.B2(n_59),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_85),
.B(n_59),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_143),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_147),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_127),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_145),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_114),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_151),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_148),
.A2(n_156),
.B1(n_131),
.B2(n_113),
.Y(n_161)
);

OAI32xp33_ASAP7_75t_L g150 ( 
.A1(n_115),
.A2(n_96),
.A3(n_102),
.B1(n_54),
.B2(n_56),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_153),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_123),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_89),
.C(n_102),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_160),
.C(n_116),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_125),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_124),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_157),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_115),
.A2(n_89),
.B1(n_107),
.B2(n_94),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_136),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_110),
.B(n_98),
.Y(n_158)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_120),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_126),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_108),
.C(n_104),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_175),
.B1(n_177),
.B2(n_138),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_169),
.C(n_148),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_120),
.C(n_122),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_117),
.B(n_119),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_170),
.A2(n_151),
.B(n_144),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_119),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_173),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_140),
.A2(n_119),
.B1(n_111),
.B2(n_135),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_172),
.A2(n_132),
.B1(n_104),
.B2(n_144),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_157),
.A2(n_118),
.B1(n_126),
.B2(n_135),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_134),
.Y(n_176)
);

OAI322xp33_ASAP7_75t_L g178 ( 
.A1(n_176),
.A2(n_158),
.A3(n_153),
.B1(n_143),
.B2(n_142),
.C1(n_141),
.C2(n_152),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_140),
.A2(n_132),
.B1(n_128),
.B2(n_134),
.Y(n_177)
);

HB1xp67_ASAP7_75t_SL g197 ( 
.A(n_178),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_179),
.A2(n_174),
.B1(n_165),
.B2(n_161),
.Y(n_199)
);

OAI21xp33_ASAP7_75t_SL g180 ( 
.A1(n_177),
.A2(n_150),
.B(n_138),
.Y(n_180)
);

HB1xp67_ASAP7_75t_SL g203 ( 
.A(n_180),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_183),
.C(n_185),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_146),
.Y(n_182)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_149),
.C(n_154),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_184),
.B(n_186),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_154),
.C(n_155),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_139),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_192),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_151),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_190),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_191),
.A2(n_174),
.B1(n_167),
.B2(n_165),
.Y(n_200)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_170),
.C(n_163),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_201),
.C(n_202),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_187),
.Y(n_206)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_200),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_171),
.C(n_167),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_176),
.C(n_144),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_6),
.C(n_10),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_189),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_208),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_203),
.A2(n_190),
.B(n_192),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_207),
.A2(n_210),
.B(n_202),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_182),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_186),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_191),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_212),
.A2(n_214),
.B1(n_211),
.B2(n_210),
.Y(n_217)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_213),
.B(n_196),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_194),
.Y(n_223)
);

NOR2xp67_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_197),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_216),
.B(n_6),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_220),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_207),
.A2(n_201),
.B1(n_198),
.B2(n_196),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_213),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_222),
.B(n_224),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_221),
.A2(n_218),
.B1(n_215),
.B2(n_13),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_226),
.B(n_10),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_223),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_227),
.A2(n_10),
.B(n_12),
.Y(n_228)
);

AO21x1_ASAP7_75t_L g232 ( 
.A1(n_228),
.A2(n_12),
.B(n_13),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_229),
.A2(n_230),
.B(n_227),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_225),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_231),
.B(n_232),
.Y(n_233)
);


endmodule