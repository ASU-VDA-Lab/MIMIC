module fake_aes_6674_n_673 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_673);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_673;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_L g77 ( .A(n_51), .Y(n_77) );
CKINVDCx16_ASAP7_75t_R g78 ( .A(n_35), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_37), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_46), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_63), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_21), .Y(n_82) );
CKINVDCx16_ASAP7_75t_R g83 ( .A(n_74), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_40), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_15), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_60), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_61), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_19), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_65), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_27), .Y(n_90) );
INVxp33_ASAP7_75t_L g91 ( .A(n_68), .Y(n_91) );
INVxp67_ASAP7_75t_SL g92 ( .A(n_32), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_59), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_17), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_16), .Y(n_95) );
NOR2xp67_ASAP7_75t_L g96 ( .A(n_50), .B(n_28), .Y(n_96) );
CKINVDCx20_ASAP7_75t_R g97 ( .A(n_56), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_42), .Y(n_98) );
OR2x2_ASAP7_75t_L g99 ( .A(n_39), .B(n_41), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_55), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_23), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_14), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_5), .Y(n_103) );
INVxp33_ASAP7_75t_SL g104 ( .A(n_15), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_76), .Y(n_105) );
NOR2xp67_ASAP7_75t_L g106 ( .A(n_47), .B(n_64), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_4), .Y(n_107) );
INVxp33_ASAP7_75t_SL g108 ( .A(n_24), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_0), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_19), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_23), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_49), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_72), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_31), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_8), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_36), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_73), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_0), .Y(n_118) );
INVxp67_ASAP7_75t_L g119 ( .A(n_3), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_30), .Y(n_120) );
CKINVDCx16_ASAP7_75t_R g121 ( .A(n_69), .Y(n_121) );
INVxp67_ASAP7_75t_SL g122 ( .A(n_34), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_62), .Y(n_123) );
INVxp67_ASAP7_75t_SL g124 ( .A(n_54), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g125 ( .A(n_91), .B(n_1), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_81), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_97), .Y(n_127) );
CKINVDCx16_ASAP7_75t_R g128 ( .A(n_78), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_116), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_79), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_111), .Y(n_131) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_79), .A2(n_75), .B(n_71), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_83), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_121), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_80), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_123), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_123), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_80), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_84), .Y(n_139) );
AND2x4_ASAP7_75t_L g140 ( .A(n_82), .B(n_1), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_104), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_116), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_108), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_77), .Y(n_144) );
OA21x2_ASAP7_75t_L g145 ( .A1(n_84), .A2(n_70), .B(n_67), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_117), .Y(n_146) );
INVxp67_ASAP7_75t_L g147 ( .A(n_82), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_119), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_86), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_100), .Y(n_150) );
BUFx3_ASAP7_75t_L g151 ( .A(n_117), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_86), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_89), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_89), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_90), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_90), .Y(n_156) );
NAND2xp33_ASAP7_75t_SL g157 ( .A(n_85), .B(n_2), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_105), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_87), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_93), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_85), .B(n_2), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_92), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_93), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_98), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_88), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_98), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_88), .B(n_3), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_140), .B(n_109), .Y(n_168) );
BUFx2_ASAP7_75t_L g169 ( .A(n_136), .Y(n_169) );
INVx4_ASAP7_75t_L g170 ( .A(n_140), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_129), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_140), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_140), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_163), .Y(n_174) );
INVx4_ASAP7_75t_L g175 ( .A(n_140), .Y(n_175) );
NAND2x1p5_ASAP7_75t_L g176 ( .A(n_161), .B(n_99), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_161), .Y(n_177) );
AND2x6_ASAP7_75t_L g178 ( .A(n_161), .B(n_112), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_147), .B(n_109), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_167), .Y(n_180) );
AO21x2_ASAP7_75t_L g181 ( .A1(n_125), .A2(n_112), .B(n_113), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_167), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_147), .B(n_120), .Y(n_183) );
CKINVDCx8_ASAP7_75t_R g184 ( .A(n_128), .Y(n_184) );
BUFx3_ASAP7_75t_L g185 ( .A(n_151), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_163), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_163), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_130), .B(n_94), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_144), .B(n_120), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_167), .Y(n_190) );
AND2x4_ASAP7_75t_L g191 ( .A(n_166), .B(n_94), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_139), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_166), .B(n_95), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_139), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_130), .B(n_114), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_139), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_137), .B(n_114), .Y(n_197) );
AND2x2_ASAP7_75t_SL g198 ( .A(n_128), .B(n_99), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_133), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_165), .A2(n_107), .B1(n_102), .B2(n_103), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_150), .B(n_113), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_159), .B(n_124), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_139), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_152), .Y(n_204) );
BUFx3_ASAP7_75t_L g205 ( .A(n_151), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_152), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_163), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_135), .B(n_95), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g209 ( .A1(n_148), .A2(n_115), .B1(n_118), .B2(n_110), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_163), .Y(n_210) );
BUFx2_ASAP7_75t_L g211 ( .A(n_134), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_129), .Y(n_212) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_129), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_163), .Y(n_214) );
OR2x2_ASAP7_75t_L g215 ( .A(n_135), .B(n_101), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_138), .B(n_118), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_152), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_129), .Y(n_218) );
BUFx2_ASAP7_75t_L g219 ( .A(n_131), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_156), .Y(n_220) );
OR2x2_ASAP7_75t_SL g221 ( .A(n_132), .B(n_101), .Y(n_221) );
INVx3_ASAP7_75t_L g222 ( .A(n_163), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_156), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_138), .B(n_110), .Y(n_224) );
NOR2x1p5_ASAP7_75t_L g225 ( .A(n_126), .B(n_122), .Y(n_225) );
NOR2x1p5_ASAP7_75t_L g226 ( .A(n_127), .B(n_4), .Y(n_226) );
BUFx2_ASAP7_75t_L g227 ( .A(n_141), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_129), .Y(n_228) );
AO22x2_ASAP7_75t_L g229 ( .A1(n_149), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_229) );
NOR3xp33_ASAP7_75t_SL g230 ( .A(n_199), .B(n_143), .C(n_157), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_192), .Y(n_231) );
NAND3xp33_ASAP7_75t_SL g232 ( .A(n_199), .B(n_162), .C(n_158), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_194), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_227), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_179), .B(n_164), .Y(n_235) );
NAND3xp33_ASAP7_75t_SL g236 ( .A(n_184), .B(n_157), .C(n_125), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_177), .B(n_164), .Y(n_237) );
INVx3_ASAP7_75t_L g238 ( .A(n_170), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_179), .B(n_155), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_179), .B(n_155), .Y(n_240) );
NAND3xp33_ASAP7_75t_SL g241 ( .A(n_184), .B(n_154), .C(n_153), .Y(n_241) );
OR2x2_ASAP7_75t_L g242 ( .A(n_227), .B(n_149), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_196), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_203), .Y(n_244) );
INVxp67_ASAP7_75t_L g245 ( .A(n_169), .Y(n_245) );
NAND2xp33_ASAP7_75t_SL g246 ( .A(n_169), .B(n_225), .Y(n_246) );
AND2x4_ASAP7_75t_L g247 ( .A(n_180), .B(n_154), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_204), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_206), .Y(n_249) );
AO22x1_ASAP7_75t_L g250 ( .A1(n_178), .A2(n_153), .B1(n_156), .B2(n_160), .Y(n_250) );
BUFx3_ASAP7_75t_L g251 ( .A(n_178), .Y(n_251) );
BUFx3_ASAP7_75t_L g252 ( .A(n_185), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_176), .B(n_160), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_178), .A2(n_151), .B1(n_160), .B2(n_146), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_217), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_176), .B(n_146), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_220), .Y(n_257) );
AOI211xp5_ASAP7_75t_L g258 ( .A1(n_182), .A2(n_146), .B(n_142), .C(n_129), .Y(n_258) );
INVx3_ASAP7_75t_L g259 ( .A(n_170), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_223), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_172), .Y(n_261) );
BUFx3_ASAP7_75t_L g262 ( .A(n_185), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_219), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_170), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_176), .B(n_142), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g266 ( .A1(n_198), .A2(n_142), .B1(n_129), .B2(n_106), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_178), .B(n_145), .Y(n_267) );
INVx8_ASAP7_75t_L g268 ( .A(n_178), .Y(n_268) );
OAI21xp33_ASAP7_75t_L g269 ( .A1(n_173), .A2(n_96), .B(n_145), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_175), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_175), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_175), .B(n_168), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_171), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_168), .B(n_145), .Y(n_274) );
INVxp67_ASAP7_75t_L g275 ( .A(n_219), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_205), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_212), .Y(n_277) );
INVx1_ASAP7_75t_SL g278 ( .A(n_178), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_183), .B(n_132), .Y(n_279) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_205), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_168), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_188), .Y(n_282) );
NAND3xp33_ASAP7_75t_SL g283 ( .A(n_200), .B(n_6), .C(n_7), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_188), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_188), .B(n_132), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_190), .B(n_145), .Y(n_286) );
NOR3xp33_ASAP7_75t_SL g287 ( .A(n_197), .B(n_8), .C(n_9), .Y(n_287) );
INVx4_ASAP7_75t_L g288 ( .A(n_191), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_216), .B(n_145), .Y(n_289) );
INVxp67_ASAP7_75t_L g290 ( .A(n_211), .Y(n_290) );
AND2x4_ASAP7_75t_L g291 ( .A(n_216), .B(n_9), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_191), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_171), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_218), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_191), .B(n_132), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_242), .B(n_193), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_243), .Y(n_297) );
OR2x2_ASAP7_75t_L g298 ( .A(n_242), .B(n_211), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_231), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_231), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_291), .B(n_208), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_233), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_268), .Y(n_303) );
INVxp67_ASAP7_75t_L g304 ( .A(n_234), .Y(n_304) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_268), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_285), .A2(n_201), .B(n_181), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_243), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g308 ( .A1(n_288), .A2(n_198), .B1(n_193), .B2(n_208), .Y(n_308) );
INVx2_ASAP7_75t_SL g309 ( .A(n_268), .Y(n_309) );
BUFx12f_ASAP7_75t_L g310 ( .A(n_234), .Y(n_310) );
OR2x6_ASAP7_75t_L g311 ( .A(n_268), .B(n_229), .Y(n_311) );
INVx2_ASAP7_75t_SL g312 ( .A(n_268), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_251), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_291), .B(n_193), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_233), .Y(n_315) );
CKINVDCx11_ASAP7_75t_R g316 ( .A(n_263), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_288), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_264), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g319 ( .A(n_288), .B(n_208), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_244), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_244), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_255), .Y(n_322) );
INVx3_ASAP7_75t_L g323 ( .A(n_288), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_255), .Y(n_324) );
OR2x2_ASAP7_75t_L g325 ( .A(n_245), .B(n_215), .Y(n_325) );
INVx3_ASAP7_75t_L g326 ( .A(n_238), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g327 ( .A1(n_291), .A2(n_229), .B1(n_181), .B2(n_195), .Y(n_327) );
BUFx3_ASAP7_75t_L g328 ( .A(n_251), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_291), .B(n_215), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_257), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_295), .A2(n_181), .B(n_189), .Y(n_331) );
INVx3_ASAP7_75t_L g332 ( .A(n_238), .Y(n_332) );
NOR2x1_ASAP7_75t_SL g333 ( .A(n_251), .B(n_224), .Y(n_333) );
O2A1O1Ixp33_ASAP7_75t_L g334 ( .A1(n_253), .A2(n_202), .B(n_226), .C(n_187), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_279), .A2(n_132), .B(n_214), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_275), .B(n_209), .Y(n_336) );
BUFx4_ASAP7_75t_SL g337 ( .A(n_282), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_290), .B(n_221), .Y(n_338) );
A2O1A1Ixp33_ASAP7_75t_L g339 ( .A1(n_261), .A2(n_284), .B(n_292), .C(n_282), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_257), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_241), .B(n_221), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_256), .B(n_10), .Y(n_342) );
AOI21x1_ASAP7_75t_L g343 ( .A1(n_274), .A2(n_174), .B(n_186), .Y(n_343) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_252), .Y(n_344) );
AOI21xp5_ASAP7_75t_L g345 ( .A1(n_267), .A2(n_174), .B(n_207), .Y(n_345) );
CKINVDCx6p67_ASAP7_75t_R g346 ( .A(n_265), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_322), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_336), .A2(n_236), .B1(n_232), .B2(n_266), .Y(n_348) );
INVx4_ASAP7_75t_L g349 ( .A(n_303), .Y(n_349) );
AO21x2_ASAP7_75t_L g350 ( .A1(n_327), .A2(n_269), .B(n_286), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_308), .A2(n_283), .B1(n_229), .B2(n_237), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_311), .A2(n_281), .B1(n_246), .B2(n_292), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_327), .A2(n_261), .B1(n_260), .B2(n_284), .Y(n_353) );
NAND3xp33_ASAP7_75t_L g354 ( .A(n_334), .B(n_258), .C(n_287), .Y(n_354) );
OAI21xp5_ASAP7_75t_L g355 ( .A1(n_331), .A2(n_289), .B(n_269), .Y(n_355) );
BUFx2_ASAP7_75t_SL g356 ( .A(n_303), .Y(n_356) );
OAI21x1_ASAP7_75t_L g357 ( .A1(n_335), .A2(n_289), .B(n_254), .Y(n_357) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_301), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_311), .A2(n_281), .B1(n_247), .B2(n_237), .Y(n_359) );
BUFx2_ASAP7_75t_SL g360 ( .A(n_303), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_311), .A2(n_260), .B1(n_278), .B2(n_235), .Y(n_361) );
AOI22xp33_ASAP7_75t_SL g362 ( .A1(n_311), .A2(n_229), .B1(n_237), .B2(n_247), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_329), .B(n_247), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_311), .A2(n_237), .B1(n_247), .B2(n_272), .Y(n_364) );
AOI22xp33_ASAP7_75t_SL g365 ( .A1(n_329), .A2(n_278), .B1(n_239), .B2(n_240), .Y(n_365) );
AOI21xp5_ASAP7_75t_SL g366 ( .A1(n_301), .A2(n_250), .B(n_252), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_322), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_314), .B(n_249), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_324), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_299), .B(n_250), .Y(n_370) );
OAI22xp5_ASAP7_75t_L g371 ( .A1(n_324), .A2(n_248), .B1(n_249), .B2(n_258), .Y(n_371) );
AO21x2_ASAP7_75t_L g372 ( .A1(n_306), .A2(n_343), .B(n_341), .Y(n_372) );
BUFx3_ASAP7_75t_L g373 ( .A(n_303), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_338), .A2(n_264), .B1(n_270), .B2(n_271), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_299), .B(n_248), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_330), .Y(n_376) );
BUFx4_ASAP7_75t_R g377 ( .A(n_337), .Y(n_377) );
AOI21xp33_ASAP7_75t_L g378 ( .A1(n_342), .A2(n_276), .B(n_280), .Y(n_378) );
INVx2_ASAP7_75t_SL g379 ( .A(n_368), .Y(n_379) );
AND2x6_ASAP7_75t_SL g380 ( .A(n_377), .B(n_316), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_347), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_348), .A2(n_296), .B1(n_298), .B2(n_304), .C(n_325), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_363), .B(n_296), .Y(n_383) );
AO221x1_ASAP7_75t_L g384 ( .A1(n_361), .A2(n_353), .B1(n_371), .B2(n_362), .C(n_366), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_363), .B(n_314), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_363), .B(n_298), .Y(n_386) );
AOI21xp5_ASAP7_75t_L g387 ( .A1(n_355), .A2(n_345), .B(n_339), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_362), .A2(n_342), .B1(n_346), .B2(n_340), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_358), .B(n_325), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_368), .B(n_330), .Y(n_390) );
BUFx3_ASAP7_75t_L g391 ( .A(n_373), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_359), .A2(n_310), .B1(n_340), .B2(n_302), .Y(n_392) );
AOI21xp5_ASAP7_75t_L g393 ( .A1(n_355), .A2(n_300), .B(n_320), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_368), .Y(n_394) );
OAI22xp5_ASAP7_75t_SL g395 ( .A1(n_352), .A2(n_310), .B1(n_321), .B2(n_300), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_364), .A2(n_302), .B1(n_315), .B2(n_320), .Y(n_396) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_373), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_347), .B(n_315), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_367), .B(n_321), .Y(n_399) );
OAI22xp33_ASAP7_75t_L g400 ( .A1(n_351), .A2(n_307), .B1(n_297), .B2(n_303), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_367), .B(n_297), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_351), .A2(n_319), .B1(n_317), .B2(n_323), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_369), .Y(n_403) );
AO31x2_ASAP7_75t_L g404 ( .A1(n_353), .A2(n_307), .A3(n_333), .B(n_228), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_365), .A2(n_313), .B1(n_328), .B2(n_344), .Y(n_405) );
OAI221xp5_ASAP7_75t_SL g406 ( .A1(n_382), .A2(n_365), .B1(n_369), .B2(n_376), .C(n_354), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_404), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_404), .Y(n_408) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_404), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_381), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_384), .A2(n_354), .B1(n_378), .B2(n_376), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_381), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_380), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_403), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_403), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_399), .Y(n_416) );
AOI222xp33_ASAP7_75t_L g417 ( .A1(n_386), .A2(n_361), .B1(n_375), .B2(n_371), .C1(n_370), .C2(n_374), .Y(n_417) );
NOR4xp25_ASAP7_75t_SL g418 ( .A(n_384), .B(n_378), .C(n_350), .D(n_230), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_404), .Y(n_419) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_397), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_394), .B(n_401), .Y(n_421) );
BUFx3_ASAP7_75t_L g422 ( .A(n_391), .Y(n_422) );
INVx2_ASAP7_75t_SL g423 ( .A(n_397), .Y(n_423) );
BUFx2_ASAP7_75t_L g424 ( .A(n_404), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_390), .B(n_350), .Y(n_425) );
OAI21xp33_ASAP7_75t_L g426 ( .A1(n_388), .A2(n_375), .B(n_370), .Y(n_426) );
NAND3xp33_ASAP7_75t_L g427 ( .A(n_387), .B(n_344), .C(n_349), .Y(n_427) );
INVx3_ASAP7_75t_L g428 ( .A(n_397), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_395), .A2(n_350), .B1(n_372), .B2(n_357), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_399), .Y(n_430) );
OAI22xp33_ASAP7_75t_L g431 ( .A1(n_379), .A2(n_349), .B1(n_373), .B2(n_313), .Y(n_431) );
AOI222xp33_ASAP7_75t_L g432 ( .A1(n_395), .A2(n_333), .B1(n_318), .B2(n_276), .C1(n_349), .C2(n_323), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_401), .Y(n_433) );
INVx4_ASAP7_75t_L g434 ( .A(n_397), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_398), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_397), .Y(n_436) );
NOR2x1p5_ASAP7_75t_L g437 ( .A(n_391), .B(n_349), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_390), .B(n_350), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_390), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_379), .B(n_372), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_421), .Y(n_441) );
AND2x2_ASAP7_75t_SL g442 ( .A(n_424), .B(n_402), .Y(n_442) );
INVx4_ASAP7_75t_L g443 ( .A(n_422), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_417), .A2(n_385), .B1(n_396), .B2(n_392), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_414), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_425), .B(n_372), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_440), .B(n_389), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_414), .Y(n_448) );
AOI211xp5_ASAP7_75t_L g449 ( .A1(n_406), .A2(n_400), .B(n_405), .C(n_383), .Y(n_449) );
OAI22xp5_ASAP7_75t_SL g450 ( .A1(n_413), .A2(n_360), .B1(n_356), .B2(n_312), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_425), .B(n_372), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_408), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_425), .B(n_393), .Y(n_453) );
AOI33xp33_ASAP7_75t_L g454 ( .A1(n_411), .A2(n_385), .A3(n_228), .B1(n_214), .B2(n_207), .B3(n_187), .Y(n_454) );
AOI322xp5_ASAP7_75t_L g455 ( .A1(n_435), .A2(n_10), .A3(n_11), .B1(n_12), .B2(n_13), .C1(n_14), .C2(n_16), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_438), .B(n_357), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_414), .Y(n_457) );
AOI21xp5_ASAP7_75t_SL g458 ( .A1(n_437), .A2(n_305), .B(n_328), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_410), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_410), .Y(n_460) );
INVxp67_ASAP7_75t_L g461 ( .A(n_421), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_440), .B(n_11), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_408), .Y(n_463) );
AOI33xp33_ASAP7_75t_L g464 ( .A1(n_411), .A2(n_186), .A3(n_218), .B1(n_17), .B2(n_18), .B3(n_20), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_412), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_421), .Y(n_466) );
INVx6_ASAP7_75t_L g467 ( .A(n_434), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_433), .Y(n_468) );
OAI31xp33_ASAP7_75t_L g469 ( .A1(n_406), .A2(n_323), .A3(n_317), .B(n_326), .Y(n_469) );
BUFx2_ASAP7_75t_L g470 ( .A(n_434), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_438), .B(n_12), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_438), .B(n_13), .Y(n_472) );
INVx1_ASAP7_75t_SL g473 ( .A(n_422), .Y(n_473) );
INVx1_ASAP7_75t_SL g474 ( .A(n_422), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_416), .B(n_318), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_412), .B(n_18), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_433), .B(n_20), .Y(n_477) );
NAND2xp33_ASAP7_75t_SL g478 ( .A(n_418), .B(n_305), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_434), .B(n_343), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_417), .A2(n_360), .B1(n_356), .B2(n_317), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_415), .Y(n_481) );
INVx2_ASAP7_75t_SL g482 ( .A(n_422), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_426), .A2(n_344), .B1(n_326), .B2(n_332), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_415), .B(n_21), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_439), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_408), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_408), .Y(n_487) );
OAI22xp33_ASAP7_75t_L g488 ( .A1(n_435), .A2(n_344), .B1(n_305), .B2(n_328), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_420), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_459), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_459), .Y(n_491) );
CKINVDCx16_ASAP7_75t_R g492 ( .A(n_443), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_460), .Y(n_493) );
CKINVDCx16_ASAP7_75t_R g494 ( .A(n_443), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_447), .B(n_424), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_452), .Y(n_496) );
CKINVDCx16_ASAP7_75t_R g497 ( .A(n_443), .Y(n_497) );
INVx1_ASAP7_75t_SL g498 ( .A(n_473), .Y(n_498) );
BUFx2_ASAP7_75t_L g499 ( .A(n_443), .Y(n_499) );
NAND2xp33_ASAP7_75t_R g500 ( .A(n_470), .B(n_418), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_465), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_447), .B(n_424), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_441), .B(n_407), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_466), .B(n_430), .Y(n_504) );
INVx1_ASAP7_75t_SL g505 ( .A(n_474), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_465), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_444), .A2(n_439), .B1(n_430), .B2(n_431), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_481), .Y(n_508) );
BUFx2_ASAP7_75t_L g509 ( .A(n_482), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_481), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_452), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_446), .B(n_407), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_446), .B(n_409), .Y(n_513) );
NAND2xp33_ASAP7_75t_R g514 ( .A(n_470), .B(n_22), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_468), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_461), .B(n_439), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_451), .B(n_409), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_471), .B(n_439), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_451), .B(n_419), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_458), .Y(n_520) );
INVxp33_ASAP7_75t_L g521 ( .A(n_458), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_471), .B(n_426), .Y(n_522) );
NAND4xp25_ASAP7_75t_SL g523 ( .A(n_455), .B(n_432), .C(n_429), .D(n_427), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_452), .Y(n_524) );
INVx2_ASAP7_75t_SL g525 ( .A(n_467), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_453), .B(n_429), .Y(n_526) );
BUFx2_ASAP7_75t_L g527 ( .A(n_482), .Y(n_527) );
NOR4xp25_ASAP7_75t_SL g528 ( .A(n_478), .B(n_432), .C(n_431), .D(n_25), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_445), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_469), .B(n_434), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_477), .B(n_22), .Y(n_531) );
INVx1_ASAP7_75t_SL g532 ( .A(n_467), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_445), .Y(n_533) );
INVx3_ASAP7_75t_L g534 ( .A(n_467), .Y(n_534) );
OAI322xp33_ASAP7_75t_L g535 ( .A1(n_477), .A2(n_427), .A3(n_25), .B1(n_24), .B2(n_423), .C1(n_213), .C2(n_212), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_472), .B(n_423), .Y(n_536) );
INVx1_ASAP7_75t_SL g537 ( .A(n_467), .Y(n_537) );
OAI31xp33_ASAP7_75t_SL g538 ( .A1(n_476), .A2(n_436), .A3(n_428), .B(n_33), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_444), .B(n_428), .Y(n_539) );
INVxp67_ASAP7_75t_SL g540 ( .A(n_463), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_448), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_448), .Y(n_542) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_450), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_456), .B(n_436), .Y(n_544) );
NOR3xp33_ASAP7_75t_L g545 ( .A(n_464), .B(n_428), .C(n_436), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_523), .A2(n_469), .B1(n_442), .B2(n_453), .Y(n_546) );
OAI21xp33_ASAP7_75t_L g547 ( .A1(n_538), .A2(n_455), .B(n_480), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_515), .B(n_472), .Y(n_548) );
OAI211xp5_ASAP7_75t_SL g549 ( .A1(n_531), .A2(n_480), .B(n_449), .C(n_462), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_490), .Y(n_550) );
NOR2xp33_ASAP7_75t_SL g551 ( .A(n_492), .B(n_450), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_504), .B(n_484), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_514), .A2(n_442), .B1(n_484), .B2(n_476), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_499), .Y(n_554) );
O2A1O1Ixp33_ASAP7_75t_L g555 ( .A1(n_535), .A2(n_475), .B(n_449), .C(n_488), .Y(n_555) );
NAND2x1p5_ASAP7_75t_L g556 ( .A(n_499), .B(n_457), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_517), .B(n_457), .Y(n_557) );
NOR3xp33_ASAP7_75t_L g558 ( .A(n_545), .B(n_454), .C(n_428), .Y(n_558) );
OAI32xp33_ASAP7_75t_L g559 ( .A1(n_494), .A2(n_487), .A3(n_486), .B1(n_463), .B2(n_485), .Y(n_559) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_527), .Y(n_560) );
AOI222xp33_ASAP7_75t_L g561 ( .A1(n_507), .A2(n_442), .B1(n_486), .B2(n_483), .C1(n_479), .C2(n_489), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_497), .A2(n_486), .B1(n_479), .B2(n_428), .Y(n_562) );
OAI22xp33_ASAP7_75t_L g563 ( .A1(n_543), .A2(n_489), .B1(n_420), .B2(n_479), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_491), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_512), .B(n_479), .Y(n_565) );
INVxp67_ASAP7_75t_L g566 ( .A(n_509), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_539), .A2(n_489), .B1(n_420), .B2(n_344), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_517), .B(n_420), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_512), .B(n_420), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_493), .Y(n_570) );
AOI221xp5_ASAP7_75t_L g571 ( .A1(n_522), .A2(n_516), .B1(n_519), .B2(n_513), .C(n_526), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_530), .A2(n_420), .B(n_313), .Y(n_572) );
XNOR2x1_ASAP7_75t_L g573 ( .A(n_526), .B(n_26), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_501), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_513), .B(n_420), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_496), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_506), .Y(n_577) );
OAI31xp33_ASAP7_75t_L g578 ( .A1(n_521), .A2(n_312), .A3(n_309), .B(n_326), .Y(n_578) );
AO22x1_ASAP7_75t_L g579 ( .A1(n_520), .A2(n_305), .B1(n_309), .B2(n_332), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_495), .B(n_212), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_519), .B(n_212), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_530), .A2(n_262), .B(n_305), .Y(n_582) );
INVxp67_ASAP7_75t_L g583 ( .A(n_527), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_540), .A2(n_262), .B(n_332), .Y(n_584) );
OAI31xp33_ASAP7_75t_L g585 ( .A1(n_532), .A2(n_332), .A3(n_259), .B(n_238), .Y(n_585) );
OAI22xp33_ASAP7_75t_L g586 ( .A1(n_520), .A2(n_259), .B1(n_270), .B2(n_271), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_498), .B(n_29), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_505), .B(n_38), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_525), .B(n_213), .Y(n_589) );
INVxp67_ASAP7_75t_L g590 ( .A(n_525), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_495), .A2(n_259), .B1(n_213), .B2(n_45), .Y(n_591) );
OAI221xp5_ASAP7_75t_L g592 ( .A1(n_500), .A2(n_213), .B1(n_222), .B2(n_210), .C(n_52), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_502), .B(n_43), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_571), .B(n_502), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_571), .B(n_503), .Y(n_595) );
INVx1_ASAP7_75t_SL g596 ( .A(n_557), .Y(n_596) );
INVxp67_ASAP7_75t_SL g597 ( .A(n_554), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_576), .Y(n_598) );
NAND3xp33_ASAP7_75t_L g599 ( .A(n_561), .B(n_528), .C(n_503), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_575), .B(n_544), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_550), .Y(n_601) );
BUFx2_ASAP7_75t_L g602 ( .A(n_556), .Y(n_602) );
NOR2xp33_ASAP7_75t_R g603 ( .A(n_551), .B(n_534), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_565), .B(n_544), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_556), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_548), .B(n_518), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_569), .B(n_496), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_564), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_570), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_552), .B(n_508), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_574), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_577), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_560), .Y(n_613) );
INVxp33_ASAP7_75t_L g614 ( .A(n_573), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_566), .B(n_510), .Y(n_615) );
NAND4xp25_ASAP7_75t_L g616 ( .A(n_553), .B(n_536), .C(n_537), .D(n_534), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_583), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_568), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_581), .Y(n_619) );
O2A1O1Ixp33_ASAP7_75t_L g620 ( .A1(n_549), .A2(n_542), .B(n_541), .C(n_533), .Y(n_620) );
INVxp67_ASAP7_75t_L g621 ( .A(n_590), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_559), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_580), .Y(n_623) );
NAND2xp33_ASAP7_75t_SL g624 ( .A(n_546), .B(n_529), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_547), .B(n_524), .Y(n_625) );
INVx1_ASAP7_75t_SL g626 ( .A(n_588), .Y(n_626) );
O2A1O1Ixp33_ASAP7_75t_SL g627 ( .A1(n_614), .A2(n_592), .B(n_563), .C(n_562), .Y(n_627) );
AOI31xp33_ASAP7_75t_L g628 ( .A1(n_622), .A2(n_593), .A3(n_572), .B(n_582), .Y(n_628) );
AO21x1_ASAP7_75t_L g629 ( .A1(n_624), .A2(n_578), .B(n_582), .Y(n_629) );
OAI221xp5_ASAP7_75t_L g630 ( .A1(n_624), .A2(n_592), .B1(n_558), .B2(n_555), .C(n_585), .Y(n_630) );
AOI21xp33_ASAP7_75t_L g631 ( .A1(n_599), .A2(n_587), .B(n_586), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_596), .B(n_511), .Y(n_632) );
OAI211xp5_ASAP7_75t_L g633 ( .A1(n_616), .A2(n_567), .B(n_572), .C(n_589), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_625), .B(n_584), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_601), .Y(n_635) );
NAND3xp33_ASAP7_75t_L g636 ( .A(n_622), .B(n_591), .C(n_579), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_594), .A2(n_584), .B1(n_210), .B2(n_222), .Y(n_637) );
O2A1O1Ixp33_ASAP7_75t_L g638 ( .A1(n_620), .A2(n_222), .B(n_210), .C(n_53), .Y(n_638) );
NOR2xp67_ASAP7_75t_L g639 ( .A(n_605), .B(n_44), .Y(n_639) );
OA22x2_ASAP7_75t_L g640 ( .A1(n_602), .A2(n_48), .B1(n_57), .B2(n_58), .Y(n_640) );
NOR2x1p5_ASAP7_75t_L g641 ( .A(n_595), .B(n_66), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_601), .Y(n_642) );
O2A1O1Ixp33_ASAP7_75t_L g643 ( .A1(n_621), .A2(n_273), .B(n_293), .C(n_294), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_635), .Y(n_644) );
NOR2xp33_ASAP7_75t_R g645 ( .A(n_640), .B(n_602), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g646 ( .A1(n_627), .A2(n_617), .B1(n_613), .B2(n_615), .C(n_610), .Y(n_646) );
INVx1_ASAP7_75t_SL g647 ( .A(n_632), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_634), .B(n_604), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_629), .B(n_603), .Y(n_649) );
AOI222xp33_ASAP7_75t_L g650 ( .A1(n_630), .A2(n_597), .B1(n_608), .B2(n_609), .C1(n_619), .C2(n_612), .Y(n_650) );
CKINVDCx5p33_ASAP7_75t_R g651 ( .A(n_641), .Y(n_651) );
NAND4xp75_ASAP7_75t_L g652 ( .A(n_631), .B(n_619), .C(n_623), .D(n_605), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_642), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_636), .A2(n_623), .B1(n_626), .B2(n_606), .Y(n_654) );
OAI211xp5_ASAP7_75t_SL g655 ( .A1(n_633), .A2(n_606), .B(n_612), .C(n_611), .Y(n_655) );
NAND4xp75_ASAP7_75t_L g656 ( .A(n_639), .B(n_607), .C(n_618), .D(n_600), .Y(n_656) );
AOI211xp5_ASAP7_75t_SL g657 ( .A1(n_628), .A2(n_600), .B(n_598), .C(n_277), .Y(n_657) );
OAI211xp5_ASAP7_75t_L g658 ( .A1(n_638), .A2(n_277), .B(n_598), .C(n_637), .Y(n_658) );
AOI21xp33_ASAP7_75t_SL g659 ( .A1(n_628), .A2(n_640), .B(n_643), .Y(n_659) );
INVxp67_ASAP7_75t_L g660 ( .A(n_636), .Y(n_660) );
A2O1A1Ixp33_ASAP7_75t_L g661 ( .A1(n_628), .A2(n_614), .B(n_624), .C(n_630), .Y(n_661) );
OR3x2_ASAP7_75t_L g662 ( .A(n_661), .B(n_660), .C(n_649), .Y(n_662) );
CKINVDCx20_ASAP7_75t_R g663 ( .A(n_651), .Y(n_663) );
AOI32xp33_ASAP7_75t_L g664 ( .A1(n_646), .A2(n_655), .A3(n_657), .B1(n_654), .B2(n_661), .Y(n_664) );
CKINVDCx5p33_ASAP7_75t_R g665 ( .A(n_654), .Y(n_665) );
OR3x2_ASAP7_75t_L g666 ( .A(n_662), .B(n_659), .C(n_645), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_665), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_663), .A2(n_650), .B1(n_652), .B2(n_656), .Y(n_668) );
INVx2_ASAP7_75t_SL g669 ( .A(n_667), .Y(n_669) );
OR3x1_ASAP7_75t_L g670 ( .A(n_666), .B(n_664), .C(n_645), .Y(n_670) );
AO22x2_ASAP7_75t_L g671 ( .A1(n_669), .A2(n_668), .B1(n_647), .B2(n_658), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_671), .A2(n_669), .B1(n_670), .B2(n_648), .Y(n_672) );
AOI21xp33_ASAP7_75t_SL g673 ( .A1(n_672), .A2(n_644), .B(n_653), .Y(n_673) );
endmodule