module fake_jpeg_26538_n_205 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_205);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_SL g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_11),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_0),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_20),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_26),
.Y(n_32)
);

BUFx2_ASAP7_75t_SL g47 ( 
.A(n_32),
.Y(n_47)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_23),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_37),
.B1(n_41),
.B2(n_18),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_24),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_24),
.A2(n_25),
.B1(n_23),
.B2(n_31),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_42),
.Y(n_48)
);

CKINVDCx12_ASAP7_75t_R g43 ( 
.A(n_42),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_53),
.B1(n_18),
.B2(n_31),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_54),
.B1(n_25),
.B2(n_32),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_35),
.B(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_51),
.Y(n_65)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_56),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_18),
.B1(n_20),
.B2(n_19),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_31),
.B1(n_29),
.B2(n_28),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_27),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_55),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_66),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_35),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_71),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_68),
.B1(n_69),
.B2(n_32),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_48),
.C(n_41),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_30),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_51),
.A2(n_39),
.B1(n_41),
.B2(n_31),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_33),
.B1(n_32),
.B2(n_38),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_33),
.B1(n_32),
.B2(n_38),
.Y(n_69)
);

AOI32xp33_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_39),
.A3(n_56),
.B1(n_25),
.B2(n_47),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_72),
.B(n_47),
.Y(n_77)
);

OAI32xp33_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_56),
.A3(n_39),
.B1(n_25),
.B2(n_27),
.Y(n_74)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_71),
.B(n_26),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_78),
.A2(n_84),
.B(n_14),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_73),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_79),
.B(n_80),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_73),
.B(n_29),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_82),
.A2(n_87),
.B1(n_61),
.B2(n_50),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_64),
.B1(n_68),
.B2(n_72),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_0),
.B(n_1),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_30),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_38),
.B1(n_33),
.B2(n_14),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_65),
.B(n_28),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_59),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_89),
.A2(n_91),
.B1(n_101),
.B2(n_82),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_83),
.A2(n_69),
.B1(n_62),
.B2(n_49),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_59),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_103),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_75),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_98),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_61),
.B(n_1),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_95),
.A2(n_102),
.B(n_77),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_84),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_21),
.Y(n_103)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_78),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_104),
.B(n_110),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_112),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_115),
.B1(n_46),
.B2(n_50),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_81),
.C(n_85),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_113),
.C(n_101),
.Y(n_121)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_75),
.Y(n_109)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_100),
.B(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_119),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_99),
.B(n_74),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_70),
.C(n_60),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_88),
.B1(n_70),
.B2(n_60),
.Y(n_115)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_26),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_30),
.B1(n_14),
.B2(n_22),
.Y(n_126)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_21),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_97),
.C(n_102),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_113),
.C(n_115),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_119),
.A2(n_90),
.B1(n_88),
.B2(n_57),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_126),
.B1(n_128),
.B2(n_133),
.Y(n_144)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_111),
.A2(n_14),
.B1(n_22),
.B2(n_17),
.Y(n_128)
);

XNOR2x1_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_21),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_130),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_114),
.B(n_21),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_0),
.B(n_1),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_22),
.B1(n_17),
.B2(n_30),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_134),
.A2(n_116),
.B(n_112),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_137),
.B(n_140),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_114),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_139),
.Y(n_159)
);

AOI322xp5_ASAP7_75t_L g140 ( 
.A1(n_129),
.A2(n_104),
.A3(n_117),
.B1(n_110),
.B2(n_118),
.C1(n_108),
.C2(n_40),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_117),
.C(n_108),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_142),
.C(n_139),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_12),
.C(n_40),
.Y(n_142)
);

BUFx12f_ASAP7_75t_SL g145 ( 
.A(n_122),
.Y(n_145)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_124),
.A2(n_17),
.B1(n_20),
.B2(n_19),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_146),
.B(n_150),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_132),
.Y(n_162)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

BUFx12_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

NOR3xp33_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_12),
.C(n_19),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_120),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_160),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_156),
.C(n_158),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_135),
.C(n_131),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_136),
.B(n_135),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_127),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_147),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_162),
.B(n_153),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_166),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_154),
.A2(n_143),
.B1(n_125),
.B2(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_152),
.B(n_156),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_169),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_163),
.A2(n_133),
.B1(n_136),
.B2(n_149),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_172),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_155),
.A2(n_149),
.B(n_128),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_11),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_174),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_10),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_167),
.A2(n_158),
.B1(n_159),
.B2(n_3),
.Y(n_175)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_168),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_12),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_159),
.C(n_12),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_179),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_12),
.C(n_40),
.Y(n_179)
);

BUFx24_ASAP7_75t_SL g184 ( 
.A(n_180),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_184),
.B(n_191),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_177),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_185)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_185),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_181),
.A2(n_9),
.B(n_12),
.Y(n_186)
);

AOI21xp33_ASAP7_75t_L g197 ( 
.A1(n_186),
.A2(n_188),
.B(n_2),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_183),
.A2(n_9),
.B(n_3),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_189),
.B(n_2),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_2),
.Y(n_191)
);

AOI322xp5_ASAP7_75t_L g201 ( 
.A1(n_192),
.A2(n_195),
.A3(n_197),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_201)
);

AOI21x1_ASAP7_75t_L g195 ( 
.A1(n_190),
.A2(n_175),
.B(n_179),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_187),
.A2(n_178),
.B1(n_176),
.B2(n_4),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_196),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_185),
.C(n_4),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_199),
.C(n_200),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_194),
.A2(n_3),
.B(n_4),
.Y(n_199)
);

OAI21x1_ASAP7_75t_L g203 ( 
.A1(n_201),
.A2(n_5),
.B(n_8),
.Y(n_203)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_8),
.C(n_202),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_8),
.Y(n_205)
);


endmodule