module fake_jpeg_10929_n_134 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_13),
.B(n_3),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_0),
.C(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_0),
.Y(n_50)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_38),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_36),
.A2(n_32),
.B1(n_30),
.B2(n_35),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_39),
.A2(n_46),
.B1(n_14),
.B2(n_19),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_21),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_54),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_32),
.A2(n_20),
.B1(n_21),
.B2(n_25),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_25),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_49),
.A2(n_29),
.B(n_33),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_50),
.B(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_29),
.B(n_17),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_26),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_62),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_26),
.B1(n_24),
.B2(n_27),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_45),
.B1(n_52),
.B2(n_41),
.Y(n_80)
);

O2A1O1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_54),
.A2(n_24),
.B(n_27),
.C(n_17),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_49),
.B(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_14),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_68),
.B1(n_71),
.B2(n_15),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_51),
.Y(n_65)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_22),
.B1(n_19),
.B2(n_18),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_70),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_49),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_22),
.B1(n_18),
.B2(n_15),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_72),
.B(n_75),
.Y(n_92)
);

AND2x6_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_11),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_76),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_64),
.A2(n_48),
.B1(n_41),
.B2(n_47),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_65),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_45),
.C(n_2),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_57),
.C(n_64),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_2),
.B1(n_10),
.B2(n_11),
.Y(n_86)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_87),
.Y(n_109)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_74),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_98),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_55),
.B(n_68),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_90),
.A2(n_80),
.B(n_82),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_84),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_91),
.B(n_94),
.Y(n_103)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

AOI221xp5_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_99),
.B1(n_89),
.B2(n_92),
.C(n_90),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_107),
.B(n_95),
.Y(n_115)
);

A2O1A1O1Ixp25_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_75),
.B(n_86),
.C(n_77),
.D(n_65),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_73),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_88),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_99),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_111),
.C(n_116),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_73),
.C(n_97),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_95),
.B1(n_97),
.B2(n_100),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_113),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_104),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_59),
.C(n_66),
.Y(n_116)
);

NOR2x1_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_114),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_108),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_120),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_109),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_122),
.B(n_121),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_127),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_114),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_128),
.A2(n_126),
.B1(n_124),
.B2(n_87),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_69),
.Y(n_129)
);

BUFx24_ASAP7_75t_SL g132 ( 
.A(n_129),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_130),
.C(n_61),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_132),
.Y(n_134)
);


endmodule