module real_aes_5688_n_422 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_421, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_401, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_399, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_415, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_400, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_408, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_409, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_398, n_89, n_277, n_331, n_93, n_182, n_363, n_417, n_323, n_199, n_350, n_142, n_223, n_67, n_405, n_368, n_250, n_85, n_406, n_45, n_5, n_244, n_118, n_139, n_402, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_416, n_410, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_412, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_404, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_413, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_407, n_217, n_419, n_55, n_62, n_411, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_420, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_418, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_414, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_403, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_422);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_421;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_401;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_399;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_415;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_400;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_408;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_409;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_398;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_417;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_405;
input n_368;
input n_250;
input n_85;
input n_406;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_402;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_416;
input n_410;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_412;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_404;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_413;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_407;
input n_217;
input n_419;
input n_55;
input n_62;
input n_411;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_420;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_418;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_414;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_403;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_422;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_786;
wire n_512;
wire n_795;
wire n_1379;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1317;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_527;
wire n_1342;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_1380;
wire n_488;
wire n_501;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1209;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_591;
wire n_1366;
wire n_678;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_1368;
wire n_994;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_617;
wire n_1404;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_895;
wire n_799;
wire n_490;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_1026;
wire n_492;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1194;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_943;
wire n_977;
wire n_905;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_816;
wire n_625;
wire n_953;
wire n_1373;
wire n_716;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_1207;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_561;
wire n_437;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_563;
wire n_891;
wire n_568;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_1083;
wire n_727;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_1139;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1127;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_1355;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1164;
wire n_433;
wire n_627;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_559;
wire n_1049;
wire n_466;
wire n_1277;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_924;
wire n_1264;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_425;
wire n_879;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_1183;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_1390;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1352;
wire n_729;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_1236;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_0), .A2(n_117), .B1(n_612), .B2(n_702), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_1), .A2(n_401), .B1(n_797), .B2(n_933), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_2), .A2(n_162), .B1(n_648), .B2(n_654), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g1358 ( .A1(n_3), .A2(n_332), .B1(n_485), .B2(n_782), .Y(n_1358) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_4), .A2(n_268), .B1(n_656), .B2(n_657), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_5), .B(n_569), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_6), .A2(n_210), .B1(n_496), .B2(n_500), .Y(n_615) );
CKINVDCx5p33_ASAP7_75t_R g690 ( .A(n_7), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_8), .A2(n_379), .B1(n_631), .B2(n_856), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_9), .A2(n_380), .B1(n_516), .B2(n_1066), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1385 ( .A1(n_10), .A2(n_324), .B1(n_1386), .B2(n_1387), .Y(n_1385) );
AO22x1_ASAP7_75t_L g835 ( .A1(n_11), .A2(n_214), .B1(n_836), .B2(n_837), .Y(n_835) );
INVx1_ASAP7_75t_L g1366 ( .A(n_12), .Y(n_1366) );
AOI221xp5_ASAP7_75t_L g803 ( .A1(n_13), .A2(n_343), .B1(n_804), .B2(n_805), .C(n_806), .Y(n_803) );
INVx1_ASAP7_75t_SL g1218 ( .A(n_14), .Y(n_1218) );
AOI22xp5_ASAP7_75t_L g1062 ( .A1(n_15), .A2(n_98), .B1(n_998), .B2(n_1063), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_16), .A2(n_250), .B1(n_444), .B2(n_701), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_17), .A2(n_231), .B1(n_656), .B2(n_657), .Y(n_975) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_18), .B(n_451), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_19), .A2(n_355), .B1(n_481), .B2(n_485), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g1125 ( .A(n_20), .Y(n_1125) );
AOI22xp33_ASAP7_75t_L g1020 ( .A1(n_21), .A2(n_224), .B1(n_612), .B2(n_613), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_22), .A2(n_319), .B1(n_506), .B2(n_687), .Y(n_810) );
AOI22xp33_ASAP7_75t_SL g1007 ( .A1(n_23), .A2(n_194), .B1(n_612), .B2(n_613), .Y(n_1007) );
AOI22xp5_ASAP7_75t_L g1355 ( .A1(n_24), .A2(n_406), .B1(n_444), .B2(n_773), .Y(n_1355) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_25), .A2(n_106), .B1(n_496), .B2(n_556), .Y(n_820) );
INVx1_ASAP7_75t_SL g759 ( .A(n_26), .Y(n_759) );
INVx1_ASAP7_75t_L g860 ( .A(n_27), .Y(n_860) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_28), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g1158 ( .A1(n_29), .A2(n_103), .B1(n_1112), .B2(n_1134), .Y(n_1158) );
INVx1_ASAP7_75t_L g929 ( .A(n_30), .Y(n_929) );
AOI22xp5_ASAP7_75t_L g1069 ( .A1(n_31), .A2(n_394), .B1(n_492), .B2(n_797), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_32), .A2(n_145), .B1(n_513), .B2(n_516), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_33), .A2(n_43), .B1(n_653), .B2(n_654), .Y(n_652) );
INVx1_ASAP7_75t_L g1050 ( .A(n_34), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_35), .A2(n_160), .B1(n_496), .B2(n_500), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_36), .A2(n_263), .B1(n_593), .B2(n_594), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_37), .A2(n_76), .B1(n_555), .B2(n_556), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_38), .B(n_660), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_39), .A2(n_342), .B1(n_1025), .B2(n_1026), .Y(n_1024) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_40), .A2(n_182), .B1(n_559), .B2(n_613), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_41), .A2(n_206), .B1(n_556), .B2(n_801), .Y(n_800) );
AOI221xp5_ASAP7_75t_L g916 ( .A1(n_42), .A2(n_397), .B1(n_591), .B2(n_662), .C(n_917), .Y(n_916) );
AOI21xp33_ASAP7_75t_L g873 ( .A1(n_44), .A2(n_660), .B(n_874), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_45), .A2(n_67), .B1(n_566), .B2(n_567), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g954 ( .A1(n_46), .A2(n_955), .B(n_957), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g1220 ( .A1(n_47), .A2(n_279), .B1(n_1152), .B2(n_1155), .Y(n_1220) );
INVx1_ASAP7_75t_L g972 ( .A(n_48), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_49), .A2(n_120), .B1(n_481), .B2(n_598), .Y(n_1043) );
AOI22xp5_ASAP7_75t_L g878 ( .A1(n_50), .A2(n_395), .B1(n_585), .B2(n_879), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_51), .A2(n_248), .B1(n_540), .B2(n_687), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_52), .A2(n_110), .B1(n_594), .B2(n_668), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_53), .A2(n_62), .B1(n_687), .B2(n_872), .Y(n_1055) );
AOI22xp33_ASAP7_75t_SL g1008 ( .A1(n_54), .A2(n_300), .B1(n_481), .B2(n_485), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_55), .A2(n_183), .B1(n_445), .B2(n_563), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_56), .A2(n_403), .B1(n_650), .B2(n_651), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_57), .A2(n_153), .B1(n_485), .B2(n_492), .Y(n_817) );
INVx1_ASAP7_75t_L g1121 ( .A(n_58), .Y(n_1121) );
AOI22x1_ASAP7_75t_L g1350 ( .A1(n_58), .A2(n_1121), .B1(n_1351), .B2(n_1352), .Y(n_1350) );
AOI22xp33_ASAP7_75t_L g1372 ( .A1(n_58), .A2(n_1373), .B1(n_1402), .B2(n_1404), .Y(n_1372) );
AO22x1_ASAP7_75t_L g917 ( .A1(n_59), .A2(n_81), .B1(n_594), .B2(n_602), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_60), .A2(n_289), .B1(n_566), .B2(n_863), .Y(n_926) );
CKINVDCx20_ASAP7_75t_R g580 ( .A(n_61), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_63), .A2(n_350), .B1(n_591), .B2(n_594), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g1394 ( .A(n_64), .B(n_688), .Y(n_1394) );
NAND2xp5_ASAP7_75t_L g1035 ( .A(n_65), .B(n_1036), .Y(n_1035) );
OA22x2_ASAP7_75t_L g457 ( .A1(n_66), .A2(n_172), .B1(n_451), .B2(n_455), .Y(n_457) );
INVx1_ASAP7_75t_L g477 ( .A(n_66), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_68), .A2(n_140), .B1(n_612), .B2(n_613), .Y(n_611) );
AOI221xp5_ASAP7_75t_L g822 ( .A1(n_69), .A2(n_78), .B1(n_569), .B2(n_823), .C(n_824), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_70), .A2(n_356), .B1(n_556), .B2(n_801), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1017 ( .A1(n_71), .A2(n_364), .B1(n_481), .B2(n_485), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_72), .A2(n_329), .B1(n_528), .B2(n_626), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_73), .A2(n_388), .B1(n_716), .B2(n_718), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_74), .A2(n_158), .B1(n_492), .B2(n_552), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_75), .A2(n_382), .B1(n_591), .B2(n_594), .Y(n_968) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_77), .B(n_196), .Y(n_432) );
INVx1_ASAP7_75t_L g454 ( .A(n_77), .Y(n_454) );
OAI21xp33_ASAP7_75t_L g478 ( .A1(n_77), .A2(n_172), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g883 ( .A(n_79), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g1086 ( .A1(n_80), .A2(n_203), .B1(n_509), .B2(n_863), .Y(n_1086) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_82), .A2(n_114), .B1(n_445), .B2(n_563), .Y(n_1070) );
INVx1_ASAP7_75t_L g944 ( .A(n_83), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g1395 ( .A1(n_84), .A2(n_187), .B1(n_692), .B2(n_1396), .Y(n_1395) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_85), .A2(n_244), .B1(n_647), .B2(n_653), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g1354 ( .A1(n_86), .A2(n_373), .B1(n_708), .B2(n_711), .Y(n_1354) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_87), .A2(n_271), .B1(n_647), .B2(n_648), .Y(n_646) );
INVx1_ASAP7_75t_SL g779 ( .A(n_88), .Y(n_779) );
INVx1_ASAP7_75t_L g992 ( .A(n_89), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_90), .A2(n_178), .B1(n_656), .B2(n_657), .Y(n_655) );
AOI21xp33_ASAP7_75t_L g663 ( .A1(n_91), .A2(n_593), .B(n_664), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_92), .A2(n_94), .B1(n_559), .B2(n_705), .Y(n_1042) );
INVx1_ASAP7_75t_L g1114 ( .A(n_93), .Y(n_1114) );
AND2x4_ASAP7_75t_L g1124 ( .A(n_93), .B(n_317), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_95), .A2(n_105), .B1(n_630), .B2(n_631), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_96), .A2(n_235), .B1(n_559), .B2(n_937), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_97), .A2(n_102), .B1(n_650), .B2(n_651), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_99), .A2(n_272), .B1(n_516), .B2(n_804), .Y(n_953) );
AOI21xp33_ASAP7_75t_L g970 ( .A1(n_100), .A2(n_602), .B(n_971), .Y(n_970) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_101), .A2(n_620), .B(n_621), .Y(n_619) );
XOR2xp5_ASAP7_75t_L g1039 ( .A(n_103), .B(n_1040), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_104), .A2(n_124), .B1(n_653), .B2(n_654), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_107), .A2(n_167), .B1(n_496), .B2(n_733), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_108), .A2(n_173), .B1(n_567), .B2(n_591), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_109), .A2(n_265), .B1(n_489), .B2(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g891 ( .A(n_111), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g1357 ( .A1(n_112), .A2(n_189), .B1(n_489), .B2(n_702), .Y(n_1357) );
INVx1_ASAP7_75t_SL g754 ( .A(n_113), .Y(n_754) );
INVx1_ASAP7_75t_L g578 ( .A(n_115), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g947 ( .A1(n_116), .A2(n_294), .B1(n_496), .B2(n_500), .Y(n_947) );
INVx1_ASAP7_75t_SL g761 ( .A(n_118), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_119), .A2(n_146), .B1(n_559), .B2(n_560), .Y(n_558) );
INVx1_ASAP7_75t_SL g1115 ( .A(n_121), .Y(n_1115) );
AND2x4_ASAP7_75t_L g1118 ( .A(n_121), .B(n_428), .Y(n_1118) );
INVx1_ASAP7_75t_L g1129 ( .A(n_121), .Y(n_1129) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_122), .A2(n_412), .B1(n_555), .B2(n_556), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_123), .A2(n_126), .B1(n_445), .B2(n_563), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g1362 ( .A1(n_125), .A2(n_128), .B1(n_630), .B2(n_631), .Y(n_1362) );
INVx1_ASAP7_75t_L g985 ( .A(n_127), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_129), .A2(n_390), .B1(n_506), .B2(n_509), .Y(n_505) );
CKINVDCx16_ASAP7_75t_R g938 ( .A(n_130), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g1179 ( .A1(n_131), .A2(n_157), .B1(n_1142), .B2(n_1180), .Y(n_1179) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_132), .A2(n_308), .B1(n_687), .B2(n_688), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_133), .A2(n_353), .B1(n_591), .B2(n_662), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_134), .A2(n_168), .B1(n_444), .B2(n_470), .Y(n_443) );
XNOR2x1_ASAP7_75t_L g964 ( .A(n_135), .B(n_965), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_136), .B(n_804), .Y(n_869) );
INVx1_ASAP7_75t_L g1116 ( .A(n_137), .Y(n_1116) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_138), .A2(n_266), .B1(n_585), .B2(n_587), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_139), .A2(n_322), .B1(n_630), .B2(n_631), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_141), .A2(n_361), .B1(n_506), .B2(n_626), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_142), .A2(n_177), .B1(n_492), .B2(n_559), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g976 ( .A1(n_143), .A2(n_184), .B1(n_651), .B2(n_653), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g1382 ( .A1(n_144), .A2(n_396), .B1(n_1383), .B2(n_1384), .Y(n_1382) );
INVx1_ASAP7_75t_L g1392 ( .A(n_147), .Y(n_1392) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_148), .B(n_857), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_149), .A2(n_400), .B1(n_688), .B2(n_1000), .Y(n_999) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_150), .A2(n_407), .B1(n_489), .B2(n_492), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_151), .A2(n_311), .B1(n_708), .B2(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g849 ( .A(n_152), .Y(n_849) );
INVx1_ASAP7_75t_L g753 ( .A(n_154), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_155), .A2(n_190), .B1(n_445), .B2(n_589), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_156), .A2(n_197), .B1(n_562), .B2(n_563), .Y(n_561) );
INVxp67_ASAP7_75t_SL g1013 ( .A(n_157), .Y(n_1013) );
AOI22xp5_ASAP7_75t_L g1379 ( .A1(n_159), .A2(n_262), .B1(n_773), .B2(n_1380), .Y(n_1379) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_161), .A2(n_415), .B1(n_489), .B2(n_492), .Y(n_1018) );
INVx1_ASAP7_75t_L g665 ( .A(n_163), .Y(n_665) );
XNOR2x1_ASAP7_75t_L g440 ( .A(n_164), .B(n_441), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_165), .A2(n_304), .B1(n_492), .B2(n_559), .Y(n_798) );
INVx1_ASAP7_75t_L g958 ( .A(n_166), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_169), .A2(n_188), .B1(n_496), .B2(n_1005), .Y(n_1019) );
CKINVDCx6p67_ASAP7_75t_R g1148 ( .A(n_170), .Y(n_1148) );
INVx1_ASAP7_75t_L g469 ( .A(n_171), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_171), .B(n_245), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_171), .B(n_475), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_172), .B(n_337), .Y(n_431) );
AOI22xp33_ASAP7_75t_SL g1003 ( .A1(n_174), .A2(n_216), .B1(n_489), .B2(n_782), .Y(n_1003) );
AOI22xp33_ASAP7_75t_SL g888 ( .A1(n_175), .A2(n_347), .B1(n_593), .B2(n_662), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_176), .A2(n_181), .B1(n_509), .B2(n_528), .Y(n_828) );
AOI21xp33_ASAP7_75t_L g1048 ( .A1(n_179), .A2(n_857), .B(n_1049), .Y(n_1048) );
XNOR2x1_ASAP7_75t_L g581 ( .A(n_180), .B(n_582), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_185), .A2(n_320), .B1(n_509), .B2(n_739), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g1135 ( .A1(n_186), .A2(n_387), .B1(n_1123), .B2(n_1127), .Y(n_1135) );
NAND2xp5_ASAP7_75t_L g1089 ( .A(n_191), .B(n_569), .Y(n_1089) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_192), .A2(n_419), .B1(n_506), .B2(n_631), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g961 ( .A(n_193), .B(n_688), .Y(n_961) );
AOI22xp5_ASAP7_75t_L g1052 ( .A1(n_195), .A2(n_234), .B1(n_555), .B2(n_556), .Y(n_1052) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_196), .B(n_461), .Y(n_460) );
AOI22xp33_ASAP7_75t_SL g881 ( .A1(n_198), .A2(n_385), .B1(n_555), .B2(n_840), .Y(n_881) );
AOI22xp5_ASAP7_75t_L g880 ( .A1(n_199), .A2(n_392), .B1(n_562), .B2(n_597), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_200), .A2(n_236), .B1(n_516), .B2(n_925), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_201), .B(n_628), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g877 ( .A1(n_202), .A2(n_358), .B1(n_598), .B2(n_705), .Y(n_877) );
AOI22xp5_ASAP7_75t_L g1004 ( .A1(n_204), .A2(n_297), .B1(n_708), .B2(n_1005), .Y(n_1004) );
AOI22xp5_ASAP7_75t_L g1159 ( .A1(n_205), .A2(n_344), .B1(n_1123), .B2(n_1127), .Y(n_1159) );
INVx1_ASAP7_75t_L g1045 ( .A(n_207), .Y(n_1045) );
INVx1_ASAP7_75t_L g526 ( .A(n_208), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_209), .A2(n_313), .B1(n_597), .B2(n_598), .Y(n_596) );
AOI21xp33_ASAP7_75t_SL g576 ( .A1(n_211), .A2(n_506), .B(n_577), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_212), .A2(n_368), .B1(n_445), .B2(n_589), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_213), .A2(n_301), .B1(n_566), .B2(n_863), .Y(n_1067) );
XNOR2x1_ASAP7_75t_L g981 ( .A(n_215), .B(n_982), .Y(n_981) );
INVx1_ASAP7_75t_L g1150 ( .A(n_217), .Y(n_1150) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_218), .A2(n_416), .B1(n_559), .B2(n_933), .Y(n_1087) );
INVx1_ASAP7_75t_L g990 ( .A(n_219), .Y(n_990) );
AOI22xp5_ASAP7_75t_L g1093 ( .A1(n_220), .A2(n_278), .B1(n_575), .B2(n_693), .Y(n_1093) );
INVx1_ASAP7_75t_SL g764 ( .A(n_221), .Y(n_764) );
INVx1_ASAP7_75t_L g669 ( .A(n_222), .Y(n_669) );
OA22x2_ASAP7_75t_L g906 ( .A1(n_223), .A2(n_907), .B1(n_918), .B2(n_919), .Y(n_906) );
INVx1_ASAP7_75t_L g919 ( .A(n_223), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g1141 ( .A1(n_223), .A2(n_359), .B1(n_1142), .B2(n_1143), .Y(n_1141) );
INVx1_ASAP7_75t_L g751 ( .A(n_225), .Y(n_751) );
AOI21xp33_ASAP7_75t_SL g1090 ( .A1(n_226), .A2(n_506), .B(n_1091), .Y(n_1090) );
INVx1_ASAP7_75t_L g996 ( .A(n_227), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_228), .A2(n_393), .B1(n_489), .B2(n_492), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_229), .A2(n_417), .B1(n_566), .B2(n_863), .Y(n_870) );
INVx1_ASAP7_75t_L g854 ( .A(n_230), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g1381 ( .A1(n_232), .A2(n_292), .B1(n_704), .B2(n_845), .Y(n_1381) );
AOI21xp33_ASAP7_75t_L g889 ( .A1(n_233), .A2(n_668), .B(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g1059 ( .A(n_237), .Y(n_1059) );
AOI22xp5_ASAP7_75t_L g1133 ( .A1(n_237), .A2(n_399), .B1(n_1112), .B2(n_1134), .Y(n_1133) );
AOI22xp33_ASAP7_75t_L g1178 ( .A1(n_238), .A2(n_331), .B1(n_1139), .B2(n_1155), .Y(n_1178) );
AOI22xp5_ASAP7_75t_L g772 ( .A1(n_239), .A2(n_351), .B1(n_773), .B2(n_775), .Y(n_772) );
INVx1_ASAP7_75t_L g850 ( .A(n_240), .Y(n_850) );
AOI221xp5_ASAP7_75t_L g1363 ( .A1(n_241), .A2(n_402), .B1(n_620), .B2(n_1364), .C(n_1365), .Y(n_1363) );
AOI21x1_ASAP7_75t_SL g519 ( .A1(n_242), .A2(n_520), .B(n_525), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_243), .A2(n_299), .B1(n_573), .B2(n_575), .Y(n_572) );
INVx1_ASAP7_75t_L g452 ( .A(n_245), .Y(n_452) );
OAI22x1_ASAP7_75t_L g608 ( .A1(n_246), .A2(n_609), .B1(n_616), .B2(n_632), .Y(n_608) );
NAND5xp2_ASAP7_75t_SL g609 ( .A(n_246), .B(n_610), .C(n_611), .D(n_614), .E(n_615), .Y(n_609) );
INVx1_ASAP7_75t_L g683 ( .A(n_247), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g1028 ( .A1(n_249), .A2(n_1029), .B(n_1031), .Y(n_1028) );
AOI22xp5_ASAP7_75t_L g769 ( .A1(n_251), .A2(n_298), .B1(n_613), .B2(n_770), .Y(n_769) );
AOI22xp5_ASAP7_75t_L g909 ( .A1(n_252), .A2(n_418), .B1(n_650), .B2(n_651), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_253), .A2(n_374), .B1(n_697), .B2(n_872), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_254), .A2(n_276), .B1(n_1139), .B2(n_1140), .Y(n_1138) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_255), .A2(n_409), .B1(n_489), .B2(n_492), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_256), .A2(n_264), .B1(n_540), .B2(n_687), .Y(n_766) );
INVx1_ASAP7_75t_L g694 ( .A(n_257), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_258), .A2(n_286), .B1(n_656), .B2(n_657), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_259), .A2(n_303), .B1(n_481), .B2(n_485), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g1053 ( .A1(n_260), .A2(n_383), .B1(n_562), .B2(n_702), .Y(n_1053) );
INVx1_ASAP7_75t_L g538 ( .A(n_261), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_267), .A2(n_410), .B1(n_647), .B2(n_648), .Y(n_893) );
AOI22xp5_ASAP7_75t_L g912 ( .A1(n_269), .A2(n_372), .B1(n_648), .B2(n_654), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_270), .A2(n_280), .B1(n_827), .B2(n_863), .Y(n_862) );
XNOR2x1_ASAP7_75t_L g866 ( .A(n_273), .B(n_867), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_274), .A2(n_275), .B1(n_496), .B2(n_500), .Y(n_1082) );
XOR2x2_ASAP7_75t_L g832 ( .A(n_277), .B(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g825 ( .A(n_281), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_282), .A2(n_291), .B1(n_647), .B2(n_662), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_283), .A2(n_411), .B1(n_708), .B2(n_711), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g1083 ( .A1(n_284), .A2(n_321), .B1(n_481), .B2(n_1084), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_285), .A2(n_404), .B1(n_566), .B2(n_575), .Y(n_1056) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_287), .A2(n_377), .B1(n_516), .B2(n_812), .Y(n_811) );
XNOR2xp5_ASAP7_75t_L g1079 ( .A(n_288), .B(n_1080), .Y(n_1079) );
AOI22xp33_ASAP7_75t_L g1164 ( .A1(n_288), .A2(n_314), .B1(n_1142), .B2(n_1143), .Y(n_1164) );
INVx1_ASAP7_75t_SL g787 ( .A(n_290), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_293), .A2(n_318), .B1(n_563), .B2(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g604 ( .A(n_295), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_296), .B(n_569), .Y(n_568) );
AOI221xp5_ASAP7_75t_SL g913 ( .A1(n_302), .A2(n_365), .B1(n_593), .B2(n_857), .C(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g726 ( .A(n_305), .Y(n_726) );
INVx1_ASAP7_75t_L g846 ( .A(n_306), .Y(n_846) );
AOI22xp5_ASAP7_75t_L g1072 ( .A1(n_307), .A2(n_413), .B1(n_559), .B2(n_1073), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_309), .A2(n_330), .B1(n_481), .B2(n_485), .Y(n_948) );
INVx1_ASAP7_75t_L g721 ( .A(n_310), .Y(n_721) );
CKINVDCx5p33_ASAP7_75t_R g679 ( .A(n_312), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g1163 ( .A1(n_315), .A2(n_346), .B1(n_1140), .B2(n_1152), .Y(n_1163) );
AOI22xp33_ASAP7_75t_SL g1397 ( .A1(n_316), .A2(n_352), .B1(n_1398), .B2(n_1399), .Y(n_1397) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_317), .Y(n_433) );
AND2x4_ASAP7_75t_L g1113 ( .A(n_317), .B(n_1114), .Y(n_1113) );
CKINVDCx5p33_ASAP7_75t_R g677 ( .A(n_323), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_325), .A2(n_345), .B1(n_485), .B2(n_563), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g1360 ( .A1(n_326), .A2(n_384), .B1(n_852), .B2(n_1361), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_327), .B(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g843 ( .A(n_328), .Y(n_843) );
INVx1_ASAP7_75t_L g858 ( .A(n_333), .Y(n_858) );
AOI22xp5_ASAP7_75t_L g1094 ( .A1(n_334), .A2(n_366), .B1(n_445), .B2(n_937), .Y(n_1094) );
INVx1_ASAP7_75t_L g807 ( .A(n_335), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_336), .A2(n_340), .B1(n_444), .B2(n_470), .Y(n_841) );
INVx1_ASAP7_75t_L g467 ( .A(n_337), .Y(n_467) );
INVxp67_ASAP7_75t_L g537 ( .A(n_337), .Y(n_537) );
INVx1_ASAP7_75t_L g1092 ( .A(n_338), .Y(n_1092) );
AOI22xp33_ASAP7_75t_SL g1374 ( .A1(n_339), .A2(n_1375), .B1(n_1376), .B2(n_1401), .Y(n_1374) );
INVx1_ASAP7_75t_L g1401 ( .A(n_339), .Y(n_1401) );
NAND2xp5_ASAP7_75t_L g1064 ( .A(n_341), .B(n_823), .Y(n_1064) );
INVxp67_ASAP7_75t_R g1153 ( .A(n_348), .Y(n_1153) );
INVx2_ASAP7_75t_L g428 ( .A(n_349), .Y(n_428) );
INVx1_ASAP7_75t_L g875 ( .A(n_354), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_357), .A2(n_370), .B1(n_612), .B2(n_937), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_360), .A2(n_398), .B1(n_556), .B2(n_801), .Y(n_935) );
AOI221xp5_ASAP7_75t_L g599 ( .A1(n_362), .A2(n_386), .B1(n_573), .B2(n_600), .C(n_603), .Y(n_599) );
INVx1_ASAP7_75t_SL g780 ( .A(n_363), .Y(n_780) );
CKINVDCx5p33_ASAP7_75t_R g915 ( .A(n_367), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_369), .B(n_743), .Y(n_886) );
INVx1_ASAP7_75t_L g814 ( .A(n_371), .Y(n_814) );
INVx1_ASAP7_75t_L g1034 ( .A(n_375), .Y(n_1034) );
AOI21xp33_ASAP7_75t_SL g1389 ( .A1(n_376), .A2(n_1390), .B(n_1391), .Y(n_1389) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_378), .A2(n_414), .B1(n_593), .B2(n_650), .Y(n_974) );
INVx1_ASAP7_75t_L g622 ( .A(n_381), .Y(n_622) );
INVx1_ASAP7_75t_L g1119 ( .A(n_389), .Y(n_1119) );
INVx1_ASAP7_75t_L g987 ( .A(n_391), .Y(n_987) );
CKINVDCx5p33_ASAP7_75t_R g784 ( .A(n_405), .Y(n_784) );
INVx1_ASAP7_75t_L g1219 ( .A(n_408), .Y(n_1219) );
XNOR2x1_ASAP7_75t_L g793 ( .A(n_420), .B(n_794), .Y(n_793) );
AOI21xp33_ASAP7_75t_L g927 ( .A1(n_421), .A2(n_739), .B(n_928), .Y(n_927) );
AOI21xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_434), .B(n_1100), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
BUFx4_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
NAND3xp33_ASAP7_75t_L g425 ( .A(n_426), .B(n_429), .C(n_433), .Y(n_425) );
AND2x2_ASAP7_75t_L g1369 ( .A(n_426), .B(n_1370), .Y(n_1369) );
AND2x2_ASAP7_75t_L g1403 ( .A(n_426), .B(n_1371), .Y(n_1403) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OA21x2_ASAP7_75t_L g1405 ( .A1(n_427), .A2(n_1115), .B(n_1406), .Y(n_1405) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND3x4_ASAP7_75t_L g1112 ( .A(n_428), .B(n_1113), .C(n_1115), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_428), .B(n_1129), .Y(n_1128) );
NOR2xp33_ASAP7_75t_L g1370 ( .A(n_429), .B(n_1371), .Y(n_1370) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AO21x2_ASAP7_75t_L g542 ( .A1(n_430), .A2(n_543), .B(n_544), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx1_ASAP7_75t_L g1371 ( .A(n_433), .Y(n_1371) );
XNOR2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_901), .Y(n_434) );
XNOR2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_722), .Y(n_435) );
XOR2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_639), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_546), .B1(n_636), .B2(n_637), .Y(n_437) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx3_ASAP7_75t_L g638 ( .A(n_440), .Y(n_638) );
NAND4xp75_ASAP7_75t_SL g441 ( .A(n_442), .B(n_487), .C(n_504), .D(n_519), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_480), .Y(n_442) );
BUFx12f_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g771 ( .A(n_445), .Y(n_771) );
BUFx6f_ASAP7_75t_L g1386 ( .A(n_445), .Y(n_1386) );
BUFx12f_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_446), .Y(n_562) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_446), .Y(n_612) );
AND2x4_ASAP7_75t_L g446 ( .A(n_447), .B(n_458), .Y(n_446) );
AND2x4_ASAP7_75t_L g482 ( .A(n_447), .B(n_483), .Y(n_482) );
AND2x4_ASAP7_75t_L g497 ( .A(n_447), .B(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g501 ( .A(n_447), .B(n_502), .Y(n_501) );
AND2x4_ASAP7_75t_L g647 ( .A(n_447), .B(n_494), .Y(n_647) );
AND2x4_ASAP7_75t_L g653 ( .A(n_447), .B(n_458), .Y(n_653) );
AND2x4_ASAP7_75t_L g656 ( .A(n_447), .B(n_498), .Y(n_656) );
AND2x4_ASAP7_75t_L g657 ( .A(n_447), .B(n_502), .Y(n_657) );
AND2x4_ASAP7_75t_L g447 ( .A(n_448), .B(n_456), .Y(n_447) );
AND2x2_ASAP7_75t_L g508 ( .A(n_448), .B(n_457), .Y(n_508) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g491 ( .A(n_449), .B(n_457), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_453), .Y(n_449) );
NAND2xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
INVx2_ASAP7_75t_L g455 ( .A(n_451), .Y(n_455) );
INVx3_ASAP7_75t_L g461 ( .A(n_451), .Y(n_461) );
NAND2xp33_ASAP7_75t_L g468 ( .A(n_451), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g479 ( .A(n_451), .Y(n_479) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_451), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_452), .B(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
OAI21xp5_ASAP7_75t_L g536 ( .A1(n_454), .A2(n_479), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g535 ( .A(n_457), .B(n_536), .Y(n_535) );
AND2x4_ASAP7_75t_L g472 ( .A(n_458), .B(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g490 ( .A(n_458), .B(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g586 ( .A(n_458), .B(n_491), .Y(n_586) );
AND2x4_ASAP7_75t_L g650 ( .A(n_458), .B(n_491), .Y(n_650) );
AND2x4_ASAP7_75t_L g654 ( .A(n_458), .B(n_473), .Y(n_654) );
AND2x4_ASAP7_75t_L g458 ( .A(n_459), .B(n_463), .Y(n_458) );
OR2x2_ASAP7_75t_L g484 ( .A(n_459), .B(n_464), .Y(n_484) );
AND2x4_ASAP7_75t_L g498 ( .A(n_459), .B(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g503 ( .A(n_459), .Y(n_503) );
AND2x2_ASAP7_75t_L g531 ( .A(n_459), .B(n_532), .Y(n_531) );
AND2x4_ASAP7_75t_L g459 ( .A(n_460), .B(n_462), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_461), .B(n_467), .Y(n_466) );
INVxp67_ASAP7_75t_L g475 ( .A(n_461), .Y(n_475) );
NAND3xp33_ASAP7_75t_L g544 ( .A(n_462), .B(n_474), .C(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g499 ( .A(n_465), .Y(n_499) );
AND2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_468), .Y(n_465) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g560 ( .A(n_471), .Y(n_560) );
INVx2_ASAP7_75t_SL g589 ( .A(n_471), .Y(n_589) );
INVx4_ASAP7_75t_L g613 ( .A(n_471), .Y(n_613) );
INVx4_ASAP7_75t_L g702 ( .A(n_471), .Y(n_702) );
INVx2_ASAP7_75t_L g879 ( .A(n_471), .Y(n_879) );
INVx4_ASAP7_75t_L g937 ( .A(n_471), .Y(n_937) );
INVx2_ASAP7_75t_L g1073 ( .A(n_471), .Y(n_1073) );
INVx8_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x4_ASAP7_75t_L g486 ( .A(n_473), .B(n_483), .Y(n_486) );
AND2x4_ASAP7_75t_L g518 ( .A(n_473), .B(n_502), .Y(n_518) );
AND2x4_ASAP7_75t_L g594 ( .A(n_473), .B(n_502), .Y(n_594) );
AND2x4_ASAP7_75t_L g648 ( .A(n_473), .B(n_483), .Y(n_648) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_478), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
BUFx6f_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_482), .Y(n_563) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_482), .Y(n_597) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_482), .Y(n_717) );
AND2x4_ASAP7_75t_L g651 ( .A(n_483), .B(n_491), .Y(n_651) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g494 ( .A(n_484), .Y(n_494) );
BUFx3_ASAP7_75t_L g1380 ( .A(n_485), .Y(n_1380) );
BUFx12f_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx6_ASAP7_75t_L g553 ( .A(n_486), .Y(n_553) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_495), .Y(n_487) );
BUFx8_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_490), .Y(n_559) );
AND2x4_ASAP7_75t_L g493 ( .A(n_491), .B(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g511 ( .A(n_491), .B(n_498), .Y(n_511) );
AND2x2_ASAP7_75t_L g524 ( .A(n_491), .B(n_502), .Y(n_524) );
AND2x4_ASAP7_75t_L g591 ( .A(n_491), .B(n_498), .Y(n_591) );
AND2x2_ASAP7_75t_L g602 ( .A(n_491), .B(n_502), .Y(n_602) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_493), .Y(n_587) );
BUFx12f_ASAP7_75t_L g705 ( .A(n_493), .Y(n_705) );
BUFx3_ASAP7_75t_L g782 ( .A(n_493), .Y(n_782) );
BUFx6f_ASAP7_75t_L g933 ( .A(n_493), .Y(n_933) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx12f_ASAP7_75t_L g555 ( .A(n_497), .Y(n_555) );
INVx3_ASAP7_75t_L g710 ( .A(n_497), .Y(n_710) );
AND2x4_ASAP7_75t_L g507 ( .A(n_498), .B(n_508), .Y(n_507) );
AND2x4_ASAP7_75t_L g593 ( .A(n_498), .B(n_508), .Y(n_593) );
AND2x4_ASAP7_75t_L g502 ( .A(n_499), .B(n_503), .Y(n_502) );
BUFx5_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_501), .Y(n_556) );
INVx1_ASAP7_75t_L g714 ( .A(n_501), .Y(n_714) );
BUFx3_ASAP7_75t_L g840 ( .A(n_501), .Y(n_840) );
AND2x4_ASAP7_75t_L g515 ( .A(n_502), .B(n_508), .Y(n_515) );
AND2x2_ASAP7_75t_L g668 ( .A(n_502), .B(n_508), .Y(n_668) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_512), .Y(n_504) );
INVx4_ASAP7_75t_L g678 ( .A(n_506), .Y(n_678) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
BUFx3_ASAP7_75t_L g620 ( .A(n_507), .Y(n_620) );
INVx1_ASAP7_75t_L g740 ( .A(n_507), .Y(n_740) );
BUFx3_ASAP7_75t_L g872 ( .A(n_507), .Y(n_872) );
INVx2_ASAP7_75t_L g988 ( .A(n_509), .Y(n_988) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
BUFx6f_ASAP7_75t_L g757 ( .A(n_510), .Y(n_757) );
INVx2_ASAP7_75t_L g1027 ( .A(n_510), .Y(n_1027) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_511), .Y(n_566) );
BUFx3_ASAP7_75t_L g626 ( .A(n_511), .Y(n_626) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx3_ASAP7_75t_L g823 ( .A(n_514), .Y(n_823) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g574 ( .A(n_515), .Y(n_574) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_515), .Y(n_693) );
BUFx8_ASAP7_75t_SL g804 ( .A(n_515), .Y(n_804) );
BUFx6f_ASAP7_75t_L g857 ( .A(n_515), .Y(n_857) );
BUFx3_ASAP7_75t_L g925 ( .A(n_515), .Y(n_925) );
INVx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g575 ( .A(n_517), .Y(n_575) );
INVx2_ASAP7_75t_L g994 ( .A(n_517), .Y(n_994) );
INVx3_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_518), .Y(n_631) );
BUFx6f_ASAP7_75t_L g697 ( .A(n_518), .Y(n_697) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g628 ( .A(n_522), .Y(n_628) );
INVx2_ASAP7_75t_L g685 ( .A(n_522), .Y(n_685) );
INVx2_ASAP7_75t_L g1047 ( .A(n_522), .Y(n_1047) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g743 ( .A(n_523), .Y(n_743) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx3_ASAP7_75t_L g570 ( .A(n_524), .Y(n_570) );
BUFx3_ASAP7_75t_L g660 ( .A(n_524), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_527), .B1(n_538), .B2(n_539), .Y(n_525) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g567 ( .A(n_529), .Y(n_567) );
INVx4_ASAP7_75t_L g687 ( .A(n_529), .Y(n_687) );
INVx3_ASAP7_75t_L g1361 ( .A(n_529), .Y(n_1361) );
INVx5_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx2_ASAP7_75t_L g863 ( .A(n_530), .Y(n_863) );
BUFx4f_ASAP7_75t_L g1000 ( .A(n_530), .Y(n_1000) );
BUFx2_ASAP7_75t_L g1033 ( .A(n_530), .Y(n_1033) );
AND2x4_ASAP7_75t_L g530 ( .A(n_531), .B(n_535), .Y(n_530) );
AND2x2_ASAP7_75t_L g662 ( .A(n_531), .B(n_535), .Y(n_662) );
AND2x4_ASAP7_75t_L g960 ( .A(n_531), .B(n_535), .Y(n_960) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
INVx1_ASAP7_75t_L g543 ( .A(n_533), .Y(n_543) );
INVx2_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
BUFx6f_ASAP7_75t_L g579 ( .A(n_541), .Y(n_579) );
BUFx6f_ASAP7_75t_L g605 ( .A(n_541), .Y(n_605) );
INVx2_ASAP7_75t_L g809 ( .A(n_541), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g914 ( .A(n_541), .B(n_915), .Y(n_914) );
INVx1_ASAP7_75t_L g1063 ( .A(n_541), .Y(n_1063) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx3_ASAP7_75t_L g624 ( .A(n_542), .Y(n_624) );
INVx2_ASAP7_75t_L g636 ( .A(n_546), .Y(n_636) );
XNOR2x1_ASAP7_75t_L g546 ( .A(n_547), .B(n_607), .Y(n_546) );
XNOR2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_581), .Y(n_547) );
XNOR2x1_ASAP7_75t_L g548 ( .A(n_549), .B(n_580), .Y(n_548) );
NOR4xp75_ASAP7_75t_L g549 ( .A(n_550), .B(n_557), .C(n_564), .D(n_571), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_554), .Y(n_550) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx5_ASAP7_75t_L g598 ( .A(n_553), .Y(n_598) );
INVx2_ASAP7_75t_L g720 ( .A(n_553), .Y(n_720) );
INVx3_ASAP7_75t_L g797 ( .A(n_553), .Y(n_797) );
INVx1_ASAP7_75t_L g1084 ( .A(n_553), .Y(n_1084) );
HB1xp67_ASAP7_75t_L g786 ( .A(n_555), .Y(n_786) );
INVx1_ASAP7_75t_L g788 ( .A(n_556), .Y(n_788) );
BUFx2_ASAP7_75t_SL g1384 ( .A(n_556), .Y(n_1384) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_561), .Y(n_557) );
BUFx3_ASAP7_75t_L g778 ( .A(n_559), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_568), .Y(n_564) );
INVx1_ASAP7_75t_L g861 ( .A(n_569), .Y(n_861) );
INVx3_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g805 ( .A(n_570), .Y(n_805) );
INVx2_ASAP7_75t_L g998 ( .A(n_570), .Y(n_998) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_572), .B(n_576), .Y(n_571) );
INVx2_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_SL g630 ( .A(n_574), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
INVx2_ASAP7_75t_L g1036 ( .A(n_579), .Y(n_1036) );
OA22x2_ASAP7_75t_L g642 ( .A1(n_581), .A2(n_643), .B1(n_670), .B2(n_671), .Y(n_642) );
INVx1_ASAP7_75t_L g670 ( .A(n_581), .Y(n_670) );
NOR2x1_ASAP7_75t_L g582 ( .A(n_583), .B(n_595), .Y(n_582) );
NAND4xp25_ASAP7_75t_L g583 ( .A(n_584), .B(n_588), .C(n_590), .D(n_592), .Y(n_583) );
BUFx4f_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
BUFx6f_ASAP7_75t_L g845 ( .A(n_586), .Y(n_845) );
NAND3xp33_ASAP7_75t_L g595 ( .A(n_596), .B(n_599), .C(n_606), .Y(n_595) );
BUFx3_ASAP7_75t_L g836 ( .A(n_597), .Y(n_836) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g874 ( .A(n_605), .B(n_875), .Y(n_874) );
BUFx3_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND4xp25_ASAP7_75t_L g633 ( .A(n_610), .B(n_611), .C(n_615), .D(n_627), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_614), .B(n_629), .Y(n_635) );
NAND3xp33_ASAP7_75t_L g616 ( .A(n_617), .B(n_627), .C(n_629), .Y(n_616) );
INVxp67_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g634 ( .A(n_618), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_625), .Y(n_618) );
INVx2_ASAP7_75t_L g986 ( .A(n_620), .Y(n_986) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx4_ASAP7_75t_L g827 ( .A(n_623), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g890 ( .A(n_623), .B(n_891), .Y(n_890) );
NOR2xp33_ASAP7_75t_L g928 ( .A(n_623), .B(n_929), .Y(n_928) );
NOR2xp33_ASAP7_75t_L g971 ( .A(n_623), .B(n_972), .Y(n_971) );
INVx4_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx3_ASAP7_75t_L g666 ( .A(n_624), .Y(n_666) );
BUFx2_ASAP7_75t_L g681 ( .A(n_626), .Y(n_681) );
INVx2_ASAP7_75t_L g1400 ( .A(n_626), .Y(n_1400) );
INVx1_ASAP7_75t_L g765 ( .A(n_628), .Y(n_765) );
INVx2_ASAP7_75t_L g760 ( .A(n_630), .Y(n_760) );
INVx4_ASAP7_75t_L g762 ( .A(n_631), .Y(n_762) );
BUFx3_ASAP7_75t_L g1396 ( .A(n_631), .Y(n_1396) );
NOR2x1_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OA22x2_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B1(n_672), .B2(n_673), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g671 ( .A(n_643), .Y(n_671) );
XOR2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_669), .Y(n_643) );
NOR2xp67_ASAP7_75t_L g644 ( .A(n_645), .B(n_658), .Y(n_644) );
NAND4xp25_ASAP7_75t_L g645 ( .A(n_646), .B(n_649), .C(n_652), .D(n_655), .Y(n_645) );
NAND4xp25_ASAP7_75t_L g658 ( .A(n_659), .B(n_661), .C(n_663), .D(n_667), .Y(n_658) );
INVx2_ASAP7_75t_L g956 ( .A(n_660), .Y(n_956) );
INVx1_ASAP7_75t_L g1030 ( .A(n_660), .Y(n_1030) );
BUFx3_ASAP7_75t_L g1364 ( .A(n_660), .Y(n_1364) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
INVx4_ASAP7_75t_L g688 ( .A(n_666), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g1091 ( .A(n_666), .B(n_1092), .Y(n_1091) );
NOR2xp33_ASAP7_75t_L g1365 ( .A(n_666), .B(n_1366), .Y(n_1365) );
INVx2_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
XOR2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_721), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_698), .Y(n_674) );
NOR3xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_682), .C(n_689), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_678), .B1(n_679), .B2(n_680), .Y(n_676) );
OAI22xp33_ASAP7_75t_L g752 ( .A1(n_678), .A2(n_753), .B1(n_754), .B2(n_755), .Y(n_752) );
OAI22xp5_ASAP7_75t_L g848 ( .A1(n_678), .A2(n_849), .B1(n_850), .B2(n_851), .Y(n_848) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OAI21xp33_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_684), .B(n_686), .Y(n_682) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_691), .B1(n_694), .B2(n_695), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
BUFx3_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
BUFx3_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NOR2xp67_ASAP7_75t_L g698 ( .A(n_699), .B(n_706), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_700), .B(n_703), .Y(n_699) );
BUFx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
BUFx3_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_715), .Y(n_706) );
BUFx4f_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g801 ( .A(n_710), .Y(n_801) );
INVx1_ASAP7_75t_L g1383 ( .A(n_710), .Y(n_1383) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g733 ( .A(n_712), .Y(n_733) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
BUFx6f_ASAP7_75t_L g1005 ( .A(n_713), .Y(n_1005) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
BUFx3_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g774 ( .A(n_717), .Y(n_774) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g775 ( .A(n_719), .Y(n_775) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
HB1xp67_ASAP7_75t_L g837 ( .A(n_720), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_830), .B1(n_899), .B2(n_900), .Y(n_722) );
INVx1_ASAP7_75t_L g899 ( .A(n_723), .Y(n_899) );
XNOR2x1_ASAP7_75t_L g723 ( .A(n_724), .B(n_746), .Y(n_723) );
BUFx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AO21x2_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_727), .B(n_745), .Y(n_725) );
NOR3xp33_ASAP7_75t_SL g745 ( .A(n_726), .B(n_729), .C(n_736), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_735), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NAND4xp25_ASAP7_75t_SL g729 ( .A(n_730), .B(n_731), .C(n_732), .D(n_734), .Y(n_729) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
NAND4xp25_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .C(n_741), .D(n_744), .Y(n_736) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g1066 ( .A(n_740), .Y(n_1066) );
BUFx3_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
OA22x2_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_748), .B1(n_791), .B2(n_792), .Y(n_746) );
INVx4_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
AO22x2_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_750), .B1(n_767), .B2(n_789), .Y(n_748) );
NOR4xp25_ASAP7_75t_L g749 ( .A(n_750), .B(n_752), .C(n_758), .D(n_763), .Y(n_749) );
CKINVDCx5p33_ASAP7_75t_R g750 ( .A(n_751), .Y(n_750) );
NOR3xp33_ASAP7_75t_SL g790 ( .A(n_752), .B(n_758), .C(n_763), .Y(n_790) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g812 ( .A(n_757), .Y(n_812) );
INVx2_ASAP7_75t_L g852 ( .A(n_757), .Y(n_852) );
OAI22xp33_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_760), .B1(n_761), .B2(n_762), .Y(n_758) );
OAI22xp5_ASAP7_75t_L g853 ( .A1(n_762), .A2(n_854), .B1(n_855), .B2(n_858), .Y(n_853) );
OAI21xp33_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_765), .B(n_766), .Y(n_763) );
NAND2xp5_ASAP7_75t_SL g789 ( .A(n_767), .B(n_790), .Y(n_789) );
NOR3xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_776), .C(n_783), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_772), .Y(n_768) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_779), .B1(n_780), .B2(n_781), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
OAI22xp5_ASAP7_75t_L g842 ( .A1(n_781), .A2(n_843), .B1(n_844), .B2(n_846), .Y(n_842) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
OAI22x1_ASAP7_75t_SL g783 ( .A1(n_784), .A2(n_785), .B1(n_787), .B2(n_788), .Y(n_783) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_SL g791 ( .A(n_792), .Y(n_791) );
XNOR2xp5_ASAP7_75t_L g792 ( .A(n_793), .B(n_813), .Y(n_792) );
NOR2x1_ASAP7_75t_L g794 ( .A(n_795), .B(n_802), .Y(n_794) );
NAND4xp25_ASAP7_75t_L g795 ( .A(n_796), .B(n_798), .C(n_799), .D(n_800), .Y(n_795) );
NAND3xp33_ASAP7_75t_L g802 ( .A(n_803), .B(n_810), .C(n_811), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
NOR2xp33_ASAP7_75t_L g1049 ( .A(n_808), .B(n_1050), .Y(n_1049) );
INVx3_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
XNOR2x1_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .Y(n_813) );
NOR2x1_ASAP7_75t_L g815 ( .A(n_816), .B(n_821), .Y(n_815) );
NAND4xp25_ASAP7_75t_L g816 ( .A(n_817), .B(n_818), .C(n_819), .D(n_820), .Y(n_816) );
NAND3xp33_ASAP7_75t_L g821 ( .A(n_822), .B(n_828), .C(n_829), .Y(n_821) );
INVx2_ASAP7_75t_L g991 ( .A(n_823), .Y(n_991) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_825), .B(n_826), .Y(n_824) );
INVx2_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g900 ( .A(n_830), .Y(n_900) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
XNOR2x1_ASAP7_75t_L g831 ( .A(n_832), .B(n_864), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_834), .B(n_847), .Y(n_833) );
NOR3xp33_ASAP7_75t_L g834 ( .A(n_835), .B(n_838), .C(n_842), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_839), .B(n_841), .Y(n_838) );
INVxp67_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
NOR3xp33_ASAP7_75t_L g847 ( .A(n_848), .B(n_853), .C(n_859), .Y(n_847) );
INVxp67_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
BUFx3_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
OAI21xp33_ASAP7_75t_L g859 ( .A1(n_860), .A2(n_861), .B(n_862), .Y(n_859) );
OA22x2_ASAP7_75t_L g864 ( .A1(n_865), .A2(n_866), .B1(n_882), .B2(n_898), .Y(n_864) );
INVx2_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
NOR2x1_ASAP7_75t_L g867 ( .A(n_868), .B(n_876), .Y(n_867) );
NAND4xp25_ASAP7_75t_L g868 ( .A(n_869), .B(n_870), .C(n_871), .D(n_873), .Y(n_868) );
BUFx2_ASAP7_75t_L g1398 ( .A(n_872), .Y(n_1398) );
NAND4xp25_ASAP7_75t_L g876 ( .A(n_877), .B(n_878), .C(n_880), .D(n_881), .Y(n_876) );
BUFx2_ASAP7_75t_SL g1387 ( .A(n_879), .Y(n_1387) );
INVx2_ASAP7_75t_L g898 ( .A(n_882), .Y(n_898) );
AO21x2_ASAP7_75t_L g882 ( .A1(n_883), .A2(n_884), .B(n_897), .Y(n_882) );
NOR3xp33_ASAP7_75t_SL g897 ( .A(n_883), .B(n_885), .C(n_892), .Y(n_897) );
OR2x2_ASAP7_75t_L g884 ( .A(n_885), .B(n_892), .Y(n_884) );
NAND4xp75_ASAP7_75t_L g885 ( .A(n_886), .B(n_887), .C(n_888), .D(n_889), .Y(n_885) );
NAND4xp25_ASAP7_75t_L g892 ( .A(n_893), .B(n_894), .C(n_895), .D(n_896), .Y(n_892) );
AOI22xp5_ASAP7_75t_L g901 ( .A1(n_902), .A2(n_1009), .B1(n_1010), .B2(n_1099), .Y(n_901) );
INVx2_ASAP7_75t_L g1099 ( .A(n_902), .Y(n_1099) );
XNOR2x1_ASAP7_75t_L g902 ( .A(n_903), .B(n_940), .Y(n_902) );
BUFx2_ASAP7_75t_SL g903 ( .A(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
OA22x2_ASAP7_75t_L g905 ( .A1(n_906), .A2(n_920), .B1(n_921), .B2(n_939), .Y(n_905) );
INVx2_ASAP7_75t_L g939 ( .A(n_906), .Y(n_939) );
OAI22xp5_ASAP7_75t_L g1078 ( .A1(n_906), .A2(n_939), .B1(n_1079), .B2(n_1095), .Y(n_1078) );
INVx1_ASAP7_75t_L g918 ( .A(n_907), .Y(n_918) );
NAND3xp33_ASAP7_75t_L g907 ( .A(n_908), .B(n_913), .C(n_916), .Y(n_907) );
AND4x1_ASAP7_75t_L g908 ( .A(n_909), .B(n_910), .C(n_911), .D(n_912), .Y(n_908) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
XNOR2x1_ASAP7_75t_L g921 ( .A(n_922), .B(n_938), .Y(n_921) );
OR2x2_ASAP7_75t_L g922 ( .A(n_923), .B(n_931), .Y(n_922) );
NAND4xp25_ASAP7_75t_L g923 ( .A(n_924), .B(n_926), .C(n_927), .D(n_930), .Y(n_923) );
NAND4xp25_ASAP7_75t_L g931 ( .A(n_932), .B(n_934), .C(n_935), .D(n_936), .Y(n_931) );
OAI22xp5_ASAP7_75t_L g1146 ( .A1(n_938), .A2(n_1117), .B1(n_1147), .B2(n_1148), .Y(n_1146) );
OA22x2_ASAP7_75t_L g940 ( .A1(n_941), .A2(n_942), .B1(n_979), .B2(n_980), .Y(n_940) );
INVx2_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
OA22x2_ASAP7_75t_L g942 ( .A1(n_943), .A2(n_962), .B1(n_963), .B2(n_978), .Y(n_942) );
INVx1_ASAP7_75t_L g978 ( .A(n_943), .Y(n_978) );
XNOR2x1_ASAP7_75t_L g943 ( .A(n_944), .B(n_945), .Y(n_943) );
NOR2x1_ASAP7_75t_L g945 ( .A(n_946), .B(n_951), .Y(n_945) );
NAND4xp25_ASAP7_75t_L g946 ( .A(n_947), .B(n_948), .C(n_949), .D(n_950), .Y(n_946) );
NAND3xp33_ASAP7_75t_L g951 ( .A(n_952), .B(n_953), .C(n_954), .Y(n_951) );
INVx2_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
OAI21xp5_ASAP7_75t_L g957 ( .A1(n_958), .A2(n_959), .B(n_961), .Y(n_957) );
INVx4_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
INVx1_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
INVx1_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
NOR2x1_ASAP7_75t_L g965 ( .A(n_966), .B(n_973), .Y(n_965) );
NAND4xp25_ASAP7_75t_L g966 ( .A(n_967), .B(n_968), .C(n_969), .D(n_970), .Y(n_966) );
NAND4xp25_ASAP7_75t_L g973 ( .A(n_974), .B(n_975), .C(n_976), .D(n_977), .Y(n_973) );
INVx2_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
INVx2_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
AND2x2_ASAP7_75t_L g982 ( .A(n_983), .B(n_1001), .Y(n_982) );
NOR3xp33_ASAP7_75t_L g983 ( .A(n_984), .B(n_989), .C(n_995), .Y(n_983) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_985), .A2(n_986), .B1(n_987), .B2(n_988), .Y(n_984) );
INVx2_ASAP7_75t_L g1025 ( .A(n_986), .Y(n_1025) );
OAI22xp5_ASAP7_75t_L g989 ( .A1(n_990), .A2(n_991), .B1(n_992), .B2(n_993), .Y(n_989) );
INVx1_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
OAI21xp33_ASAP7_75t_L g995 ( .A1(n_996), .A2(n_997), .B(n_999), .Y(n_995) );
INVx2_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
INVx2_ASAP7_75t_SL g1393 ( .A(n_1000), .Y(n_1393) );
NOR2xp33_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1006), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1004), .Y(n_1002) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_1007), .B(n_1008), .Y(n_1006) );
INVx1_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
AO22x1_ASAP7_75t_L g1010 ( .A1(n_1011), .A2(n_1076), .B1(n_1097), .B2(n_1098), .Y(n_1010) );
INVx2_ASAP7_75t_L g1098 ( .A(n_1011), .Y(n_1098) );
OA22x2_ASAP7_75t_L g1011 ( .A1(n_1012), .A2(n_1038), .B1(n_1074), .B2(n_1075), .Y(n_1011) );
INVx2_ASAP7_75t_L g1075 ( .A(n_1012), .Y(n_1075) );
AO21x2_ASAP7_75t_L g1012 ( .A1(n_1013), .A2(n_1014), .B(n_1037), .Y(n_1012) );
NOR3xp33_ASAP7_75t_L g1037 ( .A(n_1013), .B(n_1016), .C(n_1022), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_1015), .B(n_1021), .Y(n_1014) );
INVx1_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
NAND4xp25_ASAP7_75t_SL g1016 ( .A(n_1017), .B(n_1018), .C(n_1019), .D(n_1020), .Y(n_1016) );
INVx1_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
NAND3xp33_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1024), .C(n_1028), .Y(n_1022) );
BUFx3_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
INVx2_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
OAI21xp5_ASAP7_75t_SL g1031 ( .A1(n_1032), .A2(n_1034), .B(n_1035), .Y(n_1031) );
INVxp67_ASAP7_75t_L g1032 ( .A(n_1033), .Y(n_1032) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1038), .Y(n_1074) );
XNOR2xp5_ASAP7_75t_L g1038 ( .A(n_1039), .B(n_1057), .Y(n_1038) );
NAND4xp75_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1044), .C(n_1051), .D(n_1054), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1043), .Y(n_1041) );
OA21x2_ASAP7_75t_L g1044 ( .A1(n_1045), .A2(n_1046), .B(n_1048), .Y(n_1044) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_1052), .B(n_1053), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1056), .Y(n_1054) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1057), .Y(n_1096) );
XNOR2xp5_ASAP7_75t_L g1057 ( .A(n_1058), .B(n_1060), .Y(n_1057) );
CKINVDCx5p33_ASAP7_75t_R g1058 ( .A(n_1059), .Y(n_1058) );
NOR2x1_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1068), .Y(n_1060) );
NAND4xp25_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1064), .C(n_1065), .D(n_1067), .Y(n_1061) );
NAND4xp25_ASAP7_75t_L g1068 ( .A(n_1069), .B(n_1070), .C(n_1071), .D(n_1072), .Y(n_1068) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
HB1xp67_ASAP7_75t_L g1097 ( .A(n_1077), .Y(n_1097) );
XOR2x2_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1096), .Y(n_1077) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1079), .Y(n_1095) );
NOR3xp33_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1085), .C(n_1088), .Y(n_1080) );
NAND2xp5_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1083), .Y(n_1081) );
NAND2xp5_ASAP7_75t_SL g1085 ( .A(n_1086), .B(n_1087), .Y(n_1085) );
NAND4xp25_ASAP7_75t_SL g1088 ( .A(n_1089), .B(n_1090), .C(n_1093), .D(n_1094), .Y(n_1088) );
OAI221xp5_ASAP7_75t_SL g1100 ( .A1(n_1101), .A2(n_1344), .B1(n_1346), .B2(n_1367), .C(n_1372), .Y(n_1100) );
AOI21x1_ASAP7_75t_L g1101 ( .A1(n_1102), .A2(n_1259), .B(n_1308), .Y(n_1101) );
NAND5xp2_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1192), .C(n_1222), .D(n_1234), .E(n_1246), .Y(n_1102) );
AOI221xp5_ASAP7_75t_SL g1103 ( .A1(n_1104), .A2(n_1172), .B1(n_1182), .B2(n_1186), .C(n_1187), .Y(n_1103) );
A2O1A1Ixp33_ASAP7_75t_L g1104 ( .A1(n_1105), .A2(n_1156), .B(n_1160), .C(n_1165), .Y(n_1104) );
INVxp67_ASAP7_75t_SL g1342 ( .A(n_1105), .Y(n_1342) );
NAND2xp5_ASAP7_75t_L g1105 ( .A(n_1106), .B(n_1144), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
AOI211xp5_ASAP7_75t_L g1230 ( .A1(n_1107), .A2(n_1223), .B(n_1231), .C(n_1233), .Y(n_1230) );
OAI21xp33_ASAP7_75t_L g1249 ( .A1(n_1107), .A2(n_1250), .B(n_1252), .Y(n_1249) );
NAND2xp5_ASAP7_75t_L g1107 ( .A(n_1108), .B(n_1130), .Y(n_1107) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1108), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1108), .B(n_1184), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1108), .B(n_1199), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1236 ( .A(n_1108), .B(n_1237), .Y(n_1236) );
NOR2xp33_ASAP7_75t_L g1240 ( .A(n_1108), .B(n_1207), .Y(n_1240) );
NAND2xp5_ASAP7_75t_L g1269 ( .A(n_1108), .B(n_1171), .Y(n_1269) );
NAND2xp5_ASAP7_75t_L g1273 ( .A(n_1108), .B(n_1209), .Y(n_1273) );
NAND2xp5_ASAP7_75t_L g1321 ( .A(n_1108), .B(n_1160), .Y(n_1321) );
CKINVDCx6p67_ASAP7_75t_R g1108 ( .A(n_1109), .Y(n_1108) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1109), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1109), .B(n_1130), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_1109), .B(n_1144), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1109), .B(n_1209), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1109), .B(n_1262), .Y(n_1261) );
NAND2xp5_ASAP7_75t_L g1265 ( .A(n_1109), .B(n_1184), .Y(n_1265) );
NOR2xp33_ASAP7_75t_L g1287 ( .A(n_1109), .B(n_1144), .Y(n_1287) );
NOR2xp33_ASAP7_75t_L g1293 ( .A(n_1109), .B(n_1145), .Y(n_1293) );
NAND2xp5_ASAP7_75t_L g1299 ( .A(n_1109), .B(n_1300), .Y(n_1299) );
NOR2xp33_ASAP7_75t_L g1305 ( .A(n_1109), .B(n_1285), .Y(n_1305) );
OR2x6_ASAP7_75t_SL g1109 ( .A(n_1110), .B(n_1120), .Y(n_1109) );
OAI22xp5_ASAP7_75t_L g1110 ( .A1(n_1111), .A2(n_1116), .B1(n_1117), .B2(n_1119), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_1113), .B(n_1118), .Y(n_1117) );
AND2x4_ASAP7_75t_L g1134 ( .A(n_1113), .B(n_1118), .Y(n_1134) );
AND2x4_ASAP7_75t_L g1142 ( .A(n_1113), .B(n_1128), .Y(n_1142) );
AND2x4_ASAP7_75t_L g1143 ( .A(n_1113), .B(n_1118), .Y(n_1143) );
OAI221xp5_ASAP7_75t_L g1217 ( .A1(n_1117), .A2(n_1147), .B1(n_1218), .B2(n_1219), .C(n_1220), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1123 ( .A(n_1118), .B(n_1124), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1118), .B(n_1124), .Y(n_1140) );
AND2x4_ASAP7_75t_L g1155 ( .A(n_1118), .B(n_1124), .Y(n_1155) );
OAI22xp5_ASAP7_75t_L g1120 ( .A1(n_1121), .A2(n_1122), .B1(n_1125), .B2(n_1126), .Y(n_1120) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_1124), .B(n_1128), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1124), .B(n_1128), .Y(n_1139) );
AND2x4_ASAP7_75t_L g1152 ( .A(n_1124), .B(n_1128), .Y(n_1152) );
CKINVDCx5p33_ASAP7_75t_R g1406 ( .A(n_1124), .Y(n_1406) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
NAND2xp5_ASAP7_75t_L g1156 ( .A(n_1130), .B(n_1157), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1196 ( .A(n_1130), .B(n_1184), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1226 ( .A(n_1130), .B(n_1227), .Y(n_1226) );
NAND2xp5_ASAP7_75t_L g1318 ( .A(n_1130), .B(n_1210), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_1131), .B(n_1136), .Y(n_1130) );
NOR2xp33_ASAP7_75t_L g1166 ( .A(n_1131), .B(n_1157), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1131), .B(n_1137), .Y(n_1191) );
CKINVDCx5p33_ASAP7_75t_R g1131 ( .A(n_1132), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1132), .B(n_1137), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1132), .B(n_1136), .Y(n_1238) );
NAND2xp5_ASAP7_75t_L g1276 ( .A(n_1132), .B(n_1157), .Y(n_1276) );
OR2x2_ASAP7_75t_L g1316 ( .A(n_1132), .B(n_1157), .Y(n_1316) );
AND2x4_ASAP7_75t_SL g1132 ( .A(n_1133), .B(n_1135), .Y(n_1132) );
INVx2_ASAP7_75t_SL g1181 ( .A(n_1134), .Y(n_1181) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1136), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1136), .B(n_1199), .Y(n_1243) );
NOR2xp33_ASAP7_75t_L g1300 ( .A(n_1136), .B(n_1199), .Y(n_1300) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1137), .Y(n_1136) );
NAND2xp5_ASAP7_75t_L g1137 ( .A(n_1138), .B(n_1141), .Y(n_1137) );
INVx3_ASAP7_75t_L g1147 ( .A(n_1142), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1144), .B(n_1162), .Y(n_1186) );
NOR2xp33_ASAP7_75t_L g1245 ( .A(n_1144), .B(n_1201), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_1144), .B(n_1176), .Y(n_1248) );
NAND2xp5_ASAP7_75t_L g1267 ( .A(n_1144), .B(n_1175), .Y(n_1267) );
INVx3_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1145), .B(n_1161), .Y(n_1171) );
OR2x2_ASAP7_75t_L g1207 ( .A(n_1145), .B(n_1162), .Y(n_1207) );
INVx2_ASAP7_75t_L g1225 ( .A(n_1145), .Y(n_1225) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1145), .B(n_1162), .Y(n_1281) );
OR2x2_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1149), .Y(n_1145) );
OAI22xp5_ASAP7_75t_L g1149 ( .A1(n_1150), .A2(n_1151), .B1(n_1153), .B2(n_1154), .Y(n_1149) );
INVx3_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
INVx2_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
BUFx2_ASAP7_75t_L g1345 ( .A(n_1155), .Y(n_1345) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1156), .Y(n_1338) );
CKINVDCx6p67_ASAP7_75t_R g1184 ( .A(n_1157), .Y(n_1184) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1157), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1157), .B(n_1238), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1157), .B(n_1191), .Y(n_1262) );
OAI322xp33_ASAP7_75t_L g1268 ( .A1(n_1157), .A2(n_1174), .A3(n_1269), .B1(n_1270), .B2(n_1273), .C1(n_1274), .C2(n_1276), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1158), .B(n_1159), .Y(n_1157) );
AOI221xp5_ASAP7_75t_L g1246 ( .A1(n_1160), .A2(n_1247), .B1(n_1248), .B2(n_1249), .C(n_1253), .Y(n_1246) );
INVx3_ASAP7_75t_L g1288 ( .A(n_1160), .Y(n_1288) );
OAI21xp5_ASAP7_75t_L g1289 ( .A1(n_1160), .A2(n_1290), .B(n_1291), .Y(n_1289) );
INVx3_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
OR2x2_ASAP7_75t_L g1201 ( .A(n_1161), .B(n_1177), .Y(n_1201) );
NAND2xp5_ASAP7_75t_L g1212 ( .A(n_1161), .B(n_1177), .Y(n_1212) );
INVx2_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1162), .B(n_1177), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1163), .B(n_1164), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_1166), .B(n_1167), .Y(n_1165) );
NAND2xp5_ASAP7_75t_L g1292 ( .A(n_1166), .B(n_1293), .Y(n_1292) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
NOR2xp33_ASAP7_75t_L g1221 ( .A(n_1168), .B(n_1197), .Y(n_1221) );
NOR2xp33_ASAP7_75t_L g1228 ( .A(n_1168), .B(n_1229), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1171), .Y(n_1168) );
NAND2xp5_ASAP7_75t_L g1213 ( .A(n_1169), .B(n_1191), .Y(n_1213) );
NOR2xp33_ASAP7_75t_L g1304 ( .A(n_1169), .B(n_1177), .Y(n_1304) );
NOR2xp33_ASAP7_75t_L g1333 ( .A(n_1169), .B(n_1334), .Y(n_1333) );
O2A1O1Ixp33_ASAP7_75t_L g1343 ( .A1(n_1169), .A2(n_1204), .B(n_1213), .C(n_1257), .Y(n_1343) );
INVx3_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1297 ( .A(n_1171), .B(n_1174), .Y(n_1297) );
NAND3xp33_ASAP7_75t_L g1340 ( .A(n_1171), .B(n_1243), .C(n_1304), .Y(n_1340) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1172), .Y(n_1326) );
INVx3_ASAP7_75t_L g1172 ( .A(n_1173), .Y(n_1172) );
INVx3_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
NOR2xp33_ASAP7_75t_L g1187 ( .A(n_1174), .B(n_1188), .Y(n_1187) );
INVx3_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
INVx2_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
NAND2xp5_ASAP7_75t_L g1214 ( .A(n_1176), .B(n_1215), .Y(n_1214) );
A2O1A1Ixp33_ASAP7_75t_L g1337 ( .A1(n_1176), .A2(n_1206), .B(n_1338), .C(n_1339), .Y(n_1337) );
INVx3_ASAP7_75t_L g1176 ( .A(n_1177), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1177), .B(n_1206), .Y(n_1205) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1177), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1313 ( .A(n_1177), .B(n_1281), .Y(n_1313) );
AND2x4_ASAP7_75t_L g1177 ( .A(n_1178), .B(n_1179), .Y(n_1177) );
INVx2_ASAP7_75t_L g1180 ( .A(n_1181), .Y(n_1180) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1184), .B(n_1185), .Y(n_1183) );
AND2x2_ASAP7_75t_SL g1190 ( .A(n_1184), .B(n_1191), .Y(n_1190) );
NOR2xp33_ASAP7_75t_L g1232 ( .A(n_1184), .B(n_1229), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1184), .B(n_1238), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1329 ( .A(n_1184), .B(n_1209), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1185), .B(n_1199), .Y(n_1290) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1185), .Y(n_1315) );
AOI322xp5_ASAP7_75t_L g1311 ( .A1(n_1186), .A2(n_1235), .A3(n_1275), .B1(n_1312), .B2(n_1314), .C1(n_1316), .C2(n_1317), .Y(n_1311) );
INVxp67_ASAP7_75t_SL g1278 ( .A(n_1188), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1190), .Y(n_1188) );
INVxp67_ASAP7_75t_L g1256 ( .A(n_1189), .Y(n_1256) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1190), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1191), .B(n_1210), .Y(n_1215) );
AOI222xp33_ASAP7_75t_L g1234 ( .A1(n_1191), .A2(n_1235), .B1(n_1239), .B2(n_1240), .C1(n_1241), .C2(n_1245), .Y(n_1234) );
OR2x2_ASAP7_75t_L g1303 ( .A(n_1191), .B(n_1238), .Y(n_1303) );
INVxp33_ASAP7_75t_L g1334 ( .A(n_1191), .Y(n_1334) );
NOR3xp33_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1211), .C(n_1221), .Y(n_1192) );
OAI32xp33_ASAP7_75t_L g1193 ( .A1(n_1194), .A2(n_1201), .A3(n_1202), .B1(n_1204), .B2(n_1208), .Y(n_1193) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
NAND2xp5_ASAP7_75t_L g1195 ( .A(n_1196), .B(n_1197), .Y(n_1195) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1196), .Y(n_1295) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1197), .Y(n_1322) );
NAND2xp5_ASAP7_75t_L g1197 ( .A(n_1198), .B(n_1199), .Y(n_1197) );
AOI321xp33_ASAP7_75t_L g1302 ( .A1(n_1199), .A2(n_1248), .A3(n_1303), .B1(n_1304), .B2(n_1305), .C(n_1306), .Y(n_1302) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1201), .Y(n_1239) );
OAI211xp5_ASAP7_75t_L g1336 ( .A1(n_1201), .A2(n_1292), .B(n_1337), .C(n_1340), .Y(n_1336) );
CKINVDCx14_ASAP7_75t_R g1202 ( .A(n_1203), .Y(n_1202) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
OAI221xp5_ASAP7_75t_L g1279 ( .A1(n_1207), .A2(n_1280), .B1(n_1282), .B2(n_1283), .C(n_1286), .Y(n_1279) );
NAND2xp5_ASAP7_75t_L g1208 ( .A(n_1209), .B(n_1210), .Y(n_1208) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1209), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_1209), .B(n_1264), .Y(n_1263) );
NAND3xp33_ASAP7_75t_L g1286 ( .A(n_1209), .B(n_1287), .C(n_1288), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1209), .B(n_1227), .Y(n_1325) );
OAI211xp5_ASAP7_75t_L g1211 ( .A1(n_1212), .A2(n_1213), .B(n_1214), .C(n_1216), .Y(n_1211) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1212), .Y(n_1233) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1214), .Y(n_1339) );
INVx2_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
BUFx3_ASAP7_75t_L g1307 ( .A(n_1217), .Y(n_1307) );
AOI211xp5_ASAP7_75t_L g1222 ( .A1(n_1223), .A2(n_1226), .B(n_1228), .C(n_1230), .Y(n_1222) );
INVx2_ASAP7_75t_L g1223 ( .A(n_1224), .Y(n_1223) );
BUFx2_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1225), .Y(n_1251) );
NOR2xp33_ASAP7_75t_L g1271 ( .A(n_1225), .B(n_1272), .Y(n_1271) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1226), .Y(n_1252) );
NOR2xp33_ASAP7_75t_L g1301 ( .A(n_1231), .B(n_1270), .Y(n_1301) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1233), .B(n_1251), .Y(n_1275) );
AOI221xp5_ASAP7_75t_L g1294 ( .A1(n_1233), .A2(n_1295), .B1(n_1296), .B2(n_1298), .C(n_1301), .Y(n_1294) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1236), .Y(n_1235) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1238), .Y(n_1285) );
AOI21xp5_ASAP7_75t_L g1277 ( .A1(n_1239), .A2(n_1278), .B(n_1279), .Y(n_1277) );
NAND2xp5_ASAP7_75t_L g1241 ( .A(n_1242), .B(n_1244), .Y(n_1241) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1245), .Y(n_1335) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g1324 ( .A(n_1251), .B(n_1325), .Y(n_1324) );
AOI21xp5_ASAP7_75t_L g1253 ( .A1(n_1254), .A2(n_1256), .B(n_1257), .Y(n_1253) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
O2A1O1Ixp33_ASAP7_75t_L g1341 ( .A1(n_1255), .A2(n_1263), .B(n_1342), .C(n_1343), .Y(n_1341) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
NAND5xp2_ASAP7_75t_L g1259 ( .A(n_1260), .B(n_1277), .C(n_1289), .D(n_1294), .E(n_1302), .Y(n_1259) );
O2A1O1Ixp33_ASAP7_75t_L g1260 ( .A1(n_1261), .A2(n_1263), .B(n_1266), .C(n_1268), .Y(n_1260) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1262), .Y(n_1331) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1263), .Y(n_1282) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
NOR2xp33_ASAP7_75t_L g1284 ( .A(n_1265), .B(n_1285), .Y(n_1284) );
NAND2xp5_ASAP7_75t_SL g1314 ( .A(n_1265), .B(n_1315), .Y(n_1314) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1281), .Y(n_1280) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
INVxp67_ASAP7_75t_SL g1291 ( .A(n_1292), .Y(n_1291) );
AOI21xp33_ASAP7_75t_L g1327 ( .A1(n_1296), .A2(n_1328), .B(n_1330), .Y(n_1327) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1297), .Y(n_1296) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1299), .Y(n_1298) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1307), .Y(n_1306) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1309), .B(n_1341), .Y(n_1308) );
NOR2xp33_ASAP7_75t_L g1309 ( .A(n_1310), .B(n_1336), .Y(n_1309) );
NAND3xp33_ASAP7_75t_L g1310 ( .A(n_1311), .B(n_1319), .C(n_1327), .Y(n_1310) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1318), .Y(n_1317) );
A2O1A1Ixp33_ASAP7_75t_L g1319 ( .A1(n_1320), .A2(n_1322), .B(n_1323), .C(n_1326), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
AOI21xp33_ASAP7_75t_L g1330 ( .A1(n_1331), .A2(n_1332), .B(n_1335), .Y(n_1330) );
INVxp33_ASAP7_75t_L g1332 ( .A(n_1333), .Y(n_1332) );
CKINVDCx5p33_ASAP7_75t_R g1344 ( .A(n_1345), .Y(n_1344) );
INVxp67_ASAP7_75t_L g1346 ( .A(n_1347), .Y(n_1346) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1349), .Y(n_1348) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1350), .Y(n_1349) );
INVx2_ASAP7_75t_L g1351 ( .A(n_1352), .Y(n_1351) );
NAND4xp75_ASAP7_75t_L g1352 ( .A(n_1353), .B(n_1356), .C(n_1359), .D(n_1363), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1354), .B(n_1355), .Y(n_1353) );
AND2x2_ASAP7_75t_L g1356 ( .A(n_1357), .B(n_1358), .Y(n_1356) );
AND2x2_ASAP7_75t_L g1359 ( .A(n_1360), .B(n_1362), .Y(n_1359) );
HB1xp67_ASAP7_75t_L g1390 ( .A(n_1364), .Y(n_1390) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1368), .Y(n_1367) );
HB1xp67_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
INVxp67_ASAP7_75t_SL g1375 ( .A(n_1376), .Y(n_1375) );
BUFx2_ASAP7_75t_L g1376 ( .A(n_1377), .Y(n_1376) );
OR2x2_ASAP7_75t_L g1377 ( .A(n_1378), .B(n_1388), .Y(n_1377) );
NAND4xp25_ASAP7_75t_SL g1378 ( .A(n_1379), .B(n_1381), .C(n_1382), .D(n_1385), .Y(n_1378) );
NAND3xp33_ASAP7_75t_L g1388 ( .A(n_1389), .B(n_1395), .C(n_1397), .Y(n_1388) );
OAI21xp33_ASAP7_75t_L g1391 ( .A1(n_1392), .A2(n_1393), .B(n_1394), .Y(n_1391) );
INVx2_ASAP7_75t_L g1399 ( .A(n_1400), .Y(n_1399) );
BUFx3_ASAP7_75t_L g1402 ( .A(n_1403), .Y(n_1402) );
BUFx2_ASAP7_75t_L g1404 ( .A(n_1405), .Y(n_1404) );
endmodule