module fake_netlist_1_2297_n_1263 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_225, n_39, n_1263);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1263;
wire n_963;
wire n_1034;
wire n_949;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_830;
wire n_1112;
wire n_517;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_268;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_271;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_409;
wire n_315;
wire n_295;
wire n_677;
wire n_1242;
wire n_283;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_272;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_281;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_280;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_275;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1117;
wire n_1007;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_287;
wire n_606;
wire n_332;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_366;
wire n_596;
wire n_1215;
wire n_286;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_282;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_427;
wire n_703;
wire n_415;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_270;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_285;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_269;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_288;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1204;
wire n_1094;
wire n_392;
wire n_1169;
wire n_975;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_274;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_276;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_948;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_335;
wire n_700;
wire n_534;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_491;
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_48), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_262), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_173), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_249), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_13), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_186), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_81), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_77), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_78), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_121), .Y(n_277) );
BUFx3_ASAP7_75t_L g278 ( .A(n_232), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g279 ( .A(n_181), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_102), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_123), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_118), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_25), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_263), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_23), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_216), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_227), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_163), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_104), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_195), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_211), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_72), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_68), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_39), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_110), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_138), .Y(n_296) );
BUFx3_ASAP7_75t_L g297 ( .A(n_124), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_55), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_209), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_246), .Y(n_300) );
CKINVDCx16_ASAP7_75t_R g301 ( .A(n_45), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_237), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_142), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_114), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_20), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_44), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_241), .Y(n_307) );
BUFx3_ASAP7_75t_L g308 ( .A(n_127), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_115), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_185), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_117), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_153), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_252), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_76), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_156), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_92), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_116), .Y(n_317) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_217), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_133), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_58), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_139), .Y(n_321) );
CKINVDCx20_ASAP7_75t_R g322 ( .A(n_251), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_79), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_245), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_120), .Y(n_325) );
CKINVDCx16_ASAP7_75t_R g326 ( .A(n_37), .Y(n_326) );
BUFx3_ASAP7_75t_L g327 ( .A(n_144), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_49), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_193), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_43), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_264), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_48), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_257), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_51), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_1), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_239), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_134), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_31), .Y(n_338) );
BUFx3_ASAP7_75t_L g339 ( .A(n_1), .Y(n_339) );
INVxp67_ASAP7_75t_SL g340 ( .A(n_255), .Y(n_340) );
BUFx3_ASAP7_75t_L g341 ( .A(n_51), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_97), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_10), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_187), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_30), .Y(n_345) );
BUFx3_ASAP7_75t_L g346 ( .A(n_100), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_190), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_184), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_183), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_179), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_182), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_212), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_5), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_90), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_145), .Y(n_355) );
CKINVDCx14_ASAP7_75t_R g356 ( .A(n_59), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_170), .Y(n_357) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_126), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_207), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_106), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_218), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_46), .Y(n_362) );
INVxp33_ASAP7_75t_L g363 ( .A(n_157), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_265), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_98), .Y(n_365) );
NOR2xp67_ASAP7_75t_L g366 ( .A(n_149), .B(n_161), .Y(n_366) );
INVxp67_ASAP7_75t_SL g367 ( .A(n_101), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_107), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_36), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_111), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_151), .Y(n_371) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_228), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_40), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_162), .Y(n_374) );
BUFx12f_ASAP7_75t_L g375 ( .A(n_75), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_84), .Y(n_376) );
CKINVDCx14_ASAP7_75t_R g377 ( .A(n_12), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_78), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_131), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_88), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_6), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_152), .Y(n_382) );
CKINVDCx16_ASAP7_75t_R g383 ( .A(n_196), .Y(n_383) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_229), .Y(n_384) );
BUFx3_ASAP7_75t_L g385 ( .A(n_201), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_76), .Y(n_386) );
INVxp33_ASAP7_75t_L g387 ( .A(n_168), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_17), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_166), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_36), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_267), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_41), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_21), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_33), .Y(n_394) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_167), .Y(n_395) );
CKINVDCx20_ASAP7_75t_R g396 ( .A(n_18), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_113), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_84), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_213), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_109), .Y(n_400) );
BUFx3_ASAP7_75t_L g401 ( .A(n_112), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_231), .Y(n_402) );
BUFx3_ASAP7_75t_L g403 ( .A(n_158), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_238), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_258), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_208), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_214), .B(n_192), .Y(n_407) );
BUFx3_ASAP7_75t_L g408 ( .A(n_52), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_230), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_38), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_86), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_75), .Y(n_412) );
INVx4_ASAP7_75t_R g413 ( .A(n_73), .Y(n_413) );
CKINVDCx20_ASAP7_75t_R g414 ( .A(n_108), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_339), .B(n_0), .Y(n_415) );
INVx3_ASAP7_75t_L g416 ( .A(n_339), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_283), .Y(n_417) );
INVx1_ASAP7_75t_SL g418 ( .A(n_279), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_358), .B(n_0), .Y(n_419) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_303), .Y(n_420) );
INVx6_ASAP7_75t_L g421 ( .A(n_278), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_303), .Y(n_422) );
CKINVDCx6p67_ASAP7_75t_R g423 ( .A(n_383), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_283), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_303), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_338), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_303), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_363), .B(n_387), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_363), .B(n_2), .Y(n_429) );
INVx3_ASAP7_75t_L g430 ( .A(n_341), .Y(n_430) );
BUFx8_ASAP7_75t_L g431 ( .A(n_318), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_272), .B(n_2), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_338), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_388), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_274), .B(n_3), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_388), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_356), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_275), .B(n_4), .Y(n_438) );
INVxp67_ASAP7_75t_L g439 ( .A(n_341), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_318), .Y(n_440) );
INVx3_ASAP7_75t_L g441 ( .A(n_408), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_276), .B(n_6), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_412), .Y(n_443) );
AND2x6_ASAP7_75t_L g444 ( .A(n_278), .B(n_87), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_387), .B(n_7), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_292), .B(n_7), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_412), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_408), .Y(n_448) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_318), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_318), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_269), .Y(n_451) );
BUFx2_ASAP7_75t_L g452 ( .A(n_423), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_428), .B(n_273), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_429), .B(n_377), .Y(n_454) );
INVx4_ASAP7_75t_L g455 ( .A(n_444), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_415), .Y(n_456) );
OR2x6_ASAP7_75t_L g457 ( .A(n_419), .B(n_375), .Y(n_457) );
INVx2_ASAP7_75t_SL g458 ( .A(n_429), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_439), .B(n_273), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_423), .Y(n_460) );
NAND2x1p5_ASAP7_75t_L g461 ( .A(n_415), .B(n_270), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_439), .B(n_271), .Y(n_462) );
NAND3xp33_ASAP7_75t_L g463 ( .A(n_451), .B(n_281), .C(n_280), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_451), .B(n_277), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_445), .B(n_268), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_416), .Y(n_466) );
OR2x6_ASAP7_75t_L g467 ( .A(n_419), .B(n_375), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_445), .B(n_268), .Y(n_468) );
OAI22xp33_ASAP7_75t_L g469 ( .A1(n_437), .A2(n_326), .B1(n_301), .B2(n_285), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_418), .B(n_285), .Y(n_470) );
INVx3_ASAP7_75t_L g471 ( .A(n_415), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_416), .B(n_293), .Y(n_472) );
INVx3_ASAP7_75t_L g473 ( .A(n_416), .Y(n_473) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_418), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g475 ( .A(n_431), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_420), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_420), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_416), .B(n_293), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_432), .A2(n_298), .B1(n_314), .B2(n_305), .Y(n_479) );
NAND2xp33_ASAP7_75t_SL g480 ( .A(n_432), .B(n_279), .Y(n_480) );
BUFx2_ASAP7_75t_L g481 ( .A(n_431), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_430), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_435), .A2(n_323), .B1(n_330), .B2(n_328), .Y(n_483) );
BUFx3_ASAP7_75t_L g484 ( .A(n_431), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_448), .B(n_282), .Y(n_485) );
INVx1_ASAP7_75t_SL g486 ( .A(n_421), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_430), .Y(n_487) );
CKINVDCx5p33_ASAP7_75t_R g488 ( .A(n_431), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_420), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_420), .Y(n_490) );
AND2x6_ASAP7_75t_L g491 ( .A(n_430), .B(n_297), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_420), .Y(n_492) );
NAND3x1_ASAP7_75t_L g493 ( .A(n_437), .B(n_335), .C(n_332), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_441), .Y(n_494) );
INVx4_ASAP7_75t_L g495 ( .A(n_444), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_441), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_458), .A2(n_384), .B1(n_414), .B2(n_322), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_474), .B(n_435), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_458), .B(n_438), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_453), .B(n_438), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_454), .B(n_442), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_454), .B(n_442), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_452), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_484), .B(n_288), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_484), .B(n_290), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_456), .B(n_446), .Y(n_506) );
BUFx2_ASAP7_75t_L g507 ( .A(n_452), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_484), .B(n_290), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_456), .A2(n_446), .B1(n_444), .B2(n_421), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_473), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_473), .Y(n_511) );
NAND2xp33_ASAP7_75t_L g512 ( .A(n_461), .B(n_444), .Y(n_512) );
AND2x4_ASAP7_75t_L g513 ( .A(n_457), .B(n_322), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_466), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_473), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_456), .A2(n_444), .B1(n_421), .B2(n_343), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_470), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_480), .A2(n_414), .B1(n_384), .B2(n_294), .Y(n_518) );
BUFx5_ASAP7_75t_L g519 ( .A(n_491), .Y(n_519) );
NAND2x1p5_ASAP7_75t_L g520 ( .A(n_481), .B(n_345), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_482), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_465), .B(n_300), .Y(n_522) );
BUFx8_ASAP7_75t_L g523 ( .A(n_470), .Y(n_523) );
AOI22xp33_ASAP7_75t_SL g524 ( .A1(n_460), .A2(n_396), .B1(n_334), .B2(n_362), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_482), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_456), .B(n_300), .Y(n_526) );
AOI22x1_ASAP7_75t_L g527 ( .A1(n_455), .A2(n_350), .B1(n_352), .B2(n_324), .Y(n_527) );
AND2x4_ASAP7_75t_L g528 ( .A(n_457), .B(n_467), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_481), .B(n_302), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_487), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_468), .B(n_302), .Y(n_531) );
INVxp67_ASAP7_75t_L g532 ( .A(n_457), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_472), .B(n_310), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_487), .Y(n_534) );
INVx5_ASAP7_75t_L g535 ( .A(n_491), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_475), .B(n_310), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_478), .B(n_311), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_457), .B(n_306), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_494), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_494), .Y(n_540) );
CKINVDCx5p33_ASAP7_75t_R g541 ( .A(n_457), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_459), .B(n_312), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_496), .Y(n_543) );
AND2x2_ASAP7_75t_SL g544 ( .A(n_479), .B(n_353), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_467), .A2(n_334), .B1(n_362), .B2(n_306), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_496), .Y(n_546) );
AND2x4_ASAP7_75t_L g547 ( .A(n_467), .B(n_417), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_462), .B(n_325), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_493), .A2(n_396), .B1(n_369), .B2(n_376), .Y(n_549) );
NAND2x1p5_ASAP7_75t_L g550 ( .A(n_471), .B(n_373), .Y(n_550) );
NAND3xp33_ASAP7_75t_SL g551 ( .A(n_483), .B(n_392), .C(n_378), .Y(n_551) );
NAND3xp33_ASAP7_75t_SL g552 ( .A(n_461), .B(n_392), .C(n_378), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_467), .B(n_417), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_488), .B(n_325), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_464), .B(n_329), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_471), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_461), .B(n_329), .Y(n_557) );
BUFx3_ASAP7_75t_L g558 ( .A(n_467), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_485), .B(n_424), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_463), .B(n_348), .Y(n_560) );
INVx1_ASAP7_75t_SL g561 ( .A(n_491), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_469), .A2(n_386), .B1(n_390), .B2(n_381), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_463), .B(n_359), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_491), .A2(n_444), .B1(n_421), .B2(n_393), .Y(n_564) );
INVx5_ASAP7_75t_L g565 ( .A(n_491), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_486), .B(n_359), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_493), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_455), .B(n_371), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_455), .B(n_371), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_455), .A2(n_444), .B1(n_421), .B2(n_394), .Y(n_570) );
INVx8_ASAP7_75t_L g571 ( .A(n_495), .Y(n_571) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_495), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_495), .B(n_389), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_486), .B(n_391), .Y(n_574) );
OAI21xp5_ASAP7_75t_L g575 ( .A1(n_476), .A2(n_444), .B(n_286), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_492), .B(n_391), .Y(n_576) );
INVx2_ASAP7_75t_SL g577 ( .A(n_476), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_476), .B(n_397), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_477), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g580 ( .A(n_477), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_477), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_489), .B(n_397), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_492), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_489), .B(n_402), .Y(n_584) );
OAI22xp33_ASAP7_75t_SL g585 ( .A1(n_489), .A2(n_410), .B1(n_411), .B2(n_398), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_490), .A2(n_404), .B1(n_406), .B2(n_402), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_528), .B(n_404), .Y(n_587) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_503), .Y(n_588) );
AND2x4_ASAP7_75t_L g589 ( .A(n_528), .B(n_424), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_553), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_517), .B(n_426), .Y(n_591) );
A2O1A1Ixp33_ASAP7_75t_L g592 ( .A1(n_500), .A2(n_433), .B(n_434), .C(n_426), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_501), .B(n_406), .Y(n_593) );
INVx5_ASAP7_75t_L g594 ( .A(n_547), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_532), .B(n_409), .Y(n_595) );
INVx1_ASAP7_75t_SL g596 ( .A(n_507), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_520), .B(n_409), .Y(n_597) );
O2A1O1Ixp33_ASAP7_75t_L g598 ( .A1(n_501), .A2(n_434), .B(n_436), .C(n_433), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_543), .Y(n_599) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_520), .B(n_317), .Y(n_600) );
OA22x2_ASAP7_75t_L g601 ( .A1(n_497), .A2(n_436), .B1(n_447), .B2(n_443), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_502), .B(n_443), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_498), .B(n_340), .Y(n_603) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_571), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_502), .B(n_447), .Y(n_605) );
BUFx2_ASAP7_75t_L g606 ( .A(n_513), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_513), .A2(n_367), .B1(n_320), .B2(n_287), .Y(n_607) );
A2O1A1Ixp33_ASAP7_75t_L g608 ( .A1(n_506), .A2(n_289), .B(n_291), .C(n_284), .Y(n_608) );
A2O1A1Ixp33_ASAP7_75t_L g609 ( .A1(n_506), .A2(n_296), .B(n_299), .C(n_295), .Y(n_609) );
NAND2xp5_ASAP7_75t_SL g610 ( .A(n_547), .B(n_304), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_538), .B(n_524), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_556), .Y(n_612) );
AOI21xp5_ASAP7_75t_L g613 ( .A1(n_512), .A2(n_309), .B(n_307), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_550), .Y(n_614) );
OA21x2_ASAP7_75t_L g615 ( .A1(n_575), .A2(n_357), .B(n_352), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_499), .B(n_444), .Y(n_616) );
A2O1A1Ixp33_ASAP7_75t_L g617 ( .A1(n_499), .A2(n_313), .B(n_316), .C(n_315), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_558), .B(n_319), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_526), .A2(n_333), .B(n_331), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_550), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_557), .A2(n_320), .B1(n_337), .B2(n_336), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_541), .A2(n_320), .B1(n_344), .B2(n_342), .Y(n_622) );
NOR3xp33_ASAP7_75t_SL g623 ( .A(n_549), .B(n_349), .C(n_347), .Y(n_623) );
INVxp67_ASAP7_75t_SL g624 ( .A(n_523), .Y(n_624) );
OR2x6_ASAP7_75t_L g625 ( .A(n_567), .B(n_366), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_545), .B(n_351), .Y(n_626) );
NOR2xp67_ASAP7_75t_L g627 ( .A(n_535), .B(n_89), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_514), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_522), .B(n_354), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_526), .A2(n_360), .B(n_355), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_531), .B(n_361), .Y(n_631) );
NOR2xp33_ASAP7_75t_R g632 ( .A(n_552), .B(n_8), .Y(n_632) );
NOR3xp33_ASAP7_75t_SL g633 ( .A(n_549), .B(n_365), .C(n_364), .Y(n_633) );
A2O1A1Ixp33_ASAP7_75t_L g634 ( .A1(n_521), .A2(n_368), .B(n_374), .C(n_370), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_518), .A2(n_379), .B1(n_382), .B2(n_380), .Y(n_635) );
O2A1O1Ixp33_ASAP7_75t_L g636 ( .A1(n_585), .A2(n_400), .B(n_405), .C(n_399), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_525), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_568), .A2(n_490), .B(n_407), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_544), .A2(n_321), .B1(n_327), .B2(n_308), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_530), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_551), .B(n_8), .Y(n_641) );
AND2x4_ASAP7_75t_L g642 ( .A(n_559), .B(n_346), .Y(n_642) );
INVx3_ASAP7_75t_L g643 ( .A(n_510), .Y(n_643) );
A2O1A1Ixp33_ASAP7_75t_L g644 ( .A1(n_534), .A2(n_385), .B(n_403), .C(n_401), .Y(n_644) );
A2O1A1Ixp33_ASAP7_75t_L g645 ( .A1(n_539), .A2(n_403), .B(n_401), .C(n_422), .Y(n_645) );
A2O1A1Ixp33_ASAP7_75t_L g646 ( .A1(n_540), .A2(n_425), .B(n_427), .C(n_422), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_548), .B(n_9), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_546), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_511), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_515), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_536), .B(n_9), .Y(n_651) );
INVx2_ASAP7_75t_SL g652 ( .A(n_523), .Y(n_652) );
INVx5_ASAP7_75t_L g653 ( .A(n_565), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_574), .A2(n_450), .B1(n_440), .B2(n_395), .Y(n_654) );
OR2x2_ASAP7_75t_L g655 ( .A(n_562), .B(n_10), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_578), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_571), .A2(n_450), .B(n_395), .Y(n_657) );
BUFx3_ASAP7_75t_L g658 ( .A(n_555), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_527), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_571), .A2(n_395), .B(n_372), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g661 ( .A1(n_533), .A2(n_395), .B(n_372), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_537), .A2(n_372), .B(n_420), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_554), .B(n_11), .Y(n_663) );
A2O1A1Ixp33_ASAP7_75t_L g664 ( .A1(n_560), .A2(n_372), .B(n_449), .C(n_413), .Y(n_664) );
O2A1O1Ixp33_ASAP7_75t_L g665 ( .A1(n_574), .A2(n_12), .B(n_13), .C(n_14), .Y(n_665) );
OA22x2_ASAP7_75t_L g666 ( .A1(n_586), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_563), .B(n_15), .Y(n_667) );
OAI21x1_ASAP7_75t_L g668 ( .A1(n_509), .A2(n_93), .B(n_91), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_542), .B(n_16), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_582), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_584), .Y(n_671) );
NAND2x1_ASAP7_75t_L g672 ( .A(n_564), .B(n_449), .Y(n_672) );
BUFx6f_ASAP7_75t_L g673 ( .A(n_565), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_573), .A2(n_449), .B(n_95), .Y(n_674) );
OAI22x1_ASAP7_75t_L g675 ( .A1(n_529), .A2(n_17), .B1(n_18), .B2(n_19), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_566), .B(n_19), .Y(n_676) );
AND2x4_ASAP7_75t_L g677 ( .A(n_565), .B(n_20), .Y(n_677) );
OAI21x1_ASAP7_75t_L g678 ( .A1(n_516), .A2(n_96), .B(n_94), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_504), .B(n_22), .Y(n_679) );
INVx4_ASAP7_75t_L g680 ( .A(n_519), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_505), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_508), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_580), .Y(n_683) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_572), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_572), .A2(n_449), .B(n_99), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_561), .A2(n_449), .B1(n_24), .B2(n_25), .Y(n_686) );
NOR3xp33_ASAP7_75t_SL g687 ( .A(n_576), .B(n_581), .C(n_579), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_583), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_519), .B(n_23), .Y(n_689) );
INVx4_ASAP7_75t_L g690 ( .A(n_519), .Y(n_690) );
OR2x6_ASAP7_75t_L g691 ( .A(n_572), .B(n_26), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_570), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_577), .B(n_26), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_528), .A2(n_27), .B1(n_28), .B2(n_29), .Y(n_694) );
INVxp67_ASAP7_75t_L g695 ( .A(n_507), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_517), .B(n_27), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_528), .A2(n_28), .B1(n_29), .B2(n_30), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_528), .B(n_31), .Y(n_698) );
CKINVDCx5p33_ASAP7_75t_R g699 ( .A(n_503), .Y(n_699) );
BUFx6f_ASAP7_75t_L g700 ( .A(n_571), .Y(n_700) );
OAI22xp5_ASAP7_75t_SL g701 ( .A1(n_549), .A2(n_32), .B1(n_33), .B2(n_34), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_553), .Y(n_702) );
BUFx2_ASAP7_75t_L g703 ( .A(n_528), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_501), .B(n_32), .Y(n_704) );
AO32x2_ASAP7_75t_L g705 ( .A1(n_549), .A2(n_34), .A3(n_35), .B1(n_37), .B2(n_38), .Y(n_705) );
BUFx6f_ASAP7_75t_SL g706 ( .A(n_528), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_501), .B(n_35), .Y(n_707) );
NOR3xp33_ASAP7_75t_L g708 ( .A(n_549), .B(n_39), .C(n_40), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_543), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_543), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_501), .B(n_41), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_501), .B(n_42), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_528), .A2(n_42), .B1(n_43), .B2(n_44), .Y(n_713) );
INVx5_ASAP7_75t_L g714 ( .A(n_528), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_553), .Y(n_715) );
O2A1O1Ixp5_ASAP7_75t_L g716 ( .A1(n_569), .A2(n_174), .B(n_261), .C(n_260), .Y(n_716) );
AND2x4_ASAP7_75t_L g717 ( .A(n_528), .B(n_45), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_590), .B(n_46), .Y(n_718) );
CKINVDCx6p67_ASAP7_75t_R g719 ( .A(n_706), .Y(n_719) );
NAND3xp33_ASAP7_75t_L g720 ( .A(n_664), .B(n_47), .C(n_49), .Y(n_720) );
OR2x2_ASAP7_75t_L g721 ( .A(n_596), .B(n_47), .Y(n_721) );
AND2x4_ASAP7_75t_L g722 ( .A(n_614), .B(n_50), .Y(n_722) );
O2A1O1Ixp5_ASAP7_75t_L g723 ( .A1(n_661), .A2(n_175), .B(n_259), .C(n_256), .Y(n_723) );
OAI21x1_ASAP7_75t_L g724 ( .A1(n_668), .A2(n_678), .B(n_662), .Y(n_724) );
AOI221xp5_ASAP7_75t_L g725 ( .A1(n_635), .A2(n_50), .B1(n_52), .B2(n_53), .C(n_54), .Y(n_725) );
O2A1O1Ixp33_ASAP7_75t_L g726 ( .A1(n_617), .A2(n_53), .B(n_54), .C(n_55), .Y(n_726) );
OAI22x1_ASAP7_75t_L g727 ( .A1(n_717), .A2(n_56), .B1(n_57), .B2(n_58), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_602), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_628), .Y(n_729) );
AO31x2_ASAP7_75t_L g730 ( .A1(n_659), .A2(n_56), .A3(n_57), .B(n_59), .Y(n_730) );
OAI21x1_ASAP7_75t_L g731 ( .A1(n_674), .A2(n_105), .B(n_103), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_605), .Y(n_732) );
OAI21x1_ASAP7_75t_L g733 ( .A1(n_638), .A2(n_180), .B(n_254), .Y(n_733) );
AO31x2_ASAP7_75t_L g734 ( .A1(n_644), .A2(n_60), .A3(n_61), .B(n_62), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_691), .A2(n_60), .B1(n_61), .B2(n_62), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_596), .A2(n_63), .B1(n_64), .B2(n_65), .Y(n_736) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_604), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_702), .B(n_63), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_704), .Y(n_739) );
OAI22xp33_ASAP7_75t_L g740 ( .A1(n_691), .A2(n_64), .B1(n_65), .B2(n_66), .Y(n_740) );
OAI21xp33_ASAP7_75t_L g741 ( .A1(n_603), .A2(n_66), .B(n_67), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_707), .Y(n_742) );
NOR2x1_ASAP7_75t_L g743 ( .A(n_597), .B(n_67), .Y(n_743) );
A2O1A1Ixp33_ASAP7_75t_L g744 ( .A1(n_619), .A2(n_68), .B(n_69), .C(n_70), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g745 ( .A1(n_616), .A2(n_188), .B(n_253), .Y(n_745) );
A2O1A1Ixp33_ASAP7_75t_L g746 ( .A1(n_630), .A2(n_69), .B(n_70), .C(n_71), .Y(n_746) );
AO32x2_ASAP7_75t_L g747 ( .A1(n_701), .A2(n_71), .A3(n_72), .B1(n_73), .B2(n_74), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_711), .Y(n_748) );
A2O1A1Ixp33_ASAP7_75t_L g749 ( .A1(n_598), .A2(n_74), .B(n_77), .C(n_79), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_637), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_611), .A2(n_80), .B1(n_81), .B2(n_82), .Y(n_751) );
INVx5_ASAP7_75t_L g752 ( .A(n_691), .Y(n_752) );
BUFx6f_ASAP7_75t_L g753 ( .A(n_604), .Y(n_753) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_695), .Y(n_754) );
AOI21xp5_ASAP7_75t_L g755 ( .A1(n_656), .A2(n_194), .B(n_250), .Y(n_755) );
AO31x2_ASAP7_75t_L g756 ( .A1(n_645), .A2(n_80), .A3(n_82), .B(n_83), .Y(n_756) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_717), .Y(n_757) );
OAI22xp33_ASAP7_75t_L g758 ( .A1(n_655), .A2(n_83), .B1(n_85), .B2(n_86), .Y(n_758) );
INVx3_ASAP7_75t_L g759 ( .A(n_604), .Y(n_759) );
NOR2xp33_ASAP7_75t_SL g760 ( .A(n_588), .B(n_85), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_712), .Y(n_761) );
HB1xp67_ASAP7_75t_L g762 ( .A(n_699), .Y(n_762) );
AO31x2_ASAP7_75t_L g763 ( .A1(n_592), .A2(n_119), .A3(n_122), .B(n_125), .Y(n_763) );
OAI21xp5_ASAP7_75t_L g764 ( .A1(n_670), .A2(n_128), .B(n_129), .Y(n_764) );
INVx2_ASAP7_75t_SL g765 ( .A(n_652), .Y(n_765) );
INVx2_ASAP7_75t_SL g766 ( .A(n_589), .Y(n_766) );
OAI21xp5_ASAP7_75t_L g767 ( .A1(n_671), .A2(n_130), .B(n_132), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_589), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g769 ( .A1(n_606), .A2(n_135), .B1(n_136), .B2(n_137), .Y(n_769) );
NOR2xp33_ASAP7_75t_L g770 ( .A(n_703), .B(n_140), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_640), .Y(n_771) );
O2A1O1Ixp33_ASAP7_75t_L g772 ( .A1(n_608), .A2(n_141), .B(n_143), .C(n_146), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_591), .Y(n_773) );
OAI22xp5_ASAP7_75t_L g774 ( .A1(n_594), .A2(n_147), .B1(n_148), .B2(n_150), .Y(n_774) );
INVxp67_ASAP7_75t_L g775 ( .A(n_696), .Y(n_775) );
INVx2_ASAP7_75t_SL g776 ( .A(n_714), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_648), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_599), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_601), .Y(n_779) );
INVx3_ASAP7_75t_L g780 ( .A(n_700), .Y(n_780) );
O2A1O1Ixp33_ASAP7_75t_L g781 ( .A1(n_609), .A2(n_154), .B(n_155), .C(n_159), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_642), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_642), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_715), .Y(n_784) );
OAI22xp33_ASAP7_75t_L g785 ( .A1(n_624), .A2(n_160), .B1(n_164), .B2(n_165), .Y(n_785) );
AND2x4_ASAP7_75t_L g786 ( .A(n_620), .B(n_169), .Y(n_786) );
AOI22xp5_ASAP7_75t_L g787 ( .A1(n_698), .A2(n_171), .B1(n_172), .B2(n_176), .Y(n_787) );
OR2x6_ASAP7_75t_L g788 ( .A(n_701), .B(n_177), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_666), .Y(n_789) );
NOR2xp67_ASAP7_75t_L g790 ( .A(n_675), .B(n_178), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_612), .Y(n_791) );
AO31x2_ASAP7_75t_L g792 ( .A1(n_639), .A2(n_189), .A3(n_191), .B(n_197), .Y(n_792) );
BUFx3_ASAP7_75t_L g793 ( .A(n_700), .Y(n_793) );
O2A1O1Ixp33_ASAP7_75t_SL g794 ( .A1(n_646), .A2(n_198), .B(n_199), .C(n_200), .Y(n_794) );
INVx2_ASAP7_75t_L g795 ( .A(n_709), .Y(n_795) );
OR2x2_ASAP7_75t_L g796 ( .A(n_593), .B(n_202), .Y(n_796) );
INVx2_ASAP7_75t_L g797 ( .A(n_710), .Y(n_797) );
INVx1_ASAP7_75t_SL g798 ( .A(n_677), .Y(n_798) );
AOI21xp5_ASAP7_75t_L g799 ( .A1(n_613), .A2(n_203), .B(n_204), .Y(n_799) );
OAI21x1_ASAP7_75t_L g800 ( .A1(n_615), .A2(n_205), .B(n_206), .Y(n_800) );
AO32x2_ASAP7_75t_L g801 ( .A1(n_694), .A2(n_210), .A3(n_215), .B1(n_219), .B2(n_220), .Y(n_801) );
A2O1A1Ixp33_ASAP7_75t_L g802 ( .A1(n_636), .A2(n_221), .B(n_222), .C(n_223), .Y(n_802) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_681), .Y(n_803) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_594), .A2(n_224), .B1(n_225), .B2(n_226), .Y(n_804) );
A2O1A1Ixp33_ASAP7_75t_L g805 ( .A1(n_641), .A2(n_233), .B(n_234), .C(n_235), .Y(n_805) );
NAND3xp33_ASAP7_75t_L g806 ( .A(n_623), .B(n_236), .C(n_240), .Y(n_806) );
O2A1O1Ixp33_ASAP7_75t_L g807 ( .A1(n_634), .A2(n_242), .B(n_243), .C(n_244), .Y(n_807) );
CKINVDCx16_ASAP7_75t_R g808 ( .A(n_632), .Y(n_808) );
AOI21xp5_ASAP7_75t_L g809 ( .A1(n_631), .A2(n_247), .B(n_248), .Y(n_809) );
A2O1A1Ixp33_ASAP7_75t_L g810 ( .A1(n_665), .A2(n_266), .B(n_647), .C(n_676), .Y(n_810) );
AOI21xp5_ASAP7_75t_L g811 ( .A1(n_692), .A2(n_629), .B(n_688), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_679), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_626), .B(n_633), .Y(n_813) );
BUFx2_ASAP7_75t_L g814 ( .A(n_714), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_708), .A2(n_714), .B1(n_607), .B2(n_683), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_595), .A2(n_610), .B1(n_587), .B2(n_663), .Y(n_816) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_594), .A2(n_713), .B1(n_669), .B2(n_618), .Y(n_817) );
NAND3xp33_ASAP7_75t_L g818 ( .A(n_687), .B(n_651), .C(n_625), .Y(n_818) );
O2A1O1Ixp33_ASAP7_75t_L g819 ( .A1(n_697), .A2(n_621), .B(n_622), .C(n_693), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_682), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_658), .A2(n_600), .B1(n_650), .B2(n_649), .Y(n_821) );
AND2x2_ASAP7_75t_L g822 ( .A(n_625), .B(n_705), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_705), .Y(n_823) );
BUFx3_ASAP7_75t_L g824 ( .A(n_653), .Y(n_824) );
A2O1A1Ixp33_ASAP7_75t_L g825 ( .A1(n_716), .A2(n_657), .B(n_643), .C(n_660), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g826 ( .A1(n_684), .A2(n_680), .B1(n_690), .B2(n_653), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_684), .Y(n_827) );
A2O1A1Ixp33_ASAP7_75t_L g828 ( .A1(n_654), .A2(n_685), .B(n_627), .C(n_686), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_705), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_625), .Y(n_830) );
OAI221xp5_ASAP7_75t_L g831 ( .A1(n_673), .A2(n_517), .B1(n_524), .B2(n_562), .C(n_623), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_673), .Y(n_832) );
NAND2x1p5_ASAP7_75t_L g833 ( .A(n_714), .B(n_594), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_602), .Y(n_834) );
AOI21xp5_ASAP7_75t_L g835 ( .A1(n_616), .A2(n_512), .B(n_506), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_590), .B(n_501), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_611), .A2(n_513), .B1(n_567), .B2(n_528), .Y(n_837) );
O2A1O1Ixp33_ASAP7_75t_SL g838 ( .A1(n_664), .A2(n_689), .B(n_667), .C(n_592), .Y(n_838) );
A2O1A1Ixp33_ASAP7_75t_L g839 ( .A1(n_619), .A2(n_630), .B(n_598), .C(n_656), .Y(n_839) );
AOI21xp5_ASAP7_75t_L g840 ( .A1(n_616), .A2(n_512), .B(n_506), .Y(n_840) );
AND2x4_ASAP7_75t_L g841 ( .A(n_614), .B(n_528), .Y(n_841) );
CKINVDCx20_ASAP7_75t_R g842 ( .A(n_588), .Y(n_842) );
AND2x4_ASAP7_75t_L g843 ( .A(n_614), .B(n_528), .Y(n_843) );
CKINVDCx5p33_ASAP7_75t_R g844 ( .A(n_588), .Y(n_844) );
AND2x4_ASAP7_75t_L g845 ( .A(n_614), .B(n_528), .Y(n_845) );
BUFx2_ASAP7_75t_L g846 ( .A(n_596), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_590), .B(n_501), .Y(n_847) );
AND2x2_ASAP7_75t_L g848 ( .A(n_596), .B(n_517), .Y(n_848) );
OAI22xp5_ASAP7_75t_L g849 ( .A1(n_691), .A2(n_461), .B1(n_717), .B2(n_550), .Y(n_849) );
OAI21xp5_ASAP7_75t_L g850 ( .A1(n_656), .A2(n_616), .B(n_619), .Y(n_850) );
CKINVDCx20_ASAP7_75t_R g851 ( .A(n_588), .Y(n_851) );
OR2x2_ASAP7_75t_L g852 ( .A(n_596), .B(n_418), .Y(n_852) );
NAND2xp33_ASAP7_75t_L g853 ( .A(n_604), .B(n_571), .Y(n_853) );
INVx5_ASAP7_75t_L g854 ( .A(n_691), .Y(n_854) );
BUFx6f_ASAP7_75t_L g855 ( .A(n_604), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_602), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_602), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_590), .B(n_501), .Y(n_858) );
O2A1O1Ixp5_ASAP7_75t_L g859 ( .A1(n_661), .A2(n_672), .B(n_667), .C(n_664), .Y(n_859) );
INVxp67_ASAP7_75t_L g860 ( .A(n_596), .Y(n_860) );
OAI21xp5_ASAP7_75t_L g861 ( .A1(n_656), .A2(n_616), .B(n_619), .Y(n_861) );
AOI21xp5_ASAP7_75t_L g862 ( .A1(n_838), .A2(n_840), .B(n_835), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_728), .B(n_732), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_834), .B(n_856), .Y(n_864) );
OAI22xp33_ASAP7_75t_L g865 ( .A1(n_788), .A2(n_849), .B1(n_831), .B2(n_760), .Y(n_865) );
AND2x2_ASAP7_75t_L g866 ( .A(n_848), .B(n_846), .Y(n_866) );
AOI22xp33_ASAP7_75t_SL g867 ( .A1(n_788), .A2(n_752), .B1(n_854), .B2(n_722), .Y(n_867) );
AND2x2_ASAP7_75t_L g868 ( .A(n_860), .B(n_836), .Y(n_868) );
A2O1A1Ixp33_ASAP7_75t_L g869 ( .A1(n_790), .A2(n_819), .B(n_839), .C(n_857), .Y(n_869) );
OA21x2_ASAP7_75t_L g870 ( .A1(n_823), .A2(n_829), .B(n_800), .Y(n_870) );
AOI21xp5_ASAP7_75t_L g871 ( .A1(n_825), .A2(n_811), .B(n_850), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_813), .A2(n_789), .B1(n_837), .B2(n_779), .Y(n_872) );
NOR2xp33_ASAP7_75t_L g873 ( .A(n_852), .B(n_841), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_739), .A2(n_742), .B1(n_748), .B2(n_761), .Y(n_874) );
O2A1O1Ixp33_ASAP7_75t_L g875 ( .A1(n_758), .A2(n_749), .B(n_746), .C(n_744), .Y(n_875) );
OAI221xp5_ASAP7_75t_L g876 ( .A1(n_815), .A2(n_775), .B1(n_816), .B2(n_812), .C(n_847), .Y(n_876) );
NOR2xp33_ASAP7_75t_L g877 ( .A(n_841), .B(n_843), .Y(n_877) );
AOI21xp5_ASAP7_75t_L g878 ( .A1(n_861), .A2(n_859), .B(n_828), .Y(n_878) );
OA21x2_ASAP7_75t_L g879 ( .A1(n_810), .A2(n_733), .B(n_767), .Y(n_879) );
INVx4_ASAP7_75t_L g880 ( .A(n_752), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_777), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_750), .Y(n_882) );
O2A1O1Ixp33_ASAP7_75t_L g883 ( .A1(n_817), .A2(n_726), .B(n_740), .C(n_735), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_858), .B(n_773), .Y(n_884) );
HB1xp67_ASAP7_75t_L g885 ( .A(n_754), .Y(n_885) );
NOR2xp33_ASAP7_75t_L g886 ( .A(n_843), .B(n_845), .Y(n_886) );
OR2x2_ASAP7_75t_L g887 ( .A(n_721), .B(n_762), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_771), .Y(n_888) );
AND2x2_ASAP7_75t_L g889 ( .A(n_722), .B(n_845), .Y(n_889) );
OR2x6_ASAP7_75t_L g890 ( .A(n_786), .B(n_833), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_784), .Y(n_891) );
AO21x2_ASAP7_75t_L g892 ( .A1(n_822), .A2(n_720), .B(n_764), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_791), .Y(n_893) );
AOI21xp5_ASAP7_75t_L g894 ( .A1(n_745), .A2(n_796), .B(n_794), .Y(n_894) );
INVx1_ASAP7_75t_SL g895 ( .A(n_798), .Y(n_895) );
AOI221xp5_ASAP7_75t_L g896 ( .A1(n_782), .A2(n_783), .B1(n_830), .B2(n_768), .C(n_741), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_757), .A2(n_752), .B1(n_854), .B2(n_818), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_820), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_854), .A2(n_766), .B1(n_727), .B2(n_743), .Y(n_899) );
INVx2_ASAP7_75t_L g900 ( .A(n_778), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_795), .B(n_797), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_718), .Y(n_902) );
A2O1A1Ixp33_ASAP7_75t_L g903 ( .A1(n_772), .A2(n_781), .B(n_806), .C(n_807), .Y(n_903) );
HB1xp67_ASAP7_75t_L g904 ( .A(n_851), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_738), .B(n_821), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_786), .B(n_770), .Y(n_906) );
BUFx12f_ASAP7_75t_L g907 ( .A(n_844), .Y(n_907) );
AOI21xp5_ASAP7_75t_L g908 ( .A1(n_809), .A2(n_802), .B(n_755), .Y(n_908) );
AO31x2_ASAP7_75t_L g909 ( .A1(n_805), .A2(n_799), .A3(n_804), .B(n_774), .Y(n_909) );
OAI22xp5_ASAP7_75t_L g910 ( .A1(n_751), .A2(n_736), .B1(n_725), .B2(n_787), .Y(n_910) );
OR2x6_ASAP7_75t_L g911 ( .A(n_765), .B(n_855), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_808), .A2(n_719), .B1(n_814), .B2(n_776), .Y(n_912) );
BUFx6f_ASAP7_75t_L g913 ( .A(n_737), .Y(n_913) );
INVx2_ASAP7_75t_L g914 ( .A(n_827), .Y(n_914) );
NOR2xp33_ASAP7_75t_L g915 ( .A(n_803), .B(n_793), .Y(n_915) );
A2O1A1Ixp33_ASAP7_75t_L g916 ( .A1(n_769), .A2(n_723), .B(n_731), .C(n_853), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_832), .B(n_855), .Y(n_917) );
O2A1O1Ixp33_ASAP7_75t_L g918 ( .A1(n_785), .A2(n_780), .B(n_759), .C(n_826), .Y(n_918) );
AO31x2_ASAP7_75t_L g919 ( .A1(n_763), .A2(n_792), .A3(n_734), .B(n_756), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_753), .B(n_855), .Y(n_920) );
AO21x2_ASAP7_75t_L g921 ( .A1(n_792), .A2(n_763), .B(n_801), .Y(n_921) );
BUFx3_ASAP7_75t_L g922 ( .A(n_824), .Y(n_922) );
OAI221xp5_ASAP7_75t_L g923 ( .A1(n_780), .A2(n_747), .B1(n_801), .B2(n_734), .C(n_792), .Y(n_923) );
OR2x2_ASAP7_75t_L g924 ( .A(n_734), .B(n_756), .Y(n_924) );
OAI22xp5_ASAP7_75t_L g925 ( .A1(n_801), .A2(n_756), .B1(n_730), .B2(n_763), .Y(n_925) );
BUFx2_ASAP7_75t_L g926 ( .A(n_730), .Y(n_926) );
XOR2xp5_ASAP7_75t_L g927 ( .A(n_842), .B(n_851), .Y(n_927) );
A2O1A1Ixp33_ASAP7_75t_L g928 ( .A1(n_790), .A2(n_819), .B(n_839), .C(n_732), .Y(n_928) );
O2A1O1Ixp33_ASAP7_75t_L g929 ( .A1(n_831), .A2(n_813), .B(n_469), .C(n_758), .Y(n_929) );
AND2x4_ASAP7_75t_L g930 ( .A(n_728), .B(n_732), .Y(n_930) );
OA21x2_ASAP7_75t_L g931 ( .A1(n_724), .A2(n_829), .B(n_823), .Y(n_931) );
HB1xp67_ASAP7_75t_L g932 ( .A(n_846), .Y(n_932) );
AND2x2_ASAP7_75t_L g933 ( .A(n_848), .B(n_517), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_728), .B(n_856), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_777), .Y(n_935) );
INVx2_ASAP7_75t_SL g936 ( .A(n_846), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_777), .Y(n_937) );
OAI21xp5_ASAP7_75t_L g938 ( .A1(n_811), .A2(n_839), .B(n_835), .Y(n_938) );
OAI222xp33_ASAP7_75t_L g939 ( .A1(n_788), .A2(n_849), .B1(n_831), .B2(n_666), .C1(n_691), .C2(n_497), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_728), .B(n_732), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_777), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_777), .Y(n_942) );
AND2x4_ASAP7_75t_L g943 ( .A(n_728), .B(n_732), .Y(n_943) );
AO31x2_ASAP7_75t_L g944 ( .A1(n_823), .A2(n_829), .A3(n_828), .B(n_810), .Y(n_944) );
INVx1_ASAP7_75t_L g945 ( .A(n_777), .Y(n_945) );
AND2x4_ASAP7_75t_L g946 ( .A(n_728), .B(n_732), .Y(n_946) );
INVx1_ASAP7_75t_L g947 ( .A(n_777), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_777), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_728), .B(n_856), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_728), .B(n_856), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g951 ( .A(n_728), .B(n_856), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_728), .B(n_856), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_788), .A2(n_831), .B1(n_813), .B2(n_611), .Y(n_953) );
AOI21xp33_ASAP7_75t_L g954 ( .A1(n_817), .A2(n_849), .B(n_789), .Y(n_954) );
NAND2xp5_ASAP7_75t_SL g955 ( .A(n_752), .B(n_854), .Y(n_955) );
NAND2x1p5_ASAP7_75t_L g956 ( .A(n_752), .B(n_854), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_777), .Y(n_957) );
INVx1_ASAP7_75t_L g958 ( .A(n_777), .Y(n_958) );
INVx2_ASAP7_75t_L g959 ( .A(n_729), .Y(n_959) );
OA21x2_ASAP7_75t_L g960 ( .A1(n_724), .A2(n_829), .B(n_823), .Y(n_960) );
HB1xp67_ASAP7_75t_L g961 ( .A(n_846), .Y(n_961) );
O2A1O1Ixp5_ASAP7_75t_SL g962 ( .A1(n_823), .A2(n_829), .B(n_789), .C(n_830), .Y(n_962) );
OA21x2_ASAP7_75t_L g963 ( .A1(n_724), .A2(n_829), .B(n_823), .Y(n_963) );
OAI21x1_ASAP7_75t_SL g964 ( .A1(n_849), .A2(n_767), .B(n_764), .Y(n_964) );
NOR2xp33_ASAP7_75t_L g965 ( .A(n_813), .B(n_513), .Y(n_965) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_728), .B(n_856), .Y(n_966) );
AOI21xp33_ASAP7_75t_SL g967 ( .A1(n_808), .A2(n_788), .B(n_701), .Y(n_967) );
AOI221xp5_ASAP7_75t_L g968 ( .A1(n_773), .A2(n_469), .B1(n_549), .B2(n_517), .C(n_831), .Y(n_968) );
INVx2_ASAP7_75t_L g969 ( .A(n_729), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_728), .B(n_856), .Y(n_970) );
OAI21x1_ASAP7_75t_SL g971 ( .A1(n_849), .A2(n_767), .B(n_764), .Y(n_971) );
INVx3_ASAP7_75t_L g972 ( .A(n_737), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_891), .Y(n_973) );
AO21x2_ASAP7_75t_L g974 ( .A1(n_878), .A2(n_871), .B(n_938), .Y(n_974) );
AOI221xp5_ASAP7_75t_L g975 ( .A1(n_967), .A2(n_968), .B1(n_929), .B2(n_965), .C(n_876), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_881), .Y(n_976) );
BUFx2_ASAP7_75t_L g977 ( .A(n_890), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_893), .Y(n_978) );
OAI211xp5_ASAP7_75t_SL g979 ( .A1(n_912), .A2(n_887), .B(n_953), .C(n_884), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_935), .Y(n_980) );
INVx2_ASAP7_75t_L g981 ( .A(n_931), .Y(n_981) );
BUFx3_ASAP7_75t_L g982 ( .A(n_922), .Y(n_982) );
OR2x2_ASAP7_75t_L g983 ( .A(n_863), .B(n_864), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_933), .B(n_868), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_937), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_941), .Y(n_986) );
INVx3_ASAP7_75t_L g987 ( .A(n_913), .Y(n_987) );
INVx1_ASAP7_75t_L g988 ( .A(n_942), .Y(n_988) );
OR2x2_ASAP7_75t_L g989 ( .A(n_863), .B(n_864), .Y(n_989) );
HB1xp67_ASAP7_75t_L g990 ( .A(n_885), .Y(n_990) );
OR2x6_ASAP7_75t_L g991 ( .A(n_890), .B(n_956), .Y(n_991) );
AND2x2_ASAP7_75t_L g992 ( .A(n_930), .B(n_943), .Y(n_992) );
OA21x2_ASAP7_75t_L g993 ( .A1(n_938), .A2(n_925), .B(n_862), .Y(n_993) );
OAI21xp33_ASAP7_75t_L g994 ( .A1(n_869), .A2(n_928), .B(n_867), .Y(n_994) );
OA21x2_ASAP7_75t_L g995 ( .A1(n_925), .A2(n_926), .B(n_924), .Y(n_995) );
INVxp67_ASAP7_75t_SL g996 ( .A(n_934), .Y(n_996) );
INVx2_ASAP7_75t_SL g997 ( .A(n_890), .Y(n_997) );
BUFx2_ASAP7_75t_L g998 ( .A(n_946), .Y(n_998) );
INVxp67_ASAP7_75t_SL g999 ( .A(n_934), .Y(n_999) );
AOI21xp5_ASAP7_75t_SL g1000 ( .A1(n_865), .A2(n_906), .B(n_916), .Y(n_1000) );
AO21x2_ASAP7_75t_L g1001 ( .A1(n_923), .A2(n_964), .B(n_971), .Y(n_1001) );
BUFx6f_ASAP7_75t_L g1002 ( .A(n_913), .Y(n_1002) );
OR2x2_ASAP7_75t_L g1003 ( .A(n_949), .B(n_950), .Y(n_1003) );
OAI222xp33_ASAP7_75t_L g1004 ( .A1(n_906), .A2(n_899), .B1(n_910), .B2(n_883), .C1(n_956), .C2(n_872), .Y(n_1004) );
INVx3_ASAP7_75t_L g1005 ( .A(n_946), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_945), .Y(n_1006) );
OR2x6_ASAP7_75t_L g1007 ( .A(n_880), .B(n_955), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_947), .Y(n_1008) );
BUFx3_ASAP7_75t_L g1009 ( .A(n_911), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_949), .B(n_950), .Y(n_1010) );
INVx3_ASAP7_75t_L g1011 ( .A(n_880), .Y(n_1011) );
OR2x6_ASAP7_75t_L g1012 ( .A(n_918), .B(n_889), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_948), .Y(n_1013) );
AOI221xp5_ASAP7_75t_L g1014 ( .A1(n_939), .A2(n_874), .B1(n_954), .B2(n_884), .C(n_966), .Y(n_1014) );
OAI21xp5_ASAP7_75t_L g1015 ( .A1(n_910), .A2(n_875), .B(n_905), .Y(n_1015) );
AOI21xp33_ASAP7_75t_SL g1016 ( .A1(n_927), .A2(n_904), .B(n_915), .Y(n_1016) );
BUFx4f_ASAP7_75t_L g1017 ( .A(n_911), .Y(n_1017) );
HB1xp67_ASAP7_75t_L g1018 ( .A(n_866), .Y(n_1018) );
BUFx2_ASAP7_75t_R g1019 ( .A(n_951), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_957), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_958), .Y(n_1021) );
INVx1_ASAP7_75t_L g1022 ( .A(n_882), .Y(n_1022) );
AOI22xp33_ASAP7_75t_SL g1023 ( .A1(n_932), .A2(n_961), .B1(n_936), .B2(n_952), .Y(n_1023) );
OA21x2_ASAP7_75t_L g1024 ( .A1(n_894), .A2(n_908), .B(n_903), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_888), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_951), .Y(n_1026) );
BUFx2_ASAP7_75t_SL g1027 ( .A(n_959), .Y(n_1027) );
OA21x2_ASAP7_75t_L g1028 ( .A1(n_954), .A2(n_896), .B(n_905), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_952), .Y(n_1029) );
OAI21xp5_ASAP7_75t_L g1030 ( .A1(n_962), .A2(n_902), .B(n_970), .Y(n_1030) );
OR2x6_ASAP7_75t_L g1031 ( .A(n_911), .B(n_920), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_969), .B(n_966), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_970), .B(n_900), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_873), .A2(n_940), .B1(n_898), .B2(n_877), .Y(n_1034) );
BUFx6f_ASAP7_75t_L g1035 ( .A(n_920), .Y(n_1035) );
INVx2_ASAP7_75t_L g1036 ( .A(n_960), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g1037 ( .A1(n_886), .A2(n_895), .B1(n_921), .B2(n_897), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_895), .B(n_901), .Y(n_1038) );
OR2x2_ASAP7_75t_L g1039 ( .A(n_917), .B(n_919), .Y(n_1039) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_914), .B(n_919), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_919), .B(n_972), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_963), .Y(n_1042) );
OA21x2_ASAP7_75t_L g1043 ( .A1(n_921), .A2(n_944), .B(n_892), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_963), .Y(n_1044) );
INVx2_ASAP7_75t_L g1045 ( .A(n_870), .Y(n_1045) );
BUFx2_ASAP7_75t_L g1046 ( .A(n_907), .Y(n_1046) );
OA21x2_ASAP7_75t_L g1047 ( .A1(n_944), .A2(n_892), .B(n_879), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_944), .Y(n_1048) );
AOI21xp5_ASAP7_75t_SL g1049 ( .A1(n_909), .A2(n_849), .B(n_691), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_909), .B(n_930), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_909), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_891), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_891), .Y(n_1053) );
INVx2_ASAP7_75t_SL g1054 ( .A(n_890), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_891), .Y(n_1055) );
HB1xp67_ASAP7_75t_L g1056 ( .A(n_1039), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_1050), .B(n_1040), .Y(n_1057) );
HB1xp67_ASAP7_75t_L g1058 ( .A(n_1039), .Y(n_1058) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_1015), .B(n_1026), .Y(n_1059) );
AND2x4_ASAP7_75t_L g1060 ( .A(n_1050), .B(n_1041), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1040), .Y(n_1061) );
INVx5_ASAP7_75t_L g1062 ( .A(n_991), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_1032), .B(n_1033), .Y(n_1063) );
INVxp67_ASAP7_75t_SL g1064 ( .A(n_996), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1042), .Y(n_1065) );
NAND2xp5_ASAP7_75t_L g1066 ( .A(n_1029), .B(n_999), .Y(n_1066) );
OAI321xp33_ASAP7_75t_L g1067 ( .A1(n_994), .A2(n_975), .A3(n_979), .B1(n_1014), .B2(n_1037), .C(n_1030), .Y(n_1067) );
BUFx3_ASAP7_75t_L g1068 ( .A(n_1017), .Y(n_1068) );
INVx1_ASAP7_75t_L g1069 ( .A(n_1044), .Y(n_1069) );
AND2x4_ASAP7_75t_L g1070 ( .A(n_1051), .B(n_1001), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_981), .Y(n_1071) );
OR2x2_ASAP7_75t_L g1072 ( .A(n_983), .B(n_989), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_1032), .B(n_1033), .Y(n_1073) );
INVxp67_ASAP7_75t_L g1074 ( .A(n_1027), .Y(n_1074) );
BUFx3_ASAP7_75t_L g1075 ( .A(n_1017), .Y(n_1075) );
OR2x2_ASAP7_75t_L g1076 ( .A(n_1003), .B(n_1038), .Y(n_1076) );
OAI221xp5_ASAP7_75t_L g1077 ( .A1(n_1034), .A2(n_1023), .B1(n_1010), .B2(n_991), .C(n_1049), .Y(n_1077) );
HB1xp67_ASAP7_75t_L g1078 ( .A(n_1035), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_1048), .B(n_974), .Y(n_1079) );
BUFx3_ASAP7_75t_L g1080 ( .A(n_1017), .Y(n_1080) );
AO21x2_ASAP7_75t_L g1081 ( .A1(n_974), .A2(n_1045), .B(n_1036), .Y(n_1081) );
NAND2xp5_ASAP7_75t_L g1082 ( .A(n_1028), .B(n_973), .Y(n_1082) );
OR2x2_ASAP7_75t_L g1083 ( .A(n_1018), .B(n_984), .Y(n_1083) );
AND2x4_ASAP7_75t_L g1084 ( .A(n_1001), .B(n_1035), .Y(n_1084) );
OR2x2_ASAP7_75t_L g1085 ( .A(n_990), .B(n_998), .Y(n_1085) );
OR2x2_ASAP7_75t_L g1086 ( .A(n_1005), .B(n_1034), .Y(n_1086) );
HB1xp67_ASAP7_75t_L g1087 ( .A(n_1035), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_1012), .A2(n_992), .B1(n_1005), .B2(n_991), .Y(n_1088) );
OR2x2_ASAP7_75t_L g1089 ( .A(n_1005), .B(n_1012), .Y(n_1089) );
AO21x2_ASAP7_75t_L g1090 ( .A1(n_1000), .A2(n_1001), .B(n_1004), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_992), .B(n_1055), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_976), .B(n_1013), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_978), .B(n_1006), .Y(n_1093) );
HB1xp67_ASAP7_75t_L g1094 ( .A(n_1031), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_995), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_995), .Y(n_1096) );
INVx1_ASAP7_75t_L g1097 ( .A(n_995), .Y(n_1097) );
INVx1_ASAP7_75t_L g1098 ( .A(n_980), .Y(n_1098) );
INVx2_ASAP7_75t_L g1099 ( .A(n_993), .Y(n_1099) );
AND2x4_ASAP7_75t_L g1100 ( .A(n_1012), .B(n_987), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1057), .B(n_1043), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_1057), .B(n_1043), .Y(n_1102) );
HB1xp67_ASAP7_75t_L g1103 ( .A(n_1064), .Y(n_1103) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1065), .Y(n_1104) );
BUFx3_ASAP7_75t_L g1105 ( .A(n_1084), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_1061), .B(n_1043), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_1061), .B(n_1047), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1060), .B(n_1047), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_1060), .B(n_1047), .Y(n_1109) );
OR2x2_ASAP7_75t_L g1110 ( .A(n_1056), .B(n_1037), .Y(n_1110) );
NOR2x1_ASAP7_75t_L g1111 ( .A(n_1077), .B(n_1011), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_1060), .B(n_1024), .Y(n_1112) );
NOR2x1_ASAP7_75t_L g1113 ( .A(n_1077), .B(n_1011), .Y(n_1113) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1059), .B(n_1028), .Y(n_1114) );
NAND2xp5_ASAP7_75t_L g1115 ( .A(n_1059), .B(n_1028), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1079), .B(n_1024), .Y(n_1116) );
AND2x4_ASAP7_75t_L g1117 ( .A(n_1084), .B(n_1002), .Y(n_1117) );
NAND2x1p5_ASAP7_75t_L g1118 ( .A(n_1062), .B(n_987), .Y(n_1118) );
NOR2xp33_ASAP7_75t_L g1119 ( .A(n_1074), .B(n_1019), .Y(n_1119) );
NOR2xp67_ASAP7_75t_L g1120 ( .A(n_1062), .B(n_1011), .Y(n_1120) );
INVx2_ASAP7_75t_L g1121 ( .A(n_1081), .Y(n_1121) );
OR2x2_ASAP7_75t_L g1122 ( .A(n_1056), .B(n_1012), .Y(n_1122) );
AND2x2_ASAP7_75t_L g1123 ( .A(n_1079), .B(n_1024), .Y(n_1123) );
INVxp67_ASAP7_75t_L g1124 ( .A(n_1064), .Y(n_1124) );
NAND2xp5_ASAP7_75t_L g1125 ( .A(n_1066), .B(n_1020), .Y(n_1125) );
INVx1_ASAP7_75t_SL g1126 ( .A(n_1085), .Y(n_1126) );
NAND2xp5_ASAP7_75t_L g1127 ( .A(n_1066), .B(n_1021), .Y(n_1127) );
HB1xp67_ASAP7_75t_L g1128 ( .A(n_1058), .Y(n_1128) );
HB1xp67_ASAP7_75t_L g1129 ( .A(n_1058), .Y(n_1129) );
NAND2xp5_ASAP7_75t_L g1130 ( .A(n_1063), .B(n_1008), .Y(n_1130) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1069), .Y(n_1131) );
HB1xp67_ASAP7_75t_L g1132 ( .A(n_1071), .Y(n_1132) );
OR2x2_ASAP7_75t_L g1133 ( .A(n_1082), .B(n_1053), .Y(n_1133) );
AND2x4_ASAP7_75t_SL g1134 ( .A(n_1100), .B(n_991), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_1099), .B(n_1000), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1101), .B(n_1070), .Y(n_1136) );
INVx1_ASAP7_75t_SL g1137 ( .A(n_1103), .Y(n_1137) );
NAND2xp5_ASAP7_75t_L g1138 ( .A(n_1106), .B(n_1082), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1101), .B(n_1070), .Y(n_1139) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1104), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1101), .B(n_1070), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1102), .B(n_1070), .Y(n_1142) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1104), .Y(n_1143) );
OR2x2_ASAP7_75t_L g1144 ( .A(n_1126), .B(n_1076), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1102), .B(n_1063), .Y(n_1145) );
NAND2xp5_ASAP7_75t_L g1146 ( .A(n_1126), .B(n_1073), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_1102), .B(n_1073), .Y(n_1147) );
NAND2xp5_ASAP7_75t_L g1148 ( .A(n_1106), .B(n_1098), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1108), .B(n_1095), .Y(n_1149) );
OR2x2_ASAP7_75t_L g1150 ( .A(n_1128), .B(n_1076), .Y(n_1150) );
NAND2xp5_ASAP7_75t_L g1151 ( .A(n_1106), .B(n_1098), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_1108), .B(n_1095), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1153 ( .A(n_1133), .B(n_1092), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1131), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1131), .Y(n_1155) );
NAND2xp5_ASAP7_75t_L g1156 ( .A(n_1130), .B(n_1092), .Y(n_1156) );
OR2x2_ASAP7_75t_L g1157 ( .A(n_1128), .B(n_1083), .Y(n_1157) );
OR2x2_ASAP7_75t_L g1158 ( .A(n_1129), .B(n_1083), .Y(n_1158) );
OAI22xp5_ASAP7_75t_L g1159 ( .A1(n_1111), .A2(n_1088), .B1(n_1062), .B2(n_1074), .Y(n_1159) );
INVx2_ASAP7_75t_SL g1160 ( .A(n_1103), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1108), .B(n_1096), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1109), .B(n_1096), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g1163 ( .A(n_1133), .B(n_1093), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1109), .B(n_1097), .Y(n_1164) );
NOR2xp33_ASAP7_75t_L g1165 ( .A(n_1119), .B(n_1016), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1109), .B(n_1097), .Y(n_1166) );
HB1xp67_ASAP7_75t_L g1167 ( .A(n_1129), .Y(n_1167) );
INVxp67_ASAP7_75t_L g1168 ( .A(n_1125), .Y(n_1168) );
HB1xp67_ASAP7_75t_L g1169 ( .A(n_1124), .Y(n_1169) );
AND2x4_ASAP7_75t_SL g1170 ( .A(n_1117), .B(n_1100), .Y(n_1170) );
INVx2_ASAP7_75t_L g1171 ( .A(n_1121), .Y(n_1171) );
NAND5xp2_ASAP7_75t_L g1172 ( .A(n_1165), .B(n_1088), .C(n_1067), .D(n_1118), .E(n_1135), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1140), .Y(n_1173) );
INVx3_ASAP7_75t_L g1174 ( .A(n_1171), .Y(n_1174) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1157), .Y(n_1175) );
OR2x2_ASAP7_75t_L g1176 ( .A(n_1144), .B(n_1110), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1145), .B(n_1112), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1145), .B(n_1112), .Y(n_1178) );
AOI22xp5_ASAP7_75t_L g1179 ( .A1(n_1159), .A2(n_1113), .B1(n_1112), .B2(n_1134), .Y(n_1179) );
OAI21xp5_ASAP7_75t_L g1180 ( .A1(n_1159), .A2(n_1120), .B(n_1067), .Y(n_1180) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1157), .Y(n_1181) );
NAND2xp5_ASAP7_75t_SL g1182 ( .A(n_1160), .B(n_1062), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1147), .B(n_1116), .Y(n_1183) );
AND2x4_ASAP7_75t_L g1184 ( .A(n_1136), .B(n_1105), .Y(n_1184) );
OR2x2_ASAP7_75t_L g1185 ( .A(n_1144), .B(n_1110), .Y(n_1185) );
NAND2xp5_ASAP7_75t_L g1186 ( .A(n_1168), .B(n_1130), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1147), .B(n_1116), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1140), .Y(n_1188) );
NAND2xp5_ASAP7_75t_L g1189 ( .A(n_1148), .B(n_1107), .Y(n_1189) );
AOI22xp5_ASAP7_75t_L g1190 ( .A1(n_1153), .A2(n_1134), .B1(n_1090), .B2(n_1086), .Y(n_1190) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1148), .B(n_1107), .Y(n_1191) );
OR2x2_ASAP7_75t_L g1192 ( .A(n_1158), .B(n_1110), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1143), .Y(n_1193) );
A2O1A1Ixp33_ASAP7_75t_L g1194 ( .A1(n_1170), .A2(n_1134), .B(n_1062), .C(n_982), .Y(n_1194) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1136), .B(n_1116), .Y(n_1195) );
INVx2_ASAP7_75t_SL g1196 ( .A(n_1160), .Y(n_1196) );
INVx1_ASAP7_75t_SL g1197 ( .A(n_1146), .Y(n_1197) );
INVx1_ASAP7_75t_SL g1198 ( .A(n_1150), .Y(n_1198) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1175), .Y(n_1199) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1181), .Y(n_1200) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1173), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1173), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1195), .B(n_1139), .Y(n_1203) );
AOI22x1_ASAP7_75t_SL g1204 ( .A1(n_1198), .A2(n_1137), .B1(n_1046), .B2(n_1062), .Y(n_1204) );
AOI332xp33_ASAP7_75t_L g1205 ( .A1(n_1190), .A2(n_1156), .A3(n_1153), .B1(n_1163), .B2(n_1091), .B3(n_1149), .C1(n_1152), .C2(n_1166), .Y(n_1205) );
NOR2xp33_ASAP7_75t_L g1206 ( .A(n_1186), .B(n_1163), .Y(n_1206) );
OR2x2_ASAP7_75t_L g1207 ( .A(n_1192), .B(n_1138), .Y(n_1207) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1188), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1188), .Y(n_1209) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1193), .Y(n_1210) );
OR2x2_ASAP7_75t_L g1211 ( .A(n_1192), .B(n_1138), .Y(n_1211) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1193), .Y(n_1212) );
OAI22xp5_ASAP7_75t_L g1213 ( .A1(n_1194), .A2(n_1122), .B1(n_1139), .B2(n_1141), .Y(n_1213) );
A2O1A1Ixp33_ASAP7_75t_L g1214 ( .A1(n_1180), .A2(n_1170), .B(n_1080), .C(n_1075), .Y(n_1214) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1176), .Y(n_1215) );
AOI21xp33_ASAP7_75t_SL g1216 ( .A1(n_1179), .A2(n_1169), .B(n_1167), .Y(n_1216) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1176), .Y(n_1217) );
NOR2xp33_ASAP7_75t_L g1218 ( .A(n_1196), .B(n_1151), .Y(n_1218) );
AOI22xp5_ASAP7_75t_L g1219 ( .A1(n_1197), .A2(n_1149), .B1(n_1152), .B2(n_1166), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1215), .Y(n_1220) );
AOI322xp5_ASAP7_75t_L g1221 ( .A1(n_1206), .A2(n_1183), .A3(n_1187), .B1(n_1177), .B2(n_1178), .C1(n_1195), .C2(n_1189), .Y(n_1221) );
OAI21xp33_ASAP7_75t_L g1222 ( .A1(n_1216), .A2(n_1172), .B(n_1185), .Y(n_1222) );
AOI22xp5_ASAP7_75t_L g1223 ( .A1(n_1213), .A2(n_1164), .B1(n_1162), .B2(n_1161), .Y(n_1223) );
OAI22xp33_ASAP7_75t_SL g1224 ( .A1(n_1219), .A2(n_1182), .B1(n_1196), .B2(n_1185), .Y(n_1224) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1217), .Y(n_1225) );
AOI32xp33_ASAP7_75t_L g1226 ( .A1(n_1218), .A2(n_1184), .A3(n_1187), .B1(n_1183), .B2(n_1177), .Y(n_1226) );
NAND2xp5_ASAP7_75t_L g1227 ( .A(n_1206), .B(n_1178), .Y(n_1227) );
INVx1_ASAP7_75t_SL g1228 ( .A(n_1204), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1201), .Y(n_1229) );
OA21x2_ASAP7_75t_SL g1230 ( .A1(n_1205), .A2(n_1184), .B(n_1137), .Y(n_1230) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1202), .Y(n_1231) );
AOI211xp5_ASAP7_75t_L g1232 ( .A1(n_1228), .A2(n_1214), .B(n_1086), .C(n_1200), .Y(n_1232) );
AOI321xp33_ASAP7_75t_L g1233 ( .A1(n_1222), .A2(n_1199), .A3(n_1127), .B1(n_1125), .B2(n_1123), .C(n_1091), .Y(n_1233) );
OAI211xp5_ASAP7_75t_L g1234 ( .A1(n_1226), .A2(n_982), .B(n_977), .C(n_1127), .Y(n_1234) );
OAI22xp5_ASAP7_75t_L g1235 ( .A1(n_1223), .A2(n_1211), .B1(n_1207), .B2(n_1203), .Y(n_1235) );
INVx2_ASAP7_75t_L g1236 ( .A(n_1229), .Y(n_1236) );
AOI21xp33_ASAP7_75t_SL g1237 ( .A1(n_1224), .A2(n_1090), .B(n_1118), .Y(n_1237) );
AOI221xp5_ASAP7_75t_L g1238 ( .A1(n_1230), .A2(n_1212), .B1(n_1210), .B2(n_1209), .C(n_1208), .Y(n_1238) );
OAI211xp5_ASAP7_75t_SL g1239 ( .A1(n_1221), .A2(n_1191), .B(n_1054), .C(n_997), .Y(n_1239) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1220), .Y(n_1240) );
NOR2xp33_ASAP7_75t_L g1241 ( .A(n_1227), .B(n_1142), .Y(n_1241) );
NAND2xp33_ASAP7_75t_L g1242 ( .A(n_1238), .B(n_1225), .Y(n_1242) );
NAND3xp33_ASAP7_75t_L g1243 ( .A(n_1237), .B(n_1231), .C(n_986), .Y(n_1243) );
NAND4xp75_ASAP7_75t_L g1244 ( .A(n_1240), .B(n_1054), .C(n_997), .D(n_1135), .Y(n_1244) );
NAND5xp2_ASAP7_75t_L g1245 ( .A(n_1233), .B(n_1118), .C(n_1135), .D(n_1115), .E(n_1114), .Y(n_1245) );
O2A1O1Ixp33_ASAP7_75t_L g1246 ( .A1(n_1239), .A2(n_985), .B(n_1052), .C(n_988), .Y(n_1246) );
NAND4xp25_ASAP7_75t_SL g1247 ( .A(n_1232), .B(n_1122), .C(n_1089), .D(n_1072), .Y(n_1247) );
AND5x1_ASAP7_75t_L g1248 ( .A(n_1246), .B(n_1241), .C(n_1234), .D(n_1235), .E(n_1236), .Y(n_1248) );
NOR5xp2_ASAP7_75t_L g1249 ( .A(n_1243), .B(n_1094), .C(n_1132), .D(n_1078), .E(n_1087), .Y(n_1249) );
NAND3x1_ASAP7_75t_L g1250 ( .A(n_1242), .B(n_1247), .C(n_1245), .Y(n_1250) );
BUFx2_ASAP7_75t_L g1251 ( .A(n_1244), .Y(n_1251) );
INVxp33_ASAP7_75t_SL g1252 ( .A(n_1251), .Y(n_1252) );
NAND3xp33_ASAP7_75t_SL g1253 ( .A(n_1249), .B(n_1118), .C(n_1089), .Y(n_1253) );
INVx2_ASAP7_75t_L g1254 ( .A(n_1250), .Y(n_1254) );
A2O1A1Ixp33_ASAP7_75t_L g1255 ( .A1(n_1254), .A2(n_1248), .B(n_1075), .C(n_1068), .Y(n_1255) );
INVx4_ASAP7_75t_L g1256 ( .A(n_1254), .Y(n_1256) );
OAI22xp33_ASAP7_75t_SL g1257 ( .A1(n_1256), .A2(n_1252), .B1(n_1253), .B2(n_1007), .Y(n_1257) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1256), .Y(n_1258) );
OAI22xp5_ASAP7_75t_SL g1259 ( .A1(n_1258), .A2(n_1255), .B1(n_1068), .B2(n_1080), .Y(n_1259) );
A2O1A1O1Ixp25_ASAP7_75t_L g1260 ( .A1(n_1257), .A2(n_1025), .B(n_1022), .C(n_1155), .D(n_1154), .Y(n_1260) );
AOI21xp33_ASAP7_75t_L g1261 ( .A1(n_1259), .A2(n_1007), .B(n_1009), .Y(n_1261) );
OA21x2_ASAP7_75t_L g1262 ( .A1(n_1261), .A2(n_1260), .B(n_1093), .Y(n_1262) );
AOI22xp33_ASAP7_75t_L g1263 ( .A1(n_1262), .A2(n_1174), .B1(n_1105), .B2(n_1090), .Y(n_1263) );
endmodule