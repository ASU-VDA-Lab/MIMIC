module real_jpeg_31724_n_17 (n_8, n_0, n_141, n_2, n_132, n_139, n_10, n_137, n_9, n_12, n_135, n_134, n_6, n_136, n_133, n_11, n_14, n_131, n_138, n_7, n_3, n_5, n_4, n_1, n_140, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_141;
input n_2;
input n_132;
input n_139;
input n_10;
input n_137;
input n_9;
input n_12;
input n_135;
input n_134;
input n_6;
input n_136;
input n_133;
input n_11;
input n_14;
input n_131;
input n_138;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_140;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_0),
.Y(n_99)
);

AOI322xp5_ASAP7_75t_L g122 ( 
.A1(n_0),
.A2(n_94),
.A3(n_96),
.B1(n_101),
.B2(n_123),
.C1(n_125),
.C2(n_141),
.Y(n_122)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_1),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_2),
.B(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_2),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_3),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_3),
.B(n_113),
.Y(n_124)
);

AOI221xp5_ASAP7_75t_L g53 ( 
.A1(n_4),
.A2(n_10),
.B1(n_54),
.B2(n_61),
.C(n_65),
.Y(n_53)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_6),
.B(n_21),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_7),
.B(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_8),
.A2(n_19),
.B1(n_20),
.B2(n_25),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_9),
.B(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_10),
.B(n_54),
.C(n_61),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_11),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_11),
.B(n_103),
.Y(n_121)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_12),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_13),
.B(n_40),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_14),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_14),
.B(n_109),
.Y(n_120)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_26),
.Y(n_17)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_37),
.B(n_129),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_36),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_29),
.B(n_36),
.Y(n_129)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_33),
.B(n_110),
.Y(n_109)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

AOI21x1_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_45),
.B(n_128),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_44),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI31xp33_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_86),
.A3(n_111),
.B(n_118),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_78),
.C(n_79),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_69),
.B(n_77),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_53),
.B1(n_67),
.B2(n_68),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_55),
.B(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_133),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_70),
.B(n_76),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_76),
.Y(n_77)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NOR3xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_100),
.C(n_108),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_119),
.B(n_122),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_94),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NOR3xp33_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_108),
.C(n_124),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_99),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_137),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OA21x2_ASAP7_75t_SL g119 ( 
.A1(n_100),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_107),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_117),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_131),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_132),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_134),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_135),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_136),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_138),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_139),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_140),
.Y(n_114)
);


endmodule