module fake_jpeg_22891_n_29 (n_3, n_2, n_1, n_0, n_4, n_5, n_29);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_29;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_3),
.Y(n_8)
);

INVxp67_ASAP7_75t_SL g9 ( 
.A(n_3),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx4f_ASAP7_75t_SL g11 ( 
.A(n_4),
.Y(n_11)
);

INVx13_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_15),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g14 ( 
.A1(n_11),
.A2(n_5),
.B1(n_0),
.B2(n_2),
.Y(n_14)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

OAI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_10),
.A2(n_9),
.B1(n_11),
.B2(n_8),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_6),
.B(n_7),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_6),
.A2(n_10),
.B1(n_11),
.B2(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_17),
.B(n_18),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

OAI22x1_ASAP7_75t_L g23 ( 
.A1(n_22),
.A2(n_17),
.B1(n_16),
.B2(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_21),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_12),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_25),
.A2(n_22),
.B1(n_20),
.B2(n_23),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_19),
.Y(n_29)
);


endmodule