module real_aes_7104_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g111 ( .A(n_0), .Y(n_111) );
INVx1_ASAP7_75t_L g528 ( .A(n_1), .Y(n_528) );
INVx1_ASAP7_75t_L g150 ( .A(n_2), .Y(n_150) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_3), .A2(n_39), .B1(n_175), .B2(n_474), .Y(n_497) );
AOI21xp33_ASAP7_75t_L g182 ( .A1(n_4), .A2(n_166), .B(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_5), .B(n_164), .Y(n_540) );
AND2x6_ASAP7_75t_L g143 ( .A(n_6), .B(n_144), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_7), .A2(n_253), .B(n_254), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_8), .B(n_40), .Y(n_112) );
INVx1_ASAP7_75t_L g188 ( .A(n_9), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_10), .B(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g135 ( .A(n_11), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_12), .B(n_156), .Y(n_483) );
INVx1_ASAP7_75t_L g259 ( .A(n_13), .Y(n_259) );
INVx1_ASAP7_75t_L g522 ( .A(n_14), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_15), .B(n_131), .Y(n_511) );
AO32x2_ASAP7_75t_L g495 ( .A1(n_16), .A2(n_130), .A3(n_164), .B1(n_476), .B2(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_17), .B(n_175), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_18), .A2(n_102), .B1(n_113), .B2(n_736), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_19), .B(n_171), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_20), .B(n_131), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_21), .A2(n_50), .B1(n_175), .B2(n_474), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_22), .B(n_166), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_23), .A2(n_97), .B1(n_728), .B2(n_729), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_23), .Y(n_729) );
AOI22xp33_ASAP7_75t_SL g475 ( .A1(n_24), .A2(n_75), .B1(n_156), .B2(n_175), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_25), .B(n_175), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_26), .B(n_178), .Y(n_177) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_27), .A2(n_257), .B(n_258), .C(n_260), .Y(n_256) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_28), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_29), .B(n_161), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_30), .B(n_154), .Y(n_153) );
OAI22xp5_ASAP7_75t_SL g120 ( .A1(n_31), .A2(n_87), .B1(n_121), .B2(n_122), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_31), .Y(n_121) );
INVx1_ASAP7_75t_L g203 ( .A(n_32), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_33), .B(n_161), .Y(n_467) );
AOI222xp33_ASAP7_75t_L g440 ( .A1(n_34), .A2(n_441), .B1(n_726), .B2(n_727), .C1(n_730), .C2(n_732), .Y(n_440) );
INVx2_ASAP7_75t_L g141 ( .A(n_35), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_36), .B(n_175), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_37), .B(n_161), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_38), .A2(n_143), .B(n_146), .C(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g201 ( .A(n_41), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_42), .B(n_154), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_43), .B(n_175), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_44), .A2(n_85), .B1(n_223), .B2(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_45), .B(n_175), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_46), .B(n_175), .Y(n_523) );
CKINVDCx16_ASAP7_75t_R g204 ( .A(n_47), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_48), .B(n_527), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_49), .B(n_166), .Y(n_247) );
AOI22xp33_ASAP7_75t_SL g515 ( .A1(n_51), .A2(n_60), .B1(n_156), .B2(n_175), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_52), .A2(n_146), .B1(n_156), .B2(n_199), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_53), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_54), .B(n_175), .Y(n_482) );
CKINVDCx16_ASAP7_75t_R g137 ( .A(n_55), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_56), .B(n_175), .Y(n_548) );
A2O1A1Ixp33_ASAP7_75t_L g185 ( .A1(n_57), .A2(n_174), .B(n_186), .C(n_187), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_58), .Y(n_236) );
INVx1_ASAP7_75t_L g184 ( .A(n_59), .Y(n_184) );
INVx1_ASAP7_75t_L g144 ( .A(n_61), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g437 ( .A(n_62), .B(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_63), .B(n_175), .Y(n_529) );
INVx1_ASAP7_75t_L g134 ( .A(n_64), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_65), .Y(n_117) );
AO32x2_ASAP7_75t_L g471 ( .A1(n_66), .A2(n_164), .A3(n_239), .B1(n_472), .B2(n_476), .Y(n_471) );
INVx1_ASAP7_75t_L g547 ( .A(n_67), .Y(n_547) );
INVx1_ASAP7_75t_L g462 ( .A(n_68), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_SL g170 ( .A1(n_69), .A2(n_171), .B(n_172), .C(n_174), .Y(n_170) );
INVxp67_ASAP7_75t_L g173 ( .A(n_70), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_71), .B(n_156), .Y(n_463) );
INVx1_ASAP7_75t_L g106 ( .A(n_72), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g206 ( .A(n_73), .Y(n_206) );
INVx1_ASAP7_75t_L g229 ( .A(n_74), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_76), .A2(n_143), .B(n_146), .C(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_77), .B(n_474), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_78), .B(n_156), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_79), .B(n_151), .Y(n_219) );
INVx2_ASAP7_75t_L g132 ( .A(n_80), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_81), .B(n_171), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_82), .B(n_156), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_L g145 ( .A1(n_83), .A2(n_143), .B(n_146), .C(n_149), .Y(n_145) );
OR2x2_ASAP7_75t_L g108 ( .A(n_84), .B(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g444 ( .A(n_84), .B(n_110), .Y(n_444) );
INVx2_ASAP7_75t_L g449 ( .A(n_84), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_86), .A2(n_100), .B1(n_156), .B2(n_157), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_87), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_88), .B(n_161), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_89), .Y(n_159) );
A2O1A1Ixp33_ASAP7_75t_L g241 ( .A1(n_90), .A2(n_143), .B(n_146), .C(n_242), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_91), .Y(n_249) );
INVx1_ASAP7_75t_L g169 ( .A(n_92), .Y(n_169) );
CKINVDCx16_ASAP7_75t_R g255 ( .A(n_93), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_94), .B(n_151), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_95), .B(n_156), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_96), .B(n_164), .Y(n_261) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_97), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_98), .B(n_106), .Y(n_105) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_99), .A2(n_166), .B(n_167), .Y(n_165) );
CKINVDCx6p67_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
BUFx2_ASAP7_75t_L g736 ( .A(n_103), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_107), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_108), .Y(n_436) );
INVx2_ASAP7_75t_L g438 ( .A(n_108), .Y(n_438) );
NOR2x2_ASAP7_75t_L g734 ( .A(n_109), .B(n_449), .Y(n_734) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g448 ( .A(n_110), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
AO21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_118), .B(n_439), .Y(n_113) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx3_ASAP7_75t_L g735 ( .A(n_115), .Y(n_735) );
INVx2_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI21xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_435), .B(n_437), .Y(n_118) );
XNOR2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_123), .Y(n_119) );
INVx1_ASAP7_75t_L g445 ( .A(n_123), .Y(n_445) );
OAI22xp5_ASAP7_75t_SL g730 ( .A1(n_123), .A2(n_446), .B1(n_451), .B2(n_731), .Y(n_730) );
NAND2x1_ASAP7_75t_L g123 ( .A(n_124), .B(n_351), .Y(n_123) );
NOR5xp2_ASAP7_75t_L g124 ( .A(n_125), .B(n_274), .C(n_306), .D(n_321), .E(n_338), .Y(n_124) );
A2O1A1Ixp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_190), .B(n_211), .C(n_262), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_162), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_127), .B(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_127), .B(n_326), .Y(n_389) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_128), .B(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_128), .B(n_208), .Y(n_275) );
AND2x2_ASAP7_75t_L g316 ( .A(n_128), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_128), .B(n_285), .Y(n_320) );
OR2x2_ASAP7_75t_L g357 ( .A(n_128), .B(n_196), .Y(n_357) );
INVx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g195 ( .A(n_129), .B(n_196), .Y(n_195) );
INVx3_ASAP7_75t_L g265 ( .A(n_129), .Y(n_265) );
OR2x2_ASAP7_75t_L g428 ( .A(n_129), .B(n_268), .Y(n_428) );
AO21x2_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_136), .B(n_158), .Y(n_129) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_130), .A2(n_197), .B(n_205), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_130), .B(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g224 ( .A(n_130), .Y(n_224) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_131), .Y(n_164) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
AND2x2_ASAP7_75t_SL g161 ( .A(n_132), .B(n_133), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
OAI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_138), .B(n_145), .Y(n_136) );
OAI22xp33_ASAP7_75t_L g197 ( .A1(n_138), .A2(n_176), .B1(n_198), .B2(n_204), .Y(n_197) );
OAI21xp5_ASAP7_75t_L g228 ( .A1(n_138), .A2(n_229), .B(n_230), .Y(n_228) );
NAND2x1p5_ASAP7_75t_L g138 ( .A(n_139), .B(n_143), .Y(n_138) );
AND2x4_ASAP7_75t_L g166 ( .A(n_139), .B(n_143), .Y(n_166) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
INVx1_ASAP7_75t_L g527 ( .A(n_140), .Y(n_527) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g147 ( .A(n_141), .Y(n_147) );
INVx1_ASAP7_75t_L g157 ( .A(n_141), .Y(n_157) );
INVx1_ASAP7_75t_L g148 ( .A(n_142), .Y(n_148) );
INVx3_ASAP7_75t_L g152 ( .A(n_142), .Y(n_152) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_142), .Y(n_154) );
INVx1_ASAP7_75t_L g171 ( .A(n_142), .Y(n_171) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_142), .Y(n_200) );
INVx4_ASAP7_75t_SL g176 ( .A(n_143), .Y(n_176) );
OAI21xp5_ASAP7_75t_L g460 ( .A1(n_143), .A2(n_461), .B(n_464), .Y(n_460) );
BUFx3_ASAP7_75t_L g476 ( .A(n_143), .Y(n_476) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_143), .A2(n_481), .B(n_485), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_143), .A2(n_521), .B(n_525), .Y(n_520) );
OAI21xp5_ASAP7_75t_L g533 ( .A1(n_143), .A2(n_534), .B(n_537), .Y(n_533) );
INVx5_ASAP7_75t_L g168 ( .A(n_146), .Y(n_168) );
AND2x6_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_147), .Y(n_175) );
BUFx3_ASAP7_75t_L g223 ( .A(n_147), .Y(n_223) );
INVx1_ASAP7_75t_L g474 ( .A(n_147), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_153), .C(n_155), .Y(n_149) );
O2A1O1Ixp5_ASAP7_75t_SL g461 ( .A1(n_151), .A2(n_174), .B(n_462), .C(n_463), .Y(n_461) );
INVx2_ASAP7_75t_L g498 ( .A(n_151), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_151), .A2(n_535), .B(n_536), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_151), .A2(n_544), .B(n_545), .Y(n_543) );
INVx5_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_152), .B(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_152), .B(n_188), .Y(n_187) );
OAI22xp5_ASAP7_75t_SL g472 ( .A1(n_152), .A2(n_154), .B1(n_473), .B2(n_475), .Y(n_472) );
INVx2_ASAP7_75t_L g186 ( .A(n_154), .Y(n_186) );
INVx4_ASAP7_75t_L g245 ( .A(n_154), .Y(n_245) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_154), .A2(n_497), .B1(n_498), .B2(n_499), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_154), .A2(n_498), .B1(n_514), .B2(n_515), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g521 ( .A1(n_155), .A2(n_522), .B(n_523), .C(n_524), .Y(n_521) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_160), .B(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_160), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g239 ( .A(n_161), .Y(n_239) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_161), .A2(n_252), .B(n_261), .Y(n_251) );
OA21x2_ASAP7_75t_L g459 ( .A1(n_161), .A2(n_460), .B(n_467), .Y(n_459) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_161), .A2(n_480), .B(n_488), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g330 ( .A1(n_162), .A2(n_331), .B1(n_332), .B2(n_335), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_162), .B(n_265), .Y(n_414) );
AND2x2_ASAP7_75t_L g162 ( .A(n_163), .B(n_180), .Y(n_162) );
AND2x2_ASAP7_75t_L g210 ( .A(n_163), .B(n_196), .Y(n_210) );
AND2x2_ASAP7_75t_L g267 ( .A(n_163), .B(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g272 ( .A(n_163), .Y(n_272) );
INVx3_ASAP7_75t_L g285 ( .A(n_163), .Y(n_285) );
OR2x2_ASAP7_75t_L g305 ( .A(n_163), .B(n_268), .Y(n_305) );
AND2x2_ASAP7_75t_L g324 ( .A(n_163), .B(n_181), .Y(n_324) );
BUFx2_ASAP7_75t_L g356 ( .A(n_163), .Y(n_356) );
OA21x2_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_165), .B(n_177), .Y(n_163) );
INVx4_ASAP7_75t_L g179 ( .A(n_164), .Y(n_179) );
OA21x2_ASAP7_75t_L g532 ( .A1(n_164), .A2(n_533), .B(n_540), .Y(n_532) );
BUFx2_ASAP7_75t_L g253 ( .A(n_166), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_170), .C(n_176), .Y(n_167) );
O2A1O1Ixp33_ASAP7_75t_L g183 ( .A1(n_168), .A2(n_176), .B(n_184), .C(n_185), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_168), .A2(n_176), .B(n_255), .C(n_256), .Y(n_254) );
INVx1_ASAP7_75t_L g484 ( .A(n_171), .Y(n_484) );
INVx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_175), .Y(n_246) );
OA21x2_ASAP7_75t_L g181 ( .A1(n_178), .A2(n_182), .B(n_189), .Y(n_181) );
INVx3_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_SL g225 ( .A(n_179), .B(n_226), .Y(n_225) );
NAND3xp33_ASAP7_75t_L g512 ( .A(n_179), .B(n_476), .C(n_513), .Y(n_512) );
AO21x1_ASAP7_75t_L g602 ( .A1(n_179), .A2(n_513), .B(n_603), .Y(n_602) );
AND2x4_ASAP7_75t_L g271 ( .A(n_180), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_SL g180 ( .A(n_181), .Y(n_180) );
BUFx2_ASAP7_75t_L g194 ( .A(n_181), .Y(n_194) );
INVx2_ASAP7_75t_L g209 ( .A(n_181), .Y(n_209) );
OR2x2_ASAP7_75t_L g287 ( .A(n_181), .B(n_268), .Y(n_287) );
AND2x2_ASAP7_75t_L g317 ( .A(n_181), .B(n_196), .Y(n_317) );
AND2x2_ASAP7_75t_L g334 ( .A(n_181), .B(n_265), .Y(n_334) );
AND2x2_ASAP7_75t_L g374 ( .A(n_181), .B(n_285), .Y(n_374) );
AND2x2_ASAP7_75t_SL g410 ( .A(n_181), .B(n_210), .Y(n_410) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_186), .A2(n_486), .B(n_487), .Y(n_485) );
O2A1O1Ixp5_ASAP7_75t_L g546 ( .A1(n_186), .A2(n_526), .B(n_547), .C(n_548), .Y(n_546) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NAND2xp33_ASAP7_75t_SL g191 ( .A(n_192), .B(n_207), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_193), .B(n_195), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_193), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_SL g193 ( .A(n_194), .Y(n_193) );
OAI21xp33_ASAP7_75t_L g348 ( .A1(n_194), .A2(n_210), .B(n_349), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_194), .B(n_196), .Y(n_404) );
AND2x2_ASAP7_75t_L g340 ( .A(n_195), .B(n_341), .Y(n_340) );
INVx3_ASAP7_75t_L g268 ( .A(n_196), .Y(n_268) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_196), .Y(n_366) );
OAI22xp5_ASAP7_75t_SL g199 ( .A1(n_200), .A2(n_201), .B1(n_202), .B2(n_203), .Y(n_199) );
INVx2_ASAP7_75t_L g202 ( .A(n_200), .Y(n_202) );
INVx4_ASAP7_75t_L g257 ( .A(n_200), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_207), .B(n_265), .Y(n_433) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_208), .A2(n_376), .B1(n_377), .B2(n_382), .Y(n_375) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
AND2x2_ASAP7_75t_L g266 ( .A(n_209), .B(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g304 ( .A(n_209), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_SL g341 ( .A(n_209), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_210), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g395 ( .A(n_210), .Y(n_395) );
CKINVDCx16_ASAP7_75t_R g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_237), .Y(n_212) );
INVx4_ASAP7_75t_L g281 ( .A(n_213), .Y(n_281) );
AND2x2_ASAP7_75t_L g359 ( .A(n_213), .B(n_326), .Y(n_359) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_227), .Y(n_213) );
INVx3_ASAP7_75t_L g278 ( .A(n_214), .Y(n_278) );
AND2x2_ASAP7_75t_L g292 ( .A(n_214), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g296 ( .A(n_214), .Y(n_296) );
INVx2_ASAP7_75t_L g310 ( .A(n_214), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_214), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g367 ( .A(n_214), .B(n_362), .Y(n_367) );
AND2x2_ASAP7_75t_L g432 ( .A(n_214), .B(n_402), .Y(n_432) );
OR2x6_ASAP7_75t_L g214 ( .A(n_215), .B(n_225), .Y(n_214) );
AOI21xp5_ASAP7_75t_SL g215 ( .A1(n_216), .A2(n_217), .B(n_224), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_221), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_221), .A2(n_232), .B(n_233), .Y(n_231) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g260 ( .A(n_223), .Y(n_260) );
INVx1_ASAP7_75t_L g234 ( .A(n_224), .Y(n_234) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_224), .A2(n_520), .B(n_530), .Y(n_519) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_224), .A2(n_542), .B(n_549), .Y(n_541) );
AND2x2_ASAP7_75t_L g273 ( .A(n_227), .B(n_251), .Y(n_273) );
INVx2_ASAP7_75t_L g293 ( .A(n_227), .Y(n_293) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_234), .B(n_235), .Y(n_227) );
INVx1_ASAP7_75t_L g298 ( .A(n_237), .Y(n_298) );
AND2x2_ASAP7_75t_L g344 ( .A(n_237), .B(n_292), .Y(n_344) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_250), .Y(n_237) );
INVx2_ASAP7_75t_L g283 ( .A(n_238), .Y(n_283) );
INVx1_ASAP7_75t_L g291 ( .A(n_238), .Y(n_291) );
AND2x2_ASAP7_75t_L g309 ( .A(n_238), .B(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_238), .B(n_293), .Y(n_347) );
AO21x2_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_248), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_241), .B(n_247), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_246), .Y(n_242) );
AND2x2_ASAP7_75t_L g326 ( .A(n_250), .B(n_283), .Y(n_326) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g279 ( .A(n_251), .Y(n_279) );
AND2x2_ASAP7_75t_L g362 ( .A(n_251), .B(n_293), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_257), .B(n_259), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_257), .A2(n_465), .B(n_466), .Y(n_464) );
INVx1_ASAP7_75t_L g524 ( .A(n_257), .Y(n_524) );
OAI21xp5_ASAP7_75t_SL g262 ( .A1(n_263), .A2(n_269), .B(n_273), .Y(n_262) );
INVx1_ASAP7_75t_SL g307 ( .A(n_263), .Y(n_307) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_264), .B(n_271), .Y(n_364) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g313 ( .A(n_265), .B(n_268), .Y(n_313) );
AND2x2_ASAP7_75t_L g342 ( .A(n_265), .B(n_286), .Y(n_342) );
OR2x2_ASAP7_75t_L g345 ( .A(n_265), .B(n_305), .Y(n_345) );
AOI222xp33_ASAP7_75t_L g409 ( .A1(n_266), .A2(n_358), .B1(n_410), .B2(n_411), .C1(n_413), .C2(n_415), .Y(n_409) );
BUFx2_ASAP7_75t_L g323 ( .A(n_268), .Y(n_323) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g312 ( .A(n_271), .B(n_313), .Y(n_312) );
INVx3_ASAP7_75t_SL g329 ( .A(n_271), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_271), .B(n_323), .Y(n_383) );
AND2x2_ASAP7_75t_L g318 ( .A(n_273), .B(n_278), .Y(n_318) );
INVx1_ASAP7_75t_L g337 ( .A(n_273), .Y(n_337) );
OAI221xp5_ASAP7_75t_SL g274 ( .A1(n_275), .A2(n_276), .B1(n_280), .B2(n_284), .C(n_288), .Y(n_274) );
OR2x2_ASAP7_75t_L g346 ( .A(n_276), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AND2x2_ASAP7_75t_L g331 ( .A(n_278), .B(n_301), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_278), .B(n_291), .Y(n_371) );
AND2x2_ASAP7_75t_L g376 ( .A(n_278), .B(n_326), .Y(n_376) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_278), .Y(n_386) );
NAND2x1_ASAP7_75t_SL g397 ( .A(n_278), .B(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g282 ( .A(n_279), .B(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g302 ( .A(n_279), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_279), .B(n_297), .Y(n_328) );
INVx1_ASAP7_75t_L g394 ( .A(n_279), .Y(n_394) );
INVx1_ASAP7_75t_L g369 ( .A(n_280), .Y(n_369) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx1_ASAP7_75t_L g381 ( .A(n_281), .Y(n_381) );
NOR2xp67_ASAP7_75t_L g393 ( .A(n_281), .B(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g398 ( .A(n_282), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_282), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g301 ( .A(n_283), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_283), .B(n_293), .Y(n_314) );
INVx1_ASAP7_75t_L g380 ( .A(n_283), .Y(n_380) );
INVx1_ASAP7_75t_L g401 ( .A(n_284), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OAI21xp5_ASAP7_75t_SL g288 ( .A1(n_289), .A2(n_294), .B(n_303), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
AND2x2_ASAP7_75t_L g434 ( .A(n_290), .B(n_367), .Y(n_434) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g402 ( .A(n_291), .B(n_362), .Y(n_402) );
AOI32xp33_ASAP7_75t_L g315 ( .A1(n_292), .A2(n_298), .A3(n_316), .B1(n_318), .B2(n_319), .Y(n_315) );
AOI322xp5_ASAP7_75t_L g417 ( .A1(n_292), .A2(n_324), .A3(n_407), .B1(n_418), .B2(n_419), .C1(n_420), .C2(n_422), .Y(n_417) );
INVx2_ASAP7_75t_L g297 ( .A(n_293), .Y(n_297) );
INVx1_ASAP7_75t_L g407 ( .A(n_293), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_298), .B1(n_299), .B2(n_300), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_295), .B(n_301), .Y(n_350) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_296), .B(n_362), .Y(n_412) );
INVx1_ASAP7_75t_L g299 ( .A(n_297), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_297), .B(n_326), .Y(n_416) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_305), .B(n_400), .Y(n_399) );
OAI221xp5_ASAP7_75t_SL g306 ( .A1(n_307), .A2(n_308), .B1(n_311), .B2(n_314), .C(n_315), .Y(n_306) );
OR2x2_ASAP7_75t_L g327 ( .A(n_308), .B(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g336 ( .A(n_308), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g361 ( .A(n_309), .B(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g365 ( .A(n_319), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
OAI221xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_325), .B1(n_327), .B2(n_329), .C(n_330), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g353 ( .A1(n_323), .A2(n_354), .B1(n_358), .B2(n_359), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_324), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g429 ( .A(n_324), .Y(n_429) );
INVx1_ASAP7_75t_L g423 ( .A(n_326), .Y(n_423) );
INVx1_ASAP7_75t_SL g358 ( .A(n_327), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_329), .B(n_357), .Y(n_419) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_334), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_SL g400 ( .A(n_334), .Y(n_400) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
OAI221xp5_ASAP7_75t_SL g338 ( .A1(n_339), .A2(n_343), .B1(n_345), .B2(n_346), .C(n_348), .Y(n_338) );
NOR2xp33_ASAP7_75t_SL g339 ( .A(n_340), .B(n_342), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_340), .A2(n_358), .B1(n_404), .B2(n_405), .Y(n_403) );
CKINVDCx14_ASAP7_75t_R g343 ( .A(n_344), .Y(n_343) );
OAI21xp33_ASAP7_75t_L g422 ( .A1(n_345), .A2(n_423), .B(n_424), .Y(n_422) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NOR3xp33_ASAP7_75t_SL g351 ( .A(n_352), .B(n_384), .C(n_408), .Y(n_351) );
NAND4xp25_ASAP7_75t_L g352 ( .A(n_353), .B(n_360), .C(n_368), .D(n_375), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g431 ( .A(n_356), .Y(n_431) );
INVx3_ASAP7_75t_SL g425 ( .A(n_357), .Y(n_425) );
OR2x2_ASAP7_75t_L g430 ( .A(n_357), .B(n_431), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_363), .B1(n_365), .B2(n_367), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_362), .B(n_380), .Y(n_421) );
INVxp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OAI21xp5_ASAP7_75t_SL g368 ( .A1(n_369), .A2(n_370), .B(n_372), .Y(n_368) );
INVxp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_381), .Y(n_378) );
INVxp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI211xp5_ASAP7_75t_SL g384 ( .A1(n_385), .A2(n_387), .B(n_390), .C(n_403), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g418 ( .A(n_389), .Y(n_418) );
AOI222xp33_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_395), .B1(n_396), .B2(n_399), .C1(n_401), .C2(n_402), .Y(n_390) );
INVxp67_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND4xp25_ASAP7_75t_SL g427 ( .A(n_400), .B(n_428), .C(n_429), .D(n_430), .Y(n_427) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND3xp33_ASAP7_75t_SL g408 ( .A(n_409), .B(n_417), .C(n_426), .Y(n_408) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_432), .B1(n_433), .B2(n_434), .Y(n_426) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AOI21xp33_ASAP7_75t_L g439 ( .A1(n_437), .A2(n_440), .B(n_735), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_445), .B1(n_446), .B2(n_450), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g731 ( .A(n_443), .Y(n_731) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_647), .Y(n_451) );
NAND3xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_596), .C(n_638), .Y(n_452) );
AOI211xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_505), .B(n_550), .C(n_572), .Y(n_453) );
OAI211xp5_ASAP7_75t_SL g454 ( .A1(n_455), .A2(n_468), .B(n_489), .C(n_500), .Y(n_454) );
INVxp67_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_456), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g659 ( .A(n_456), .B(n_576), .Y(n_659) );
BUFx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g561 ( .A(n_457), .B(n_492), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_457), .B(n_479), .Y(n_678) );
INVx1_ASAP7_75t_L g696 ( .A(n_457), .Y(n_696) );
AND2x2_ASAP7_75t_L g705 ( .A(n_457), .B(n_593), .Y(n_705) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g588 ( .A(n_458), .B(n_479), .Y(n_588) );
AND2x2_ASAP7_75t_L g646 ( .A(n_458), .B(n_593), .Y(n_646) );
INVx1_ASAP7_75t_L g690 ( .A(n_458), .Y(n_690) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g567 ( .A(n_459), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g575 ( .A(n_459), .Y(n_575) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_459), .Y(n_615) );
INVxp67_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_477), .Y(n_469) );
AND2x2_ASAP7_75t_L g554 ( .A(n_470), .B(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g587 ( .A(n_470), .Y(n_587) );
OR2x2_ASAP7_75t_L g713 ( .A(n_470), .B(n_714), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_470), .B(n_479), .Y(n_717) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g492 ( .A(n_471), .Y(n_492) );
INVx1_ASAP7_75t_L g503 ( .A(n_471), .Y(n_503) );
AND2x2_ASAP7_75t_L g576 ( .A(n_471), .B(n_494), .Y(n_576) );
AND2x2_ASAP7_75t_L g616 ( .A(n_471), .B(n_495), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g542 ( .A1(n_476), .A2(n_543), .B(n_546), .Y(n_542) );
INVxp67_ASAP7_75t_L g658 ( .A(n_477), .Y(n_658) );
AND2x4_ASAP7_75t_L g683 ( .A(n_477), .B(n_576), .Y(n_683) );
BUFx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_SL g574 ( .A(n_478), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g493 ( .A(n_479), .B(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g562 ( .A(n_479), .B(n_495), .Y(n_562) );
INVx1_ASAP7_75t_L g568 ( .A(n_479), .Y(n_568) );
INVx2_ASAP7_75t_L g594 ( .A(n_479), .Y(n_594) );
AND2x2_ASAP7_75t_L g610 ( .A(n_479), .B(n_611), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .B(n_484), .Y(n_481) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_490), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_493), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx2_ASAP7_75t_L g565 ( .A(n_492), .Y(n_565) );
AND2x2_ASAP7_75t_L g673 ( .A(n_492), .B(n_494), .Y(n_673) );
AND2x2_ASAP7_75t_L g590 ( .A(n_493), .B(n_575), .Y(n_590) );
AND2x2_ASAP7_75t_L g689 ( .A(n_493), .B(n_690), .Y(n_689) );
NOR2xp67_ASAP7_75t_L g611 ( .A(n_494), .B(n_612), .Y(n_611) );
OR2x2_ASAP7_75t_L g714 ( .A(n_494), .B(n_575), .Y(n_714) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx2_ASAP7_75t_L g504 ( .A(n_495), .Y(n_504) );
AND2x2_ASAP7_75t_L g593 ( .A(n_495), .B(n_594), .Y(n_593) );
O2A1O1Ixp33_ASAP7_75t_L g525 ( .A1(n_498), .A2(n_526), .B(n_528), .C(n_529), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_498), .A2(n_538), .B(n_539), .Y(n_537) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_504), .Y(n_501) );
AND2x2_ASAP7_75t_L g639 ( .A(n_502), .B(n_574), .Y(n_639) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_503), .B(n_575), .Y(n_624) );
INVx2_ASAP7_75t_L g623 ( .A(n_504), .Y(n_623) );
OAI222xp33_ASAP7_75t_L g627 ( .A1(n_504), .A2(n_567), .B1(n_628), .B2(n_630), .C1(n_631), .C2(n_634), .Y(n_627) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_516), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g552 ( .A(n_509), .Y(n_552) );
OR2x2_ASAP7_75t_L g663 ( .A(n_509), .B(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx3_ASAP7_75t_L g585 ( .A(n_510), .Y(n_585) );
NOR2x1_ASAP7_75t_L g636 ( .A(n_510), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g642 ( .A(n_510), .B(n_556), .Y(n_642) );
AND2x4_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
INVx1_ASAP7_75t_L g603 ( .A(n_511), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_516), .A2(n_606), .B1(n_645), .B2(n_646), .Y(n_644) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_531), .Y(n_516) );
INVx3_ASAP7_75t_L g578 ( .A(n_517), .Y(n_578) );
OR2x2_ASAP7_75t_L g711 ( .A(n_517), .B(n_587), .Y(n_711) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g584 ( .A(n_518), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g600 ( .A(n_518), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g608 ( .A(n_518), .B(n_556), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_518), .B(n_532), .Y(n_664) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g555 ( .A(n_519), .B(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g559 ( .A(n_519), .B(n_532), .Y(n_559) );
AND2x2_ASAP7_75t_L g635 ( .A(n_519), .B(n_582), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_519), .B(n_541), .Y(n_675) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_531), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g591 ( .A(n_531), .B(n_552), .Y(n_591) );
AND2x2_ASAP7_75t_L g595 ( .A(n_531), .B(n_585), .Y(n_595) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_541), .Y(n_531) );
INVx3_ASAP7_75t_L g556 ( .A(n_532), .Y(n_556) );
AND2x2_ASAP7_75t_L g581 ( .A(n_532), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g716 ( .A(n_532), .B(n_699), .Y(n_716) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_541), .Y(n_570) );
INVx2_ASAP7_75t_L g582 ( .A(n_541), .Y(n_582) );
AND2x2_ASAP7_75t_L g626 ( .A(n_541), .B(n_602), .Y(n_626) );
INVx1_ASAP7_75t_L g669 ( .A(n_541), .Y(n_669) );
OR2x2_ASAP7_75t_L g700 ( .A(n_541), .B(n_602), .Y(n_700) );
AND2x2_ASAP7_75t_L g720 ( .A(n_541), .B(n_556), .Y(n_720) );
OAI21xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_553), .B(n_557), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g558 ( .A(n_552), .B(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_552), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g677 ( .A(n_554), .Y(n_677) );
INVx2_ASAP7_75t_SL g571 ( .A(n_555), .Y(n_571) );
AND2x2_ASAP7_75t_L g691 ( .A(n_555), .B(n_585), .Y(n_691) );
INVx2_ASAP7_75t_L g637 ( .A(n_556), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_556), .B(n_669), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_560), .B1(n_563), .B2(n_569), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_559), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_SL g725 ( .A(n_559), .Y(n_725) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
INVx1_ASAP7_75t_L g650 ( .A(n_561), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_561), .B(n_593), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_562), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g666 ( .A(n_562), .B(n_615), .Y(n_666) );
INVx2_ASAP7_75t_L g722 ( .A(n_562), .Y(n_722) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
AND2x2_ASAP7_75t_L g592 ( .A(n_565), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_565), .B(n_610), .Y(n_643) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_567), .B(n_587), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
INVx1_ASAP7_75t_L g704 ( .A(n_570), .Y(n_704) );
O2A1O1Ixp33_ASAP7_75t_SL g654 ( .A1(n_571), .A2(n_655), .B(n_657), .C(n_660), .Y(n_654) );
OR2x2_ASAP7_75t_L g681 ( .A(n_571), .B(n_585), .Y(n_681) );
OAI221xp5_ASAP7_75t_SL g572 ( .A1(n_573), .A2(n_577), .B1(n_579), .B2(n_586), .C(n_589), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_574), .B(n_576), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_574), .B(n_623), .Y(n_630) );
AND2x2_ASAP7_75t_L g672 ( .A(n_574), .B(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g708 ( .A(n_574), .Y(n_708) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_575), .Y(n_599) );
INVx1_ASAP7_75t_L g612 ( .A(n_575), .Y(n_612) );
NOR2xp67_ASAP7_75t_L g632 ( .A(n_578), .B(n_633), .Y(n_632) );
INVxp67_ASAP7_75t_L g686 ( .A(n_578), .Y(n_686) );
NAND2xp5_ASAP7_75t_SL g702 ( .A(n_578), .B(n_626), .Y(n_702) );
INVx2_ASAP7_75t_L g688 ( .A(n_579), .Y(n_688) );
OR2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_583), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g629 ( .A(n_581), .B(n_600), .Y(n_629) );
O2A1O1Ixp33_ASAP7_75t_L g638 ( .A1(n_581), .A2(n_597), .B(n_639), .C(n_640), .Y(n_638) );
AND2x2_ASAP7_75t_L g607 ( .A(n_582), .B(n_602), .Y(n_607) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_586), .B(n_685), .Y(n_684) );
OR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
OR2x2_ASAP7_75t_L g655 ( .A(n_587), .B(n_656), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B1(n_592), .B2(n_595), .Y(n_589) );
INVx1_ASAP7_75t_L g709 ( .A(n_591), .Y(n_709) );
INVx1_ASAP7_75t_L g656 ( .A(n_593), .Y(n_656) );
INVx1_ASAP7_75t_L g707 ( .A(n_595), .Y(n_707) );
AOI211xp5_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_600), .B(n_604), .C(n_627), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g619 ( .A(n_599), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g670 ( .A(n_600), .Y(n_670) );
AND2x2_ASAP7_75t_L g719 ( .A(n_600), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OAI21xp33_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_609), .B(n_617), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
INVx2_ASAP7_75t_L g633 ( .A(n_607), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_607), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g625 ( .A(n_608), .B(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g701 ( .A(n_608), .Y(n_701) );
OAI32xp33_ASAP7_75t_L g712 ( .A1(n_608), .A2(n_660), .A3(n_667), .B1(n_708), .B2(n_713), .Y(n_712) );
NOR2xp33_ASAP7_75t_SL g609 ( .A(n_610), .B(n_613), .Y(n_609) );
INVx1_ASAP7_75t_SL g680 ( .A(n_610), .Y(n_680) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_SL g620 ( .A(n_616), .Y(n_620) );
OAI21xp33_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_621), .B(n_625), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OAI22xp33_ASAP7_75t_L g692 ( .A1(n_619), .A2(n_667), .B1(n_693), .B2(n_695), .Y(n_692) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_623), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g660 ( .A(n_626), .Y(n_660) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2x1p5_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g653 ( .A(n_637), .Y(n_653) );
OAI21xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_643), .B(n_644), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_646), .A2(n_688), .B1(n_689), .B2(n_691), .C(n_692), .Y(n_687) );
NAND5xp2_ASAP7_75t_L g647 ( .A(n_648), .B(n_671), .C(n_687), .D(n_697), .E(n_715), .Y(n_647) );
AOI211xp5_ASAP7_75t_SL g648 ( .A1(n_649), .A2(n_651), .B(n_654), .C(n_661), .Y(n_648) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g718 ( .A(n_655), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
OAI22xp33_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_663), .B1(n_665), .B2(n_667), .Y(n_661) );
INVx1_ASAP7_75t_SL g694 ( .A(n_664), .Y(n_694) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OAI322xp33_ASAP7_75t_L g676 ( .A1(n_667), .A2(n_677), .A3(n_678), .B1(n_679), .B2(n_680), .C1(n_681), .C2(n_682), .Y(n_676) );
OR2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_670), .Y(n_667) );
INVx1_ASAP7_75t_L g679 ( .A(n_669), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_669), .B(n_694), .Y(n_693) );
AOI211xp5_ASAP7_75t_SL g671 ( .A1(n_672), .A2(n_674), .B(n_676), .C(n_684), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
OAI22xp33_ASAP7_75t_L g706 ( .A1(n_680), .A2(n_707), .B1(n_708), .B2(n_709), .Y(n_706) );
INVx1_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g723 ( .A(n_690), .Y(n_723) );
AOI221xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_705), .B1(n_706), .B2(n_710), .C(n_712), .Y(n_697) );
OAI211xp5_ASAP7_75t_SL g698 ( .A1(n_699), .A2(n_701), .B(n_702), .C(n_703), .Y(n_698) );
INVx1_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
OR2x2_ASAP7_75t_L g724 ( .A(n_700), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AOI221xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_717), .B1(n_718), .B2(n_719), .C(n_721), .Y(n_715) );
AOI21xp33_ASAP7_75t_SL g721 ( .A1(n_722), .A2(n_723), .B(n_724), .Y(n_721) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
INVx3_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
endmodule