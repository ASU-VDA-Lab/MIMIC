module fake_jpeg_12618_n_129 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_129);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx6_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_23),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_4),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_7),
.B(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_45),
.A2(n_49),
.B1(n_52),
.B2(n_48),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_58),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_52),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_62),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_53),
.B(n_1),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

AOI21xp33_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_4),
.B(n_7),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_8),
.Y(n_68)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_73),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2x1_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_46),
.B(n_43),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_50),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_83),
.B(n_89),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_51),
.B1(n_42),
.B2(n_40),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_87),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_67),
.A2(n_9),
.B(n_55),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_91),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_70),
.A2(n_40),
.B1(n_51),
.B2(n_55),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_9),
.B(n_39),
.C(n_11),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_10),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_38),
.B1(n_14),
.B2(n_16),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_90),
.B(n_92),
.Y(n_95)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_12),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_18),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_102),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_19),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_84),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_20),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_80),
.B(n_21),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_105),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_22),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_28),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_93),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_110),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_112),
.B(n_117),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_115),
.B1(n_96),
.B2(n_106),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_98),
.A2(n_33),
.B(n_34),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_114),
.A2(n_95),
.B(n_107),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_96),
.B1(n_94),
.B2(n_100),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_108),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_109),
.C(n_101),
.Y(n_123)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_123),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_116),
.C(n_110),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_124),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_126),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_127),
.Y(n_128)
);

AOI221xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_122),
.B1(n_118),
.B2(n_111),
.C(n_120),
.Y(n_129)
);


endmodule