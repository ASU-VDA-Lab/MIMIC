module real_jpeg_6007_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_1),
.A2(n_134),
.B1(n_154),
.B2(n_157),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_1),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_1),
.A2(n_157),
.B1(n_211),
.B2(n_213),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_1),
.A2(n_157),
.B1(n_280),
.B2(n_282),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_1),
.A2(n_157),
.B1(n_332),
.B2(n_335),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_3),
.A2(n_65),
.B1(n_70),
.B2(n_71),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_3),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_3),
.A2(n_51),
.B1(n_60),
.B2(n_70),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_4),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_4),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_5),
.A2(n_49),
.B1(n_51),
.B2(n_53),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_5),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_5),
.A2(n_53),
.B1(n_122),
.B2(n_125),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g345 ( 
.A1(n_5),
.A2(n_53),
.B1(n_84),
.B2(n_346),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_6),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_6),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_6),
.A2(n_133),
.B1(n_268),
.B2(n_291),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_6),
.A2(n_133),
.B1(n_203),
.B2(n_308),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_6),
.A2(n_133),
.B1(n_353),
.B2(n_371),
.Y(n_370)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_7),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_8),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_8),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_8),
.Y(n_206)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_8),
.Y(n_229)
);

INVx8_ASAP7_75t_L g320 ( 
.A(n_8),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_9),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_9),
.A2(n_195),
.B1(n_254),
.B2(n_257),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_9),
.B(n_270),
.C(n_274),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_9),
.B(n_108),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_9),
.B(n_89),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_9),
.B(n_55),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_9),
.B(n_341),
.Y(n_340)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_10),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_10),
.Y(n_146)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_10),
.Y(n_149)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_11),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_12),
.Y(n_132)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_12),
.Y(n_137)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_12),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_12),
.Y(n_144)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_12),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_12),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_12),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_13),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_13),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_13),
.A2(n_85),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_14),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_14),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_14),
.A2(n_59),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_14),
.A2(n_59),
.B1(n_236),
.B2(n_240),
.Y(n_235)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_15),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_16),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_16),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_16),
.A2(n_118),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_16),
.A2(n_118),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_16),
.A2(n_67),
.B1(n_118),
.B2(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_244),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_243),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_217),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_21),
.B(n_217),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_160),
.C(n_173),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_22),
.A2(n_23),
.B1(n_160),
.B2(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_90),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_24),
.B(n_91),
.C(n_159),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_63),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_25),
.B(n_63),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_48),
.B1(n_54),
.B2(n_56),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_26),
.A2(n_253),
.B(n_260),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_26),
.A2(n_54),
.B1(n_290),
.B2(n_331),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_26),
.A2(n_260),
.B(n_331),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_27),
.A2(n_55),
.B1(n_57),
.B2(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_27),
.A2(n_55),
.B1(n_162),
.B2(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_27),
.B(n_261),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_38),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_28)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_32),
.Y(n_335)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_33),
.Y(n_112)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_33),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_33),
.Y(n_268)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_34),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_37),
.Y(n_226)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_38),
.A2(n_290),
.B(n_294),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_44),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_44),
.Y(n_286)
);

BUFx5_ASAP7_75t_L g347 ( 
.A(n_44),
.Y(n_347)
);

INVx8_ASAP7_75t_L g302 ( 
.A(n_45),
.Y(n_302)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_48),
.A2(n_54),
.B(n_294),
.Y(n_396)
);

INVx5_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_52),
.Y(n_223)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_52),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_52),
.Y(n_293)
);

INVx6_ASAP7_75t_L g334 ( 
.A(n_52),
.Y(n_334)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_55),
.B(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AO22x2_ASAP7_75t_L g108 ( 
.A1(n_61),
.A2(n_109),
.B1(n_112),
.B2(n_113),
.Y(n_108)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_74),
.B1(n_82),
.B2(n_88),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_64),
.Y(n_207)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_68),
.Y(n_169)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_68),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_69),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_74),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_74),
.B(n_285),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_74),
.A2(n_315),
.B1(n_316),
.B2(n_317),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_74),
.A2(n_199),
.B1(n_345),
.B2(n_377),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_81),
.Y(n_200)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_81),
.Y(n_309)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_83),
.A2(n_164),
.B1(n_165),
.B2(n_167),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_89),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_129),
.B1(n_158),
.B2(n_159),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_91),
.Y(n_158)
);

AOI22x1_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_108),
.B1(n_114),
.B2(n_120),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_92),
.A2(n_209),
.B(n_215),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_92),
.A2(n_215),
.B(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_92),
.B(n_114),
.Y(n_373)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_93),
.A2(n_121),
.B1(n_216),
.B2(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_93),
.A2(n_210),
.B1(n_216),
.B2(n_370),
.Y(n_395)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_108),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_99),
.B1(n_104),
.B2(n_105),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_99),
.Y(n_341)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_102),
.Y(n_186)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_103),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_103),
.Y(n_214)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_103),
.Y(n_239)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_108),
.Y(n_216)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx8_ASAP7_75t_L g356 ( 
.A(n_110),
.Y(n_356)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_112),
.Y(n_264)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_115),
.B(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_116),
.B(n_193),
.Y(n_192)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_128),
.Y(n_353)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_138),
.B1(n_147),
.B2(n_153),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_130),
.A2(n_176),
.B(n_178),
.Y(n_175)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_138),
.A2(n_153),
.B(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_179),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_139),
.A2(n_392),
.B(n_393),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_147),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_140)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_142),
.Y(n_191)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_147),
.B(n_195),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_147)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_149),
.Y(n_152)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_160),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_161),
.B(n_163),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_164),
.A2(n_198),
.B1(n_204),
.B2(n_207),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_164),
.A2(n_167),
.B(n_228),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_164),
.A2(n_279),
.B(n_284),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_164),
.A2(n_195),
.B(n_284),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_173),
.B(n_411),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_182),
.C(n_208),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_174),
.A2(n_175),
.B1(n_208),
.B2(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_177),
.B(n_179),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_182),
.B(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_196),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_183),
.A2(n_196),
.B1(n_197),
.B2(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_183),
.Y(n_385)
);

OAI32xp33_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_187),
.A3(n_191),
.B1(n_192),
.B2(n_194),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_SL g392 ( 
.A1(n_188),
.A2(n_194),
.B(n_195),
.Y(n_392)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_SL g338 ( 
.A1(n_195),
.A2(n_213),
.B(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_200),
.Y(n_283)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_205),
.B(n_285),
.Y(n_284)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_208),
.Y(n_406)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx6_ASAP7_75t_SL g213 ( 
.A(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_216),
.A2(n_370),
.B(n_373),
.Y(n_369)
);

BUFx24_ASAP7_75t_SL g422 ( 
.A(n_217),
.Y(n_422)
);

FAx1_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_219),
.CI(n_231),
.CON(n_217),
.SN(n_217)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_227),
.B2(n_230),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_223),
.Y(n_354)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx4_ASAP7_75t_SL g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_227),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_228),
.A2(n_307),
.B(n_310),
.Y(n_306)
);

INVx5_ASAP7_75t_L g377 ( 
.A(n_228),
.Y(n_377)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_241),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_239),
.Y(n_240)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_239),
.Y(n_372)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_242),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_399),
.B(n_418),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

AOI21x1_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_380),
.B(n_398),
.Y(n_246)
);

AO21x1_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_361),
.B(n_379),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_325),
.B(n_360),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_297),
.B(n_324),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_277),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_251),
.B(n_277),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_265),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_252),
.A2(n_265),
.B1(n_266),
.B2(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_252),
.Y(n_322)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_269),
.Y(n_266)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_287),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_278),
.B(n_288),
.C(n_296),
.Y(n_326)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_279),
.Y(n_316)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_295),
.B2(n_296),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_313),
.B(n_323),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_305),
.B(n_312),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_304),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_311),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_311),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_307),
.Y(n_315)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_310),
.A2(n_344),
.B(n_348),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_321),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_321),
.Y(n_323)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx8_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_320),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_327),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_342),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_330),
.B1(n_336),
.B2(n_337),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_330),
.B(n_336),
.C(n_342),
.Y(n_362)
);

INVx3_ASAP7_75t_SL g332 ( 
.A(n_333),
.Y(n_332)
);

INVx8_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_334),
.Y(n_359)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVxp33_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

AOI32xp33_ASAP7_75t_L g351 ( 
.A1(n_340),
.A2(n_352),
.A3(n_354),
.B1(n_355),
.B2(n_357),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_351),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_343),
.B(n_351),
.Y(n_367)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx5_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx5_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

NAND2xp33_ASAP7_75t_SL g357 ( 
.A(n_356),
.B(n_358),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_362),
.B(n_363),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_364),
.A2(n_365),
.B1(n_368),
.B2(n_378),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_366),
.B(n_367),
.C(n_378),
.Y(n_381)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_368),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_369),
.B(n_374),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_369),
.B(n_375),
.C(n_376),
.Y(n_386)
);

INVx8_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_381),
.B(n_382),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_389),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_384),
.A2(n_386),
.B1(n_387),
.B2(n_388),
.Y(n_383)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_384),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_386),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_386),
.B(n_387),
.C(n_389),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_390),
.A2(n_391),
.B1(n_394),
.B2(n_397),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_390),
.B(n_395),
.C(n_396),
.Y(n_409)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_394),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_395),
.B(n_396),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_401),
.B(n_413),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_402),
.A2(n_419),
.B(n_420),
.Y(n_418)
);

NOR2x1_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_410),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_403),
.B(n_410),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_407),
.C(n_409),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_404),
.B(n_416),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_407),
.A2(n_408),
.B1(n_409),
.B2(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_409),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_415),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_414),
.B(n_415),
.Y(n_419)
);


endmodule