module fake_jpeg_15437_n_125 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_125);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx2_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_28),
.B(n_39),
.Y(n_53)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_33),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_40),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_1),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_42),
.Y(n_66)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_1),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_26),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_19),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_45),
.B(n_8),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_29),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_51),
.B1(n_61),
.B2(n_65),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_49),
.B(n_55),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_22),
.B1(n_26),
.B2(n_12),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_2),
.B(n_4),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_18),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_58),
.B(n_62),
.Y(n_80)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_64),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_30),
.A2(n_25),
.B1(n_14),
.B2(n_18),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_32),
.B(n_12),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_25),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_28),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_73),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_79),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_9),
.Y(n_92)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_8),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_53),
.Y(n_90)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_63),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_77),
.B1(n_82),
.B2(n_67),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_70),
.B1(n_56),
.B2(n_78),
.Y(n_101)
);

OAI221xp5_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_57),
.B1(n_49),
.B2(n_50),
.C(n_44),
.Y(n_87)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_92),
.Y(n_98)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_67),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_81),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_94),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_106),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_101),
.A2(n_97),
.B1(n_103),
.B2(n_100),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_68),
.C(n_70),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_104),
.C(n_89),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_SL g107 ( 
.A1(n_103),
.A2(n_97),
.B(n_89),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_80),
.C(n_73),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_107),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_88),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_108),
.A2(n_92),
.B(n_98),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_105),
.A2(n_91),
.B1(n_85),
.B2(n_83),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_93),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_109),
.C(n_98),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_107),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_118),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

OAI31xp33_ASAP7_75t_L g122 ( 
.A1(n_119),
.A2(n_121),
.A3(n_114),
.B(n_115),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_118),
.B(n_92),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_122),
.A2(n_123),
.B(n_47),
.Y(n_124)
);

OAI311xp33_ASAP7_75t_L g123 ( 
.A1(n_120),
.A2(n_117),
.A3(n_74),
.B1(n_84),
.C1(n_73),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_59),
.Y(n_125)
);


endmodule