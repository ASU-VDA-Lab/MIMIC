module real_jpeg_27903_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_164;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_0),
.B(n_50),
.Y(n_49)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_0),
.Y(n_152)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_24)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_2),
.A2(n_28),
.B1(n_87),
.B2(n_109),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_2),
.A2(n_28),
.B1(n_37),
.B2(n_38),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_2),
.A2(n_28),
.B1(n_50),
.B2(n_53),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_4),
.B(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_4),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_SL g86 ( 
.A1(n_4),
.A2(n_26),
.B(n_46),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_4),
.A2(n_74),
.B1(n_87),
.B2(n_109),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_4),
.A2(n_37),
.B(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_4),
.B(n_37),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_4),
.B(n_42),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_4),
.A2(n_78),
.B1(n_148),
.B2(n_152),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_4),
.A2(n_25),
.B(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_5),
.A2(n_50),
.B1(n_53),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_5),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_6),
.A2(n_37),
.B1(n_38),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_6),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_6),
.A2(n_50),
.B1(n_53),
.B2(n_69),
.Y(n_79)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_7),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_8),
.A2(n_50),
.B1(n_53),
.B2(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_8),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_9),
.A2(n_37),
.B1(n_38),
.B2(n_41),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_9),
.A2(n_41),
.B1(n_50),
.B2(n_53),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_10),
.A2(n_50),
.B1(n_53),
.B2(n_62),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_11),
.A2(n_37),
.B1(n_38),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_11),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_67),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_11),
.A2(n_50),
.B1(n_53),
.B2(n_67),
.Y(n_137)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_14),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_15),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_15),
.A2(n_37),
.B1(n_38),
.B2(n_54),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_115),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_113),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_82),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_19),
.B(n_82),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_59),
.C(n_70),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_20),
.A2(n_21),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_43),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_22),
.B(n_44),
.C(n_48),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_29),
.B1(n_40),
.B2(n_42),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_24),
.A2(n_30),
.B1(n_34),
.B2(n_163),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_31),
.B(n_33),
.C(n_34),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_31),
.Y(n_33)
);

AO22x1_ASAP7_75t_L g45 ( 
.A1(n_25),
.A2(n_26),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

OAI32xp33_ASAP7_75t_L g72 ( 
.A1(n_25),
.A2(n_35),
.A3(n_38),
.B1(n_73),
.B2(n_75),
.Y(n_72)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_26),
.B(n_74),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_30),
.A2(n_34),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_34)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_37),
.A2(n_38),
.B1(n_62),
.B2(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_37),
.B(n_76),
.Y(n_75)
);

OAI32xp33_ASAP7_75t_L g126 ( 
.A1(n_37),
.A2(n_53),
.A3(n_64),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_40),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_48),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_45),
.A2(n_108),
.B1(n_111),
.B2(n_112),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_45),
.A2(n_46),
.B(n_109),
.C(n_110),
.Y(n_108)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

NAND2xp33_ASAP7_75t_SL g110 ( 
.A(n_46),
.B(n_109),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_74),
.B(n_86),
.C(n_87),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_52),
.B1(n_55),
.B2(n_57),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_49),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_49),
.A2(n_55),
.B1(n_57),
.B2(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_49),
.A2(n_55),
.B1(n_141),
.B2(n_143),
.Y(n_140)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_50),
.B(n_62),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_50),
.B(n_154),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_52),
.Y(n_81)
);

INVx5_ASAP7_75t_SL g80 ( 
.A(n_55),
.Y(n_80)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_56),
.A2(n_78),
.B1(n_142),
.B2(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_56),
.B(n_74),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_59),
.A2(n_70),
.B1(n_71),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_59),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_65),
.B2(n_68),
.Y(n_59)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_60),
.A2(n_61),
.B1(n_122),
.B2(n_124),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_60),
.A2(n_61),
.B1(n_124),
.B2(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_63),
.Y(n_60)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_61),
.B(n_74),
.Y(n_149)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_66),
.A2(n_104),
.B1(n_106),
.B2(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_68),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_77),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_72),
.B(n_77),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_73),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_137),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_95),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_84),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_89),
.Y(n_84)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_107),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_101),
.B2(n_102),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_173),
.B(n_179),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_158),
.B(n_172),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_138),
.B(n_157),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_129),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_119),
.B(n_129),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_125),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_120),
.A2(n_121),
.B1(n_125),
.B2(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_123),
.Y(n_127)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_136),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_134),
.C(n_136),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_135),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_137),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_145),
.B(n_156),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_140),
.B(n_144),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_150),
.B(n_155),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_147),
.B(n_149),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_153),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_159),
.B(n_160),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_160)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_161)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_165),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_168),
.C(n_171),
.Y(n_174)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_169),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_174),
.B(n_175),
.Y(n_179)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);


endmodule