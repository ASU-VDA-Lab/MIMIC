module fake_jpeg_1926_n_570 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_570);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_570;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_3),
.B(n_18),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_53),
.B(n_56),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_20),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_29),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_58),
.B(n_72),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_39),
.B(n_16),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_103),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_60),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_63),
.Y(n_165)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_21),
.B(n_16),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_70),
.B(n_89),
.Y(n_131)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_71),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_29),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_74),
.B(n_80),
.Y(n_162)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_75),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_26),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_84),
.Y(n_168)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_34),
.B(n_0),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_90),
.Y(n_147)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

INVx3_ASAP7_75t_SL g92 ( 
.A(n_31),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_92),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_28),
.B(n_0),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_93),
.B(n_50),
.Y(n_142)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

INVx4_ASAP7_75t_SL g95 ( 
.A(n_39),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_95),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_97),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_19),
.Y(n_98)
);

NAND2xp33_ASAP7_75t_SL g122 ( 
.A(n_98),
.B(n_101),
.Y(n_122)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_26),
.Y(n_100)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

INVx5_ASAP7_75t_SL g101 ( 
.A(n_36),
.Y(n_101)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_24),
.Y(n_102)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_27),
.Y(n_121)
);

BUFx4f_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

BUFx8_ASAP7_75t_L g106 ( 
.A(n_24),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_L g161 ( 
.A1(n_106),
.A2(n_42),
.B(n_33),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_27),
.B1(n_37),
.B2(n_38),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_108),
.A2(n_115),
.B1(n_128),
.B2(n_129),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_L g115 ( 
.A1(n_84),
.A2(n_37),
.B1(n_36),
.B2(n_46),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_121),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_54),
.A2(n_46),
.B1(n_38),
.B2(n_36),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_59),
.A2(n_27),
.B1(n_38),
.B2(n_46),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_60),
.A2(n_27),
.B1(n_46),
.B2(n_38),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_132),
.A2(n_139),
.B1(n_144),
.B2(n_154),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_57),
.B(n_48),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_133),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_61),
.A2(n_34),
.B1(n_49),
.B2(n_47),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_78),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_140),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_142),
.B(n_170),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_63),
.A2(n_73),
.B1(n_100),
.B2(n_87),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_106),
.A2(n_34),
.B(n_42),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_149),
.A2(n_161),
.B(n_41),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_79),
.A2(n_50),
.B1(n_49),
.B2(n_47),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_98),
.B(n_45),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_69),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_83),
.A2(n_45),
.B1(n_44),
.B2(n_21),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_159),
.A2(n_32),
.B1(n_23),
.B2(n_96),
.Y(n_214)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_64),
.Y(n_167)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_92),
.Y(n_169)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_95),
.B(n_44),
.Y(n_170)
);

OR2x2_ASAP7_75t_SL g171 ( 
.A(n_107),
.B(n_106),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_171),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_111),
.Y(n_173)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_173),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g174 ( 
.A(n_114),
.Y(n_174)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_174),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_176),
.Y(n_260)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_110),
.Y(n_177)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_112),
.Y(n_178)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_178),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_180),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_131),
.B(n_42),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_181),
.B(n_195),
.Y(n_243)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_182),
.Y(n_282)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_125),
.Y(n_183)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_185),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_138),
.B(n_71),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_186),
.B(n_196),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_133),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_187),
.B(n_207),
.Y(n_249)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_113),
.Y(n_189)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_189),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_162),
.Y(n_190)
);

NAND3xp33_ASAP7_75t_L g286 ( 
.A(n_190),
.B(n_198),
.C(n_201),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_153),
.A2(n_33),
.B1(n_19),
.B2(n_76),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_191),
.A2(n_193),
.B1(n_194),
.B2(n_221),
.Y(n_238)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_116),
.Y(n_192)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_192),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_153),
.A2(n_19),
.B1(n_33),
.B2(n_77),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_107),
.A2(n_102),
.B1(n_69),
.B2(n_41),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_126),
.B(n_90),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_75),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_122),
.Y(n_197)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_197),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_146),
.B(n_62),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_199),
.B(n_200),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_156),
.B(n_55),
.Y(n_200)
);

AOI21xp33_ASAP7_75t_L g201 ( 
.A1(n_163),
.A2(n_101),
.B(n_103),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_151),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g233 ( 
.A(n_202),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_203),
.Y(n_277)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_119),
.Y(n_204)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_204),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_130),
.B(n_86),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_136),
.Y(n_208)
);

INVx13_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_141),
.Y(n_209)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_209),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_136),
.B(n_104),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_210),
.B(n_213),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_149),
.B(n_105),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_211),
.B(n_217),
.Y(n_245)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_117),
.Y(n_212)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_212),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g213 ( 
.A(n_127),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_214),
.A2(n_150),
.B1(n_165),
.B2(n_135),
.Y(n_258)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_127),
.Y(n_216)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_216),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_118),
.B(n_32),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_166),
.Y(n_218)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_218),
.Y(n_270)
);

BUFx2_ASAP7_75t_SL g219 ( 
.A(n_137),
.Y(n_219)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_219),
.Y(n_278)
);

BUFx12f_ASAP7_75t_L g220 ( 
.A(n_137),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_227),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_159),
.A2(n_23),
.B1(n_103),
.B2(n_104),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_155),
.Y(n_222)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_222),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_124),
.B(n_0),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_224),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_164),
.B(n_0),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_141),
.A2(n_43),
.B1(n_3),
.B2(n_4),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_225),
.A2(n_145),
.B1(n_119),
.B2(n_134),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_137),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_226),
.B(n_228),
.Y(n_250)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_135),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_147),
.B(n_121),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_147),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_230),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_166),
.B(n_2),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_157),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_109),
.Y(n_267)
);

AND2x4_ASAP7_75t_L g232 ( 
.A(n_148),
.B(n_43),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_157),
.C(n_128),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_235),
.B(n_10),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_179),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_236),
.B(n_241),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_179),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_184),
.A2(n_115),
.B1(n_132),
.B2(n_168),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_248),
.A2(n_264),
.B1(n_192),
.B2(n_218),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_258),
.A2(n_268),
.B1(n_271),
.B2(n_274),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_181),
.B(n_143),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_259),
.B(n_279),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_217),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_280),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_197),
.A2(n_150),
.B1(n_151),
.B2(n_160),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_223),
.B(n_148),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_266),
.B(n_276),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_267),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_184),
.A2(n_165),
.B1(n_134),
.B2(n_168),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_205),
.A2(n_203),
.B1(n_211),
.B2(n_214),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_273),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_205),
.A2(n_160),
.B1(n_120),
.B2(n_119),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_206),
.B(n_109),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_275),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_224),
.B(n_145),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_171),
.B(n_120),
.C(n_43),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_195),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_215),
.B(n_2),
.C(n_3),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_283),
.B(n_5),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_182),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_208),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_280),
.A2(n_221),
.B1(n_187),
.B2(n_172),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_289),
.B(n_316),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_246),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_290),
.B(n_295),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_238),
.A2(n_172),
.B(n_232),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_292),
.A2(n_297),
.B(n_311),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_260),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_293),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_246),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_247),
.A2(n_232),
.B(n_209),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_284),
.Y(n_298)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_298),
.Y(n_347)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_299),
.Y(n_353)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_300),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_271),
.A2(n_232),
.B1(n_227),
.B2(n_216),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_301),
.A2(n_302),
.B1(n_303),
.B2(n_306),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_263),
.A2(n_189),
.B1(n_212),
.B2(n_188),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_245),
.A2(n_188),
.B1(n_176),
.B2(n_202),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_237),
.Y(n_304)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_304),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_305),
.A2(n_321),
.B1(n_338),
.B2(n_283),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_245),
.A2(n_183),
.B1(n_175),
.B2(n_213),
.Y(n_306)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_281),
.Y(n_308)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_308),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_252),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_309),
.B(n_313),
.Y(n_345)
);

INVx4_ASAP7_75t_SL g310 ( 
.A(n_236),
.Y(n_310)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_310),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_277),
.A2(n_213),
.B(n_174),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_287),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_274),
.A2(n_204),
.B1(n_174),
.B2(n_173),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_314),
.A2(n_317),
.B1(n_318),
.B2(n_320),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_256),
.B(n_173),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_248),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_243),
.A2(n_235),
.B1(n_269),
.B2(n_276),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_287),
.B(n_220),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_319),
.B(n_324),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_243),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_266),
.A2(n_220),
.B1(n_6),
.B2(n_8),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_253),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_322),
.B(n_329),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_323),
.B(n_325),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_256),
.B(n_8),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_259),
.B(n_9),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_237),
.Y(n_326)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_326),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_247),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_327)
);

AO21x1_ASAP7_75t_L g360 ( 
.A1(n_327),
.A2(n_278),
.B(n_285),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_241),
.A2(n_9),
.B(n_10),
.Y(n_328)
);

NAND2x1_ASAP7_75t_L g344 ( 
.A(n_328),
.B(n_279),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_251),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_331),
.B(n_278),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_253),
.B(n_12),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_332),
.B(n_335),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_255),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_333),
.B(n_257),
.Y(n_367)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_239),
.Y(n_334)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_334),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_239),
.B(n_12),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_249),
.B(n_12),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_336),
.B(n_337),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_286),
.B(n_13),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_250),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_339),
.Y(n_387)
);

CKINVDCx14_ASAP7_75t_R g342 ( 
.A(n_291),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_342),
.B(n_343),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_291),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_344),
.A2(n_378),
.B(n_311),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_330),
.B(n_240),
.C(n_270),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_348),
.B(n_351),
.C(n_357),
.Y(n_385)
);

XOR2x2_ASAP7_75t_L g350 ( 
.A(n_330),
.B(n_240),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_350),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_318),
.B(n_270),
.C(n_262),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_300),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_354),
.B(n_358),
.Y(n_397)
);

CKINVDCx14_ASAP7_75t_R g356 ( 
.A(n_319),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_356),
.B(n_375),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_315),
.B(n_262),
.C(n_261),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_294),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_360),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_294),
.B(n_261),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_363),
.B(n_364),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_315),
.B(n_257),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_367),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_335),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_369),
.B(n_332),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_373),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_329),
.B(n_254),
.C(n_265),
.Y(n_375)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_310),
.B(n_242),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_377),
.B(n_383),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_297),
.B(n_292),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_304),
.Y(n_379)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_379),
.Y(n_390)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_326),
.Y(n_380)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_380),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_313),
.B(n_254),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_381),
.B(n_382),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_312),
.B(n_265),
.Y(n_382)
);

OR2x2_ASAP7_75t_SL g383 ( 
.A(n_310),
.B(n_244),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g384 ( 
.A1(n_358),
.A2(n_305),
.B1(n_309),
.B2(n_288),
.Y(n_384)
);

OAI22xp33_ASAP7_75t_SL g446 ( 
.A1(n_384),
.A2(n_402),
.B1(n_417),
.B2(n_418),
.Y(n_446)
);

CKINVDCx14_ASAP7_75t_R g443 ( 
.A(n_386),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_377),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_388),
.B(n_392),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_346),
.A2(n_296),
.B1(n_301),
.B2(n_289),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_389),
.A2(n_391),
.B1(n_393),
.B2(n_399),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_346),
.A2(n_296),
.B1(n_316),
.B2(n_307),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_343),
.B(n_324),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_370),
.A2(n_306),
.B1(n_317),
.B2(n_331),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_340),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_396),
.B(n_400),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_370),
.A2(n_331),
.B1(n_303),
.B2(n_295),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_345),
.Y(n_400)
);

XOR2x1_ASAP7_75t_L g448 ( 
.A(n_401),
.B(n_353),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_361),
.A2(n_290),
.B1(n_314),
.B2(n_321),
.Y(n_402)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_347),
.Y(n_404)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_404),
.Y(n_422)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_347),
.Y(n_405)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_405),
.Y(n_424)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_353),
.Y(n_411)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_411),
.Y(n_425)
);

OA22x2_ASAP7_75t_L g412 ( 
.A1(n_362),
.A2(n_302),
.B1(n_299),
.B2(n_298),
.Y(n_412)
);

OA21x2_ASAP7_75t_L g442 ( 
.A1(n_412),
.A2(n_368),
.B(n_380),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_369),
.B(n_325),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_413),
.B(n_415),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_378),
.A2(n_333),
.B1(n_336),
.B2(n_337),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_414),
.A2(n_372),
.B1(n_373),
.B2(n_375),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_354),
.B(n_334),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_378),
.A2(n_338),
.B1(n_328),
.B2(n_293),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_351),
.A2(n_293),
.B1(n_320),
.B2(n_308),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_362),
.A2(n_242),
.B1(n_282),
.B2(n_327),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_419),
.A2(n_349),
.B(n_360),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_352),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_420),
.B(n_368),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_341),
.B(n_323),
.Y(n_421)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_421),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_385),
.B(n_350),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_423),
.B(n_436),
.Y(n_469)
);

XNOR2x2_ASAP7_75t_SL g427 ( 
.A(n_401),
.B(n_363),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_427),
.A2(n_431),
.B(n_408),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_385),
.B(n_348),
.C(n_364),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_429),
.B(n_432),
.C(n_437),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_400),
.B(n_341),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_430),
.B(n_420),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_416),
.B(n_357),
.C(n_355),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_433),
.A2(n_419),
.B1(n_372),
.B2(n_374),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_395),
.A2(n_349),
.B(n_360),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_434),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_403),
.B(n_355),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_394),
.B(n_344),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_406),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_439),
.B(n_442),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_394),
.B(n_344),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_440),
.B(n_445),
.C(n_447),
.Y(n_464)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_444),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_396),
.B(n_415),
.C(n_387),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_413),
.B(n_383),
.C(n_379),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_448),
.B(n_449),
.Y(n_457)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_390),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_390),
.Y(n_450)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_450),
.Y(n_473)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_398),
.Y(n_451)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_451),
.Y(n_475)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_398),
.Y(n_452)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_452),
.Y(n_476)
);

AO22x1_ASAP7_75t_L g453 ( 
.A1(n_409),
.A2(n_376),
.B1(n_365),
.B2(n_371),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_453),
.A2(n_388),
.B1(n_395),
.B2(n_397),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_408),
.B(n_376),
.C(n_371),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_454),
.B(n_411),
.C(n_405),
.Y(n_468)
);

NOR2xp67_ASAP7_75t_SL g499 ( 
.A(n_455),
.B(n_433),
.Y(n_499)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_456),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_441),
.A2(n_391),
.B1(n_389),
.B2(n_397),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_459),
.A2(n_460),
.B1(n_465),
.B2(n_466),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_426),
.B(n_392),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_461),
.B(n_462),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_444),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_441),
.A2(n_402),
.B1(n_417),
.B2(n_393),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_446),
.A2(n_399),
.B1(n_410),
.B2(n_418),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_442),
.A2(n_414),
.B1(n_407),
.B2(n_386),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_467),
.A2(n_479),
.B1(n_481),
.B2(n_449),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_468),
.B(n_474),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_429),
.B(n_421),
.C(n_404),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_470),
.B(n_472),
.C(n_477),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_423),
.B(n_412),
.C(n_365),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_432),
.B(n_412),
.C(n_366),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_454),
.Y(n_478)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_478),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_442),
.A2(n_412),
.B1(n_359),
.B2(n_366),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_443),
.A2(n_412),
.B1(n_374),
.B2(n_281),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_437),
.B(n_282),
.C(n_244),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_482),
.B(n_448),
.C(n_436),
.Y(n_489)
);

BUFx12_ASAP7_75t_L g483 ( 
.A(n_479),
.Y(n_483)
);

INVxp33_ASAP7_75t_L g523 ( 
.A(n_483),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_468),
.B(n_426),
.Y(n_484)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_484),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_469),
.B(n_440),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_487),
.B(n_497),
.Y(n_513)
);

BUFx12_ASAP7_75t_L g488 ( 
.A(n_482),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_488),
.B(n_490),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_489),
.B(n_491),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_467),
.B(n_439),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_458),
.A2(n_434),
.B(n_431),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_464),
.B(n_445),
.C(n_447),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_492),
.B(n_495),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_471),
.B(n_428),
.Y(n_493)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_493),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_458),
.B(n_453),
.Y(n_494)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_494),
.Y(n_524)
);

BUFx12_ASAP7_75t_L g495 ( 
.A(n_464),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_466),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_496),
.B(n_501),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_480),
.A2(n_438),
.B(n_453),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_499),
.B(n_469),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_500),
.A2(n_465),
.B1(n_427),
.B2(n_476),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_477),
.B(n_472),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_463),
.B(n_435),
.C(n_438),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_505),
.B(n_470),
.C(n_455),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_457),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_506),
.A2(n_481),
.B1(n_480),
.B2(n_459),
.Y(n_507)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_507),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_R g508 ( 
.A(n_486),
.B(n_456),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_508),
.B(n_518),
.Y(n_530)
);

AOI22x1_ASAP7_75t_L g534 ( 
.A1(n_511),
.A2(n_483),
.B1(n_484),
.B2(n_503),
.Y(n_534)
);

NOR2xp67_ASAP7_75t_L g531 ( 
.A(n_514),
.B(n_489),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_515),
.B(n_487),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_485),
.B(n_463),
.C(n_422),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_486),
.A2(n_425),
.B(n_424),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_519),
.A2(n_497),
.B(n_494),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_498),
.A2(n_496),
.B1(n_500),
.B2(n_506),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_520),
.A2(n_523),
.B1(n_524),
.B2(n_510),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_485),
.B(n_473),
.C(n_475),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_521),
.B(n_522),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_492),
.B(n_272),
.C(n_234),
.Y(n_522)
);

FAx1_ASAP7_75t_SL g526 ( 
.A(n_508),
.B(n_499),
.CI(n_514),
.CON(n_526),
.SN(n_526)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_526),
.B(n_527),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_517),
.B(n_505),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_528),
.B(n_529),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_531),
.A2(n_532),
.B(n_515),
.Y(n_543)
);

NAND2x1p5_ASAP7_75t_L g532 ( 
.A(n_513),
.B(n_493),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_534),
.B(n_537),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_518),
.B(n_504),
.C(n_503),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_535),
.B(n_538),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_521),
.B(n_502),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_536),
.B(n_540),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_512),
.B(n_495),
.C(n_491),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_525),
.B(n_260),
.Y(n_540)
);

OAI21xp33_ASAP7_75t_L g541 ( 
.A1(n_530),
.A2(n_509),
.B(n_522),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g552 ( 
.A1(n_541),
.A2(n_542),
.B(n_543),
.Y(n_552)
);

A2O1A1Ixp33_ASAP7_75t_SL g542 ( 
.A1(n_529),
.A2(n_523),
.B(n_509),
.C(n_483),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_538),
.A2(n_513),
.B(n_516),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_544),
.A2(n_547),
.B1(n_545),
.B2(n_551),
.Y(n_556)
);

AOI221xp5_ASAP7_75t_L g549 ( 
.A1(n_533),
.A2(n_520),
.B1(n_519),
.B2(n_495),
.C(n_483),
.Y(n_549)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_549),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_535),
.B(n_233),
.Y(n_550)
);

NOR2xp67_ASAP7_75t_L g553 ( 
.A(n_550),
.B(n_539),
.Y(n_553)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_553),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_548),
.B(n_534),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_554),
.A2(n_557),
.B(n_558),
.Y(n_560)
);

NAND2xp33_ASAP7_75t_SL g562 ( 
.A(n_556),
.B(n_526),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_546),
.B(n_537),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_542),
.B(n_532),
.C(n_527),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_SL g561 ( 
.A1(n_555),
.A2(n_552),
.B(n_526),
.Y(n_561)
);

MAJx2_ASAP7_75t_L g564 ( 
.A(n_561),
.B(n_554),
.C(n_488),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_562),
.B(n_488),
.Y(n_565)
);

O2A1O1Ixp33_ASAP7_75t_SL g563 ( 
.A1(n_559),
.A2(n_542),
.B(n_558),
.C(n_557),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_563),
.A2(n_272),
.B(n_234),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_SL g566 ( 
.A1(n_564),
.A2(n_565),
.B(n_560),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g568 ( 
.A1(n_566),
.A2(n_567),
.B1(n_233),
.B2(n_15),
.Y(n_568)
);

AOI31xp67_ASAP7_75t_L g569 ( 
.A1(n_568),
.A2(n_15),
.A3(n_233),
.B(n_328),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_569),
.B(n_15),
.Y(n_570)
);


endmodule