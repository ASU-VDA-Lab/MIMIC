module fake_jpeg_13_n_256 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_107;
wire n_39;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_3),
.B(n_1),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_45),
.Y(n_118)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_23),
.B(n_14),
.Y(n_47)
);

OAI21xp33_ASAP7_75t_L g120 ( 
.A1(n_47),
.A2(n_50),
.B(n_51),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_23),
.B(n_14),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_22),
.B(n_0),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_3),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_56),
.B(n_58),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_26),
.B(n_4),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_5),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_78),
.Y(n_91)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_60),
.Y(n_94)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_67),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_69),
.Y(n_100)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_71),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_36),
.B(n_5),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_74),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_37),
.B(n_5),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_6),
.Y(n_105)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_76),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_9),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_31),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_52),
.A2(n_32),
.B1(n_28),
.B2(n_37),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_82),
.A2(n_87),
.B1(n_118),
.B2(n_88),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_58),
.B(n_41),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_84),
.B(n_106),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_40),
.B1(n_38),
.B2(n_17),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_85),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_53),
.A2(n_32),
.B1(n_40),
.B2(n_17),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_47),
.A2(n_50),
.B(n_59),
.C(n_56),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_90),
.B(n_105),
.Y(n_134)
);

AO22x1_ASAP7_75t_SL g99 ( 
.A1(n_77),
.A2(n_38),
.B1(n_41),
.B2(n_31),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_115),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_67),
.A2(n_79),
.B1(n_57),
.B2(n_43),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_101),
.B(n_107),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_48),
.B(n_39),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_62),
.B(n_39),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_64),
.B(n_6),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_94),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_6),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_113),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_60),
.B(n_8),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_45),
.B(n_8),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_9),
.Y(n_126)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_125),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_126),
.B(n_131),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_127),
.A2(n_129),
.B1(n_141),
.B2(n_93),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_100),
.A2(n_34),
.B1(n_116),
.B2(n_110),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_34),
.B1(n_81),
.B2(n_92),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_130),
.A2(n_138),
.B1(n_140),
.B2(n_132),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_117),
.Y(n_131)
);

INVx3_ASAP7_75t_SL g132 ( 
.A(n_110),
.Y(n_132)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_132),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_100),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_133),
.B(n_138),
.Y(n_171)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_140),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_80),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_142),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_95),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_90),
.B(n_86),
.Y(n_139)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_134),
.C(n_145),
.Y(n_166)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_91),
.B(n_102),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_91),
.B(n_108),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_144),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_149),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_148),
.B(n_154),
.Y(n_179)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

AND2x2_ASAP7_75t_SL g151 ( 
.A(n_118),
.B(n_103),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_144),
.C(n_155),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_103),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_153),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_87),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_155),
.Y(n_175)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_150),
.A2(n_82),
.B1(n_119),
.B2(n_88),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_168),
.B1(n_152),
.B2(n_146),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_133),
.A2(n_93),
.B(n_83),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_157),
.B(n_166),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_151),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_174),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_119),
.B(n_83),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_163),
.A2(n_157),
.B(n_177),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_128),
.A2(n_146),
.B1(n_132),
.B2(n_139),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_169),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_122),
.B(n_124),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_128),
.B(n_148),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_151),
.C(n_123),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_128),
.B(n_122),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_179),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_188),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_184),
.C(n_194),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_145),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_135),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_189),
.Y(n_210)
);

AO21x1_ASAP7_75t_L g186 ( 
.A1(n_172),
.A2(n_149),
.B(n_136),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_186),
.A2(n_196),
.B(n_169),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_178),
.A2(n_158),
.B1(n_163),
.B2(n_171),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_147),
.B1(n_125),
.B2(n_141),
.Y(n_191)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_191),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_166),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_197),
.B(n_199),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_165),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_198),
.B(n_177),
.Y(n_200)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_202),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_159),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_159),
.Y(n_204)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_204),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_186),
.Y(n_205)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_205),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_173),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_207),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_198),
.Y(n_208)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_208),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_211),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_184),
.Y(n_212)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_212),
.Y(n_222)
);

AOI21x1_ASAP7_75t_SL g213 ( 
.A1(n_196),
.A2(n_175),
.B(n_167),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_187),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_173),
.Y(n_214)
);

OAI321xp33_ASAP7_75t_L g218 ( 
.A1(n_214),
.A2(n_192),
.A3(n_195),
.B1(n_183),
.B2(n_199),
.C(n_182),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_192),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_220),
.C(n_225),
.Y(n_230)
);

OA21x2_ASAP7_75t_SL g234 ( 
.A1(n_218),
.A2(n_221),
.B(n_201),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_195),
.C(n_180),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_175),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_187),
.Y(n_229)
);

OAI321xp33_ASAP7_75t_L g227 ( 
.A1(n_215),
.A2(n_201),
.A3(n_210),
.B1(n_204),
.B2(n_202),
.C(n_200),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_231),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_209),
.Y(n_228)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_228),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_232),
.Y(n_241)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_219),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_223),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_234),
.C(n_235),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_211),
.Y(n_235)
);

AOI321xp33_ASAP7_75t_L g237 ( 
.A1(n_235),
.A2(n_224),
.A3(n_222),
.B1(n_220),
.B2(n_216),
.C(n_225),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_237),
.B(n_213),
.Y(n_246)
);

NOR2x1p5_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_201),
.Y(n_240)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_240),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_230),
.C(n_239),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_244),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_239),
.A2(n_229),
.B(n_226),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_243),
.A2(n_240),
.B(n_245),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_238),
.B(n_230),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_246),
.B(n_241),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_249),
.Y(n_252)
);

OAI221xp5_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_203),
.B1(n_193),
.B2(n_180),
.C(n_170),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_175),
.C(n_167),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_193),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_170),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_254),
.B(n_252),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_251),
.Y(n_256)
);


endmodule