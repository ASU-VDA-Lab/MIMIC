module fake_ibex_537_n_7783 (n_151, n_85, n_599, n_778, n_822, n_1042, n_507, n_743, n_1060, n_540, n_754, n_395, n_1011, n_84, n_64, n_992, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_1041, n_688, n_130, n_177, n_946, n_707, n_76, n_273, n_309, n_330, n_926, n_9, n_1031, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_947, n_972, n_981, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_956, n_790, n_920, n_452, n_86, n_70, n_664, n_1067, n_255, n_175, n_586, n_773, n_994, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_962, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_957, n_1015, n_678, n_663, n_969, n_194, n_249, n_334, n_634, n_733, n_961, n_991, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_1034, n_371, n_974, n_1036, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_959, n_258, n_861, n_1018, n_1044, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_1077, n_43, n_216, n_996, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_1045, n_753, n_645, n_500, n_747, n_963, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1061, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_1056, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_1010, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_948, n_158, n_1029, n_859, n_259, n_276, n_339, n_470, n_770, n_965, n_210, n_348, n_220, n_875, n_941, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_989, n_373, n_1051, n_854, n_1008, n_458, n_244, n_73, n_1053, n_343, n_310, n_714, n_1076, n_1032, n_936, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_967, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_1055, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_1025, n_465, n_1057, n_1068, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_1013, n_982, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_1024, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_977, n_1075, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_215, n_279, n_49, n_1037, n_374, n_235, n_464, n_538, n_669, n_838, n_987, n_750, n_1021, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_1052, n_852, n_789, n_880, n_654, n_656, n_1014, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_1023, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_944, n_1001, n_156, n_570, n_126, n_623, n_585, n_1030, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_980, n_454, n_1070, n_1074, n_777, n_1017, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_953, n_625, n_968, n_619, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_1064, n_1071, n_207, n_922, n_438, n_851, n_993, n_1012, n_1028, n_689, n_960, n_1022, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_973, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_999, n_1038, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_1009, n_635, n_979, n_844, n_1066, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_1020, n_847, n_830, n_1062, n_1004, n_473, n_1027, n_445, n_629, n_335, n_413, n_1072, n_82, n_263, n_1069, n_27, n_573, n_353, n_966, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_949, n_1007, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_954, n_363, n_1006, n_402, n_725, n_180, n_369, n_976, n_596, n_201, n_699, n_14, n_1063, n_351, n_368, n_456, n_834, n_257, n_77, n_998, n_935, n_869, n_925, n_718, n_801, n_918, n_1054, n_44, n_672, n_1039, n_722, n_401, n_1046, n_553, n_554, n_1043, n_66, n_735, n_305, n_882, n_942, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_955, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_943, n_1049, n_763, n_745, n_329, n_447, n_940, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_1065, n_592, n_986, n_495, n_762, n_410, n_905, n_308, n_975, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_512, n_615, n_950, n_685, n_1026, n_283, n_366, n_397, n_111, n_803, n_894, n_1033, n_692, n_36, n_627, n_990, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_971, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_978, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_1019, n_1059, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_951, n_511, n_23, n_734, n_468, n_223, n_381, n_1073, n_525, n_815, n_919, n_780, n_535, n_1002, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_952, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_997, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_1016, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_958, n_485, n_870, n_46, n_284, n_811, n_1047, n_808, n_80, n_172, n_250, n_945, n_493, n_460, n_609, n_1040, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_1048, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_1005, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_985, n_572, n_867, n_983, n_1003, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_970, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_1058, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_964, n_424, n_565, n_916, n_823, n_701, n_271, n_995, n_241, n_68, n_503, n_292, n_807, n_984, n_394, n_79, n_1000, n_81, n_35, n_364, n_687, n_895, n_988, n_159, n_202, n_231, n_298, n_587, n_1035, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_1050, n_7783);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_1042;
input n_507;
input n_743;
input n_1060;
input n_540;
input n_754;
input n_395;
input n_1011;
input n_84;
input n_64;
input n_992;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_1041;
input n_688;
input n_130;
input n_177;
input n_946;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_9;
input n_1031;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_947;
input n_972;
input n_981;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_956;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_1067;
input n_255;
input n_175;
input n_586;
input n_773;
input n_994;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_962;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_957;
input n_1015;
input n_678;
input n_663;
input n_969;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_961;
input n_991;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_1034;
input n_371;
input n_974;
input n_1036;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_959;
input n_258;
input n_861;
input n_1018;
input n_1044;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_1077;
input n_43;
input n_216;
input n_996;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_1045;
input n_753;
input n_645;
input n_500;
input n_747;
input n_963;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1061;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_1056;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_1010;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_948;
input n_158;
input n_1029;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_965;
input n_210;
input n_348;
input n_220;
input n_875;
input n_941;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_989;
input n_373;
input n_1051;
input n_854;
input n_1008;
input n_458;
input n_244;
input n_73;
input n_1053;
input n_343;
input n_310;
input n_714;
input n_1076;
input n_1032;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_967;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_1055;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_1025;
input n_465;
input n_1057;
input n_1068;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_1013;
input n_982;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_1024;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_977;
input n_1075;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_215;
input n_279;
input n_49;
input n_1037;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_987;
input n_750;
input n_1021;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_1052;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_1014;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_1023;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_944;
input n_1001;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_1030;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_980;
input n_454;
input n_1070;
input n_1074;
input n_777;
input n_1017;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_953;
input n_625;
input n_968;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_1064;
input n_1071;
input n_207;
input n_922;
input n_438;
input n_851;
input n_993;
input n_1012;
input n_1028;
input n_689;
input n_960;
input n_1022;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_973;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_999;
input n_1038;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_1009;
input n_635;
input n_979;
input n_844;
input n_1066;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_1020;
input n_847;
input n_830;
input n_1062;
input n_1004;
input n_473;
input n_1027;
input n_445;
input n_629;
input n_335;
input n_413;
input n_1072;
input n_82;
input n_263;
input n_1069;
input n_27;
input n_573;
input n_353;
input n_966;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_949;
input n_1007;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_954;
input n_363;
input n_1006;
input n_402;
input n_725;
input n_180;
input n_369;
input n_976;
input n_596;
input n_201;
input n_699;
input n_14;
input n_1063;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_998;
input n_935;
input n_869;
input n_925;
input n_718;
input n_801;
input n_918;
input n_1054;
input n_44;
input n_672;
input n_1039;
input n_722;
input n_401;
input n_1046;
input n_553;
input n_554;
input n_1043;
input n_66;
input n_735;
input n_305;
input n_882;
input n_942;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_955;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_943;
input n_1049;
input n_763;
input n_745;
input n_329;
input n_447;
input n_940;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_1065;
input n_592;
input n_986;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_975;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_512;
input n_615;
input n_950;
input n_685;
input n_1026;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_1033;
input n_692;
input n_36;
input n_627;
input n_990;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_971;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_978;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_1019;
input n_1059;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_951;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_1073;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_1002;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_952;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_997;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_1016;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_958;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_1047;
input n_808;
input n_80;
input n_172;
input n_250;
input n_945;
input n_493;
input n_460;
input n_609;
input n_1040;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_1048;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_1005;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_985;
input n_572;
input n_867;
input n_983;
input n_1003;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_970;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_1058;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_964;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_995;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_984;
input n_394;
input n_79;
input n_1000;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_988;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_1035;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;
input n_1050;

output n_7783;

wire n_4557;
wire n_6873;
wire n_6210;
wire n_5285;
wire n_6516;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_4983;
wire n_3548;
wire n_5647;
wire n_7170;
wire n_1382;
wire n_2949;
wire n_2840;
wire n_6537;
wire n_3319;
wire n_3915;
wire n_5002;
wire n_5155;
wire n_5130;
wire n_7029;
wire n_4204;
wire n_5899;
wire n_6259;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_3817;
wire n_2038;
wire n_2504;
wire n_7042;
wire n_4607;
wire n_4514;
wire n_3674;
wire n_4249;
wire n_4931;
wire n_1859;
wire n_5827;
wire n_4805;
wire n_1765;
wire n_2392;
wire n_5008;
wire n_6183;
wire n_3280;
wire n_7262;
wire n_7551;
wire n_6616;
wire n_6848;
wire n_4371;
wire n_7766;
wire n_4601;
wire n_6035;
wire n_5858;
wire n_5879;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1782;
wire n_2889;
wire n_6567;
wire n_7063;
wire n_2391;
wire n_4585;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_4169;
wire n_6744;
wire n_7707;
wire n_3570;
wire n_5760;
wire n_4875;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2506;
wire n_7589;
wire n_6229;
wire n_7643;
wire n_3598;
wire n_1752;
wire n_4172;
wire n_6639;
wire n_1730;
wire n_5243;
wire n_3479;
wire n_5587;
wire n_3751;
wire n_3262;
wire n_4673;
wire n_3537;
wire n_5667;
wire n_2343;
wire n_5615;
wire n_1480;
wire n_7147;
wire n_6327;
wire n_1463;
wire n_1823;
wire n_4781;
wire n_6256;
wire n_4423;
wire n_5517;
wire n_1766;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_7067;
wire n_5962;
wire n_3347;
wire n_3395;
wire n_4808;
wire n_6658;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_6842;
wire n_4526;
wire n_6286;
wire n_3472;
wire n_7485;
wire n_5922;
wire n_1981;
wire n_7636;
wire n_3976;
wire n_4348;
wire n_5931;
wire n_7450;
wire n_7492;
wire n_6760;
wire n_7396;
wire n_3807;
wire n_2998;
wire n_3845;
wire n_7082;
wire n_2163;
wire n_4450;
wire n_4467;
wire n_6159;
wire n_6517;
wire n_7313;
wire n_7305;
wire n_4801;
wire n_6005;
wire n_3639;
wire n_5809;
wire n_7332;
wire n_1664;
wire n_4144;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4955;
wire n_3208;
wire n_5588;
wire n_4569;
wire n_5404;
wire n_3671;
wire n_7673;
wire n_1778;
wire n_7151;
wire n_2839;
wire n_7013;
wire n_4998;
wire n_1698;
wire n_1496;
wire n_2333;
wire n_2705;
wire n_5505;
wire n_1214;
wire n_1274;
wire n_1595;
wire n_6530;
wire n_4510;
wire n_5658;
wire n_4567;
wire n_7672;
wire n_5151;
wire n_2362;
wire n_5478;
wire n_2822;
wire n_1306;
wire n_5994;
wire n_1493;
wire n_2597;
wire n_2774;
wire n_7776;
wire n_6602;
wire n_7753;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_5037;
wire n_5878;
wire n_5716;
wire n_1960;
wire n_6562;
wire n_7397;
wire n_7324;
wire n_3979;
wire n_3714;
wire n_6534;
wire n_6629;
wire n_7105;
wire n_2844;
wire n_6192;
wire n_3565;
wire n_7560;
wire n_5304;
wire n_3883;
wire n_5866;
wire n_5941;
wire n_3943;
wire n_4563;
wire n_1309;
wire n_5882;
wire n_1316;
wire n_1562;
wire n_6102;
wire n_7187;
wire n_4854;
wire n_6732;
wire n_3769;
wire n_6456;
wire n_1445;
wire n_6026;
wire n_2147;
wire n_5591;
wire n_6083;
wire n_7229;
wire n_2253;
wire n_4479;
wire n_5381;
wire n_3858;
wire n_4173;
wire n_6674;
wire n_6486;
wire n_5261;
wire n_5895;
wire n_7099;
wire n_5944;
wire n_6328;
wire n_5673;
wire n_7251;
wire n_7189;
wire n_1078;
wire n_4422;
wire n_5743;
wire n_6868;
wire n_1865;
wire n_5033;
wire n_6491;
wire n_4786;
wire n_4842;
wire n_1170;
wire n_3842;
wire n_2980;
wire n_7706;
wire n_6219;
wire n_5075;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_6241;
wire n_7507;
wire n_1305;
wire n_2088;
wire n_6724;
wire n_1248;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_7097;
wire n_3780;
wire n_5571;
wire n_1653;
wire n_1375;
wire n_6254;
wire n_1118;
wire n_6066;
wire n_7241;
wire n_1881;
wire n_3798;
wire n_5241;
wire n_4809;
wire n_3060;
wire n_5129;
wire n_4124;
wire n_4499;
wire n_1350;
wire n_3627;
wire n_5191;
wire n_7264;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_5259;
wire n_3293;
wire n_7372;
wire n_2550;
wire n_5913;
wire n_6302;
wire n_6580;
wire n_7607;
wire n_5266;
wire n_3381;
wire n_2750;
wire n_1650;
wire n_1453;
wire n_5580;
wire n_1108;
wire n_6078;
wire n_7521;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_4714;
wire n_5660;
wire n_5955;
wire n_1209;
wire n_5419;
wire n_3732;
wire n_6070;
wire n_6926;
wire n_3295;
wire n_3199;
wire n_1616;
wire n_6625;
wire n_7628;
wire n_2389;
wire n_5612;
wire n_6408;
wire n_6638;
wire n_7358;
wire n_2107;
wire n_3435;
wire n_4828;
wire n_4480;
wire n_1613;
wire n_3874;
wire n_6878;
wire n_2782;
wire n_4258;
wire n_1549;
wire n_4290;
wire n_1531;
wire n_2919;
wire n_6019;
wire n_4577;
wire n_7316;
wire n_1424;
wire n_2444;
wire n_2625;
wire n_3652;
wire n_4913;
wire n_2199;
wire n_1610;
wire n_4398;
wire n_7207;
wire n_1298;
wire n_1844;
wire n_6485;
wire n_4055;
wire n_3194;
wire n_4692;
wire n_7112;
wire n_7083;
wire n_5987;
wire n_6421;
wire n_6009;
wire n_2431;
wire n_2084;
wire n_1243;
wire n_7026;
wire n_3572;
wire n_6114;
wire n_6996;
wire n_1121;
wire n_4823;
wire n_7366;
wire n_5195;
wire n_7657;
wire n_5541;
wire n_7033;
wire n_6081;
wire n_3951;
wire n_4927;
wire n_3355;
wire n_2019;
wire n_1407;
wire n_4680;
wire n_1821;
wire n_7103;
wire n_5609;
wire n_5904;
wire n_4757;
wire n_5254;
wire n_6334;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_5423;
wire n_4653;
wire n_3466;
wire n_3370;
wire n_6606;
wire n_1504;
wire n_6864;
wire n_1781;
wire n_4331;
wire n_7733;
wire n_2028;
wire n_3678;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_5732;
wire n_5141;
wire n_1293;
wire n_7711;
wire n_3968;
wire n_4825;
wire n_6178;
wire n_3950;
wire n_5252;
wire n_6209;
wire n_7445;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_4623;
wire n_4523;
wire n_4411;
wire n_3811;
wire n_6941;
wire n_1271;
wire n_6011;
wire n_7667;
wire n_3416;
wire n_6824;
wire n_3147;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_7140;
wire n_4225;
wire n_7169;
wire n_5238;
wire n_6533;
wire n_3859;
wire n_6540;
wire n_4489;
wire n_6912;
wire n_3455;
wire n_6940;
wire n_1591;
wire n_7048;
wire n_2289;
wire n_2841;
wire n_4271;
wire n_7303;
wire n_1409;
wire n_2744;
wire n_3524;
wire n_6085;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_4404;
wire n_1521;
wire n_5502;
wire n_3054;
wire n_2456;
wire n_2924;
wire n_5288;
wire n_2264;
wire n_1987;
wire n_7192;
wire n_5749;
wire n_1129;
wire n_1244;
wire n_7639;
wire n_3365;
wire n_4974;
wire n_6802;
wire n_4725;
wire n_6691;
wire n_6431;
wire n_1932;
wire n_3775;
wire n_6196;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_7394;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_1715;
wire n_6377;
wire n_3300;
wire n_5969;
wire n_5920;
wire n_1713;
wire n_3621;
wire n_2036;
wire n_1255;
wire n_6855;
wire n_2740;
wire n_2622;
wire n_4250;
wire n_7003;
wire n_1218;
wire n_4572;
wire n_5705;
wire n_4374;
wire n_6146;
wire n_7161;
wire n_3708;
wire n_2626;
wire n_1446;
wire n_7723;
wire n_7748;
wire n_6958;
wire n_3218;
wire n_2880;
wire n_5887;
wire n_5948;
wire n_7226;
wire n_2423;
wire n_3849;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_4469;
wire n_2580;
wire n_3222;
wire n_3529;
wire n_6711;
wire n_6124;
wire n_3352;
wire n_4180;
wire n_2964;
wire n_4062;
wire n_1498;
wire n_7356;
wire n_5199;
wire n_7377;
wire n_1207;
wire n_1735;
wire n_3813;
wire n_1825;
wire n_4232;
wire n_7360;
wire n_7315;
wire n_4199;
wire n_6061;
wire n_5099;
wire n_1210;
wire n_7081;
wire n_6136;
wire n_7559;
wire n_4033;
wire n_2522;
wire n_4608;
wire n_7446;
wire n_1201;
wire n_5859;
wire n_7224;
wire n_1246;
wire n_5258;
wire n_4231;
wire n_7541;
wire n_6187;
wire n_1724;
wire n_2838;
wire n_1540;
wire n_3243;
wire n_7583;
wire n_3214;
wire n_1890;
wire n_3128;
wire n_4073;
wire n_6402;
wire n_2549;
wire n_4325;
wire n_7131;
wire n_2440;
wire n_4113;
wire n_7777;
wire n_1440;
wire n_4646;
wire n_7155;
wire n_6305;
wire n_1751;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_4819;
wire n_4261;
wire n_4884;
wire n_1083;
wire n_3205;
wire n_4490;
wire n_2358;
wire n_6971;
wire n_7553;
wire n_6128;
wire n_2361;
wire n_6804;
wire n_4128;
wire n_5213;
wire n_6469;
wire n_5354;
wire n_2062;
wire n_7700;
wire n_3932;
wire n_2339;
wire n_7338;
wire n_1963;
wire n_1418;
wire n_1137;
wire n_2552;
wire n_7221;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_3345;
wire n_6714;
wire n_4114;
wire n_6983;
wire n_1776;
wire n_6113;
wire n_3544;
wire n_5049;
wire n_1279;
wire n_6857;
wire n_4209;
wire n_3692;
wire n_5163;
wire n_1408;
wire n_5707;
wire n_3913;
wire n_3535;
wire n_6859;
wire n_2287;
wire n_3597;
wire n_4190;
wire n_7101;
wire n_2954;
wire n_6379;
wire n_6911;
wire n_6766;
wire n_2046;
wire n_6454;
wire n_4443;
wire n_4151;
wire n_4625;
wire n_4170;
wire n_7692;
wire n_7173;
wire n_4424;
wire n_6570;
wire n_1465;
wire n_6071;
wire n_4674;
wire n_6893;
wire n_6450;
wire n_1232;
wire n_2715;
wire n_6270;
wire n_4679;
wire n_6065;
wire n_7530;
wire n_1345;
wire n_4456;
wire n_5574;
wire n_1590;
wire n_7729;
wire n_7349;
wire n_2133;
wire n_3553;
wire n_5081;
wire n_6850;
wire n_6332;
wire n_6345;
wire n_1471;
wire n_5385;
wire n_3441;
wire n_4559;
wire n_5336;
wire n_2551;
wire n_4641;
wire n_4064;
wire n_5668;
wire n_4110;
wire n_4379;
wire n_3397;
wire n_5310;
wire n_4145;
wire n_6507;
wire n_1627;
wire n_3880;
wire n_7749;
wire n_5192;
wire n_4664;
wire n_3829;
wire n_7690;
wire n_1864;
wire n_6827;
wire n_5206;
wire n_2010;
wire n_2733;
wire n_6120;
wire n_7068;
wire n_3796;
wire n_5719;
wire n_6544;
wire n_5157;
wire n_1836;
wire n_6384;
wire n_4753;
wire n_1420;
wire n_2651;
wire n_1699;
wire n_6699;
wire n_4894;
wire n_5892;
wire n_5216;
wire n_6901;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_4321;
wire n_5375;
wire n_2418;
wire n_1087;
wire n_1599;
wire n_3070;
wire n_3477;
wire n_1575;
wire n_6773;
wire n_4416;
wire n_7430;
wire n_5998;
wire n_4024;
wire n_5521;
wire n_3975;
wire n_3164;
wire n_6314;
wire n_1448;
wire n_3034;
wire n_6765;
wire n_7703;
wire n_6605;
wire n_5433;
wire n_2628;
wire n_4361;
wire n_1705;
wire n_4237;
wire n_2263;
wire n_3495;
wire n_3169;
wire n_6349;
wire n_3759;
wire n_4777;
wire n_7391;
wire n_4800;
wire n_3629;
wire n_5573;
wire n_7695;
wire n_5620;
wire n_4117;
wire n_6527;
wire n_7283;
wire n_2884;
wire n_3383;
wire n_7148;
wire n_3687;
wire n_6626;
wire n_4154;
wire n_3459;
wire n_6105;
wire n_6704;
wire n_2691;
wire n_2243;
wire n_3092;
wire n_7592;
wire n_5330;
wire n_4385;
wire n_2759;
wire n_3434;
wire n_7254;
wire n_2654;
wire n_7199;
wire n_5729;
wire n_2975;
wire n_2503;
wire n_4072;
wire n_1512;
wire n_4908;
wire n_3885;
wire n_7509;
wire n_1426;
wire n_2365;
wire n_6528;
wire n_2245;
wire n_3877;
wire n_6939;
wire n_5083;
wire n_3260;
wire n_6463;
wire n_2776;
wire n_6727;
wire n_2630;
wire n_6348;
wire n_1967;
wire n_1095;
wire n_6883;
wire n_5801;
wire n_3834;
wire n_5579;
wire n_1378;
wire n_7457;
wire n_3257;
wire n_2459;
wire n_6652;
wire n_2439;
wire n_7619;
wire n_7760;
wire n_1430;
wire n_5365;
wire n_2450;
wire n_6459;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_5263;
wire n_6950;
wire n_4851;
wire n_4963;
wire n_1122;
wire n_3387;
wire n_7327;
wire n_6126;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_2728;
wire n_4685;
wire n_6915;
wire n_6115;
wire n_3428;
wire n_5959;
wire n_6282;
wire n_2427;
wire n_5017;
wire n_1127;
wire n_5938;
wire n_7025;
wire n_1845;
wire n_3835;
wire n_7645;
wire n_3723;
wire n_3389;
wire n_5292;
wire n_2422;
wire n_6277;
wire n_5190;
wire n_1679;
wire n_2342;
wire n_5926;
wire n_2755;
wire n_6531;
wire n_2301;
wire n_6922;
wire n_1578;
wire n_2712;
wire n_5316;
wire n_4314;
wire n_6731;
wire n_6502;
wire n_2788;
wire n_2089;
wire n_7090;
wire n_1857;
wire n_7587;
wire n_7574;
wire n_1997;
wire n_7174;
wire n_3314;
wire n_5135;
wire n_1349;
wire n_7250;
wire n_3891;
wire n_4704;
wire n_1777;
wire n_3409;
wire n_6646;
wire n_1546;
wire n_6394;
wire n_4003;
wire n_4775;
wire n_3420;
wire n_5840;
wire n_4192;
wire n_4633;
wire n_1950;
wire n_6439;
wire n_6084;
wire n_4593;
wire n_3914;
wire n_3289;
wire n_6902;
wire n_1834;
wire n_3372;
wire n_7641;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_4488;
wire n_3405;
wire n_6837;
wire n_1657;
wire n_1741;
wire n_4264;
wire n_4183;
wire n_4118;
wire n_4302;
wire n_2138;
wire n_4916;
wire n_6767;
wire n_7102;
wire n_4858;
wire n_6733;
wire n_1914;
wire n_3833;
wire n_5833;
wire n_6723;
wire n_3339;
wire n_7177;
wire n_6900;
wire n_3673;
wire n_5792;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_3556;
wire n_5617;
wire n_1340;
wire n_2562;
wire n_6191;
wire n_3269;
wire n_7539;
wire n_5491;
wire n_2223;
wire n_5024;
wire n_3876;
wire n_4971;
wire n_1267;
wire n_2683;
wire n_3432;
wire n_5696;
wire n_1816;
wire n_7233;
wire n_4645;
wire n_4619;
wire n_2318;
wire n_2141;
wire n_1422;
wire n_6044;
wire n_4339;
wire n_5493;
wire n_4085;
wire n_3190;
wire n_3878;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_5406;
wire n_1754;
wire n_3686;
wire n_6595;
wire n_7742;
wire n_2679;
wire n_4028;
wire n_5704;
wire n_7031;
wire n_1517;
wire n_5973;
wire n_7012;
wire n_7238;
wire n_3670;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_4289;
wire n_7030;
wire n_7110;
wire n_5555;
wire n_1895;
wire n_1860;
wire n_5727;
wire n_6856;
wire n_5770;
wire n_1763;
wire n_6976;
wire n_3912;
wire n_5169;
wire n_1607;
wire n_6682;
wire n_2959;
wire n_2380;
wire n_2420;
wire n_3265;
wire n_2221;
wire n_5274;
wire n_1774;
wire n_7517;
wire n_2516;
wire n_2031;
wire n_7121;
wire n_1348;
wire n_7317;
wire n_1191;
wire n_4099;
wire n_7190;
wire n_3899;
wire n_6153;
wire n_4729;
wire n_5957;
wire n_7429;
wire n_1617;
wire n_2639;
wire n_5323;
wire n_6777;
wire n_3099;
wire n_6412;
wire n_4745;
wire n_4057;
wire n_7390;
wire n_2410;
wire n_7145;
wire n_3206;
wire n_2633;
wire n_2049;
wire n_6245;
wire n_2113;
wire n_1690;
wire n_6553;
wire n_4466;
wire n_4132;
wire n_3361;
wire n_6543;
wire n_5566;
wire n_7561;
wire n_7529;
wire n_6185;
wire n_6706;
wire n_5342;
wire n_6884;
wire n_4603;
wire n_1135;
wire n_4300;
wire n_3277;
wire n_7533;
wire n_2758;
wire n_5787;
wire n_6745;
wire n_7210;
wire n_4417;
wire n_5967;
wire n_1550;
wire n_1169;
wire n_6224;
wire n_1938;
wire n_3452;
wire n_7563;
wire n_4022;
wire n_5843;
wire n_2194;
wire n_6072;
wire n_4320;
wire n_1173;
wire n_2736;
wire n_2845;
wire n_3886;
wire n_7191;
wire n_1901;
wire n_5332;
wire n_6073;
wire n_3096;
wire n_6097;
wire n_2059;
wire n_1278;
wire n_5553;
wire n_4730;
wire n_5763;
wire n_4616;
wire n_4760;
wire n_1710;
wire n_3021;
wire n_6881;
wire n_1603;
wire n_5864;
wire n_5227;
wire n_7136;
wire n_3404;
wire n_2072;
wire n_2963;
wire n_1489;
wire n_1993;
wire n_4859;
wire n_7213;
wire n_1455;
wire n_2182;
wire n_3115;
wire n_5352;
wire n_4583;
wire n_7034;
wire n_1502;
wire n_4923;
wire n_3920;
wire n_5370;
wire n_4082;
wire n_3273;
wire n_4367;
wire n_4282;
wire n_5600;
wire n_4475;
wire n_2286;
wire n_2563;
wire n_4893;
wire n_6990;
wire n_3650;
wire n_6948;
wire n_5014;
wire n_3513;
wire n_2677;
wire n_2531;
wire n_6591;
wire n_4029;
wire n_3212;
wire n_1321;
wire n_1779;
wire n_2489;
wire n_6816;
wire n_7512;
wire n_2950;
wire n_2272;
wire n_3574;
wire n_2608;
wire n_6712;
wire n_5824;
wire n_6280;
wire n_7682;
wire n_5472;
wire n_5950;
wire n_3739;
wire n_2825;
wire n_7098;
wire n_4338;
wire n_5546;
wire n_6222;
wire n_5972;
wire n_4985;
wire n_2742;
wire n_3604;
wire n_1740;
wire n_3540;
wire n_2680;
wire n_1343;
wire n_1371;
wire n_4198;
wire n_5924;
wire n_4529;
wire n_2861;
wire n_2976;
wire n_6656;
wire n_7323;
wire n_2366;
wire n_6318;
wire n_6200;
wire n_7149;
wire n_7219;
wire n_4919;
wire n_7320;
wire n_7175;
wire n_4111;
wire n_4200;
wire n_1659;
wire n_4575;
wire n_4847;
wire n_4803;
wire n_1878;
wire n_1374;
wire n_7357;
wire n_2851;
wire n_2973;
wire n_3651;
wire n_6637;
wire n_4666;
wire n_5752;
wire n_1242;
wire n_2810;
wire n_1119;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_5233;
wire n_3438;
wire n_4835;
wire n_3464;
wire n_4390;
wire n_5977;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_5968;
wire n_2871;
wire n_2764;
wire n_5713;
wire n_3648;
wire n_3234;
wire n_6577;
wire n_4058;
wire n_6268;
wire n_5403;
wire n_7593;
wire n_4611;
wire n_5527;
wire n_2714;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_5831;
wire n_1459;
wire n_4032;
wire n_6032;
wire n_2232;
wire n_4541;
wire n_4530;
wire n_1570;
wire n_5048;
wire n_5671;
wire n_6129;
wire n_1303;
wire n_1994;
wire n_7449;
wire n_6058;
wire n_1526;
wire n_4268;
wire n_2367;
wire n_3236;
wire n_1961;
wire n_3013;
wire n_4265;
wire n_3062;
wire n_3806;
wire n_3256;
wire n_3126;
wire n_5834;
wire n_1257;
wire n_6641;
wire n_2864;
wire n_1632;
wire n_3104;
wire n_5951;
wire n_4895;
wire n_5480;
wire n_7663;
wire n_3354;
wire n_4069;
wire n_5289;
wire n_3373;
wire n_7218;
wire n_6863;
wire n_2784;
wire n_4140;
wire n_1909;
wire n_7292;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_6556;
wire n_4778;
wire n_4789;
wire n_2703;
wire n_6152;
wire n_7582;
wire n_2574;
wire n_7659;
wire n_7142;
wire n_5492;
wire n_1887;
wire n_6106;
wire n_7428;
wire n_3504;
wire n_3511;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_3101;
wire n_6805;
wire n_5260;
wire n_6416;
wire n_7602;
wire n_5069;
wire n_2364;
wire n_7133;
wire n_2641;
wire n_7306;
wire n_7202;
wire n_6771;
wire n_4751;
wire n_7730;
wire n_5930;
wire n_5309;
wire n_6695;
wire n_3774;
wire n_2494;
wire n_3863;
wire n_5782;
wire n_2228;
wire n_4474;
wire n_5646;
wire n_7691;
wire n_1518;
wire n_4350;
wire n_5327;
wire n_4478;
wire n_2872;
wire n_2411;
wire n_3539;
wire n_2266;
wire n_4473;
wire n_6673;
wire n_7138;
wire n_7370;
wire n_3761;
wire n_2830;
wire n_4675;
wire n_3083;
wire n_6978;
wire n_7626;
wire n_5927;
wire n_3844;
wire n_4049;
wire n_2044;
wire n_2091;
wire n_4945;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_5019;
wire n_4891;
wire n_6910;
wire n_2394;
wire n_1572;
wire n_7236;
wire n_1245;
wire n_4867;
wire n_7387;
wire n_2929;
wire n_6346;
wire n_4911;
wire n_5414;
wire n_1329;
wire n_2409;
wire n_6403;
wire n_2405;
wire n_2601;
wire n_4405;
wire n_3118;
wire n_6172;
wire n_7122;
wire n_3742;
wire n_6004;
wire n_3532;
wire n_6347;
wire n_6482;
wire n_7698;
wire n_5280;
wire n_5466;
wire n_5469;
wire n_6925;
wire n_7024;
wire n_6483;
wire n_4686;
wire n_7466;
wire n_6358;
wire n_4682;
wire n_5750;
wire n_5305;
wire n_2914;
wire n_1833;
wire n_6598;
wire n_6800;
wire n_7410;
wire n_5186;
wire n_7257;
wire n_1986;
wire n_2882;
wire n_4301;
wire n_2493;
wire n_6499;
wire n_6944;
wire n_6215;
wire n_2115;
wire n_2013;
wire n_1556;
wire n_3547;
wire n_4898;
wire n_6980;
wire n_3700;
wire n_5180;
wire n_6594;
wire n_6233;
wire n_4733;
wire n_5368;
wire n_6338;
wire n_5757;
wire n_3947;
wire n_4684;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_6621;
wire n_7282;
wire n_2532;
wire n_3782;
wire n_1720;
wire n_3831;
wire n_2293;
wire n_7495;
wire n_7334;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_6053;
wire n_2734;
wire n_1166;
wire n_7346;
wire n_5267;
wire n_7649;
wire n_6020;
wire n_2310;
wire n_2674;
wire n_1284;
wire n_7532;
wire n_7740;
wire n_6432;
wire n_6426;
wire n_2689;
wire n_1992;
wire n_4493;
wire n_4962;
wire n_1082;
wire n_5397;
wire n_4797;
wire n_2596;
wire n_1488;
wire n_7401;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_3606;
wire n_5232;
wire n_7245;
wire n_1866;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_6946;
wire n_5890;
wire n_4644;
wire n_4412;
wire n_6068;
wire n_5802;
wire n_4266;
wire n_5815;
wire n_5605;
wire n_6897;
wire n_3124;
wire n_2634;
wire n_2982;
wire n_5384;
wire n_6550;
wire n_3015;
wire n_3321;
wire n_3081;
wire n_4639;
wire n_2291;
wire n_5664;
wire n_4102;
wire n_3612;
wire n_2172;
wire n_1728;
wire n_5863;
wire n_1230;
wire n_7075;
wire n_7710;
wire n_3622;
wire n_5276;
wire n_3857;
wire n_6847;
wire n_6042;
wire n_2357;
wire n_5197;
wire n_4354;
wire n_5320;
wire n_2937;
wire n_3728;
wire n_5087;
wire n_5265;
wire n_4401;
wire n_4727;
wire n_7367;
wire n_6265;
wire n_4296;
wire n_5312;
wire n_5534;
wire n_2967;
wire n_6737;
wire n_3005;
wire n_4627;
wire n_6936;
wire n_5107;
wire n_6780;
wire n_4309;
wire n_4027;
wire n_7132;
wire n_7486;
wire n_6758;
wire n_2056;
wire n_2054;
wire n_2226;
wire n_1402;
wire n_3267;
wire n_3008;
wire n_6452;
wire n_2802;
wire n_4728;
wire n_7419;
wire n_2279;
wire n_1536;
wire n_1719;
wire n_5281;
wire n_4046;
wire n_7201;
wire n_2961;
wire n_6458;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_7555;
wire n_1736;
wire n_6176;
wire n_7265;
wire n_7232;
wire n_2907;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_6092;
wire n_7023;
wire n_3675;
wire n_7227;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_4901;
wire n_3133;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_5025;
wire n_4539;
wire n_1205;
wire n_5575;
wire n_2969;
wire n_6052;
wire n_5753;
wire n_3550;
wire n_5401;
wire n_7642;
wire n_5509;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_6468;
wire n_1414;
wire n_5506;
wire n_6063;
wire n_7273;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_3275;
wire n_2645;
wire n_7623;
wire n_5417;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_7774;
wire n_5015;
wire n_5372;
wire n_1675;
wire n_6909;
wire n_1551;
wire n_1533;
wire n_3792;
wire n_2515;
wire n_3089;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_3988;
wire n_3758;
wire n_6418;
wire n_2353;
wire n_4251;
wire n_4106;
wire n_3662;
wire n_6344;
wire n_1354;
wire n_3329;
wire n_1277;
wire n_5995;
wire n_3233;
wire n_3193;
wire n_2582;
wire n_7070;
wire n_5253;
wire n_3789;
wire n_6308;
wire n_2174;
wire n_6989;
wire n_2510;
wire n_7634;
wire n_2435;
wire n_3934;
wire n_2583;
wire n_1678;
wire n_4606;
wire n_1287;
wire n_1525;
wire n_6662;
wire n_6461;
wire n_7046;
wire n_1150;
wire n_1674;
wire n_6304;
wire n_3980;
wire n_2912;
wire n_2710;
wire n_6617;
wire n_2970;
wire n_1393;
wire n_4691;
wire n_5937;
wire n_2978;
wire n_5291;
wire n_3502;
wire n_5460;
wire n_3935;
wire n_5379;
wire n_1854;
wire n_1084;
wire n_2804;
wire n_5390;
wire n_5691;
wire n_4926;
wire n_5043;
wire n_6549;
wire n_7194;
wire n_4688;
wire n_5097;
wire n_5675;
wire n_3144;
wire n_4234;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_4932;
wire n_6179;
wire n_1930;
wire n_5577;
wire n_1234;
wire n_4881;
wire n_7527;
wire n_7290;
wire n_3755;
wire n_1469;
wire n_4632;
wire n_7146;
wire n_3255;
wire n_1652;
wire n_2183;
wire n_6607;
wire n_1883;
wire n_2037;
wire n_4550;
wire n_6960;
wire n_1226;
wire n_7253;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_5181;
wire n_3105;
wire n_3146;
wire n_4892;
wire n_4343;
wire n_7615;
wire n_3931;
wire n_5745;
wire n_7434;
wire n_4421;
wire n_2322;
wire n_7477;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_7452;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_5893;
wire n_3843;
wire n_2847;
wire n_4399;
wire n_1308;
wire n_5067;
wire n_6823;
wire n_3904;
wire n_4378;
wire n_6455;
wire n_3729;
wire n_5637;
wire n_3484;
wire n_7414;
wire n_2485;
wire n_5614;
wire n_4477;
wire n_5177;
wire n_5643;
wire n_2179;
wire n_6725;
wire n_4654;
wire n_3984;
wire n_4233;
wire n_4765;
wire n_7475;
wire n_7775;
wire n_7184;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_5695;
wire n_3726;
wire n_6914;
wire n_5438;
wire n_4277;
wire n_4431;
wire n_7152;
wire n_4771;
wire n_4970;
wire n_4652;
wire n_6927;
wire n_5179;
wire n_3804;
wire n_1908;
wire n_6457;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_4285;
wire n_4928;
wire n_3251;
wire n_6916;
wire n_6973;
wire n_2921;
wire n_3724;
wire n_3192;
wire n_3753;
wire n_5683;
wire n_3566;
wire n_7554;
wire n_6564;
wire n_2820;
wire n_2311;
wire n_5701;
wire n_4403;
wire n_3242;
wire n_6566;
wire n_7114;
wire n_1654;
wire n_6428;
wire n_5774;
wire n_3330;
wire n_2707;
wire n_4746;
wire n_7354;
wire n_4382;
wire n_4002;
wire n_3631;
wire n_6808;
wire n_7609;
wire n_7037;
wire n_2537;
wire n_1130;
wire n_4545;
wire n_2643;
wire n_4246;
wire n_2336;
wire n_3987;
wire n_7709;
wire n_3969;
wire n_1081;
wire n_4437;
wire n_6747;
wire n_7335;
wire n_3856;
wire n_6496;
wire n_1155;
wire n_5394;
wire n_1292;
wire n_5462;
wire n_2432;
wire n_3043;
wire n_2273;
wire n_5428;
wire n_4491;
wire n_4672;
wire n_5001;
wire n_2421;
wire n_3237;
wire n_6095;
wire n_6787;
wire n_1970;
wire n_3946;
wire n_7183;
wire n_2953;
wire n_3949;
wire n_3507;
wire n_6150;
wire n_3926;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_2436;
wire n_1663;
wire n_6784;
wire n_4267;
wire n_5933;
wire n_4723;
wire n_7433;
wire n_2269;
wire n_6741;
wire n_2472;
wire n_2846;
wire n_3699;
wire n_4312;
wire n_5874;
wire n_5104;
wire n_2249;
wire n_3022;
wire n_4014;
wire n_3766;
wire n_3707;
wire n_7669;
wire n_4217;
wire n_3973;
wire n_5964;
wire n_5551;
wire n_5319;
wire n_4769;
wire n_4724;
wire n_2260;
wire n_5543;
wire n_4721;
wire n_2663;
wire n_3882;
wire n_6807;
wire n_2595;
wire n_5723;
wire n_5621;
wire n_6795;
wire n_7437;
wire n_6898;
wire n_5386;
wire n_4433;
wire n_5133;
wire n_5056;
wire n_6785;
wire n_7384;
wire n_7588;
wire n_6738;
wire n_3030;
wire n_5631;
wire n_6818;
wire n_5983;
wire n_7516;
wire n_5796;
wire n_4503;
wire n_6232;
wire n_3917;
wire n_3679;
wire n_7393;
wire n_4517;
wire n_6021;
wire n_3210;
wire n_3221;
wire n_4511;
wire n_6966;
wire n_1672;
wire n_4171;
wire n_3764;
wire n_5405;
wire n_6389;
wire n_3795;
wire n_6055;
wire n_4788;
wire n_4754;
wire n_1817;
wire n_5848;
wire n_5221;
wire n_1301;
wire n_5997;
wire n_4166;
wire n_2242;
wire n_4845;
wire n_1561;
wire n_5122;
wire n_2247;
wire n_3177;
wire n_3399;
wire n_5439;
wire n_6899;
wire n_4850;
wire n_1869;
wire n_7614;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_3676;
wire n_1753;
wire n_6351;
wire n_7503;
wire n_4610;
wire n_6441;
wire n_5854;
wire n_6754;
wire n_4067;
wire n_6822;
wire n_6849;
wire n_6796;
wire n_6836;
wire n_4997;
wire n_5906;
wire n_7355;
wire n_6755;
wire n_7608;
wire n_4393;
wire n_5205;
wire n_3777;
wire n_7084;
wire n_5916;
wire n_7685;
wire n_5993;
wire n_4553;
wire n_5240;
wire n_3961;
wire n_1520;
wire n_7515;
wire n_2509;
wire n_5714;
wire n_4283;
wire n_4174;
wire n_4870;
wire n_2399;
wire n_1370;
wire n_1708;
wire n_3038;
wire n_7483;
wire n_6476;
wire n_5828;
wire n_7648;
wire n_6276;
wire n_5907;
wire n_5284;
wire n_4804;
wire n_3716;
wire n_1649;
wire n_3450;
wire n_6669;
wire n_5357;
wire n_6717;
wire n_4994;
wire n_4518;
wire n_4732;
wire n_1936;
wire n_1717;
wire n_6040;
wire n_2257;
wire n_4856;
wire n_5088;
wire n_5250;
wire n_1467;
wire n_6388;
wire n_3217;
wire n_2511;
wire n_5461;
wire n_6298;
wire n_6988;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2661;
wire n_4079;
wire n_7256;
wire n_3573;
wire n_7652;
wire n_3563;
wire n_4993;
wire n_3510;
wire n_7172;
wire n_4248;
wire n_2334;
wire n_2350;
wire n_5958;
wire n_5619;
wire n_7117;
wire n_1709;
wire n_6655;
wire n_6541;
wire n_2649;
wire n_3607;
wire n_4476;
wire n_6460;
wire n_3241;
wire n_2746;
wire n_5471;
wire n_2256;
wire n_5210;
wire n_2445;
wire n_1980;
wire n_6790;
wire n_3583;
wire n_4987;
wire n_3832;
wire n_4649;
wire n_3508;
wire n_6295;
wire n_1862;
wire n_4693;
wire n_3415;
wire n_2355;
wire n_4992;
wire n_1543;
wire n_3386;
wire n_4568;
wire n_4359;
wire n_3814;
wire n_1441;
wire n_4573;
wire n_4105;
wire n_4206;
wire n_5273;
wire n_7722;
wire n_4177;
wire n_1888;
wire n_6497;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_5877;
wire n_6535;
wire n_5457;
wire n_5482;
wire n_4700;
wire n_2828;
wire n_1964;
wire n_6090;
wire n_3720;
wire n_1196;
wire n_6840;
wire n_1182;
wire n_4074;
wire n_5237;
wire n_5360;
wire n_3633;
wire n_1731;
wire n_5596;
wire n_2879;
wire n_3514;
wire n_3091;
wire n_5625;
wire n_4037;
wire n_4582;
wire n_5539;
wire n_3426;
wire n_7287;
wire n_4308;
wire n_2288;
wire n_3075;
wire n_1671;
wire n_6748;
wire n_3448;
wire n_3788;
wire n_6164;
wire n_6211;
wire n_2076;
wire n_3733;
wire n_1831;
wire n_4853;
wire n_6676;
wire n_6117;
wire n_6563;
wire n_1312;
wire n_5844;
wire n_6470;
wire n_7301;
wire n_6448;
wire n_3684;
wire n_6667;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_6018;
wire n_6094;
wire n_3970;
wire n_3291;
wire n_2454;
wire n_4008;
wire n_4973;
wire n_2829;
wire n_4966;
wire n_2968;
wire n_4494;
wire n_3473;
wire n_5362;
wire n_6236;
wire n_6208;
wire n_5294;
wire n_6197;
wire n_3263;
wire n_4501;
wire n_7156;
wire n_1772;
wire n_2858;
wire n_7780;
wire n_1283;
wire n_6552;
wire n_1421;
wire n_4922;
wire n_6237;
wire n_5089;
wire n_2424;
wire n_1793;
wire n_2573;
wire n_6993;
wire n_2390;
wire n_7544;
wire n_7203;
wire n_4402;
wire n_2793;
wire n_4813;
wire n_6653;
wire n_3098;
wire n_7732;
wire n_6449;
wire n_1711;
wire n_3069;
wire n_5465;
wire n_3107;
wire n_5488;
wire n_4134;
wire n_4131;
wire n_6539;
wire n_4330;
wire n_5832;
wire n_2176;
wire n_2805;
wire n_5165;
wire n_2319;
wire n_5678;
wire n_7658;
wire n_3757;
wire n_5811;
wire n_1933;
wire n_7408;
wire n_7605;
wire n_1842;
wire n_3364;
wire n_3429;
wire n_3306;
wire n_5234;
wire n_3787;
wire n_5140;
wire n_3445;
wire n_2080;
wire n_5655;
wire n_5514;
wire n_2554;
wire n_6130;
wire n_1676;
wire n_7476;
wire n_7624;
wire n_5020;
wire n_5225;
wire n_1136;
wire n_1918;
wire n_3642;
wire n_2461;
wire n_1229;
wire n_1490;
wire n_1179;
wire n_4818;
wire n_7566;
wire n_4462;
wire n_1153;
wire n_6560;
wire n_7307;
wire n_2787;
wire n_4540;
wire n_6987;
wire n_4187;
wire n_7684;
wire n_1273;
wire n_3821;
wire n_2930;
wire n_2616;
wire n_4979;
wire n_7409;
wire n_7087;
wire n_3503;
wire n_2441;
wire n_7280;
wire n_7680;
wire n_4063;
wire n_4362;
wire n_5318;
wire n_3312;
wire n_1848;
wire n_4009;
wire n_7107;
wire n_2650;
wire n_2888;
wire n_3614;
wire n_5946;
wire n_6131;
wire n_3394;
wire n_6207;
wire n_6984;
wire n_5942;
wire n_2530;
wire n_2792;
wire n_2372;
wire n_4191;
wire n_4965;
wire n_1522;
wire n_2523;
wire n_6701;
wire n_6326;
wire n_3488;
wire n_6365;
wire n_7288;
wire n_7248;
wire n_2832;
wire n_4991;
wire n_4525;
wire n_4011;
wire n_3526;
wire n_5242;
wire n_2142;
wire n_6519;
wire n_3703;
wire n_5116;
wire n_6635;
wire n_6907;
wire n_4554;
wire n_1260;
wire n_7038;
wire n_4097;
wire n_4861;
wire n_3239;
wire n_6155;
wire n_5953;
wire n_2600;
wire n_3952;
wire n_1171;
wire n_1126;
wire n_6151;
wire n_6074;
wire n_4596;
wire n_2434;
wire n_3578;
wire n_4734;
wire n_5947;
wire n_6661;
wire n_6730;
wire n_4492;
wire n_3470;
wire n_1738;
wire n_6370;
wire n_1729;
wire n_5563;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_7153;
wire n_5194;
wire n_7230;
wire n_4579;
wire n_5628;
wire n_6994;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_4936;
wire n_2097;
wire n_2109;
wire n_2648;
wire n_6262;
wire n_2398;
wire n_7572;
wire n_1593;
wire n_7308;
wire n_1775;
wire n_6889;
wire n_6361;
wire n_6803;
wire n_7481;
wire n_2570;
wire n_4025;
wire n_6751;
wire n_2184;
wire n_3948;
wire n_2842;
wire n_1400;
wire n_7403;
wire n_2469;
wire n_6024;
wire n_3074;
wire n_4640;
wire n_5790;
wire n_6523;
wire n_5746;
wire n_5883;
wire n_7369;
wire n_5630;
wire n_3136;
wire n_3108;
wire n_6696;
wire n_2395;
wire n_7089;
wire n_6062;
wire n_4059;
wire n_7258;
wire n_4130;
wire n_2752;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_4642;
wire n_3625;
wire n_1746;
wire n_2716;
wire n_2212;
wire n_6943;
wire n_4878;
wire n_1832;
wire n_1128;
wire n_2376;
wire n_3398;
wire n_3718;
wire n_6252;
wire n_7080;
wire n_7718;
wire n_5193;
wire n_2170;
wire n_6407;
wire n_4904;
wire n_1785;
wire n_3999;
wire n_1405;
wire n_4087;
wire n_7002;
wire n_5153;
wire n_6235;
wire n_5369;
wire n_7745;
wire n_6726;
wire n_7689;
wire n_3238;
wire n_6740;
wire n_4318;
wire n_3731;
wire n_3555;
wire n_3254;
wire n_5007;
wire n_4717;
wire n_4052;
wire n_6447;
wire n_6799;
wire n_2463;
wire n_6932;
wire n_6434;
wire n_2478;
wire n_3178;
wire n_4245;
wire n_7008;
wire n_3378;
wire n_5689;
wire n_3350;
wire n_6391;
wire n_5399;
wire n_4873;
wire n_6630;
wire n_6631;
wire n_3936;
wire n_1560;
wire n_5513;
wire n_3166;
wire n_3953;
wire n_3385;
wire n_1265;
wire n_2488;
wire n_2042;
wire n_5891;
wire n_1925;
wire n_6489;
wire n_7049;
wire n_1251;
wire n_6657;
wire n_3090;
wire n_1247;
wire n_5030;
wire n_3816;
wire n_5098;
wire n_5755;
wire n_4636;
wire n_7062;
wire n_7493;
wire n_5408;
wire n_4256;
wire n_1185;
wire n_3575;
wire n_6716;
wire n_6797;
wire n_2765;
wire n_4278;
wire n_6165;
wire n_6263;
wire n_6481;
wire n_4609;
wire n_5148;
wire n_7215;
wire n_7340;
wire n_4822;
wire n_6694;
wire n_2936;
wire n_7154;
wire n_2985;
wire n_3106;
wire n_6597;
wire n_4030;
wire n_4276;
wire n_6238;
wire n_4612;
wire n_1148;
wire n_1667;
wire n_6272;
wire n_5454;
wire n_3902;
wire n_1707;
wire n_4203;
wire n_5650;
wire n_2055;
wire n_4866;
wire n_2385;
wire n_6965;
wire n_3864;
wire n_3026;
wire n_3294;
wire n_4831;
wire n_5656;
wire n_1143;
wire n_6647;
wire n_7279;
wire n_7499;
wire n_2584;
wire n_4381;
wire n_5183;
wire n_7771;
wire n_2442;
wire n_5072;
wire n_4441;
wire n_2000;
wire n_4083;
wire n_2696;
wire n_4960;
wire n_5146;
wire n_6846;
wire n_5131;
wire n_1894;
wire n_2904;
wire n_3064;
wire n_2896;
wire n_4228;
wire n_4699;
wire n_5803;
wire n_1331;
wire n_1223;
wire n_5754;
wire n_1739;
wire n_3130;
wire n_1353;
wire n_7052;
wire n_5018;
wire n_2386;
wire n_7662;
wire n_3324;
wire n_3073;
wire n_2029;
wire n_4254;
wire n_4536;
wire n_7728;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_6931;
wire n_4924;
wire n_2238;
wire n_6398;
wire n_6700;
wire n_5786;
wire n_4138;
wire n_3100;
wire n_1727;
wire n_6366;
wire n_6853;
wire n_1294;
wire n_1351;
wire n_6679;
wire n_5035;
wire n_5425;
wire n_1380;
wire n_6036;
wire n_3336;
wire n_6104;
wire n_1291;
wire n_5742;
wire n_5901;
wire n_3763;
wire n_7158;
wire n_4284;
wire n_5943;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_6253;
wire n_7299;
wire n_1830;
wire n_6770;
wire n_3476;
wire n_3990;
wire n_2011;
wire n_4044;
wire n_5499;
wire n_7095;
wire n_7464;
wire n_1662;
wire n_7426;
wire n_3443;
wire n_5143;
wire n_3029;
wire n_4135;
wire n_7076;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_5302;
wire n_1660;
wire n_5640;
wire n_4000;
wire n_5841;
wire n_5011;
wire n_2556;
wire n_1537;
wire n_3908;
wire n_3696;
wire n_2902;
wire n_6242;
wire n_6660;
wire n_3608;
wire n_4269;
wire n_4016;
wire n_4915;
wire n_4286;
wire n_3048;
wire n_6414;
wire n_7666;
wire n_1962;
wire n_5296;
wire n_7246;
wire n_5159;
wire n_1952;
wire n_1624;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_7459;
wire n_2250;
wire n_1491;
wire n_3778;
wire n_7570;
wire n_2075;
wire n_4816;
wire n_6951;
wire n_3335;
wire n_4846;
wire n_3669;
wire n_1899;
wire n_4001;
wire n_6029;
wire n_2892;
wire n_3356;
wire n_4377;
wire n_3220;
wire n_3422;
wire n_5798;
wire n_2309;
wire n_2274;
wire n_6278;
wire n_6949;
wire n_5096;
wire n_6480;
wire n_7380;
wire n_6443;
wire n_3712;
wire n_5805;
wire n_5171;
wire n_2143;
wire n_4637;
wire n_4976;
wire n_4021;
wire n_5351;
wire n_2739;
wire n_2528;
wire n_7167;
wire n_7537;
wire n_2548;
wire n_3216;
wire n_6157;
wire n_6453;
wire n_3061;
wire n_3717;
wire n_3424;
wire n_3745;
wire n_3245;
wire n_6693;
wire n_4855;
wire n_5851;
wire n_4643;
wire n_5217;
wire n_6030;
wire n_4736;
wire n_2817;
wire n_1790;
wire n_4202;
wire n_3196;
wire n_5767;
wire n_4287;
wire n_2809;
wire n_6615;
wire n_3921;
wire n_3480;
wire n_7455;
wire n_1494;
wire n_2060;
wire n_2214;
wire n_7755;
wire n_1726;
wire n_5751;
wire n_6819;
wire n_1241;
wire n_5929;
wire n_2589;
wire n_5928;
wire n_1231;
wire n_1208;
wire n_1604;
wire n_4947;
wire n_3506;
wire n_1976;
wire n_1337;
wire n_2984;
wire n_4890;
wire n_4538;
wire n_4023;
wire n_3031;
wire n_4920;
wire n_5869;
wire n_5862;
wire n_1238;
wire n_3959;
wire n_6937;
wire n_4288;
wire n_7629;
wire n_2452;
wire n_6274;
wire n_2144;
wire n_4763;
wire n_7725;
wire n_2592;
wire n_2251;
wire n_5201;
wire n_1644;
wire n_4586;
wire n_6190;
wire n_3860;
wire n_5353;
wire n_1871;
wire n_2868;
wire n_3044;
wire n_3493;
wire n_2818;
wire n_7474;
wire n_3486;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_4034;
wire n_5444;
wire n_1149;
wire n_6860;
wire n_7739;
wire n_4905;
wire n_6100;
wire n_1457;
wire n_3172;
wire n_6833;
wire n_2159;
wire n_6865;
wire n_2700;
wire n_1222;
wire n_1630;
wire n_1959;
wire n_1198;
wire n_7135;
wire n_6794;
wire n_3637;
wire n_7216;
wire n_3393;
wire n_5772;
wire n_1261;
wire n_5520;
wire n_3327;
wire n_1114;
wire n_7487;
wire n_5277;
wire n_5900;
wire n_7421;
wire n_7694;
wire n_3647;
wire n_6240;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_1846;
wire n_1573;
wire n_7399;
wire n_1956;
wire n_7186;
wire n_5569;
wire n_5779;
wire n_4270;
wire n_2983;
wire n_4273;
wire n_7580;
wire n_7632;
wire n_6498;
wire n_6720;
wire n_1669;
wire n_7562;
wire n_6247;
wire n_5109;
wire n_1885;
wire n_1989;
wire n_5837;
wire n_5402;
wire n_1801;
wire n_3740;
wire n_3001;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_2576;
wire n_6854;
wire n_4344;
wire n_1342;
wire n_6574;
wire n_2756;
wire n_7197;
wire n_7015;
wire n_7747;
wire n_1175;
wire n_4408;
wire n_6832;
wire n_5473;
wire n_1221;
wire n_3875;
wire n_5113;
wire n_7066;
wire n_4341;
wire n_4759;
wire n_7688;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_6779;
wire n_2567;
wire n_5645;
wire n_7044;
wire n_1085;
wire n_2981;
wire n_2222;
wire n_4439;
wire n_5102;
wire n_6258;
wire n_7329;
wire n_6139;
wire n_5167;
wire n_7756;
wire n_4565;
wire n_5562;
wire n_7713;
wire n_1451;
wire n_7438;
wire n_4663;
wire n_2471;
wire n_5666;
wire n_1288;
wire n_1275;
wire n_4519;
wire n_2757;
wire n_1622;
wire n_3121;
wire n_2121;
wire n_6887;
wire n_4515;
wire n_1893;
wire n_5639;
wire n_5607;
wire n_7735;
wire n_2278;
wire n_6769;
wire n_6903;
wire n_2433;
wire n_7255;
wire n_2798;
wire n_3425;
wire n_1771;
wire n_3308;
wire n_6169;
wire n_1507;
wire n_5914;
wire n_1206;
wire n_3576;
wire n_5275;
wire n_3109;
wire n_4838;
wire n_2553;
wire n_4524;
wire n_2218;
wire n_6861;
wire n_2130;
wire n_4862;
wire n_7270;
wire n_5114;
wire n_7071;
wire n_7773;
wire n_6697;
wire n_4260;
wire n_4628;
wire n_4696;
wire n_1097;
wire n_3122;
wire n_3012;
wire n_6826;
wire n_5005;
wire n_5004;
wire n_7768;
wire n_3368;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_7235;
wire n_4597;
wire n_1812;
wire n_5090;
wire n_4574;
wire n_7129;
wire n_4242;
wire n_7243;
wire n_4949;
wire n_4748;
wire n_4959;
wire n_1747;
wire n_7342;
wire n_3400;
wire n_2508;
wire n_4243;
wire n_2540;
wire n_7547;
wire n_3820;
wire n_5395;
wire n_6494;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_2316;
wire n_5489;
wire n_5649;
wire n_7581;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_7310;
wire n_2911;
wire n_1828;
wire n_6972;
wire n_1389;
wire n_6380;
wire n_7200;
wire n_7751;
wire n_5791;
wire n_1798;
wire n_5559;
wire n_6703;
wire n_7116;
wire n_4562;
wire n_1584;
wire n_7540;
wire n_7720;
wire n_5009;
wire n_6034;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_6719;
wire n_6526;
wire n_4986;
wire n_4453;
wire n_1366;
wire n_7208;
wire n_1187;
wire n_3173;
wire n_6212;
wire n_4281;
wire n_4332;
wire n_7337;
wire n_3433;
wire n_3998;
wire n_1686;
wire n_4464;
wire n_3017;
wire n_4605;
wire n_4737;
wire n_6111;
wire n_2542;
wire n_2843;
wire n_3305;
wire n_1635;
wire n_7055;
wire n_5295;
wire n_6427;
wire n_4310;
wire n_3752;
wire n_7073;
wire n_2637;
wire n_7417;
wire n_7159;
wire n_5047;
wire n_5504;
wire n_7494;
wire n_5076;
wire n_3543;
wire n_5693;
wire n_3655;
wire n_7314;
wire n_3791;
wire n_6904;
wire n_6778;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_7294;
wire n_6520;
wire n_4906;
wire n_4257;
wire n_7016;
wire n_5712;
wire n_4516;
wire n_2913;
wire n_5028;
wire n_1381;
wire n_2254;
wire n_1597;
wire n_1486;
wire n_6444;
wire n_7422;
wire n_5622;
wire n_4196;
wire n_5255;
wire n_2371;
wire n_6362;
wire n_3898;
wire n_6749;
wire n_3366;
wire n_3453;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_6648;
wire n_2408;
wire n_6985;
wire n_4961;
wire n_6330;
wire n_5013;
wire n_2140;
wire n_6622;
wire n_2134;
wire n_2483;
wire n_2466;
wire n_3661;
wire n_5348;
wire n_6405;
wire n_2048;
wire n_2760;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_4964;
wire n_5251;
wire n_5036;
wire n_3665;
wire n_2079;
wire n_4807;
wire n_4886;
wire n_6488;
wire n_4342;
wire n_5554;
wire n_2671;
wire n_3296;
wire n_5919;
wire n_5978;
wire n_6220;
wire n_1390;
wire n_2775;
wire n_7178;
wire n_7330;
wire n_3223;
wire n_2005;
wire n_7764;
wire n_1116;
wire n_7704;
wire n_2811;
wire n_1758;
wire n_7388;
wire n_2848;
wire n_6087;
wire n_1784;
wire n_3200;
wire n_1213;
wire n_3483;
wire n_5702;
wire n_3207;
wire n_5450;
wire n_7697;
wire n_5806;
wire n_1180;
wire n_4657;
wire n_3869;
wire n_3852;
wire n_1220;
wire n_5071;
wire n_5308;
wire n_5982;
wire n_6692;
wire n_7079;
wire n_6590;
wire n_7536;
wire n_3036;
wire n_7209;
wire n_5012;
wire n_5376;
wire n_6501;
wire n_5778;
wire n_4207;
wire n_1760;
wire n_5208;
wire n_6396;
wire n_2173;
wire n_2824;
wire n_7467;
wire n_4038;
wire n_5503;
wire n_7206;
wire n_4793;
wire n_4472;
wire n_2588;
wire n_6702;
wire n_3046;
wire n_7505;
wire n_6551;
wire n_1142;
wire n_1385;
wire n_4395;
wire n_4274;
wire n_5644;
wire n_7501;
wire n_6368;
wire n_2533;
wire n_1500;
wire n_2706;
wire n_1868;
wire n_2303;
wire n_7490;
wire n_4532;
wire n_5235;
wire n_5062;
wire n_6309;
wire n_3332;
wire n_5161;
wire n_4413;
wire n_4743;
wire n_2403;
wire n_5016;
wire n_2702;
wire n_3922;
wire n_7051;
wire n_7278;
wire n_2791;
wire n_1450;
wire n_7416;
wire n_2092;
wire n_6248;
wire n_5996;
wire n_3189;
wire n_7611;
wire n_2797;
wire n_7600;
wire n_1089;
wire n_4275;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_7447;
wire n_2996;
wire n_2836;
wire n_1404;
wire n_3582;
wire n_4830;
wire n_7520;
wire n_4442;
wire n_7702;
wire n_5700;
wire n_7274;
wire n_2168;
wire n_1442;
wire n_7668;
wire n_4689;
wire n_2886;
wire n_5699;
wire n_6287;
wire n_6022;
wire n_1968;
wire n_6579;
wire n_6820;
wire n_4018;
wire n_2609;
wire n_6633;
wire n_4613;
wire n_5940;
wire n_6614;
wire n_1483;
wire n_1703;
wire n_7591;
wire n_1953;
wire n_3715;
wire n_6952;
wire n_7617;
wire n_3261;
wire n_5324;
wire n_7534;
wire n_6547;
wire n_7065;
wire n_5421;
wire n_3861;
wire n_5175;
wire n_3161;
wire n_3313;
wire n_1807;
wire n_1310;
wire n_3198;
wire n_5820;
wire n_3463;
wire n_2559;
wire n_6589;
wire n_6995;
wire n_4188;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_5340;
wire n_3738;
wire n_1640;
wire n_5694;
wire n_5022;
wire n_7461;
wire n_1145;
wire n_2307;
wire n_3546;
wire n_1511;
wire n_1651;
wire n_6297;
wire n_5245;
wire n_7326;
wire n_5651;
wire n_3944;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1696;
wire n_6367;
wire n_7761;
wire n_6198;
wire n_1355;
wire n_5364;
wire n_5459;
wire n_4534;
wire n_3635;
wire n_7423;
wire n_3270;
wire n_5168;
wire n_7443;
wire n_4590;
wire n_4602;
wire n_5510;
wire n_5329;
wire n_7746;
wire n_6251;
wire n_1335;
wire n_3213;
wire n_4394;
wire n_1900;
wire n_6583;
wire n_3418;
wire n_2614;
wire n_5581;
wire n_7556;
wire n_1780;
wire n_1091;
wire n_3865;
wire n_2769;
wire n_4220;
wire n_6879;
wire n_5812;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_2100;
wire n_4948;
wire n_3903;
wire n_3895;
wire n_1194;
wire n_3851;
wire n_4508;
wire n_4934;
wire n_7104;
wire n_7631;
wire n_3482;
wire n_2282;
wire n_3654;
wire n_4939;
wire n_4213;
wire n_2430;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_5711;
wire n_3268;
wire n_4703;
wire n_1655;
wire n_3494;
wire n_7106;
wire n_3615;
wire n_7693;
wire n_7198;
wire n_7656;
wire n_7381;
wire n_5970;
wire n_3363;
wire n_7731;
wire n_1186;
wire n_3180;
wire n_5570;
wire n_1743;
wire n_7182;
wire n_6310;
wire n_6852;
wire n_5061;
wire n_1506;
wire n_2594;
wire n_1474;
wire n_3150;
wire n_5550;
wire n_4773;
wire n_3853;
wire n_6961;
wire n_2512;
wire n_4449;
wire n_5219;
wire n_6618;
wire n_7670;
wire n_2607;
wire n_4615;
wire n_3911;
wire n_7126;
wire n_5132;
wire n_4883;
wire n_1079;
wire n_6249;
wire n_3559;
wire n_6956;
wire n_5184;
wire n_6440;
wire n_7564;
wire n_5747;
wire n_6575;
wire n_4943;
wire n_5821;
wire n_2498;
wire n_7524;
wire n_4630;
wire n_3812;
wire n_6584;
wire n_6689;
wire n_2017;
wire n_1227;
wire n_5326;
wire n_3750;
wire n_5909;
wire n_6050;
wire n_3838;
wire n_5868;
wire n_1954;
wire n_4749;
wire n_1125;
wire n_6643;
wire n_2687;
wire n_3456;
wire n_6569;
wire n_6814;
wire n_3132;
wire n_5618;
wire n_6596;
wire n_7176;
wire n_4159;
wire n_7056;
wire n_4372;
wire n_5528;
wire n_4731;
wire n_4004;
wire n_1134;
wire n_1684;
wire n_7594;
wire n_4353;
wire n_5593;
wire n_3334;
wire n_3819;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_5740;
wire n_1233;
wire n_5108;
wire n_3653;
wire n_4360;
wire n_6123;
wire n_4897;
wire n_2139;
wire n_3693;
wire n_5477;
wire n_5934;
wire n_5218;
wire n_1138;
wire n_2943;
wire n_5272;
wire n_1096;
wire n_7535;
wire n_3135;
wire n_4239;
wire n_3175;
wire n_6273;
wire n_7368;
wire n_5464;
wire n_6895;
wire n_6548;
wire n_7627;
wire n_6420;
wire n_6474;
wire n_1268;
wire n_3187;
wire n_3830;
wire n_2724;
wire n_6890;
wire n_5688;
wire n_6141;
wire n_1829;
wire n_1338;
wire n_6234;
wire n_1327;
wire n_5204;
wire n_6789;
wire n_5400;
wire n_3407;
wire n_3315;
wire n_4470;
wire n_4690;
wire n_3982;
wire n_6311;
wire n_6867;
wire n_2565;
wire n_4201;
wire n_6634;
wire n_6288;
wire n_1636;
wire n_1687;
wire n_5303;
wire n_4584;
wire n_3184;
wire n_6290;
wire n_5804;
wire n_6764;
wire n_4155;
wire n_3890;
wire n_5519;
wire n_5023;
wire n_2032;
wire n_3392;
wire n_4802;
wire n_6935;
wire n_1258;
wire n_2208;
wire n_1344;
wire n_5971;
wire n_2198;
wire n_1929;
wire n_5095;
wire n_1680;
wire n_1195;
wire n_5902;
wire n_4304;
wire n_4975;
wire n_4821;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_4910;
wire n_5064;
wire n_6478;
wire n_7382;
wire n_3641;
wire n_5203;
wire n_5065;
wire n_4887;
wire n_5436;
wire n_7579;
wire n_3996;
wire n_7130;
wire n_6942;
wire n_6056;
wire n_7647;
wire n_2873;
wire n_1576;
wire n_6772;
wire n_6466;
wire n_3049;
wire n_4015;
wire n_4211;
wire n_4119;
wire n_3620;
wire n_2558;
wire n_2347;
wire n_3884;
wire n_3103;
wire n_3770;
wire n_4591;
wire n_2527;
wire n_5314;
wire n_7469;
wire n_5044;
wire n_1509;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_6228;
wire n_1841;
wire n_6955;
wire n_5886;
wire n_2685;
wire n_5344;
wire n_1313;
wire n_4223;
wire n_2090;
wire n_5173;
wire n_5585;
wire n_3722;
wire n_5981;
wire n_3802;
wire n_5343;
wire n_5783;
wire n_2215;
wire n_1449;
wire n_1723;
wire n_3129;
wire n_5515;
wire n_4806;
wire n_2116;
wire n_5784;
wire n_5337;
wire n_3592;
wire n_5545;
wire n_1645;
wire n_3186;
wire n_6393;
wire n_7654;
wire n_6375;
wire n_7762;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_5209;
wire n_1269;
wire n_2773;
wire n_2906;
wire n_3097;
wire n_5495;
wire n_7427;
wire n_6908;
wire n_3910;
wire n_4238;
wire n_1466;
wire n_3667;
wire n_6424;
wire n_7506;
wire n_3822;
wire n_1276;
wire n_6874;
wire n_1637;
wire n_2900;
wire n_5799;
wire n_6296;
wire n_3765;
wire n_2216;
wire n_5888;
wire n_6736;
wire n_4259;
wire n_1620;
wire n_7376;
wire n_5196;
wire n_5086;
wire n_7018;
wire n_6025;
wire n_6168;
wire n_7498;
wire n_3518;
wire n_5885;
wire n_2022;
wire n_7134;
wire n_3967;
wire n_2373;
wire n_7456;
wire n_1853;
wire n_2275;
wire n_5398;
wire n_5434;
wire n_5797;
wire n_2899;
wire n_5830;
wire n_5896;
wire n_3351;
wire n_7480;
wire n_2008;
wire n_5052;
wire n_2859;
wire n_5952;
wire n_6003;
wire n_2564;
wire n_5110;
wire n_7348;
wire n_5918;
wire n_4799;
wire n_1356;
wire n_2591;
wire n_3965;
wire n_1969;
wire n_5808;
wire n_6119;
wire n_1296;
wire n_4444;
wire n_4676;
wire n_5212;
wire n_6525;
wire n_1764;
wire n_7383;
wire n_1250;
wire n_1190;
wire n_5733;
wire n_4598;
wire n_3259;
wire n_7053;
wire n_7660;
wire n_5483;
wire n_6713;
wire n_6919;
wire n_4533;
wire n_4078;
wire n_1794;
wire n_7557;
wire n_3779;
wire n_3203;
wire n_7240;
wire n_7468;
wire n_3923;
wire n_4392;
wire n_3808;
wire n_6750;
wire n_4455;
wire n_3093;
wire n_2664;
wire n_1434;
wire n_4129;
wire n_5278;
wire n_2114;
wire n_6204;
wire n_1609;
wire n_5522;
wire n_3530;
wire n_6981;
wire n_1132;
wire n_5584;
wire n_4548;
wire n_6675;
wire n_1803;
wire n_5264;
wire n_6321;
wire n_1281;
wire n_4535;
wire n_1447;
wire n_2150;
wire n_6337;
wire n_4999;
wire n_5328;
wire n_7604;
wire n_2660;
wire n_5447;
wire n_5029;
wire n_5127;
wire n_5006;
wire n_5679;
wire n_4604;
wire n_7585;
wire n_6828;
wire n_5123;
wire n_6160;
wire n_7043;
wire n_3467;
wire n_6156;
wire n_4240;
wire n_7074;
wire n_7119;
wire n_7596;
wire n_2219;
wire n_6116;
wire n_4522;
wire n_1387;
wire n_3371;
wire n_4713;
wire n_1368;
wire n_1154;
wire n_6267;
wire n_2539;
wire n_6875;
wire n_1701;
wire n_5236;
wire n_7567;
wire n_6678;
wire n_5239;
wire n_5307;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_3317;
wire n_3963;
wire n_6870;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_6561;
wire n_6715;
wire n_2529;
wire n_4103;
wire n_4126;
wire n_4710;
wire n_5576;
wire n_3282;
wire n_5144;
wire n_2708;
wire n_5164;
wire n_6557;
wire n_2748;
wire n_5359;
wire n_7386;
wire n_6503;
wire n_5925;
wire n_2224;
wire n_5526;
wire n_5810;
wire n_2233;
wire n_2499;
wire n_6333;
wire n_5172;
wire n_3888;
wire n_4549;
wire n_3309;
wire n_5126;
wire n_1924;
wire n_3024;
wire n_7701;
wire n_4767;
wire n_7007;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_7027;
wire n_5999;
wire n_5147;
wire n_7616;
wire n_5407;
wire n_7432;
wire n_1553;
wire n_3542;
wire n_5536;
wire n_1090;
wire n_6002;
wire n_3374;
wire n_3704;
wire n_7661;
wire n_2786;
wire n_1905;
wire n_4355;
wire n_2958;
wire n_7009;
wire n_6140;
wire n_5903;
wire n_7263;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_4834;
wire n_6336;
wire n_3660;
wire n_2718;
wire n_4712;
wire n_5849;
wire n_7772;
wire n_6663;
wire n_1795;
wire n_7610;
wire n_3634;
wire n_4096;
wire n_6844;
wire n_2101;
wire n_5378;
wire n_1152;
wire n_3626;
wire n_2599;
wire n_6999;
wire n_4571;
wire n_7214;
wire n_6982;
wire n_5389;
wire n_6166;
wire n_3171;
wire n_6170;
wire n_1733;
wire n_6257;
wire n_7613;
wire n_3986;
wire n_2853;
wire n_1552;
wire n_6620;
wire n_4930;
wire n_5345;
wire n_2217;
wire n_3594;
wire n_2866;
wire n_5138;
wire n_3153;
wire n_6202;
wire n_1189;
wire n_4995;
wire n_6529;
wire n_4039;
wire n_4253;
wire n_4681;
wire n_2623;
wire n_6843;
wire n_3232;
wire n_5228;
wire n_2178;
wire n_1181;
wire n_3815;
wire n_4375;
wire n_5629;
wire n_5945;
wire n_4205;
wire n_6161;
wire n_3790;
wire n_6147;
wire n_2404;
wire n_5601;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_6554;
wire n_3640;
wire n_6877;
wire n_2821;
wire n_6892;
wire n_4768;
wire n_6133;
wire n_6109;
wire n_6585;
wire n_5985;
wire n_7162;
wire n_5435;
wire n_5665;
wire n_3299;
wire n_4070;
wire n_4558;
wire n_6436;
wire n_3065;
wire n_2375;
wire n_2572;
wire n_1656;
wire n_2063;
wire n_3082;
wire n_5709;
wire n_4504;
wire n_5176;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_4864;
wire n_3855;
wire n_3357;
wire n_4485;
wire n_1510;
wire n_5003;
wire n_2852;
wire n_2132;
wire n_5567;
wire n_1236;
wire n_3412;
wire n_5765;
wire n_1712;
wire n_6409;
wire n_4537;
wire n_5771;
wire n_5271;
wire n_1184;
wire n_2585;
wire n_7510;
wire n_2220;
wire n_4005;
wire n_1364;
wire n_3183;
wire n_4323;
wire n_5068;
wire n_4184;
wire n_2468;
wire n_5078;
wire n_7268;
wire n_3248;
wire n_2606;
wire n_5980;
wire n_7465;
wire n_4337;
wire n_4826;
wire n_7398;
wire n_2152;
wire n_5073;
wire n_5420;
wire n_6386;
wire n_5599;
wire n_4952;
wire n_3785;
wire n_3525;
wire n_5508;
wire n_2779;
wire n_1117;
wire n_2547;
wire n_6473;
wire n_1748;
wire n_7304;
wire n_7036;
wire n_2935;
wire n_5084;
wire n_6651;
wire n_7462;
wire n_2490;
wire n_3127;
wire n_7171;
wire n_3496;
wire n_3568;
wire n_5789;
wire n_4876;
wire n_5322;
wire n_6490;
wire n_3841;
wire n_4626;
wire n_1334;
wire n_7678;
wire n_7597;
wire n_3879;
wire n_6558;
wire n_2402;
wire n_1200;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_6500;
wire n_5590;
wire n_5638;
wire n_4747;
wire n_5152;
wire n_3341;
wire n_4347;
wire n_1852;
wire n_3868;
wire n_4791;
wire n_5497;
wire n_2481;
wire n_4409;
wire n_5361;
wire n_7293;
wire n_1264;
wire n_6752;
wire n_2808;
wire n_5010;
wire n_6363;
wire n_3396;
wire n_6007;
wire n_2102;
wire n_7568;
wire n_3492;
wire n_3558;
wire n_2751;
wire n_1548;
wire n_4824;
wire n_5117;
wire n_2977;
wire n_1682;
wire n_6142;
wire n_3599;
wire n_7363;
wire n_6244;
wire n_1896;
wire n_1704;
wire n_2234;
wire n_6369;
wire n_6518;
wire n_5050;
wire n_5608;
wire n_5610;
wire n_4152;
wire n_6698;
wire n_1352;
wire n_5125;
wire n_2328;
wire n_6977;
wire n_6578;
wire n_4587;
wire n_6118;
wire n_6429;
wire n_6158;
wire n_2332;
wire n_7511;
wire n_7028;
wire n_1628;
wire n_6810;
wire n_1773;
wire n_7237;
wire n_3580;
wire n_2369;
wire n_5474;
wire n_3584;
wire n_4500;
wire n_5845;
wire n_1115;
wire n_1395;
wire n_7039;
wire n_4660;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_6049;
wire n_2419;
wire n_6671;
wire n_6791;
wire n_5794;
wire n_5299;
wire n_2807;
wire n_4047;
wire n_5905;
wire n_4157;
wire n_3956;
wire n_1431;
wire n_5202;
wire n_6967;
wire n_5170;
wire n_5724;
wire n_6610;
wire n_7442;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_6108;
wire n_2241;
wire n_7618;
wire n_6768;
wire n_2458;
wire n_7489;
wire n_7144;
wire n_3401;
wire n_3032;
wire n_7362;
wire n_5042;
wire n_1750;
wire n_2833;
wire n_3179;
wire n_6382;
wire n_5662;
wire n_1563;
wire n_4051;
wire n_3123;
wire n_6576;
wire n_1875;
wire n_6947;
wire n_1615;
wire n_3719;
wire n_5334;
wire n_5595;
wire n_6938;
wire n_7765;
wire n_6260;
wire n_5244;
wire n_7453;
wire n_2635;
wire n_4077;
wire n_3897;
wire n_3475;
wire n_2077;
wire n_2520;
wire n_2193;
wire n_4010;
wire n_4942;
wire n_4255;
wire n_5692;
wire n_2908;
wire n_4561;
wire n_6906;
wire n_4957;
wire n_2053;
wire n_1580;
wire n_5728;
wire n_7758;
wire n_2200;
wire n_2304;
wire n_4683;
wire n_6148;
wire n_6404;
wire n_1439;
wire n_2352;
wire n_4839;
wire n_2185;
wire n_7124;
wire n_2476;
wire n_1266;
wire n_4814;
wire n_2781;
wire n_6217;
wire n_6324;
wire n_6918;
wire n_2460;
wire n_4694;
wire n_3600;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_2308;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_4026;
wire n_7143;
wire n_2903;
wire n_3659;
wire n_5795;
wire n_4496;
wire n_6048;
wire n_1528;
wire n_3840;
wire n_5889;
wire n_5856;
wire n_7606;
wire n_3481;
wire n_4719;
wire n_4100;
wire n_3517;
wire n_5722;
wire n_1413;
wire n_2464;
wire n_6834;
wire n_5498;
wire n_2925;
wire n_2270;
wire n_5034;
wire n_5725;
wire n_6812;
wire n_1706;
wire n_1592;
wire n_6110;
wire n_1461;
wire n_2695;
wire n_6300;
wire n_5657;
wire n_3656;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_5282;
wire n_5511;
wire n_7123;
wire n_2414;
wire n_5736;
wire n_5642;
wire n_6624;
wire n_3316;
wire n_2465;
wire n_3925;
wire n_4089;
wire n_1683;
wire n_7072;
wire n_4175;
wire n_4458;
wire n_7488;
wire n_6001;
wire n_3955;
wire n_3158;
wire n_3657;
wire n_5776;
wire n_5826;
wire n_6687;
wire n_2684;
wire n_1104;
wire n_2205;
wire n_3284;
wire n_2875;
wire n_1437;
wire n_2747;
wire n_5932;
wire n_4185;
wire n_2064;
wire n_3088;
wire n_1497;
wire n_2002;
wire n_7734;
wire n_6088;
wire n_6762;
wire n_4815;
wire n_2545;
wire n_2050;
wire n_3695;
wire n_6239;
wire n_2500;
wire n_6992;
wire n_7109;
wire n_1917;
wire n_1444;
wire n_6091;
wire n_4316;
wire n_5453;
wire n_3328;
wire n_2763;
wire n_7644;
wire n_5136;
wire n_6352;
wire n_2761;
wire n_4020;
wire n_5494;
wire n_6101;
wire n_1920;
wire n_4306;
wire n_6319;
wire n_2997;
wire n_3735;
wire n_2127;
wire n_6188;
wire n_5718;
wire n_5634;
wire n_3228;
wire n_3028;
wire n_5079;
wire n_3706;
wire n_6395;
wire n_1432;
wire n_3322;
wire n_7325;
wire n_1174;
wire n_6037;
wire n_4512;
wire n_4483;
wire n_3499;
wire n_3552;
wire n_4164;
wire n_1286;
wire n_6759;
wire n_3784;
wire n_4142;
wire n_6206;
wire n_7137;
wire n_4621;
wire n_7526;
wire n_3016;
wire n_7699;
wire n_1629;
wire n_5706;
wire n_7350;
wire n_2694;
wire n_6177;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1850;
wire n_1670;
wire n_4123;
wire n_7311;
wire n_7458;
wire n_2317;
wire n_1384;
wire n_1612;
wire n_5496;
wire n_1099;
wire n_3113;
wire n_4305;
wire n_2909;
wire n_3960;
wire n_4007;
wire n_7244;
wire n_1524;
wire n_7681;
wire n_4707;
wire n_4429;
wire n_1991;
wire n_2566;
wire n_7339;
wire n_2210;
wire n_5606;
wire n_6322;
wire n_1225;
wire n_7247;
wire n_2346;
wire n_4695;
wire n_7331;
wire n_7128;
wire n_2180;
wire n_3376;
wire n_6313;
wire n_5989;
wire n_2617;
wire n_5870;
wire n_7284;
wire n_4163;
wire n_7321;
wire n_2831;
wire n_6504;
wire n_2865;
wire n_1625;
wire n_4638;
wire n_5530;
wire n_4498;
wire n_2240;
wire n_7309;
wire n_1797;
wire n_4750;
wire n_3993;
wire n_7163;
wire n_2120;
wire n_1289;
wire n_1557;
wire n_1567;
wire n_2007;
wire n_2004;
wire n_5424;
wire n_5230;
wire n_2086;
wire n_6886;
wire n_4832;
wire n_5229;
wire n_7054;
wire n_3666;
wire n_6374;
wire n_1839;
wire n_5160;
wire n_2330;
wire n_2555;
wire n_1587;
wire n_6356;
wire n_6640;
wire n_5313;
wire n_2108;
wire n_6462;
wire n_5333;
wire n_5207;
wire n_2535;
wire n_6959;
wire n_5158;
wire n_2945;
wire n_5154;
wire n_3057;
wire n_7413;
wire n_4319;
wire n_3760;
wire n_5721;
wire n_7185;
wire n_1396;
wire n_1923;
wire n_1224;
wire n_5654;
wire n_2196;
wire n_5860;
wire n_1538;
wire n_3773;
wire n_6710;
wire n_5884;
wire n_2604;
wire n_3462;
wire n_4373;
wire n_6945;
wire n_2351;
wire n_2437;
wire n_1889;
wire n_6776;
wire n_1124;
wire n_5839;
wire n_2688;
wire n_4990;
wire n_7336;
wire n_3302;
wire n_1673;
wire n_5058;
wire n_2085;
wire n_3304;
wire n_1725;
wire n_6231;
wire n_2149;
wire n_7630;
wire n_2001;
wire n_1800;
wire n_3746;
wire n_6905;
wire n_7737;
wire n_7120;
wire n_3645;
wire n_5823;
wire n_4262;
wire n_4019;
wire n_2735;
wire n_6401;
wire n_2035;
wire n_4436;
wire n_4697;
wire n_1906;
wire n_1647;
wire n_4357;
wire n_7374;
wire n_6521;
wire n_4849;
wire n_5101;
wire n_5532;
wire n_4366;
wire n_6582;
wire n_7491;
wire n_6964;
wire n_4139;
wire n_1270;
wire n_5297;
wire n_4340;
wire n_1476;
wire n_7001;
wire n_2027;
wire n_5611;
wire n_2012;
wire n_3512;
wire n_4720;
wire n_3892;
wire n_7111;
wire n_6623;
wire n_1880;
wire n_6225;
wire n_7519;
wire n_1642;
wire n_5744;
wire n_6798;
wire n_2447;
wire n_3358;
wire n_5538;
wire n_2894;
wire n_5249;
wire n_5669;
wire n_2587;
wire n_1605;
wire n_6134;
wire n_2099;
wire n_1202;
wire n_5793;
wire n_3410;
wire n_4900;
wire n_6493;
wire n_6364;
wire n_5715;
wire n_6665;
wire n_7538;
wire n_3408;
wire n_3182;
wire n_1879;
wire n_4941;
wire n_1311;
wire n_5966;
wire n_2299;
wire n_2078;
wire n_6284;
wire n_3709;
wire n_3011;
wire n_5383;
wire n_6649;
wire n_5775;
wire n_2315;
wire n_3623;
wire n_6230;
wire n_5558;
wire n_7165;
wire n_2157;
wire n_6546;
wire n_3446;
wire n_5547;
wire n_5572;
wire n_5659;
wire n_5223;
wire n_6555;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_6010;
wire n_3058;
wire n_4334;
wire n_6331;
wire n_6888;
wire n_2211;
wire n_6047;
wire n_5708;
wire n_7599;
wire n_6532;
wire n_5817;
wire n_3384;
wire n_4698;
wire n_6677;
wire n_2225;
wire n_1411;
wire n_5867;
wire n_7389;
wire n_1501;
wire n_7418;
wire n_5636;
wire n_5106;
wire n_5800;
wire n_7375;
wire n_7671;
wire n_7096;
wire n_5257;
wire n_7719;
wire n_7281;
wire n_7300;
wire n_4397;
wire n_6920;
wire n_3611;
wire n_4186;
wire n_2093;
wire n_2675;
wire n_5371;
wire n_6524;
wire n_6781;
wire n_4229;
wire n_4294;
wire n_7085;
wire n_1919;
wire n_4351;
wire n_6811;
wire n_6226;
wire n_2893;
wire n_6281;
wire n_2009;
wire n_6514;
wire n_5731;
wire n_4162;
wire n_1416;
wire n_3465;
wire n_7683;
wire n_1515;
wire n_6921;
wire n_4127;
wire n_4620;
wire n_1314;
wire n_3059;
wire n_3085;
wire n_2867;
wire n_2229;
wire n_4770;
wire n_7212;
wire n_7285;
wire n_7676;
wire n_3871;
wire n_2388;
wire n_6685;
wire n_7590;
wire n_3112;
wire n_5623;
wire n_5921;
wire n_6082;
wire n_3413;
wire n_4580;
wire n_7032;
wire n_2624;
wire n_1813;
wire n_4581;
wire n_4618;
wire n_7125;
wire n_5178;
wire n_6609;
wire n_5853;
wire n_7160;
wire n_7100;
wire n_1105;
wire n_5898;
wire n_5198;
wire n_2898;
wire n_5437;
wire n_6627;
wire n_2519;
wire n_2231;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_5053;
wire n_1256;
wire n_4670;
wire n_7319;
wire n_6162;
wire n_7638;
wire n_5592;
wire n_5484;
wire n_6650;
wire n_4982;
wire n_5418;
wire n_6079;
wire n_6013;
wire n_5432;
wire n_1769;
wire n_7635;
wire n_5270;
wire n_1372;
wire n_1847;
wire n_5166;
wire n_5358;
wire n_3805;
wire n_2406;
wire n_4017;
wire n_7504;
wire n_1586;
wire n_3497;
wire n_6722;
wire n_5156;
wire n_6592;
wire n_3382;
wire n_4236;
wire n_4313;
wire n_5548;
wire n_5687;
wire n_3561;
wire n_2543;
wire n_6512;
wire n_2992;
wire n_1541;
wire n_6008;
wire n_6522;
wire n_4907;
wire n_4659;
wire n_2128;
wire n_1697;
wire n_1872;
wire n_5822;
wire n_2690;
wire n_3942;
wire n_2020;
wire n_5758;
wire n_1939;
wire n_7767;
wire n_5366;
wire n_4053;
wire n_5392;
wire n_4279;
wire n_3937;
wire n_6400;
wire n_7371;
wire n_3303;
wire n_5115;
wire n_5046;
wire n_7361;
wire n_5139;
wire n_4555;
wire n_5829;
wire n_5686;
wire n_7440;
wire n_5735;
wire n_3549;
wire n_1481;
wire n_6613;
wire n_1928;
wire n_4235;
wire n_3972;
wire n_5674;
wire n_2314;
wire n_2126;
wire n_3403;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_1361;
wire n_5039;
wire n_6538;
wire n_1693;
wire n_2081;
wire n_5341;
wire n_2993;
wire n_7010;
wire n_5032;
wire n_3018;
wire n_4820;
wire n_2449;
wire n_2131;
wire n_7289;
wire n_2526;
wire n_4794;
wire n_1302;
wire n_5041;
wire n_6505;
wire n_3989;
wire n_6581;
wire n_5565;
wire n_7021;
wire n_7004;
wire n_6350;
wire n_4752;
wire n_4546;
wire n_7234;
wire n_3918;
wire n_6378;
wire n_3191;
wire n_3051;
wire n_6975;
wire n_7266;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_4415;
wire n_2487;
wire n_3343;
wire n_3163;
wire n_6243;
wire n_3786;
wire n_4061;
wire n_4432;
wire n_6484;
wire n_1912;
wire n_4552;
wire n_3143;
wire n_1876;
wire n_7754;
wire n_6573;
wire n_6786;
wire n_6774;
wire n_6419;
wire n_4790;
wire n_1811;
wire n_1285;
wire n_5448;
wire n_4263;
wire n_3725;
wire n_5974;
wire n_5852;
wire n_6143;
wire n_6851;
wire n_1529;
wire n_1824;
wire n_3522;
wire n_4528;
wire n_4888;
wire n_4502;
wire n_5085;
wire n_7211;
wire n_4335;
wire n_7141;
wire n_3444;
wire n_4218;
wire n_4705;
wire n_6112;
wire n_6138;
wire n_3009;
wire n_4471;
wire n_1141;
wire n_3297;
wire n_6729;
wire n_7150;
wire n_6882;
wire n_1168;
wire n_5500;
wire n_7378;
wire n_6045;
wire n_5293;
wire n_6203;
wire n_7470;
wire n_3000;
wire n_2305;
wire n_1192;
wire n_1290;
wire n_2514;
wire n_4386;
wire n_6568;
wire n_4547;
wire n_7633;
wire n_4836;
wire n_5458;
wire n_3545;
wire n_1101;
wire n_4193;
wire n_5670;
wire n_7420;
wire n_1336;
wire n_6433;
wire n_6023;
wire n_1358;
wire n_3318;
wire n_5684;
wire n_1397;
wire n_1359;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_4984;
wire n_1532;
wire n_5624;
wire n_3430;
wire n_1685;
wire n_7558;
wire n_5325;
wire n_2801;
wire n_3225;
wire n_3067;
wire n_6189;
wire n_6167;
wire n_5059;
wire n_1462;
wire n_5825;
wire n_3823;
wire n_4718;
wire n_3185;
wire n_2326;
wire n_5586;
wire n_6998;
wire n_1398;
wire n_5222;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_4634;
wire n_6335;
wire n_5741;
wire n_1692;
wire n_5875;
wire n_6721;
wire n_4796;
wire n_6312;
wire n_4560;
wire n_1240;
wire n_3285;
wire n_5045;
wire n_7640;
wire n_1814;
wire n_4882;
wire n_1808;
wire n_2768;
wire n_1658;
wire n_6611;
wire n_7484;
wire n_5038;
wire n_5769;
wire n_3837;
wire n_7708;
wire n_4841;
wire n_6213;
wire n_3076;
wire n_6264;
wire n_4954;
wire n_4635;
wire n_4521;
wire n_5703;
wire n_3893;
wire n_4272;
wire n_2148;
wire n_2104;
wire n_2653;
wire n_2855;
wire n_6301;
wire n_2618;
wire n_7598;
wire n_4448;
wire n_3359;
wire n_5501;
wire n_6216;
wire n_2331;
wire n_1600;
wire n_7271;
wire n_5894;
wire n_4701;
wire n_5248;
wire n_5872;
wire n_4088;
wire n_2136;
wire n_7322;
wire n_7549;
wire n_7022;
wire n_5443;
wire n_6193;
wire n_1913;
wire n_6885;
wire n_7217;
wire n_7166;
wire n_3056;
wire n_4208;
wire n_5363;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_6806;
wire n_4865;
wire n_2066;
wire n_7584;
wire n_1974;
wire n_1158;
wire n_6588;
wire n_4589;
wire n_3924;
wire n_6933;
wire n_1915;
wire n_2534;
wire n_5908;
wire n_4972;
wire n_5597;
wire n_4617;
wire n_3311;
wire n_1160;
wire n_4094;
wire n_4772;
wire n_4857;
wire n_7297;
wire n_7664;
wire n_3613;
wire n_1383;
wire n_7546;
wire n_2057;
wire n_7179;
wire n_5984;
wire n_6385;
wire n_7415;
wire n_5533;
wire n_1822;
wire n_6051;
wire n_1804;
wire n_1581;
wire n_7057;
wire n_5387;
wire n_4776;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_2246;
wire n_2738;
wire n_6793;
wire n_1851;
wire n_1755;
wire n_5589;
wire n_6746;
wire n_4702;
wire n_1341;
wire n_7411;
wire n_4486;
wire n_4946;
wire n_2202;
wire n_5380;
wire n_2262;
wire n_5134;
wire n_1333;
wire n_4506;
wire n_7108;
wire n_7736;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_4153;
wire n_7220;
wire n_6015;
wire n_4329;
wire n_6435;
wire n_4877;
wire n_3442;
wire n_2327;
wire n_4780;
wire n_6411;
wire n_4327;
wire n_5954;
wire n_5412;
wire n_2656;
wire n_6323;
wire n_4168;
wire n_2258;
wire n_4396;
wire n_2039;
wire n_5174;
wire n_4465;
wire n_6174;
wire n_7223;
wire n_2544;
wire n_7261;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_3266;
wire n_7092;
wire n_5468;
wire n_1843;
wire n_2030;
wire n_4576;
wire n_6728;
wire n_4075;
wire n_5429;
wire n_3593;
wire n_6586;
wire n_2536;
wire n_1399;
wire n_3685;
wire n_5269;
wire n_4833;
wire n_1903;
wire n_1849;
wire n_7275;
wire n_3768;
wire n_4224;
wire n_7272;
wire n_4868;
wire n_5124;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_7436;
wire n_3181;
wire n_7249;
wire n_3644;
wire n_5287;
wire n_4387;
wire n_5865;
wire n_2368;
wire n_6437;
wire n_4896;
wire n_1157;
wire n_7168;
wire n_2065;
wire n_2901;
wire n_5583;
wire n_3818;
wire n_4368;
wire n_1295;
wire n_1983;
wire n_4798;
wire n_2201;
wire n_1582;
wire n_7712;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_5416;
wire n_7743;
wire n_2569;
wire n_7705;
wire n_1998;
wire n_1596;
wire n_3077;
wire n_7091;
wire n_1100;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_2123;
wire n_4364;
wire n_3019;
wire n_2235;
wire n_5373;
wire n_4967;
wire n_6067;
wire n_6858;
wire n_7679;
wire n_1080;
wire n_5377;
wire n_2290;
wire n_6479;
wire n_7228;
wire n_3272;
wire n_7353;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_5350;
wire n_6279;
wire n_6841;
wire n_4668;
wire n_7696;
wire n_2383;
wire n_5632;
wire n_2640;
wire n_7687;
wire n_1492;
wire n_6425;
wire n_1478;
wire n_6896;
wire n_1796;
wire n_3569;
wire n_2374;
wire n_1614;
wire n_4648;
wire n_2598;
wire n_1722;
wire n_5290;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_4785;
wire n_5120;
wire n_2230;
wire n_5535;
wire n_3033;
wire n_2151;
wire n_5382;
wire n_6354;
wire n_4912;
wire n_6320;
wire n_1971;
wire n_5759;
wire n_2479;
wire n_4914;
wire n_6954;
wire n_2359;
wire n_2360;
wire n_4902;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_6612;
wire n_6376;
wire n_2571;
wire n_7000;
wire n_5479;
wire n_6006;
wire n_5598;
wire n_7040;
wire n_6132;
wire n_7196;
wire n_2799;
wire n_7655;
wire n_4708;
wire n_4592;
wire n_1307;
wire n_5578;
wire n_2644;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_6872;
wire n_6089;
wire n_5211;
wire n_7205;
wire n_1668;
wire n_7260;
wire n_7500;
wire n_5861;
wire n_7086;
wire n_6417;
wire n_1681;
wire n_4031;
wire n_7569;
wire n_4120;
wire n_3533;
wire n_3896;
wire n_2192;
wire n_7763;
wire n_4578;
wire n_3323;
wire n_1937;
wire n_3839;
wire n_3509;
wire n_1749;
wire n_2918;
wire n_3353;
wire n_5092;
wire n_1945;
wire n_5182;
wire n_5430;
wire n_2638;
wire n_3939;
wire n_7577;
wire n_4874;
wire n_1228;
wire n_7047;
wire n_7412;
wire n_4840;
wire n_7717;
wire n_2354;
wire n_5956;
wire n_6027;
wire n_6477;
wire n_4311;
wire n_5766;
wire n_6269;
wire n_1133;
wire n_1926;
wire n_2363;
wire n_2814;
wire n_5094;
wire n_6275;
wire n_3264;
wire n_3204;
wire n_6390;
wire n_2003;
wire n_3727;
wire n_2621;
wire n_2922;
wire n_6306;
wire n_3881;
wire n_1910;
wire n_5446;
wire n_1606;
wire n_5315;
wire n_3711;
wire n_7077;
wire n_2164;
wire n_7565;
wire n_1618;
wire n_3748;
wire n_4389;
wire n_3668;
wire n_3197;
wire n_1955;
wire n_4556;
wire n_2413;
wire n_3148;
wire n_4779;
wire n_6122;
wire n_1253;
wire n_1484;
wire n_2686;
wire n_4214;
wire n_4430;
wire n_3151;
wire n_3977;
wire n_3125;
wire n_2812;
wire n_4889;
wire n_4221;
wire n_1638;
wire n_6831;
wire n_6175;
wire n_5279;
wire n_6506;
wire n_6690;
wire n_4650;
wire n_6968;
wire n_6415;
wire n_2280;
wire n_7576;
wire n_4428;
wire n_4784;
wire n_2393;
wire n_4766;
wire n_7523;
wire n_3809;
wire n_1999;
wire n_3810;
wire n_5103;
wire n_5835;
wire n_4968;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_5311;
wire n_2283;
wire n_2806;
wire n_6184;
wire n_2813;
wire n_5268;
wire n_4295;
wire n_1716;
wire n_1412;
wire n_6285;
wire n_5773;
wire n_3310;
wire n_4182;
wire n_7750;
wire n_1401;
wire n_2951;
wire n_5451;
wire n_7578;
wire n_5452;
wire n_2145;
wire n_2122;
wire n_6644;
wire n_1588;
wire n_2579;
wire n_6688;
wire n_7402;
wire n_2876;
wire n_6670;
wire n_7473;
wire n_5321;
wire n_3301;
wire n_2370;
wire n_5215;
wire n_4600;
wire n_2025;
wire n_3451;
wire n_1219;
wire n_6680;
wire n_4513;
wire n_5635;
wire n_1252;
wire n_2730;
wire n_1927;
wire n_5356;
wire n_4735;
wire n_2767;
wire n_4667;
wire n_5150;
wire n_2826;
wire n_2112;
wire n_6180;
wire n_5613;
wire n_7405;
wire n_6137;
wire n_2762;
wire n_4774;
wire n_4711;
wire n_3023;
wire n_7343;
wire n_3224;
wire n_7721;
wire n_4481;
wire n_3762;
wire n_6410;
wire n_5063;
wire n_4671;
wire n_1326;
wire n_6046;
wire n_4981;
wire n_1799;
wire n_7252;
wire n_1689;
wire n_1304;
wire n_6465;
wire n_5653;
wire n_2541;
wire n_4879;
wire n_2987;
wire n_5788;
wire n_1702;
wire n_3916;
wire n_3630;
wire n_1558;
wire n_2722;
wire n_5057;
wire n_3618;
wire n_2727;
wire n_6991;
wire n_5560;
wire n_2719;
wire n_2213;
wire n_5476;
wire n_3521;
wire n_6121;
wire n_2723;
wire n_6077;
wire n_4054;
wire n_1569;
wire n_6000;
wire n_6205;
wire n_4012;
wire n_5582;
wire n_6705;
wire n_3567;
wire n_7601;
wire n_4352;
wire n_1988;
wire n_5935;
wire n_6201;
wire n_2401;
wire n_1787;
wire n_3094;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2631;
wire n_1867;
wire n_5697;
wire n_4252;
wire n_4505;
wire n_4219;
wire n_5119;
wire n_2292;
wire n_7451;
wire n_6471;
wire n_3560;
wire n_5813;
wire n_1742;
wire n_1818;
wire n_5100;
wire n_3847;
wire n_2203;
wire n_5427;
wire n_4909;
wire n_2693;
wire n_1159;
wire n_2281;
wire n_3202;
wire n_7603;
wire n_7575;
wire n_7188;
wire n_6913;
wire n_5467;
wire n_2646;
wire n_7525;
wire n_5346;
wire n_3887;
wire n_3800;
wire n_7528;
wire n_7113;
wire n_4435;
wire n_1235;
wire n_6329;
wire n_4755;
wire n_6355;
wire n_3827;
wire n_6145;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_5633;
wire n_7637;
wire n_1835;
wire n_2697;
wire n_3531;
wire n_2470;
wire n_5726;
wire n_2890;
wire n_6734;
wire n_4400;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_5415;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_5445;
wire n_6446;
wire n_4996;
wire n_4136;
wire n_5040;
wire n_7471;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_5031;
wire n_1360;
wire n_5814;
wire n_5374;
wire n_2070;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3039;
wire n_7296;
wire n_3900;
wire n_3478;
wire n_3701;
wire n_2766;
wire n_3756;
wire n_3754;
wire n_4156;
wire n_6057;
wire n_5818;
wire n_7781;
wire n_2416;
wire n_2962;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_6221;
wire n_5876;
wire n_5529;
wire n_3006;
wire n_3348;
wire n_4758;
wire n_2236;
wire n_5317;
wire n_3957;
wire n_2377;
wire n_2577;
wire n_3165;
wire n_4419;
wire n_2795;
wire n_7741;
wire n_5490;
wire n_3520;
wire n_2632;
wire n_4406;
wire n_7727;
wire n_6825;
wire n_5897;
wire n_5331;
wire n_6107;
wire n_6743;
wire n_1106;
wire n_4655;
wire n_6080;
wire n_1634;
wire n_5556;
wire n_1452;
wire n_4953;
wire n_7345;
wire n_7472;
wire n_6339;
wire n_4570;
wire n_5391;
wire n_5431;
wire n_3966;
wire n_4293;
wire n_6371;
wire n_6014;
wire n_1577;
wire n_1700;
wire n_4122;
wire n_4542;
wire n_5021;
wire n_2819;
wire n_5456;
wire n_5523;
wire n_1140;
wire n_1985;
wire n_4740;
wire n_3007;
wire n_1487;
wire n_6373;
wire n_1237;
wire n_4230;
wire n_7157;
wire n_1109;
wire n_2741;
wire n_4333;
wire n_7674;
wire n_5231;
wire n_6809;
wire n_5512;
wire n_6406;
wire n_3436;
wire n_6223;
wire n_4460;
wire n_2312;
wire n_2946;
wire n_4040;
wire n_7622;
wire n_7115;
wire n_1884;
wire n_6632;
wire n_2717;
wire n_1589;
wire n_5720;
wire n_7286;
wire n_4527;
wire n_2877;
wire n_5881;
wire n_1996;
wire n_5857;
wire n_5256;
wire n_3964;
wire n_3110;
wire n_5717;
wire n_1677;
wire n_4384;
wire n_2297;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_6654;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_4762;
wire n_5561;
wire n_1877;
wire n_6871;
wire n_1477;
wire n_3155;
wire n_4938;
wire n_5487;
wire n_4407;
wire n_5961;
wire n_5077;
wire n_6672;
wire n_5214;
wire n_1249;
wire n_3468;
wire n_7344;
wire n_2006;
wire n_7714;
wire n_1990;
wire n_5413;
wire n_3680;
wire n_6227;
wire n_7612;
wire n_3624;
wire n_6098;
wire n_4989;
wire n_7744;
wire n_2467;
wire n_5066;
wire n_4292;
wire n_6953;
wire n_7779;
wire n_3145;
wire n_5682;
wire n_6891;
wire n_2662;
wire n_3872;
wire n_5602;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_6163;
wire n_1566;
wire n_1464;
wire n_7127;
wire n_6601;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_6565;
wire n_2277;
wire n_1982;
wire n_2252;
wire n_1695;
wire n_3331;
wire n_2999;
wire n_2910;
wire n_4414;
wire n_6979;
wire n_2294;
wire n_2295;
wire n_4977;
wire n_4706;
wire n_1602;
wire n_2965;
wire n_6076;
wire n_7650;
wire n_5347;
wire n_2382;
wire n_2557;
wire n_2505;
wire n_7050;
wire n_3554;
wire n_7431;
wire n_6199;
wire n_3730;
wire n_4307;
wire n_4356;
wire n_6930;
wire n_1935;
wire n_7770;
wire n_5568;
wire n_3367;
wire n_1146;
wire n_2785;
wire n_7118;
wire n_7259;
wire n_5060;
wire n_4929;
wire n_5121;
wire n_1608;
wire n_3776;
wire n_4951;
wire n_5756;
wire n_5162;
wire n_5224;
wire n_2160;
wire n_2699;
wire n_2991;
wire n_6513;
wire n_6214;
wire n_1436;
wire n_6821;
wire n_4137;
wire n_1485;
wire n_7448;
wire n_2239;
wire n_6289;
wire n_3826;
wire n_4365;
wire n_1979;
wire n_3781;
wire n_6775;
wire n_4215;
wire n_4315;
wire n_6559;
wire n_2971;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_7518;
wire n_3797;
wire n_6683;
wire n_3281;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2934;
wire n_6815;
wire n_6430;
wire n_4042;
wire n_5663;
wire n_2525;
wire n_5552;
wire n_4624;
wire n_6043;
wire n_4317;
wire n_3087;
wire n_7726;
wire n_4925;
wire n_2197;
wire n_7069;
wire n_1470;
wire n_2098;
wire n_1761;
wire n_4041;
wire n_5672;
wire n_7478;
wire n_4958;
wire n_5051;
wire n_4297;
wire n_5367;
wire n_5339;
wire n_4709;
wire n_3379;
wire n_4425;
wire n_3390;
wire n_5000;
wire n_1806;
wire n_1539;
wire n_2711;
wire n_3646;
wire n_7011;
wire n_2209;
wire n_3020;
wire n_3142;
wire n_2612;
wire n_5226;
wire n_2095;
wire n_2486;
wire n_5855;
wire n_5819;
wire n_2521;
wire n_5388;
wire n_1574;
wire n_6608;
wire n_7686;
wire n_6186;
wire n_4764;
wire n_4899;
wire n_6283;
wire n_6445;
wire n_7716;
wire n_4141;
wire n_4614;
wire n_2979;
wire n_4739;
wire n_1300;
wire n_4035;
wire n_4291;
wire n_6372;
wire n_3419;
wire n_4935;
wire n_4880;
wire n_7759;
wire n_3167;
wire n_5188;
wire n_2986;
wire n_4969;
wire n_7675;
wire n_2400;
wire n_6467;
wire n_6144;
wire n_5681;
wire n_2507;
wire n_3682;
wire n_3131;
wire n_1495;
wire n_6291;
wire n_1357;
wire n_6593;
wire n_7482;
wire n_4566;
wire n_5262;
wire n_2794;
wire n_6542;
wire n_3672;
wire n_2496;
wire n_4918;
wire n_2974;
wire n_6763;
wire n_6782;
wire n_7621;
wire n_5604;
wire n_3449;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_4933;
wire n_4872;
wire n_5910;
wire n_1315;
wire n_4647;
wire n_7552;
wire n_6839;
wire n_2340;
wire n_6125;
wire n_2117;
wire n_5990;
wire n_1328;
wire n_4837;
wire n_6218;
wire n_3638;
wire n_2106;
wire n_5880;
wire n_5685;
wire n_7164;
wire n_6619;
wire n_6515;
wire n_6060;
wire n_1263;
wire n_4940;
wire n_4176;
wire n_4454;
wire n_7017;
wire n_7454;
wire n_6664;
wire n_5992;
wire n_5105;
wire n_6761;
wire n_5807;
wire n_3772;
wire n_7769;
wire n_2948;
wire n_4322;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_5449;
wire n_3867;
wire n_4956;
wire n_2045;
wire n_1535;
wire n_4227;
wire n_6599;
wire n_2190;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_3929;
wire n_6974;
wire n_1898;
wire n_1254;
wire n_7312;
wire n_6894;
wire n_2524;
wire n_3927;
wire n_7045;
wire n_1941;
wire n_5338;
wire n_5070;
wire n_3564;
wire n_3095;
wire n_1783;
wire n_5842;
wire n_3279;
wire n_1815;
wire n_3344;
wire n_6173;
wire n_4133;
wire n_6093;
wire n_3985;
wire n_7277;
wire n_6099;
wire n_5939;
wire n_7502;
wire n_5481;
wire n_5187;
wire n_5762;
wire n_3252;
wire n_1162;
wire n_2578;
wire n_5486;
wire n_5426;
wire n_2745;
wire n_2110;
wire n_6031;
wire n_6064;
wire n_6997;
wire n_3747;
wire n_1323;
wire n_6753;
wire n_5846;
wire n_6033;
wire n_3710;
wire n_1429;
wire n_6316;
wire n_3209;
wire n_2026;
wire n_5537;
wire n_3588;
wire n_7778;
wire n_5220;
wire n_6341;
wire n_2103;
wire n_4497;
wire n_4388;
wire n_7359;
wire n_3632;
wire n_5200;
wire n_7225;
wire n_1874;
wire n_7651;
wire n_4116;
wire n_3377;
wire n_5816;
wire n_1601;
wire n_3414;
wire n_2933;
wire n_7020;
wire n_3828;
wire n_1367;
wire n_3240;
wire n_2895;
wire n_1458;
wire n_1694;
wire n_7392;
wire n_2271;
wire n_2356;
wire n_5676;
wire n_5463;
wire n_2261;
wire n_4066;
wire n_2994;
wire n_4980;
wire n_2105;
wire n_2187;
wire n_5780;
wire n_2642;
wire n_6924;
wire n_5485;
wire n_5737;
wire n_6876;
wire n_7424;
wire n_1643;
wire n_1789;
wire n_7625;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_6571;
wire n_1112;
wire n_2384;
wire n_6962;
wire n_1376;
wire n_1858;
wire n_3523;
wire n_2815;
wire n_2446;
wire n_3388;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_6039;
wire n_5355;
wire n_4048;
wire n_7059;
wire n_4084;
wire n_5149;
wire n_1527;
wire n_3174;
wire n_4848;
wire n_6970;
wire n_5185;
wire n_6829;
wire n_2849;
wire n_6509;
wire n_6642;
wire n_5847;
wire n_5091;
wire n_5936;
wire n_1177;
wire n_3292;
wire n_6442;
wire n_7522;
wire n_6636;
wire n_3940;
wire n_6475;
wire n_2502;
wire n_5396;
wire n_4860;
wire n_4438;
wire n_5300;
wire n_6830;
wire n_3290;
wire n_7365;
wire n_3585;
wire n_7094;
wire n_2878;
wire n_1810;
wire n_7439;
wire n_6342;
wire n_3047;
wire n_2610;
wire n_5917;
wire n_7035;
wire n_5306;
wire n_3427;
wire n_1188;
wire n_3431;
wire n_2024;
wire n_3783;
wire n_1503;
wire n_1942;
wire n_4326;
wire n_3141;
wire n_6838;
wire n_2698;
wire n_6869;
wire n_3930;
wire n_4149;
wire n_5518;
wire n_5531;
wire n_1259;
wire n_4101;
wire n_6735;
wire n_4792;
wire n_2916;
wire n_3736;
wire n_2611;
wire n_6012;
wire n_6866;
wire n_4383;
wire n_7395;
wire n_2709;
wire n_5074;
wire n_6492;
wire n_7005;
wire n_2244;
wire n_6387;
wire n_3664;
wire n_1456;
wire n_3907;
wire n_5246;
wire n_2665;
wire n_5544;
wire n_6742;
wire n_3063;
wire n_4543;
wire n_6969;
wire n_2881;
wire n_3862;
wire n_2018;
wire n_3134;
wire n_5652;
wire n_7180;
wire n_5409;
wire n_2581;
wire n_6271;
wire n_5540;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_6929;
wire n_2255;
wire n_1820;
wire n_6986;
wire n_3906;
wire n_3474;
wire n_1946;
wire n_3111;
wire n_4212;
wire n_7752;
wire n_6709;
wire n_4827;
wire n_1639;
wire n_2154;
wire n_6149;
wire n_3162;
wire n_4599;
wire n_2732;
wire n_3004;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4783;
wire n_3276;
wire n_2956;
wire n_1415;
wire n_3743;
wire n_7724;
wire n_4068;
wire n_7385;
wire n_2153;
wire n_5777;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_6545;
wire n_4434;
wire n_2737;
wire n_5557;
wire n_1406;
wire n_3591;
wire n_6054;
wire n_2137;
wire n_7444;
wire n_6756;
wire n_5442;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_1176;
wire n_7620;
wire n_3848;
wire n_1897;
wire n_2477;
wire n_4622;
wire n_5549;
wire n_3139;
wire n_4715;
wire n_7441;
wire n_6250;
wire n_6718;
wire n_4222;
wire n_5730;
wire n_2206;
wire n_3734;
wire n_7078;
wire n_3538;
wire n_4716;
wire n_4588;
wire n_2265;
wire n_5054;
wire n_5349;
wire n_7093;
wire n_1167;
wire n_7333;
wire n_3231;
wire n_6423;
wire n_6659;
wire n_3138;
wire n_6303;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_3349;
wire n_7508;
wire n_4988;
wire n_5128;
wire n_3454;
wire n_6668;
wire n_6299;
wire n_4143;
wire n_5027;
wire n_4410;
wire n_5026;
wire n_5189;
wire n_1718;
wire n_3229;
wire n_6757;
wire n_2546;
wire n_4741;
wire n_6383;
wire n_5516;
wire n_1139;
wire n_2345;
wire n_1324;
wire n_4440;
wire n_7496;
wire n_3649;
wire n_1838;
wire n_6880;
wire n_3824;
wire n_7425;
wire n_3439;
wire n_5525;
wire n_1513;
wire n_5836;
wire n_5677;
wire n_6182;
wire n_6510;
wire n_1788;
wire n_5764;
wire n_2348;
wire n_6171;
wire n_2417;
wire n_7550;
wire n_2043;
wire n_3601;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_7715;
wire n_5768;
wire n_6353;
wire n_7302;
wire n_6472;
wire n_2248;
wire n_3500;
wire n_2850;
wire n_3962;
wire n_6360;
wire n_3846;
wire n_4328;
wire n_7548;
wire n_5142;
wire n_1433;
wire n_6934;
wire n_5082;
wire n_1907;
wire n_6686;
wire n_7019;
wire n_3994;
wire n_5911;
wire n_5118;
wire n_2135;
wire n_5781;
wire n_5739;
wire n_7595;
wire n_1088;
wire n_7088;
wire n_6666;
wire n_6075;
wire n_1102;
wire n_5145;
wire n_7542;
wire n_4487;
wire n_7204;
wire n_7014;
wire n_1165;
wire n_6708;
wire n_5111;
wire n_4148;
wire n_3066;
wire n_6135;
wire n_2869;
wire n_6422;
wire n_4829;
wire n_2455;
wire n_2874;
wire n_4937;
wire n_7665;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_7341;
wire n_7407;
wire n_6266;
wire n_5748;
wire n_1809;
wire n_7757;
wire n_3491;
wire n_4844;
wire n_3271;
wire n_5734;
wire n_2667;
wire n_7514;
wire n_6317;
wire n_7646;
wire n_7653;
wire n_6059;
wire n_5247;
wire n_1565;
wire n_2325;
wire n_6041;
wire n_3346;
wire n_5411;
wire n_5422;
wire n_3391;
wire n_6801;
wire n_1547;
wire n_1542;
wire n_5991;
wire n_1362;
wire n_6343;
wire n_4178;
wire n_4324;
wire n_7193;
wire n_3288;
wire n_2518;
wire n_6069;
wire n_3045;
wire n_3014;
wire n_5475;
wire n_6511;
wire n_1951;
wire n_1330;
wire n_5850;
wire n_6307;
wire n_7373;
wire n_5440;
wire n_1940;
wire n_3767;
wire n_1212;
wire n_1199;
wire n_4852;
wire n_1978;
wire n_1767;
wire n_1443;
wire n_5641;
wire n_1861;
wire n_1564;
wire n_7291;
wire n_2593;
wire n_1623;
wire n_6413;
wire n_6603;
wire n_1131;
wire n_6707;
wire n_3120;
wire n_1554;
wire n_4843;
wire n_7239;
wire n_6255;
wire n_4761;
wire n_6294;
wire n_2021;
wire n_6835;
wire n_7406;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_3342;
wire n_5441;
wire n_2939;
wire n_6587;
wire n_6792;
wire n_4036;
wire n_1147;
wire n_5055;
wire n_4380;
wire n_2790;
wire n_2034;
wire n_3102;
wire n_4345;
wire n_6487;
wire n_1892;
wire n_5761;
wire n_6195;
wire n_2061;
wire n_6038;
wire n_1373;
wire n_7677;
wire n_3866;
wire n_3803;
wire n_2083;
wire n_2119;
wire n_5976;
wire n_7513;
wire n_2207;
wire n_4210;
wire n_7782;
wire n_3485;
wire n_4810;
wire n_3149;
wire n_5871;
wire n_2827;
wire n_5680;
wire n_3278;
wire n_2701;
wire n_6928;
wire n_2337;
wire n_4045;
wire n_4871;
wire n_2513;
wire n_1369;
wire n_1297;
wire n_1734;
wire n_4461;
wire n_2323;
wire n_7242;
wire n_6086;
wire n_5915;
wire n_5524;
wire n_7573;
wire n_5112;
wire n_3042;
wire n_5542;
wire n_5627;
wire n_2561;
wire n_5785;
wire n_2491;
wire n_6438;
wire n_5298;
wire n_7181;
wire n_1161;
wire n_1103;
wire n_6739;
wire n_4363;
wire n_5564;
wire n_5603;
wire n_3551;
wire n_3992;
wire n_4147;
wire n_6451;
wire n_4811;
wire n_6495;
wire n_5093;
wire n_5710;
wire n_3176;
wire n_2429;
wire n_3326;
wire n_5986;
wire n_3581;
wire n_3423;
wire n_1646;
wire n_4161;
wire n_5137;
wire n_1759;
wire n_2096;
wire n_5912;
wire n_2296;
wire n_7139;
wire n_6194;
wire n_1911;
wire n_7586;
wire n_6381;
wire n_7404;
wire n_2870;
wire n_6862;
wire n_4869;
wire n_6397;
wire n_4013;
wire n_1211;
wire n_4482;
wire n_3794;
wire n_6628;
wire n_5283;
wire n_1419;
wire n_7328;
wire n_6783;
wire n_4738;
wire n_7231;
wire n_6604;
wire n_1193;
wire n_2928;
wire n_3380;
wire n_3557;
wire n_7435;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_7058;
wire n_5286;
wire n_2627;
wire n_1827;
wire n_3369;
wire n_5626;
wire n_4086;
wire n_5410;
wire n_4112;
wire n_2501;
wire n_2051;
wire n_1805;
wire n_3737;
wire n_1183;
wire n_7041;
wire n_3160;
wire n_4744;
wire n_1204;
wire n_1151;
wire n_3286;
wire n_1092;
wire n_6788;
wire n_2668;
wire n_6684;
wire n_1386;
wire n_2931;
wire n_7364;
wire n_2492;
wire n_5960;
wire n_3636;
wire n_4787;
wire n_4885;
wire n_2927;
wire n_4459;
wire n_7738;
wire n_1516;
wire n_4551;
wire n_4484;
wire n_5988;
wire n_1499;
wire n_5838;
wire n_2155;
wire n_3938;
wire n_6103;
wire n_7006;
wire n_6016;
wire n_3114;
wire n_3905;
wire n_6817;
wire n_1661;
wire n_6261;
wire n_7276;
wire n_1965;
wire n_5616;
wire n_1757;
wire n_7571;
wire n_7269;
wire n_6399;
wire n_4726;
wire n_3617;
wire n_3602;
wire n_4298;
wire n_6181;
wire n_3053;
wire n_5965;
wire n_3894;
wire n_6645;
wire n_2407;
wire n_6845;
wire n_2267;
wire n_2302;
wire n_2082;
wire n_2453;
wire n_2560;
wire n_6572;
wire n_4544;
wire n_7531;
wire n_7222;
wire n_4418;
wire n_4595;
wire n_2770;
wire n_7463;
wire n_2704;
wire n_6246;
wire n_1762;
wire n_7347;
wire n_4944;
wire n_7060;
wire n_4468;
wire n_5923;
wire n_6357;
wire n_6508;
wire n_6536;
wire n_3421;
wire n_7064;
wire n_4950;
wire n_3247;
wire n_1454;
wire n_4108;
wire n_6917;
wire n_7545;
wire n_4594;
wire n_6359;
wire n_5949;
wire n_7479;
wire n_1325;
wire n_2754;
wire n_4629;
wire n_4903;
wire n_3041;
wire n_7400;
wire n_4194;
wire n_3713;
wire n_2692;
wire n_5738;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_2324;
wire n_6096;
wire n_4921;
wire n_1111;
wire n_1819;
wire n_4863;
wire n_6813;
wire n_2670;
wire n_7379;
wire n_1745;
wire n_7352;
wire n_7318;
wire n_3941;
wire n_3516;
wire n_3933;
wire n_7295;
wire n_3562;
wire n_1916;
wire n_3873;
wire n_7267;
wire n_2073;
wire n_4093;
wire n_1947;
wire n_2165;
wire n_2016;
wire n_3793;
wire n_5080;
wire n_7497;
wire n_5975;
wire n_1791;
wire n_5301;
wire n_6464;
wire n_1113;
wire n_6963;
wire n_4817;
wire n_1468;
wire n_4917;
wire n_6017;
wire n_5507;
wire n_1164;
wire n_6340;
wire n_7543;
wire n_3749;
wire n_5470;
wire n_6315;
wire n_6923;
wire n_3691;
wire n_4452;
wire n_3501;
wire n_2538;
wire n_1559;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_6392;
wire n_4280;
wire n_2285;
wire n_5979;
wire n_1934;
wire n_2040;
wire n_3246;
wire n_2186;
wire n_5648;
wire n_1665;
wire n_5335;
wire n_5594;
wire n_3417;
wire n_2725;
wire n_6681;
wire n_1482;
wire n_5393;
wire n_4782;
wire n_5661;
wire n_4978;
wire n_6292;
wire n_5690;
wire n_2349;
wire n_1902;
wire n_2474;
wire n_6154;
wire n_7460;
wire n_5963;
wire n_6293;
wire n_1417;
wire n_5455;
wire n_7061;
wire n_7351;
wire n_3536;
wire n_1346;
wire n_5873;
wire n_2834;
wire n_6127;
wire n_1123;
wire n_1272;
wire n_7298;
wire n_2497;
wire n_7195;
wire n_3040;
wire n_6028;
wire n_6325;
wire n_1410;
wire n_6600;
wire n_3528;
wire n_3677;
wire n_2657;
wire n_6957;
wire n_2743;
wire n_5698;
wire n_4662;
wire n_2658;

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_294),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_972),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_574),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_909),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_503),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_1009),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_48),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_861),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_114),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_860),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_946),
.Y(n_1088)
);

INVx1_ASAP7_75t_SL g1089 ( 
.A(n_168),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_158),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_557),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_537),
.Y(n_1092)
);

INVx1_ASAP7_75t_SL g1093 ( 
.A(n_988),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_602),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_644),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_305),
.Y(n_1096)
);

CKINVDCx16_ASAP7_75t_R g1097 ( 
.A(n_137),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_171),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_295),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_659),
.Y(n_1100)
);

BUFx5_ASAP7_75t_L g1101 ( 
.A(n_972),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_442),
.Y(n_1102)
);

BUFx10_ASAP7_75t_L g1103 ( 
.A(n_989),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1018),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_778),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_40),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_953),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_827),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_999),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_1067),
.Y(n_1110)
);

CKINVDCx16_ASAP7_75t_R g1111 ( 
.A(n_1035),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_161),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_396),
.Y(n_1113)
);

INVx4_ASAP7_75t_R g1114 ( 
.A(n_431),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_353),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_912),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_306),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_233),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_815),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_190),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_398),
.Y(n_1121)
);

BUFx10_ASAP7_75t_L g1122 ( 
.A(n_328),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_986),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_462),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_321),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_328),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_91),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_189),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_226),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_837),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_999),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_465),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_809),
.Y(n_1133)
);

INVx1_ASAP7_75t_SL g1134 ( 
.A(n_606),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_434),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_715),
.Y(n_1136)
);

CKINVDCx20_ASAP7_75t_R g1137 ( 
.A(n_1005),
.Y(n_1137)
);

CKINVDCx20_ASAP7_75t_R g1138 ( 
.A(n_814),
.Y(n_1138)
);

CKINVDCx14_ASAP7_75t_R g1139 ( 
.A(n_983),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_218),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_928),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_458),
.Y(n_1142)
);

INVxp67_ASAP7_75t_L g1143 ( 
.A(n_674),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_780),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_1017),
.Y(n_1145)
);

CKINVDCx16_ASAP7_75t_R g1146 ( 
.A(n_577),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_695),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_378),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_737),
.Y(n_1149)
);

HB1xp67_ASAP7_75t_L g1150 ( 
.A(n_264),
.Y(n_1150)
);

INVx4_ASAP7_75t_R g1151 ( 
.A(n_999),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_571),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_350),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_314),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1025),
.Y(n_1155)
);

BUFx8_ASAP7_75t_SL g1156 ( 
.A(n_1072),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1076),
.Y(n_1157)
);

CKINVDCx20_ASAP7_75t_R g1158 ( 
.A(n_405),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_376),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_327),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_506),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_848),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_1059),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_973),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_984),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_740),
.Y(n_1166)
);

INVxp67_ASAP7_75t_L g1167 ( 
.A(n_514),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_39),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_970),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_613),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_487),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_495),
.Y(n_1172)
);

INVx1_ASAP7_75t_SL g1173 ( 
.A(n_846),
.Y(n_1173)
);

CKINVDCx14_ASAP7_75t_R g1174 ( 
.A(n_62),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_967),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_21),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_981),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_410),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_956),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_723),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_17),
.Y(n_1181)
);

INVx1_ASAP7_75t_SL g1182 ( 
.A(n_855),
.Y(n_1182)
);

CKINVDCx20_ASAP7_75t_R g1183 ( 
.A(n_295),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_118),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_183),
.Y(n_1185)
);

INVx2_ASAP7_75t_SL g1186 ( 
.A(n_809),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_607),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_667),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_207),
.Y(n_1189)
);

CKINVDCx20_ASAP7_75t_R g1190 ( 
.A(n_1013),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_829),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_1023),
.Y(n_1192)
);

INVx1_ASAP7_75t_SL g1193 ( 
.A(n_688),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_993),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_1071),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_350),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_30),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_861),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_905),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_1039),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_1074),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_407),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_531),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_611),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_224),
.Y(n_1205)
);

BUFx10_ASAP7_75t_L g1206 ( 
.A(n_156),
.Y(n_1206)
);

BUFx10_ASAP7_75t_L g1207 ( 
.A(n_935),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_28),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_94),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_354),
.Y(n_1210)
);

CKINVDCx20_ASAP7_75t_R g1211 ( 
.A(n_32),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_1010),
.Y(n_1212)
);

INVx1_ASAP7_75t_SL g1213 ( 
.A(n_269),
.Y(n_1213)
);

INVx1_ASAP7_75t_SL g1214 ( 
.A(n_47),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_30),
.Y(n_1215)
);

INVx2_ASAP7_75t_SL g1216 ( 
.A(n_698),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_127),
.Y(n_1217)
);

BUFx10_ASAP7_75t_L g1218 ( 
.A(n_1004),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_932),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_120),
.Y(n_1220)
);

CKINVDCx20_ASAP7_75t_R g1221 ( 
.A(n_244),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_894),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_240),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_107),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_171),
.Y(n_1225)
);

CKINVDCx20_ASAP7_75t_R g1226 ( 
.A(n_462),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_203),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_17),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_503),
.Y(n_1229)
);

INVx2_ASAP7_75t_SL g1230 ( 
.A(n_945),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_595),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_467),
.Y(n_1232)
);

INVx4_ASAP7_75t_R g1233 ( 
.A(n_632),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_597),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_850),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_428),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_906),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_171),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_48),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1012),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_925),
.Y(n_1241)
);

CKINVDCx20_ASAP7_75t_R g1242 ( 
.A(n_261),
.Y(n_1242)
);

CKINVDCx20_ASAP7_75t_R g1243 ( 
.A(n_213),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_73),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_285),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_1034),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_831),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_155),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_380),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_980),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_526),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_962),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_1008),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_224),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1028),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_761),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_150),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_81),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_477),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_208),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_725),
.Y(n_1261)
);

BUFx10_ASAP7_75t_L g1262 ( 
.A(n_37),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_841),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_165),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_441),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_490),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_548),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_727),
.Y(n_1268)
);

CKINVDCx20_ASAP7_75t_R g1269 ( 
.A(n_789),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_950),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_932),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_927),
.Y(n_1272)
);

CKINVDCx20_ASAP7_75t_R g1273 ( 
.A(n_329),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_510),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_395),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_1021),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_243),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_60),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_106),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_456),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_779),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_307),
.Y(n_1282)
);

CKINVDCx16_ASAP7_75t_R g1283 ( 
.A(n_635),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_21),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_83),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_675),
.Y(n_1286)
);

INVx1_ASAP7_75t_SL g1287 ( 
.A(n_330),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_344),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_31),
.Y(n_1289)
);

BUFx10_ASAP7_75t_L g1290 ( 
.A(n_321),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_466),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1000),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_804),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_463),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1041),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_1029),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_125),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_518),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_661),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_548),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_102),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_518),
.Y(n_1302)
);

CKINVDCx12_ASAP7_75t_R g1303 ( 
.A(n_217),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_340),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_280),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_958),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_589),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_960),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_798),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_30),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_1062),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1033),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_703),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_366),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_101),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_76),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_1006),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_536),
.Y(n_1318)
);

BUFx10_ASAP7_75t_L g1319 ( 
.A(n_53),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_45),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_997),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_201),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_200),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_835),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_574),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_259),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_450),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1016),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1069),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_299),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_785),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_617),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_579),
.Y(n_1333)
);

INVx2_ASAP7_75t_SL g1334 ( 
.A(n_1002),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_694),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_796),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_342),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_467),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1005),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_913),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_602),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_1036),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_511),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_981),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_885),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_395),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_987),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_29),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_94),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_183),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_593),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_916),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_279),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_456),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_670),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_525),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_848),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_620),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1040),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_871),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_279),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_238),
.Y(n_1362)
);

INVx1_ASAP7_75t_SL g1363 ( 
.A(n_421),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_659),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_844),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1022),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_977),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_807),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_497),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_971),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_609),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_441),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1011),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_390),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_777),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_902),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_358),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_923),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_1030),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_904),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_71),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_959),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_159),
.Y(n_1383)
);

CKINVDCx16_ASAP7_75t_R g1384 ( 
.A(n_549),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1020),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_663),
.Y(n_1386)
);

CKINVDCx14_ASAP7_75t_R g1387 ( 
.A(n_530),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_722),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_472),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_668),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_541),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_1056),
.Y(n_1392)
);

INVx2_ASAP7_75t_SL g1393 ( 
.A(n_499),
.Y(n_1393)
);

INVx1_ASAP7_75t_SL g1394 ( 
.A(n_362),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1002),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1003),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_658),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_519),
.Y(n_1398)
);

CKINVDCx16_ASAP7_75t_R g1399 ( 
.A(n_683),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_699),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_47),
.Y(n_1401)
);

INVx1_ASAP7_75t_SL g1402 ( 
.A(n_273),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1075),
.Y(n_1403)
);

INVxp67_ASAP7_75t_SL g1404 ( 
.A(n_871),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_843),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_264),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_691),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_948),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_300),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_1032),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_137),
.Y(n_1411)
);

CKINVDCx20_ASAP7_75t_R g1412 ( 
.A(n_772),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1011),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_408),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_808),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_222),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_474),
.Y(n_1417)
);

CKINVDCx20_ASAP7_75t_R g1418 ( 
.A(n_1033),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_93),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1002),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_151),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_162),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_153),
.Y(n_1423)
);

BUFx10_ASAP7_75t_L g1424 ( 
.A(n_17),
.Y(n_1424)
);

CKINVDCx20_ASAP7_75t_R g1425 ( 
.A(n_435),
.Y(n_1425)
);

CKINVDCx20_ASAP7_75t_R g1426 ( 
.A(n_182),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_384),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_239),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_991),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_982),
.Y(n_1430)
);

INVx2_ASAP7_75t_SL g1431 ( 
.A(n_952),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_995),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_280),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_393),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_127),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_749),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_222),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_818),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_922),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_403),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_99),
.Y(n_1441)
);

BUFx10_ASAP7_75t_L g1442 ( 
.A(n_193),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_120),
.Y(n_1443)
);

INVx2_ASAP7_75t_SL g1444 ( 
.A(n_255),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_725),
.Y(n_1445)
);

INVxp67_ASAP7_75t_L g1446 ( 
.A(n_370),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_643),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_101),
.Y(n_1448)
);

CKINVDCx16_ASAP7_75t_R g1449 ( 
.A(n_444),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_492),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_123),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_388),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_20),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_455),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_828),
.Y(n_1455)
);

INVx1_ASAP7_75t_SL g1456 ( 
.A(n_273),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_279),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_192),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_288),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_792),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_246),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_428),
.Y(n_1462)
);

BUFx8_ASAP7_75t_SL g1463 ( 
.A(n_1028),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_330),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_146),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_123),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_767),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_162),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1013),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_673),
.Y(n_1470)
);

INVx1_ASAP7_75t_SL g1471 ( 
.A(n_578),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_585),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_732),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_490),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_329),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_109),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_981),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_122),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_394),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_101),
.Y(n_1480)
);

CKINVDCx16_ASAP7_75t_R g1481 ( 
.A(n_872),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_373),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_520),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_793),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_994),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_116),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_455),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1001),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_475),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1047),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_145),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_415),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_1037),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_942),
.Y(n_1494)
);

INVx1_ASAP7_75t_SL g1495 ( 
.A(n_1041),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_256),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_392),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_1059),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_125),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_604),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_504),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_41),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_969),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_82),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_845),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_286),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_244),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_1054),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_956),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_767),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_947),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_501),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1021),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_921),
.Y(n_1514)
);

CKINVDCx20_ASAP7_75t_R g1515 ( 
.A(n_978),
.Y(n_1515)
);

CKINVDCx20_ASAP7_75t_R g1516 ( 
.A(n_995),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_868),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_842),
.Y(n_1518)
);

CKINVDCx20_ASAP7_75t_R g1519 ( 
.A(n_1049),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_950),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1059),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_682),
.Y(n_1522)
);

CKINVDCx20_ASAP7_75t_R g1523 ( 
.A(n_65),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_449),
.Y(n_1524)
);

CKINVDCx16_ASAP7_75t_R g1525 ( 
.A(n_133),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1077),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_659),
.Y(n_1527)
);

BUFx3_ASAP7_75t_L g1528 ( 
.A(n_976),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_957),
.Y(n_1529)
);

BUFx2_ASAP7_75t_SL g1530 ( 
.A(n_992),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_51),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_838),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_153),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_75),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_655),
.Y(n_1535)
);

BUFx6f_ASAP7_75t_L g1536 ( 
.A(n_577),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_178),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_404),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_710),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1015),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_810),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_55),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_1034),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_508),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_134),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_5),
.Y(n_1546)
);

BUFx10_ASAP7_75t_L g1547 ( 
.A(n_40),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_958),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_741),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_280),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_209),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_701),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_975),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_543),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_601),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_685),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_892),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_997),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_510),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_739),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_12),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_104),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_459),
.Y(n_1563)
);

CKINVDCx20_ASAP7_75t_R g1564 ( 
.A(n_142),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_626),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_506),
.Y(n_1566)
);

BUFx3_ASAP7_75t_L g1567 ( 
.A(n_565),
.Y(n_1567)
);

BUFx10_ASAP7_75t_L g1568 ( 
.A(n_1044),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_1009),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_468),
.Y(n_1570)
);

CKINVDCx20_ASAP7_75t_R g1571 ( 
.A(n_336),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_854),
.Y(n_1572)
);

BUFx3_ASAP7_75t_L g1573 ( 
.A(n_265),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_518),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_892),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_914),
.Y(n_1576)
);

BUFx3_ASAP7_75t_L g1577 ( 
.A(n_201),
.Y(n_1577)
);

BUFx6f_ASAP7_75t_L g1578 ( 
.A(n_833),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_653),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_663),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_584),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_893),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_177),
.Y(n_1583)
);

CKINVDCx20_ASAP7_75t_R g1584 ( 
.A(n_334),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1012),
.Y(n_1585)
);

CKINVDCx16_ASAP7_75t_R g1586 ( 
.A(n_1007),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_965),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_965),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_708),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_289),
.Y(n_1590)
);

BUFx10_ASAP7_75t_L g1591 ( 
.A(n_742),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_70),
.Y(n_1592)
);

CKINVDCx20_ASAP7_75t_R g1593 ( 
.A(n_399),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_785),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_749),
.Y(n_1595)
);

CKINVDCx20_ASAP7_75t_R g1596 ( 
.A(n_652),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_256),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_1014),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_681),
.Y(n_1599)
);

CKINVDCx20_ASAP7_75t_R g1600 ( 
.A(n_399),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_449),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_702),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_990),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_1027),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_66),
.Y(n_1605)
);

BUFx3_ASAP7_75t_L g1606 ( 
.A(n_45),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_217),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_955),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_433),
.Y(n_1609)
);

CKINVDCx16_ASAP7_75t_R g1610 ( 
.A(n_299),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1024),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_671),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_949),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_117),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_495),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_548),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_992),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1043),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_1054),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_1019),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_333),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_906),
.Y(n_1622)
);

INVx2_ASAP7_75t_SL g1623 ( 
.A(n_985),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_536),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_394),
.Y(n_1625)
);

BUFx3_ASAP7_75t_L g1626 ( 
.A(n_10),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_954),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_438),
.Y(n_1628)
);

INVx1_ASAP7_75t_SL g1629 ( 
.A(n_736),
.Y(n_1629)
);

INVx1_ASAP7_75t_SL g1630 ( 
.A(n_830),
.Y(n_1630)
);

INVx2_ASAP7_75t_SL g1631 ( 
.A(n_961),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_673),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_62),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_31),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_344),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_174),
.Y(n_1636)
);

CKINVDCx14_ASAP7_75t_R g1637 ( 
.A(n_299),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1038),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_344),
.Y(n_1639)
);

BUFx6f_ASAP7_75t_L g1640 ( 
.A(n_655),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_658),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_496),
.Y(n_1642)
);

BUFx3_ASAP7_75t_L g1643 ( 
.A(n_197),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_228),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1019),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_963),
.Y(n_1646)
);

BUFx10_ASAP7_75t_L g1647 ( 
.A(n_262),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_996),
.Y(n_1648)
);

INVx1_ASAP7_75t_SL g1649 ( 
.A(n_998),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_214),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_716),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_625),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_656),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_413),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_639),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_1031),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_641),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_228),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_735),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_306),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1040),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_522),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_941),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_774),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_979),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_10),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_650),
.Y(n_1667)
);

BUFx6f_ASAP7_75t_L g1668 ( 
.A(n_949),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_777),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_772),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_674),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_568),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_105),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_968),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_771),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_459),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_1026),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_252),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_353),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_964),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_594),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_951),
.Y(n_1682)
);

BUFx5_ASAP7_75t_L g1683 ( 
.A(n_338),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_594),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_735),
.Y(n_1685)
);

CKINVDCx20_ASAP7_75t_R g1686 ( 
.A(n_65),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_820),
.Y(n_1687)
);

BUFx10_ASAP7_75t_L g1688 ( 
.A(n_48),
.Y(n_1688)
);

CKINVDCx20_ASAP7_75t_R g1689 ( 
.A(n_172),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_72),
.Y(n_1690)
);

INVx1_ASAP7_75t_SL g1691 ( 
.A(n_464),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_155),
.Y(n_1692)
);

BUFx8_ASAP7_75t_SL g1693 ( 
.A(n_955),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_956),
.Y(n_1694)
);

BUFx6f_ASAP7_75t_L g1695 ( 
.A(n_976),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_194),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_966),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_994),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_805),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_259),
.Y(n_1700)
);

CKINVDCx5p33_ASAP7_75t_R g1701 ( 
.A(n_422),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_563),
.Y(n_1702)
);

CKINVDCx5p33_ASAP7_75t_R g1703 ( 
.A(n_442),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_935),
.Y(n_1704)
);

BUFx2_ASAP7_75t_L g1705 ( 
.A(n_372),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_98),
.Y(n_1706)
);

CKINVDCx16_ASAP7_75t_R g1707 ( 
.A(n_326),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_328),
.Y(n_1708)
);

CKINVDCx20_ASAP7_75t_R g1709 ( 
.A(n_35),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_542),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_441),
.Y(n_1711)
);

INVx2_ASAP7_75t_SL g1712 ( 
.A(n_974),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_569),
.Y(n_1713)
);

INVxp67_ASAP7_75t_SL g1714 ( 
.A(n_646),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_912),
.Y(n_1715)
);

INVx2_ASAP7_75t_SL g1716 ( 
.A(n_240),
.Y(n_1716)
);

CKINVDCx20_ASAP7_75t_R g1717 ( 
.A(n_64),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_59),
.Y(n_1718)
);

INVx2_ASAP7_75t_SL g1719 ( 
.A(n_392),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_473),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_219),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_315),
.Y(n_1722)
);

CKINVDCx14_ASAP7_75t_R g1723 ( 
.A(n_1139),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1262),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1262),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1262),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1424),
.Y(n_1727)
);

BUFx3_ASAP7_75t_L g1728 ( 
.A(n_1626),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_1139),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1424),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1424),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_1174),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1547),
.Y(n_1733)
);

BUFx10_ASAP7_75t_L g1734 ( 
.A(n_1181),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_1174),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1547),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1547),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1106),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1176),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_1387),
.Y(n_1740)
);

CKINVDCx20_ASAP7_75t_R g1741 ( 
.A(n_1211),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_1387),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_1637),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1197),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1208),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1348),
.Y(n_1746)
);

INVxp67_ASAP7_75t_SL g1747 ( 
.A(n_1626),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1186),
.Y(n_1748)
);

BUFx2_ASAP7_75t_L g1749 ( 
.A(n_1637),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1216),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_1156),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1393),
.Y(n_1752)
);

INVxp67_ASAP7_75t_L g1753 ( 
.A(n_1381),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1431),
.Y(n_1754)
);

INVxp67_ASAP7_75t_L g1755 ( 
.A(n_1705),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1444),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1101),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1445),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_1156),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1101),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1473),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_1463),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_1463),
.Y(n_1763)
);

CKINVDCx5p33_ASAP7_75t_R g1764 ( 
.A(n_1693),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1150),
.Y(n_1765)
);

INVxp67_ASAP7_75t_L g1766 ( 
.A(n_1618),
.Y(n_1766)
);

INVxp67_ASAP7_75t_SL g1767 ( 
.A(n_1380),
.Y(n_1767)
);

BUFx3_ASAP7_75t_L g1768 ( 
.A(n_1380),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1623),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1101),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1631),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1716),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1719),
.Y(n_1773)
);

CKINVDCx16_ASAP7_75t_R g1774 ( 
.A(n_1097),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_1693),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1380),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1403),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1403),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_1303),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_1215),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1403),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1661),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1230),
.Y(n_1783)
);

CKINVDCx20_ASAP7_75t_R g1784 ( 
.A(n_1211),
.Y(n_1784)
);

INVxp67_ASAP7_75t_SL g1785 ( 
.A(n_1102),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1230),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1311),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1101),
.Y(n_1788)
);

BUFx6f_ASAP7_75t_L g1789 ( 
.A(n_1159),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1311),
.Y(n_1790)
);

BUFx3_ASAP7_75t_L g1791 ( 
.A(n_1101),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1334),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1334),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_1284),
.Y(n_1794)
);

INVxp67_ASAP7_75t_SL g1795 ( 
.A(n_1102),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1712),
.Y(n_1796)
);

CKINVDCx20_ASAP7_75t_R g1797 ( 
.A(n_1228),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1712),
.Y(n_1798)
);

BUFx3_ASAP7_75t_L g1799 ( 
.A(n_1101),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1082),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1094),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1101),
.Y(n_1802)
);

INVx3_ASAP7_75t_L g1803 ( 
.A(n_1103),
.Y(n_1803)
);

CKINVDCx20_ASAP7_75t_R g1804 ( 
.A(n_1228),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1095),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1096),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_1289),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1104),
.Y(n_1808)
);

CKINVDCx5p33_ASAP7_75t_R g1809 ( 
.A(n_1310),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_1453),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1113),
.Y(n_1811)
);

INVxp67_ASAP7_75t_L g1812 ( 
.A(n_1124),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1115),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1683),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1117),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1119),
.Y(n_1816)
);

INVxp67_ASAP7_75t_SL g1817 ( 
.A(n_1124),
.Y(n_1817)
);

INVx1_ASAP7_75t_SL g1818 ( 
.A(n_1168),
.Y(n_1818)
);

CKINVDCx5p33_ASAP7_75t_R g1819 ( 
.A(n_1502),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1126),
.Y(n_1820)
);

NOR2xp67_ASAP7_75t_L g1821 ( 
.A(n_1128),
.B(n_0),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1683),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_1546),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1131),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1133),
.Y(n_1825)
);

CKINVDCx14_ASAP7_75t_R g1826 ( 
.A(n_1103),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1683),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1135),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1140),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_L g1830 ( 
.A(n_1111),
.B(n_0),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1142),
.Y(n_1831)
);

INVx1_ASAP7_75t_SL g1832 ( 
.A(n_1561),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1147),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1157),
.Y(n_1834)
);

CKINVDCx20_ASAP7_75t_R g1835 ( 
.A(n_1709),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1683),
.Y(n_1836)
);

INVx2_ASAP7_75t_SL g1837 ( 
.A(n_1103),
.Y(n_1837)
);

CKINVDCx16_ASAP7_75t_R g1838 ( 
.A(n_1146),
.Y(n_1838)
);

INVxp33_ASAP7_75t_L g1839 ( 
.A(n_1160),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_1634),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1683),
.Y(n_1841)
);

CKINVDCx5p33_ASAP7_75t_R g1842 ( 
.A(n_1666),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1161),
.Y(n_1843)
);

INVxp67_ASAP7_75t_SL g1844 ( 
.A(n_1220),
.Y(n_1844)
);

INVxp67_ASAP7_75t_L g1845 ( 
.A(n_1220),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1169),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1175),
.Y(n_1847)
);

CKINVDCx20_ASAP7_75t_R g1848 ( 
.A(n_1709),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1178),
.Y(n_1849)
);

INVxp67_ASAP7_75t_SL g1850 ( 
.A(n_1241),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_1283),
.Y(n_1851)
);

CKINVDCx20_ASAP7_75t_R g1852 ( 
.A(n_1105),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1179),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1184),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1185),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1188),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1189),
.Y(n_1857)
);

INVxp67_ASAP7_75t_SL g1858 ( 
.A(n_1241),
.Y(n_1858)
);

CKINVDCx20_ASAP7_75t_R g1859 ( 
.A(n_1741),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1768),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1795),
.Y(n_1861)
);

HB1xp67_ASAP7_75t_L g1862 ( 
.A(n_1818),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1795),
.Y(n_1863)
);

CKINVDCx16_ASAP7_75t_R g1864 ( 
.A(n_1826),
.Y(n_1864)
);

INVxp67_ASAP7_75t_SL g1865 ( 
.A(n_1818),
.Y(n_1865)
);

INVxp67_ASAP7_75t_L g1866 ( 
.A(n_1765),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1817),
.Y(n_1867)
);

INVxp67_ASAP7_75t_L g1868 ( 
.A(n_1749),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_1780),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_1794),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_1807),
.Y(n_1871)
);

CKINVDCx5p33_ASAP7_75t_R g1872 ( 
.A(n_1809),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1817),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1858),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1858),
.Y(n_1875)
);

CKINVDCx5p33_ASAP7_75t_R g1876 ( 
.A(n_1810),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1803),
.B(n_1384),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1728),
.Y(n_1878)
);

BUFx6f_ASAP7_75t_SL g1879 ( 
.A(n_1734),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1747),
.Y(n_1880)
);

BUFx3_ASAP7_75t_L g1881 ( 
.A(n_1734),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1767),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1812),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_1819),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_1823),
.Y(n_1885)
);

NOR2xp33_ASAP7_75t_L g1886 ( 
.A(n_1803),
.B(n_1399),
.Y(n_1886)
);

CKINVDCx20_ASAP7_75t_R g1887 ( 
.A(n_1784),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1812),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1845),
.Y(n_1889)
);

CKINVDCx20_ASAP7_75t_R g1890 ( 
.A(n_1797),
.Y(n_1890)
);

INVxp67_ASAP7_75t_SL g1891 ( 
.A(n_1766),
.Y(n_1891)
);

CKINVDCx20_ASAP7_75t_R g1892 ( 
.A(n_1804),
.Y(n_1892)
);

CKINVDCx20_ASAP7_75t_R g1893 ( 
.A(n_1835),
.Y(n_1893)
);

HB1xp67_ASAP7_75t_L g1894 ( 
.A(n_1832),
.Y(n_1894)
);

INVxp33_ASAP7_75t_SL g1895 ( 
.A(n_1840),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_1842),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1845),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1783),
.Y(n_1898)
);

NOR2xp67_ASAP7_75t_L g1899 ( 
.A(n_1753),
.B(n_1143),
.Y(n_1899)
);

INVx3_ASAP7_75t_L g1900 ( 
.A(n_1786),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1791),
.Y(n_1901)
);

CKINVDCx5p33_ASAP7_75t_R g1902 ( 
.A(n_1751),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1787),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_1759),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1790),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_1762),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1792),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_1763),
.Y(n_1908)
);

INVxp67_ASAP7_75t_SL g1909 ( 
.A(n_1766),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1793),
.Y(n_1910)
);

CKINVDCx20_ASAP7_75t_R g1911 ( 
.A(n_1848),
.Y(n_1911)
);

CKINVDCx20_ASAP7_75t_R g1912 ( 
.A(n_1852),
.Y(n_1912)
);

CKINVDCx5p33_ASAP7_75t_R g1913 ( 
.A(n_1764),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1796),
.Y(n_1914)
);

NOR2xp67_ASAP7_75t_L g1915 ( 
.A(n_1753),
.B(n_1167),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1798),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1785),
.Y(n_1917)
);

CKINVDCx5p33_ASAP7_75t_R g1918 ( 
.A(n_1775),
.Y(n_1918)
);

HB1xp67_ASAP7_75t_L g1919 ( 
.A(n_1832),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1844),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1850),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1748),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1750),
.Y(n_1923)
);

CKINVDCx20_ASAP7_75t_R g1924 ( 
.A(n_1774),
.Y(n_1924)
);

CKINVDCx5p33_ASAP7_75t_R g1925 ( 
.A(n_1838),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1755),
.B(n_1782),
.Y(n_1926)
);

CKINVDCx5p33_ASAP7_75t_R g1927 ( 
.A(n_1723),
.Y(n_1927)
);

CKINVDCx5p33_ASAP7_75t_R g1928 ( 
.A(n_1851),
.Y(n_1928)
);

NOR2xp33_ASAP7_75t_L g1929 ( 
.A(n_1837),
.B(n_1449),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1752),
.Y(n_1930)
);

CKINVDCx5p33_ASAP7_75t_R g1931 ( 
.A(n_1779),
.Y(n_1931)
);

HB1xp67_ASAP7_75t_L g1932 ( 
.A(n_1755),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1754),
.Y(n_1933)
);

CKINVDCx5p33_ASAP7_75t_R g1934 ( 
.A(n_1729),
.Y(n_1934)
);

CKINVDCx5p33_ASAP7_75t_R g1935 ( 
.A(n_1732),
.Y(n_1935)
);

CKINVDCx5p33_ASAP7_75t_R g1936 ( 
.A(n_1735),
.Y(n_1936)
);

NOR2xp33_ASAP7_75t_L g1937 ( 
.A(n_1724),
.B(n_1481),
.Y(n_1937)
);

CKINVDCx20_ASAP7_75t_R g1938 ( 
.A(n_1740),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1799),
.Y(n_1939)
);

INVxp67_ASAP7_75t_L g1940 ( 
.A(n_1725),
.Y(n_1940)
);

CKINVDCx16_ASAP7_75t_R g1941 ( 
.A(n_1830),
.Y(n_1941)
);

NOR2xp33_ASAP7_75t_L g1942 ( 
.A(n_1726),
.B(n_1525),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1756),
.Y(n_1943)
);

CKINVDCx20_ASAP7_75t_R g1944 ( 
.A(n_1742),
.Y(n_1944)
);

CKINVDCx5p33_ASAP7_75t_R g1945 ( 
.A(n_1743),
.Y(n_1945)
);

INVxp67_ASAP7_75t_L g1946 ( 
.A(n_1727),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_1730),
.Y(n_1947)
);

HB1xp67_ASAP7_75t_L g1948 ( 
.A(n_1839),
.Y(n_1948)
);

CKINVDCx5p33_ASAP7_75t_R g1949 ( 
.A(n_1731),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1733),
.B(n_1586),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1758),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1761),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1769),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_1736),
.Y(n_1954)
);

CKINVDCx20_ASAP7_75t_R g1955 ( 
.A(n_1737),
.Y(n_1955)
);

CKINVDCx20_ASAP7_75t_R g1956 ( 
.A(n_1771),
.Y(n_1956)
);

CKINVDCx5p33_ASAP7_75t_R g1957 ( 
.A(n_1772),
.Y(n_1957)
);

CKINVDCx5p33_ASAP7_75t_R g1958 ( 
.A(n_1773),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1776),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1777),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1778),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1781),
.Y(n_1962)
);

INVxp33_ASAP7_75t_SL g1963 ( 
.A(n_1738),
.Y(n_1963)
);

CKINVDCx16_ASAP7_75t_R g1964 ( 
.A(n_1739),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1744),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1745),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1746),
.Y(n_1967)
);

CKINVDCx20_ASAP7_75t_R g1968 ( 
.A(n_1800),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1801),
.Y(n_1969)
);

CKINVDCx5p33_ASAP7_75t_R g1970 ( 
.A(n_1805),
.Y(n_1970)
);

INVx1_ASAP7_75t_SL g1971 ( 
.A(n_1857),
.Y(n_1971)
);

CKINVDCx20_ASAP7_75t_R g1972 ( 
.A(n_1806),
.Y(n_1972)
);

NOR2xp67_ASAP7_75t_L g1973 ( 
.A(n_1808),
.B(n_1446),
.Y(n_1973)
);

CKINVDCx5p33_ASAP7_75t_R g1974 ( 
.A(n_1811),
.Y(n_1974)
);

CKINVDCx5p33_ASAP7_75t_R g1975 ( 
.A(n_1813),
.Y(n_1975)
);

BUFx3_ASAP7_75t_L g1976 ( 
.A(n_1757),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1760),
.Y(n_1977)
);

BUFx2_ASAP7_75t_L g1978 ( 
.A(n_1815),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1816),
.Y(n_1979)
);

INVxp67_ASAP7_75t_SL g1980 ( 
.A(n_1820),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1824),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1825),
.Y(n_1982)
);

CKINVDCx5p33_ASAP7_75t_R g1983 ( 
.A(n_1828),
.Y(n_1983)
);

NOR2xp67_ASAP7_75t_L g1984 ( 
.A(n_1829),
.B(n_1252),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1831),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1833),
.Y(n_1986)
);

CKINVDCx20_ASAP7_75t_R g1987 ( 
.A(n_1834),
.Y(n_1987)
);

CKINVDCx20_ASAP7_75t_R g1988 ( 
.A(n_1843),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1846),
.Y(n_1989)
);

CKINVDCx20_ASAP7_75t_R g1990 ( 
.A(n_1847),
.Y(n_1990)
);

CKINVDCx20_ASAP7_75t_R g1991 ( 
.A(n_1849),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1853),
.B(n_1610),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_1854),
.Y(n_1993)
);

HB1xp67_ASAP7_75t_L g1994 ( 
.A(n_1855),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1770),
.Y(n_1995)
);

CKINVDCx20_ASAP7_75t_R g1996 ( 
.A(n_1856),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1788),
.Y(n_1997)
);

CKINVDCx5p33_ASAP7_75t_R g1998 ( 
.A(n_1802),
.Y(n_1998)
);

CKINVDCx5p33_ASAP7_75t_R g1999 ( 
.A(n_1814),
.Y(n_1999)
);

CKINVDCx20_ASAP7_75t_R g2000 ( 
.A(n_1822),
.Y(n_2000)
);

CKINVDCx5p33_ASAP7_75t_R g2001 ( 
.A(n_1827),
.Y(n_2001)
);

CKINVDCx20_ASAP7_75t_R g2002 ( 
.A(n_1836),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1841),
.Y(n_2003)
);

INVxp67_ASAP7_75t_L g2004 ( 
.A(n_1821),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1789),
.Y(n_2005)
);

CKINVDCx20_ASAP7_75t_R g2006 ( 
.A(n_1789),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1789),
.Y(n_2007)
);

CKINVDCx5p33_ASAP7_75t_R g2008 ( 
.A(n_1826),
.Y(n_2008)
);

CKINVDCx5p33_ASAP7_75t_R g2009 ( 
.A(n_1826),
.Y(n_2009)
);

CKINVDCx20_ASAP7_75t_R g2010 ( 
.A(n_1741),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1768),
.Y(n_2011)
);

HB1xp67_ASAP7_75t_L g2012 ( 
.A(n_1818),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_1826),
.Y(n_2013)
);

CKINVDCx5p33_ASAP7_75t_R g2014 ( 
.A(n_1826),
.Y(n_2014)
);

BUFx10_ASAP7_75t_L g2015 ( 
.A(n_1780),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1768),
.Y(n_2016)
);

CKINVDCx5p33_ASAP7_75t_R g2017 ( 
.A(n_1826),
.Y(n_2017)
);

CKINVDCx5p33_ASAP7_75t_R g2018 ( 
.A(n_1826),
.Y(n_2018)
);

NOR2xp67_ASAP7_75t_L g2019 ( 
.A(n_1803),
.B(n_1252),
.Y(n_2019)
);

CKINVDCx5p33_ASAP7_75t_R g2020 ( 
.A(n_1826),
.Y(n_2020)
);

INVxp67_ASAP7_75t_SL g2021 ( 
.A(n_1818),
.Y(n_2021)
);

CKINVDCx5p33_ASAP7_75t_R g2022 ( 
.A(n_1826),
.Y(n_2022)
);

INVx3_ASAP7_75t_L g2023 ( 
.A(n_1768),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1768),
.Y(n_2024)
);

INVxp67_ASAP7_75t_SL g2025 ( 
.A(n_1818),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_1826),
.Y(n_2026)
);

CKINVDCx20_ASAP7_75t_R g2027 ( 
.A(n_1741),
.Y(n_2027)
);

BUFx6f_ASAP7_75t_SL g2028 ( 
.A(n_1734),
.Y(n_2028)
);

CKINVDCx5p33_ASAP7_75t_R g2029 ( 
.A(n_1826),
.Y(n_2029)
);

CKINVDCx5p33_ASAP7_75t_R g2030 ( 
.A(n_1826),
.Y(n_2030)
);

CKINVDCx5p33_ASAP7_75t_R g2031 ( 
.A(n_1826),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1768),
.Y(n_2032)
);

HB1xp67_ASAP7_75t_L g2033 ( 
.A(n_1818),
.Y(n_2033)
);

CKINVDCx5p33_ASAP7_75t_R g2034 ( 
.A(n_1826),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1768),
.Y(n_2035)
);

CKINVDCx20_ASAP7_75t_R g2036 ( 
.A(n_1741),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1768),
.Y(n_2037)
);

NOR2xp33_ASAP7_75t_L g2038 ( 
.A(n_1803),
.B(n_1707),
.Y(n_2038)
);

CKINVDCx16_ASAP7_75t_R g2039 ( 
.A(n_1826),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1768),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1768),
.Y(n_2041)
);

CKINVDCx20_ASAP7_75t_R g2042 ( 
.A(n_1741),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1768),
.Y(n_2043)
);

CKINVDCx20_ASAP7_75t_R g2044 ( 
.A(n_1741),
.Y(n_2044)
);

CKINVDCx20_ASAP7_75t_R g2045 ( 
.A(n_1741),
.Y(n_2045)
);

CKINVDCx20_ASAP7_75t_R g2046 ( 
.A(n_1741),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1768),
.Y(n_2047)
);

CKINVDCx5p33_ASAP7_75t_R g2048 ( 
.A(n_1826),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1768),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1768),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1768),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1768),
.Y(n_2052)
);

CKINVDCx5p33_ASAP7_75t_R g2053 ( 
.A(n_1826),
.Y(n_2053)
);

CKINVDCx5p33_ASAP7_75t_R g2054 ( 
.A(n_1826),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_1826),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1768),
.Y(n_2056)
);

INVxp67_ASAP7_75t_SL g2057 ( 
.A(n_1818),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1768),
.Y(n_2058)
);

CKINVDCx5p33_ASAP7_75t_R g2059 ( 
.A(n_1826),
.Y(n_2059)
);

CKINVDCx20_ASAP7_75t_R g2060 ( 
.A(n_1741),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1728),
.Y(n_2061)
);

CKINVDCx5p33_ASAP7_75t_R g2062 ( 
.A(n_1826),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1768),
.Y(n_2063)
);

CKINVDCx20_ASAP7_75t_R g2064 ( 
.A(n_1741),
.Y(n_2064)
);

CKINVDCx5p33_ASAP7_75t_R g2065 ( 
.A(n_1826),
.Y(n_2065)
);

CKINVDCx20_ASAP7_75t_R g2066 ( 
.A(n_1741),
.Y(n_2066)
);

CKINVDCx5p33_ASAP7_75t_R g2067 ( 
.A(n_1826),
.Y(n_2067)
);

BUFx6f_ASAP7_75t_L g2068 ( 
.A(n_1789),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1768),
.Y(n_2069)
);

CKINVDCx5p33_ASAP7_75t_R g2070 ( 
.A(n_1826),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1768),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1768),
.Y(n_2072)
);

CKINVDCx16_ASAP7_75t_R g2073 ( 
.A(n_1826),
.Y(n_2073)
);

CKINVDCx16_ASAP7_75t_R g2074 ( 
.A(n_1826),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1768),
.Y(n_2075)
);

INVx1_ASAP7_75t_SL g2076 ( 
.A(n_1818),
.Y(n_2076)
);

HB1xp67_ASAP7_75t_L g2077 ( 
.A(n_1818),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1768),
.Y(n_2078)
);

CKINVDCx5p33_ASAP7_75t_R g2079 ( 
.A(n_1826),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1768),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1768),
.Y(n_2081)
);

NOR2xp33_ASAP7_75t_L g2082 ( 
.A(n_1803),
.B(n_1078),
.Y(n_2082)
);

CKINVDCx20_ASAP7_75t_R g2083 ( 
.A(n_1741),
.Y(n_2083)
);

CKINVDCx20_ASAP7_75t_R g2084 ( 
.A(n_1741),
.Y(n_2084)
);

CKINVDCx20_ASAP7_75t_R g2085 ( 
.A(n_1741),
.Y(n_2085)
);

CKINVDCx5p33_ASAP7_75t_R g2086 ( 
.A(n_1826),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1768),
.Y(n_2087)
);

CKINVDCx5p33_ASAP7_75t_R g2088 ( 
.A(n_2076),
.Y(n_2088)
);

AOI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_1963),
.A2(n_1080),
.B1(n_1081),
.B2(n_1079),
.Y(n_2089)
);

BUFx6f_ASAP7_75t_L g2090 ( 
.A(n_1881),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1900),
.Y(n_2091)
);

OAI21x1_ASAP7_75t_L g2092 ( 
.A1(n_1900),
.A2(n_1155),
.B(n_1148),
.Y(n_2092)
);

AND2x4_ASAP7_75t_L g2093 ( 
.A(n_1948),
.B(n_1105),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1862),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_2012),
.B(n_1122),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2033),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2077),
.Y(n_2097)
);

BUFx2_ASAP7_75t_L g2098 ( 
.A(n_1865),
.Y(n_2098)
);

NOR2xp33_ASAP7_75t_L g2099 ( 
.A(n_1940),
.B(n_1946),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_1866),
.B(n_1122),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1971),
.B(n_1683),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_2061),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1898),
.Y(n_2103)
);

AND2x4_ASAP7_75t_L g2104 ( 
.A(n_2021),
.B(n_1404),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1903),
.Y(n_2105)
);

BUFx8_ASAP7_75t_L g2106 ( 
.A(n_1879),
.Y(n_2106)
);

BUFx3_ASAP7_75t_L g2107 ( 
.A(n_2006),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_1866),
.B(n_1122),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2025),
.B(n_1206),
.Y(n_2109)
);

NAND2xp33_ASAP7_75t_R g2110 ( 
.A(n_1925),
.B(n_1083),
.Y(n_2110)
);

CKINVDCx16_ASAP7_75t_R g2111 ( 
.A(n_1864),
.Y(n_2111)
);

CKINVDCx5p33_ASAP7_75t_R g2112 ( 
.A(n_2039),
.Y(n_2112)
);

INVx4_ASAP7_75t_L g2113 ( 
.A(n_1879),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1905),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_1980),
.B(n_1683),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_1994),
.B(n_1084),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1907),
.Y(n_2117)
);

CKINVDCx20_ASAP7_75t_R g2118 ( 
.A(n_1859),
.Y(n_2118)
);

INVx3_ASAP7_75t_L g2119 ( 
.A(n_2023),
.Y(n_2119)
);

OAI22xp5_ASAP7_75t_SL g2120 ( 
.A1(n_1887),
.A2(n_1138),
.B1(n_1158),
.B2(n_1137),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_2057),
.B(n_1085),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1910),
.Y(n_2122)
);

CKINVDCx20_ASAP7_75t_R g2123 ( 
.A(n_1890),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1914),
.Y(n_2124)
);

INVx3_ASAP7_75t_L g2125 ( 
.A(n_2023),
.Y(n_2125)
);

CKINVDCx20_ASAP7_75t_R g2126 ( 
.A(n_1892),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_1916),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1891),
.B(n_1086),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1878),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1922),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_1894),
.B(n_1919),
.Y(n_2131)
);

CKINVDCx5p33_ASAP7_75t_R g2132 ( 
.A(n_2073),
.Y(n_2132)
);

BUFx6f_ASAP7_75t_L g2133 ( 
.A(n_2015),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1909),
.B(n_1087),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_SL g2135 ( 
.A(n_1969),
.B(n_1206),
.Y(n_2135)
);

CKINVDCx5p33_ASAP7_75t_R g2136 ( 
.A(n_2074),
.Y(n_2136)
);

HB1xp67_ASAP7_75t_L g2137 ( 
.A(n_1964),
.Y(n_2137)
);

INVx2_ASAP7_75t_SL g2138 ( 
.A(n_1932),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1923),
.Y(n_2139)
);

BUFx6f_ASAP7_75t_L g2140 ( 
.A(n_2015),
.Y(n_2140)
);

NOR2x1_ASAP7_75t_L g2141 ( 
.A(n_1926),
.B(n_1270),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_1959),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1960),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1961),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_1962),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1861),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_1863),
.Y(n_2147)
);

CKINVDCx5p33_ASAP7_75t_R g2148 ( 
.A(n_2028),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_1978),
.B(n_1206),
.Y(n_2149)
);

BUFx6f_ASAP7_75t_L g2150 ( 
.A(n_2008),
.Y(n_2150)
);

AND2x4_ASAP7_75t_L g2151 ( 
.A(n_1940),
.B(n_1714),
.Y(n_2151)
);

HB1xp67_ASAP7_75t_L g2152 ( 
.A(n_1968),
.Y(n_2152)
);

AND2x4_ASAP7_75t_L g2153 ( 
.A(n_2009),
.B(n_1137),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1930),
.Y(n_2154)
);

AND2x4_ASAP7_75t_L g2155 ( 
.A(n_2013),
.B(n_1138),
.Y(n_2155)
);

BUFx2_ASAP7_75t_L g2156 ( 
.A(n_1972),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1933),
.Y(n_2157)
);

BUFx8_ASAP7_75t_L g2158 ( 
.A(n_2028),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1943),
.Y(n_2159)
);

OA21x2_ASAP7_75t_L g2160 ( 
.A1(n_1997),
.A2(n_1204),
.B(n_1191),
.Y(n_2160)
);

AOI22x1_ASAP7_75t_SL g2161 ( 
.A1(n_1893),
.A2(n_1183),
.B1(n_1190),
.B2(n_1158),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1951),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1952),
.Y(n_2163)
);

OAI22xp5_ASAP7_75t_SL g2164 ( 
.A1(n_1911),
.A2(n_2010),
.B1(n_2036),
.B2(n_2027),
.Y(n_2164)
);

CKINVDCx20_ASAP7_75t_R g2165 ( 
.A(n_2042),
.Y(n_2165)
);

BUFx2_ASAP7_75t_L g2166 ( 
.A(n_1987),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_1867),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_1883),
.B(n_1088),
.Y(n_2168)
);

AND2x4_ASAP7_75t_L g2169 ( 
.A(n_2014),
.B(n_2017),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1953),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1873),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1874),
.Y(n_2172)
);

INVx6_ASAP7_75t_L g2173 ( 
.A(n_1950),
.Y(n_2173)
);

NOR2xp33_ASAP7_75t_L g2174 ( 
.A(n_1946),
.B(n_1090),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1875),
.Y(n_2175)
);

OA21x2_ASAP7_75t_L g2176 ( 
.A1(n_2003),
.A2(n_1229),
.B(n_1222),
.Y(n_2176)
);

BUFx8_ASAP7_75t_L g2177 ( 
.A(n_1924),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_1888),
.B(n_1889),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1882),
.Y(n_2179)
);

HB1xp67_ASAP7_75t_L g2180 ( 
.A(n_1988),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1880),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1984),
.Y(n_2182)
);

BUFx6f_ASAP7_75t_L g2183 ( 
.A(n_2018),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_1897),
.B(n_1091),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_1868),
.B(n_1207),
.Y(n_2185)
);

AND2x4_ASAP7_75t_L g2186 ( 
.A(n_2020),
.B(n_1183),
.Y(n_2186)
);

CKINVDCx5p33_ASAP7_75t_R g2187 ( 
.A(n_1895),
.Y(n_2187)
);

AND2x4_ASAP7_75t_L g2188 ( 
.A(n_2022),
.B(n_1190),
.Y(n_2188)
);

INVx3_ASAP7_75t_L g2189 ( 
.A(n_2026),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1917),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1920),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_1976),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1921),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2082),
.B(n_1092),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2019),
.Y(n_2195)
);

AND2x4_ASAP7_75t_L g2196 ( 
.A(n_2029),
.B(n_1221),
.Y(n_2196)
);

OAI22xp5_ASAP7_75t_SL g2197 ( 
.A1(n_2044),
.A2(n_1223),
.B1(n_1226),
.B2(n_1221),
.Y(n_2197)
);

BUFx6f_ASAP7_75t_L g2198 ( 
.A(n_2030),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_1970),
.B(n_1098),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_1860),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_1868),
.B(n_1207),
.Y(n_2201)
);

CKINVDCx5p33_ASAP7_75t_R g2202 ( 
.A(n_2031),
.Y(n_2202)
);

INVx3_ASAP7_75t_L g2203 ( 
.A(n_2034),
.Y(n_2203)
);

CKINVDCx5p33_ASAP7_75t_R g2204 ( 
.A(n_2048),
.Y(n_2204)
);

AND2x4_ASAP7_75t_L g2205 ( 
.A(n_1973),
.B(n_2004),
.Y(n_2205)
);

INVx3_ASAP7_75t_L g2206 ( 
.A(n_2053),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2011),
.Y(n_2207)
);

CKINVDCx16_ASAP7_75t_R g2208 ( 
.A(n_1990),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1974),
.Y(n_2209)
);

BUFx8_ASAP7_75t_L g2210 ( 
.A(n_2045),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2016),
.Y(n_2211)
);

INVxp67_ASAP7_75t_L g2212 ( 
.A(n_1877),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_2024),
.Y(n_2213)
);

INVx3_ASAP7_75t_L g2214 ( 
.A(n_2054),
.Y(n_2214)
);

NOR2xp33_ASAP7_75t_L g2215 ( 
.A(n_1929),
.B(n_1099),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_1975),
.B(n_1207),
.Y(n_2216)
);

CKINVDCx20_ASAP7_75t_R g2217 ( 
.A(n_2046),
.Y(n_2217)
);

CKINVDCx20_ASAP7_75t_R g2218 ( 
.A(n_2060),
.Y(n_2218)
);

BUFx2_ASAP7_75t_L g2219 ( 
.A(n_1991),
.Y(n_2219)
);

INVx3_ASAP7_75t_L g2220 ( 
.A(n_2055),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1983),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_1993),
.B(n_1100),
.Y(n_2222)
);

CKINVDCx5p33_ASAP7_75t_R g2223 ( 
.A(n_2059),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1979),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1981),
.Y(n_2225)
);

AOI22xp5_ASAP7_75t_L g2226 ( 
.A1(n_1937),
.A2(n_1108),
.B1(n_1109),
.B2(n_1107),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_2032),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_1982),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_2035),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1985),
.Y(n_2230)
);

BUFx6f_ASAP7_75t_L g2231 ( 
.A(n_2062),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_2037),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_2040),
.Y(n_2233)
);

CKINVDCx5p33_ASAP7_75t_R g2234 ( 
.A(n_2065),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1986),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1989),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_SL g2237 ( 
.A(n_1947),
.B(n_1218),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2041),
.Y(n_2238)
);

BUFx8_ASAP7_75t_L g2239 ( 
.A(n_2064),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_1965),
.B(n_1110),
.Y(n_2240)
);

BUFx12f_ASAP7_75t_L g2241 ( 
.A(n_1931),
.Y(n_2241)
);

NAND2xp33_ASAP7_75t_L g2242 ( 
.A(n_2067),
.B(n_1159),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2043),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2047),
.Y(n_2244)
);

BUFx6f_ASAP7_75t_L g2245 ( 
.A(n_2070),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2049),
.Y(n_2246)
);

INVx3_ASAP7_75t_L g2247 ( 
.A(n_2079),
.Y(n_2247)
);

BUFx6f_ASAP7_75t_L g2248 ( 
.A(n_2086),
.Y(n_2248)
);

CKINVDCx5p33_ASAP7_75t_R g2249 ( 
.A(n_2066),
.Y(n_2249)
);

INVxp67_ASAP7_75t_L g2250 ( 
.A(n_1886),
.Y(n_2250)
);

OA21x2_ASAP7_75t_L g2251 ( 
.A1(n_1977),
.A2(n_1235),
.B(n_1232),
.Y(n_2251)
);

OAI22xp5_ASAP7_75t_L g2252 ( 
.A1(n_1992),
.A2(n_1116),
.B1(n_1118),
.B2(n_1112),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2050),
.Y(n_2253)
);

NAND2xp33_ASAP7_75t_L g2254 ( 
.A(n_1949),
.B(n_1159),
.Y(n_2254)
);

HB1xp67_ASAP7_75t_L g2255 ( 
.A(n_1996),
.Y(n_2255)
);

CKINVDCx5p33_ASAP7_75t_R g2256 ( 
.A(n_2083),
.Y(n_2256)
);

AND2x2_ASAP7_75t_L g2257 ( 
.A(n_1899),
.B(n_1218),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_2051),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2052),
.Y(n_2259)
);

AND2x4_ASAP7_75t_L g2260 ( 
.A(n_1915),
.B(n_1223),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2056),
.Y(n_2261)
);

OAI22xp5_ASAP7_75t_L g2262 ( 
.A1(n_1954),
.A2(n_1121),
.B1(n_1123),
.B2(n_1120),
.Y(n_2262)
);

INVx1_ASAP7_75t_SL g2263 ( 
.A(n_1869),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_2058),
.Y(n_2264)
);

CKINVDCx5p33_ASAP7_75t_R g2265 ( 
.A(n_2084),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2063),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2069),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_1966),
.B(n_1125),
.Y(n_2268)
);

AND2x4_ASAP7_75t_L g2269 ( 
.A(n_1956),
.B(n_1226),
.Y(n_2269)
);

OA21x2_ASAP7_75t_L g2270 ( 
.A1(n_1995),
.A2(n_1245),
.B(n_1240),
.Y(n_2270)
);

CKINVDCx20_ASAP7_75t_R g2271 ( 
.A(n_2085),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2071),
.Y(n_2272)
);

HB1xp67_ASAP7_75t_L g2273 ( 
.A(n_1870),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2072),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2075),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2078),
.Y(n_2276)
);

INVx3_ASAP7_75t_L g2277 ( 
.A(n_2080),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_1967),
.B(n_1127),
.Y(n_2278)
);

AND2x4_ASAP7_75t_L g2279 ( 
.A(n_2004),
.B(n_1270),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_2081),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2087),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_1998),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_1999),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_1957),
.Y(n_2284)
);

BUFx6f_ASAP7_75t_L g2285 ( 
.A(n_1871),
.Y(n_2285)
);

BUFx6f_ASAP7_75t_L g2286 ( 
.A(n_1872),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_2038),
.B(n_1129),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1958),
.Y(n_2288)
);

HB1xp67_ASAP7_75t_L g2289 ( 
.A(n_1876),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2000),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2002),
.Y(n_2291)
);

INVxp67_ASAP7_75t_L g2292 ( 
.A(n_1884),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1942),
.Y(n_2293)
);

AND2x4_ASAP7_75t_L g2294 ( 
.A(n_1955),
.B(n_1300),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_2001),
.B(n_1130),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_1901),
.Y(n_2296)
);

INVx4_ASAP7_75t_L g2297 ( 
.A(n_1885),
.Y(n_2297)
);

BUFx6f_ASAP7_75t_L g2298 ( 
.A(n_1896),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_2005),
.Y(n_2299)
);

AND2x4_ASAP7_75t_L g2300 ( 
.A(n_1927),
.B(n_1238),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_1939),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_1941),
.B(n_1132),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_1934),
.B(n_1136),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_1935),
.B(n_1141),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_1936),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_1945),
.B(n_1218),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2007),
.Y(n_2307)
);

AOI22xp5_ASAP7_75t_L g2308 ( 
.A1(n_1928),
.A2(n_1145),
.B1(n_1149),
.B2(n_1144),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2068),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2068),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_1938),
.B(n_1152),
.Y(n_2311)
);

INVx3_ASAP7_75t_L g2312 ( 
.A(n_1902),
.Y(n_2312)
);

CKINVDCx8_ASAP7_75t_R g2313 ( 
.A(n_1904),
.Y(n_2313)
);

BUFx6f_ASAP7_75t_L g2314 ( 
.A(n_2068),
.Y(n_2314)
);

BUFx6f_ASAP7_75t_L g2315 ( 
.A(n_2068),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_1944),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_1906),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_1908),
.Y(n_2318)
);

BUFx2_ASAP7_75t_L g2319 ( 
.A(n_1913),
.Y(n_2319)
);

NOR2xp33_ASAP7_75t_L g2320 ( 
.A(n_1918),
.B(n_1153),
.Y(n_2320)
);

INVx2_ASAP7_75t_L g2321 ( 
.A(n_1912),
.Y(n_2321)
);

CKINVDCx8_ASAP7_75t_R g2322 ( 
.A(n_1864),
.Y(n_2322)
);

BUFx2_ASAP7_75t_L g2323 ( 
.A(n_1862),
.Y(n_2323)
);

XNOR2xp5_ASAP7_75t_L g2324 ( 
.A(n_1859),
.B(n_1238),
.Y(n_2324)
);

INVx3_ASAP7_75t_L g2325 ( 
.A(n_2076),
.Y(n_2325)
);

OAI22xp5_ASAP7_75t_L g2326 ( 
.A1(n_2076),
.A2(n_1162),
.B1(n_1163),
.B2(n_1154),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_1900),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_1971),
.B(n_1165),
.Y(n_2328)
);

NOR2x1_ASAP7_75t_L g2329 ( 
.A(n_1881),
.B(n_1300),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_1900),
.Y(n_2330)
);

AOI22xp5_ASAP7_75t_L g2331 ( 
.A1(n_1963),
.A2(n_1170),
.B1(n_1171),
.B2(n_1166),
.Y(n_2331)
);

CKINVDCx5p33_ASAP7_75t_R g2332 ( 
.A(n_2076),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_1900),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_1900),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_1900),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_1900),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_1971),
.B(n_1172),
.Y(n_2337)
);

AND2x4_ASAP7_75t_L g2338 ( 
.A(n_2076),
.B(n_1304),
.Y(n_2338)
);

OA21x2_ASAP7_75t_L g2339 ( 
.A1(n_1997),
.A2(n_1255),
.B(n_1249),
.Y(n_2339)
);

BUFx6f_ASAP7_75t_L g2340 ( 
.A(n_1881),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_1900),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_1900),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_1900),
.Y(n_2343)
);

AND2x4_ASAP7_75t_L g2344 ( 
.A(n_2076),
.B(n_1304),
.Y(n_2344)
);

CKINVDCx20_ASAP7_75t_R g2345 ( 
.A(n_2076),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_1900),
.Y(n_2346)
);

INVx5_ASAP7_75t_L g2347 ( 
.A(n_2023),
.Y(n_2347)
);

CKINVDCx5p33_ASAP7_75t_R g2348 ( 
.A(n_2076),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_1900),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_1900),
.Y(n_2350)
);

AND2x4_ASAP7_75t_L g2351 ( 
.A(n_2076),
.B(n_1364),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_1900),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_1900),
.Y(n_2353)
);

CKINVDCx6p67_ASAP7_75t_R g2354 ( 
.A(n_1879),
.Y(n_2354)
);

OA21x2_ASAP7_75t_L g2355 ( 
.A1(n_1997),
.A2(n_1258),
.B(n_1257),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_1900),
.Y(n_2356)
);

CKINVDCx16_ASAP7_75t_R g2357 ( 
.A(n_1864),
.Y(n_2357)
);

HB1xp67_ASAP7_75t_L g2358 ( 
.A(n_2076),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_1900),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_1900),
.Y(n_2360)
);

CKINVDCx20_ASAP7_75t_R g2361 ( 
.A(n_2076),
.Y(n_2361)
);

AND2x4_ASAP7_75t_L g2362 ( 
.A(n_2076),
.B(n_1242),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_1900),
.Y(n_2363)
);

INVxp67_ASAP7_75t_L g2364 ( 
.A(n_1948),
.Y(n_2364)
);

NOR2xp33_ASAP7_75t_L g2365 ( 
.A(n_1963),
.B(n_1177),
.Y(n_2365)
);

BUFx6f_ASAP7_75t_L g2366 ( 
.A(n_1881),
.Y(n_2366)
);

BUFx6f_ASAP7_75t_L g2367 ( 
.A(n_1881),
.Y(n_2367)
);

CKINVDCx20_ASAP7_75t_R g2368 ( 
.A(n_2076),
.Y(n_2368)
);

BUFx6f_ASAP7_75t_L g2369 ( 
.A(n_1881),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_1900),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_1900),
.Y(n_2371)
);

CKINVDCx5p33_ASAP7_75t_R g2372 ( 
.A(n_2076),
.Y(n_2372)
);

INVx3_ASAP7_75t_L g2373 ( 
.A(n_2076),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_1900),
.Y(n_2374)
);

CKINVDCx5p33_ASAP7_75t_R g2375 ( 
.A(n_2076),
.Y(n_2375)
);

AND2x4_ASAP7_75t_L g2376 ( 
.A(n_2076),
.B(n_1364),
.Y(n_2376)
);

AND2x4_ASAP7_75t_L g2377 ( 
.A(n_2076),
.B(n_1474),
.Y(n_2377)
);

OAI22xp5_ASAP7_75t_L g2378 ( 
.A1(n_2076),
.A2(n_1187),
.B1(n_1192),
.B2(n_1180),
.Y(n_2378)
);

INVx4_ASAP7_75t_L g2379 ( 
.A(n_1881),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_1900),
.Y(n_2380)
);

INVxp33_ASAP7_75t_SL g2381 ( 
.A(n_2076),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_1900),
.Y(n_2382)
);

HB1xp67_ASAP7_75t_L g2383 ( 
.A(n_2076),
.Y(n_2383)
);

BUFx6f_ASAP7_75t_L g2384 ( 
.A(n_1881),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_1900),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_1900),
.Y(n_2386)
);

AOI22xp5_ASAP7_75t_L g2387 ( 
.A1(n_1963),
.A2(n_1195),
.B1(n_1196),
.B2(n_1194),
.Y(n_2387)
);

BUFx6f_ASAP7_75t_L g2388 ( 
.A(n_1881),
.Y(n_2388)
);

INVx3_ASAP7_75t_L g2389 ( 
.A(n_2076),
.Y(n_2389)
);

AND2x2_ASAP7_75t_L g2390 ( 
.A(n_1948),
.B(n_1290),
.Y(n_2390)
);

BUFx3_ASAP7_75t_L g2391 ( 
.A(n_2076),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_1900),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_1948),
.B(n_1290),
.Y(n_2393)
);

CKINVDCx20_ASAP7_75t_R g2394 ( 
.A(n_2076),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_1900),
.Y(n_2395)
);

CKINVDCx5p33_ASAP7_75t_R g2396 ( 
.A(n_2076),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_1900),
.Y(n_2397)
);

CKINVDCx5p33_ASAP7_75t_R g2398 ( 
.A(n_2076),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_2092),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_2327),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_2335),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_2341),
.Y(n_2402)
);

BUFx2_ASAP7_75t_L g2403 ( 
.A(n_2345),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_2099),
.B(n_1198),
.Y(n_2404)
);

INVxp33_ASAP7_75t_SL g2405 ( 
.A(n_2088),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2251),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2251),
.Y(n_2407)
);

NAND2xp33_ASAP7_75t_SL g2408 ( 
.A(n_2361),
.B(n_1242),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_SL g2409 ( 
.A(n_2391),
.B(n_1199),
.Y(n_2409)
);

NOR3xp33_ASAP7_75t_L g2410 ( 
.A(n_2208),
.B(n_1093),
.C(n_1089),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_SL g2411 ( 
.A(n_2381),
.B(n_1200),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2342),
.Y(n_2412)
);

OR2x2_ASAP7_75t_L g2413 ( 
.A(n_2358),
.B(n_1134),
.Y(n_2413)
);

AND2x2_ASAP7_75t_L g2414 ( 
.A(n_2323),
.B(n_2131),
.Y(n_2414)
);

BUFx3_ASAP7_75t_L g2415 ( 
.A(n_2368),
.Y(n_2415)
);

HB1xp67_ASAP7_75t_L g2416 ( 
.A(n_2383),
.Y(n_2416)
);

AND2x2_ASAP7_75t_L g2417 ( 
.A(n_2323),
.B(n_1243),
.Y(n_2417)
);

BUFx6f_ASAP7_75t_L g2418 ( 
.A(n_2270),
.Y(n_2418)
);

OR2x2_ASAP7_75t_SL g2419 ( 
.A(n_2111),
.B(n_2357),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2346),
.Y(n_2420)
);

INVx8_ASAP7_75t_L g2421 ( 
.A(n_2394),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_SL g2422 ( 
.A(n_2325),
.B(n_2373),
.Y(n_2422)
);

AND2x4_ASAP7_75t_L g2423 ( 
.A(n_2389),
.B(n_2133),
.Y(n_2423)
);

INVx3_ASAP7_75t_L g2424 ( 
.A(n_2347),
.Y(n_2424)
);

NOR2xp33_ASAP7_75t_L g2425 ( 
.A(n_2364),
.B(n_2212),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2352),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2359),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_SL g2428 ( 
.A(n_2332),
.B(n_1202),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_2371),
.Y(n_2429)
);

NOR2xp33_ASAP7_75t_L g2430 ( 
.A(n_2250),
.B(n_1243),
.Y(n_2430)
);

AOI21x1_ASAP7_75t_L g2431 ( 
.A1(n_2307),
.A2(n_1261),
.B(n_1260),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2385),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2151),
.B(n_1203),
.Y(n_2433)
);

INVx2_ASAP7_75t_L g2434 ( 
.A(n_2386),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2146),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2147),
.Y(n_2436)
);

CKINVDCx5p33_ASAP7_75t_R g2437 ( 
.A(n_2348),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2167),
.Y(n_2438)
);

INVx1_ASAP7_75t_SL g2439 ( 
.A(n_2372),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2270),
.Y(n_2440)
);

INVx3_ASAP7_75t_L g2441 ( 
.A(n_2347),
.Y(n_2441)
);

AOI21x1_ASAP7_75t_L g2442 ( 
.A1(n_2160),
.A2(n_1272),
.B(n_1265),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2224),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2225),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_SL g2445 ( 
.A(n_2375),
.B(n_1205),
.Y(n_2445)
);

INVxp33_ASAP7_75t_L g2446 ( 
.A(n_2137),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_2091),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_2330),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_SL g2449 ( 
.A(n_2396),
.B(n_1209),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_2333),
.Y(n_2450)
);

BUFx6f_ASAP7_75t_L g2451 ( 
.A(n_2160),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2179),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2171),
.Y(n_2453)
);

NOR2xp33_ASAP7_75t_L g2454 ( 
.A(n_2138),
.B(n_1253),
.Y(n_2454)
);

NOR2xp33_ASAP7_75t_SL g2455 ( 
.A(n_2398),
.B(n_1253),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2172),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_2334),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_SL g2458 ( 
.A(n_2098),
.B(n_1210),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2336),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2175),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_2343),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2181),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_2349),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_2151),
.B(n_1212),
.Y(n_2464)
);

BUFx3_ASAP7_75t_L g2465 ( 
.A(n_2133),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2190),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2191),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_2098),
.B(n_1217),
.Y(n_2468)
);

INVx2_ASAP7_75t_L g2469 ( 
.A(n_2350),
.Y(n_2469)
);

AND2x4_ASAP7_75t_L g2470 ( 
.A(n_2140),
.B(n_1274),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2193),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_SL g2472 ( 
.A(n_2338),
.B(n_2344),
.Y(n_2472)
);

INVx3_ASAP7_75t_L g2473 ( 
.A(n_2347),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2353),
.Y(n_2474)
);

AOI21x1_ASAP7_75t_L g2475 ( 
.A1(n_2176),
.A2(n_1282),
.B(n_1277),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2356),
.Y(n_2476)
);

AOI21x1_ASAP7_75t_L g2477 ( 
.A1(n_2176),
.A2(n_1286),
.B(n_1285),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2103),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2360),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2363),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2370),
.Y(n_2481)
);

BUFx10_ASAP7_75t_L g2482 ( 
.A(n_2140),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2105),
.Y(n_2483)
);

NOR2xp33_ASAP7_75t_L g2484 ( 
.A(n_2173),
.B(n_1269),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_2374),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2114),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2117),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2380),
.Y(n_2488)
);

NOR2x1_ASAP7_75t_L g2489 ( 
.A(n_2113),
.B(n_1269),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_2382),
.Y(n_2490)
);

NOR2xp33_ASAP7_75t_L g2491 ( 
.A(n_2173),
.B(n_1273),
.Y(n_2491)
);

AND2x2_ASAP7_75t_L g2492 ( 
.A(n_2362),
.B(n_1273),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2228),
.Y(n_2493)
);

AO22x2_ASAP7_75t_L g2494 ( 
.A1(n_2161),
.A2(n_1335),
.B1(n_1352),
.B2(n_1318),
.Y(n_2494)
);

CKINVDCx5p33_ASAP7_75t_R g2495 ( 
.A(n_2177),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2392),
.Y(n_2496)
);

OR2x6_ASAP7_75t_L g2497 ( 
.A(n_2241),
.B(n_1530),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_SL g2498 ( 
.A(n_2338),
.B(n_1219),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_2395),
.Y(n_2499)
);

INVx2_ASAP7_75t_L g2500 ( 
.A(n_2397),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2230),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2142),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2143),
.Y(n_2503)
);

CKINVDCx5p33_ASAP7_75t_R g2504 ( 
.A(n_2210),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_2144),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2235),
.Y(n_2506)
);

NOR2xp33_ASAP7_75t_L g2507 ( 
.A(n_2302),
.B(n_1318),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2145),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_2127),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2200),
.Y(n_2510)
);

INVxp33_ASAP7_75t_SL g2511 ( 
.A(n_2187),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2207),
.Y(n_2512)
);

NOR2xp33_ASAP7_75t_L g2513 ( 
.A(n_2100),
.B(n_1335),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2211),
.Y(n_2514)
);

BUFx3_ASAP7_75t_L g2515 ( 
.A(n_2106),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_SL g2516 ( 
.A(n_2344),
.B(n_1224),
.Y(n_2516)
);

INVx2_ASAP7_75t_L g2517 ( 
.A(n_2213),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2109),
.B(n_1225),
.Y(n_2518)
);

INVxp33_ASAP7_75t_SL g2519 ( 
.A(n_2324),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2236),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2227),
.Y(n_2521)
);

NAND2xp5_ASAP7_75t_SL g2522 ( 
.A(n_2351),
.B(n_1227),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2122),
.Y(n_2523)
);

INVx2_ASAP7_75t_L g2524 ( 
.A(n_2229),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2124),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2232),
.Y(n_2526)
);

INVx8_ASAP7_75t_L g2527 ( 
.A(n_2090),
.Y(n_2527)
);

INVx8_ASAP7_75t_L g2528 ( 
.A(n_2090),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_SL g2529 ( 
.A(n_2351),
.B(n_1231),
.Y(n_2529)
);

INVx2_ASAP7_75t_SL g2530 ( 
.A(n_2376),
.Y(n_2530)
);

NAND2xp33_ASAP7_75t_L g2531 ( 
.A(n_2108),
.B(n_1234),
.Y(n_2531)
);

INVx2_ASAP7_75t_SL g2532 ( 
.A(n_2376),
.Y(n_2532)
);

INVx3_ASAP7_75t_L g2533 ( 
.A(n_2192),
.Y(n_2533)
);

INVx3_ASAP7_75t_L g2534 ( 
.A(n_2119),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2130),
.Y(n_2535)
);

OR2x2_ASAP7_75t_L g2536 ( 
.A(n_2269),
.B(n_1173),
.Y(n_2536)
);

INVxp33_ASAP7_75t_L g2537 ( 
.A(n_2324),
.Y(n_2537)
);

NOR2xp33_ASAP7_75t_L g2538 ( 
.A(n_2185),
.B(n_1352),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2233),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2139),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2258),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2264),
.Y(n_2542)
);

AOI21x1_ASAP7_75t_L g2543 ( 
.A1(n_2339),
.A2(n_1309),
.B(n_1302),
.Y(n_2543)
);

AND3x2_ASAP7_75t_L g2544 ( 
.A(n_2319),
.B(n_1418),
.C(n_1412),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_L g2545 ( 
.A(n_2293),
.B(n_1236),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2280),
.Y(n_2546)
);

INVx3_ASAP7_75t_L g2547 ( 
.A(n_2125),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2104),
.B(n_1237),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2154),
.Y(n_2549)
);

BUFx2_ASAP7_75t_L g2550 ( 
.A(n_2156),
.Y(n_2550)
);

INVx2_ASAP7_75t_SL g2551 ( 
.A(n_2377),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2102),
.Y(n_2552)
);

AO21x2_ASAP7_75t_L g2553 ( 
.A1(n_2101),
.A2(n_1326),
.B(n_1314),
.Y(n_2553)
);

AND2x2_ASAP7_75t_L g2554 ( 
.A(n_2365),
.B(n_1412),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2104),
.B(n_1239),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2377),
.B(n_1244),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2157),
.Y(n_2557)
);

INVxp67_ASAP7_75t_SL g2558 ( 
.A(n_2107),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_2296),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2301),
.Y(n_2560)
);

INVx3_ASAP7_75t_L g2561 ( 
.A(n_2277),
.Y(n_2561)
);

BUFx10_ASAP7_75t_L g2562 ( 
.A(n_2169),
.Y(n_2562)
);

INVx3_ASAP7_75t_L g2563 ( 
.A(n_2129),
.Y(n_2563)
);

BUFx10_ASAP7_75t_L g2564 ( 
.A(n_2285),
.Y(n_2564)
);

INVx2_ASAP7_75t_L g2565 ( 
.A(n_2339),
.Y(n_2565)
);

INVx2_ASAP7_75t_L g2566 ( 
.A(n_2355),
.Y(n_2566)
);

CKINVDCx5p33_ASAP7_75t_R g2567 ( 
.A(n_2239),
.Y(n_2567)
);

NOR2xp33_ASAP7_75t_L g2568 ( 
.A(n_2201),
.B(n_1418),
.Y(n_2568)
);

AOI21x1_ASAP7_75t_L g2569 ( 
.A1(n_2355),
.A2(n_1332),
.B(n_1330),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2159),
.Y(n_2570)
);

BUFx6f_ASAP7_75t_L g2571 ( 
.A(n_2314),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2162),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2163),
.Y(n_2573)
);

NOR2x1p5_ASAP7_75t_L g2574 ( 
.A(n_2354),
.B(n_1246),
.Y(n_2574)
);

AND3x2_ASAP7_75t_L g2575 ( 
.A(n_2319),
.B(n_1426),
.C(n_1425),
.Y(n_2575)
);

NOR2xp33_ASAP7_75t_L g2576 ( 
.A(n_2094),
.B(n_1425),
.Y(n_2576)
);

INVx2_ASAP7_75t_L g2577 ( 
.A(n_2238),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_2243),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2095),
.B(n_1426),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2244),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2246),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_2253),
.Y(n_2582)
);

AND2x2_ASAP7_75t_L g2583 ( 
.A(n_2294),
.B(n_1432),
.Y(n_2583)
);

OR2x6_ASAP7_75t_L g2584 ( 
.A(n_2297),
.B(n_1474),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2170),
.Y(n_2585)
);

AOI21x1_ASAP7_75t_L g2586 ( 
.A1(n_2115),
.A2(n_1343),
.B(n_1333),
.Y(n_2586)
);

INVx5_ASAP7_75t_L g2587 ( 
.A(n_2340),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2259),
.Y(n_2588)
);

CKINVDCx6p67_ASAP7_75t_R g2589 ( 
.A(n_2118),
.Y(n_2589)
);

OR2x2_ASAP7_75t_L g2590 ( 
.A(n_2093),
.B(n_1182),
.Y(n_2590)
);

INVx2_ASAP7_75t_L g2591 ( 
.A(n_2261),
.Y(n_2591)
);

INVx3_ASAP7_75t_L g2592 ( 
.A(n_2266),
.Y(n_2592)
);

INVxp33_ASAP7_75t_SL g2593 ( 
.A(n_2263),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_SL g2594 ( 
.A(n_2216),
.B(n_1247),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_2267),
.Y(n_2595)
);

BUFx10_ASAP7_75t_L g2596 ( 
.A(n_2285),
.Y(n_2596)
);

OR2x2_ASAP7_75t_L g2597 ( 
.A(n_2156),
.B(n_1193),
.Y(n_2597)
);

AND2x2_ASAP7_75t_L g2598 ( 
.A(n_2294),
.B(n_1432),
.Y(n_2598)
);

INVx3_ASAP7_75t_L g2599 ( 
.A(n_2272),
.Y(n_2599)
);

INVxp33_ASAP7_75t_L g2600 ( 
.A(n_2152),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2174),
.B(n_1250),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2274),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2275),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2276),
.Y(n_2604)
);

BUFx6f_ASAP7_75t_SL g2605 ( 
.A(n_2150),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2281),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2182),
.Y(n_2607)
);

AOI21x1_ASAP7_75t_L g2608 ( 
.A1(n_2309),
.A2(n_1353),
.B(n_1350),
.Y(n_2608)
);

XOR2x2_ASAP7_75t_L g2609 ( 
.A(n_2164),
.B(n_2120),
.Y(n_2609)
);

NOR2xp33_ASAP7_75t_L g2610 ( 
.A(n_2096),
.B(n_1515),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_2195),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_2299),
.Y(n_2612)
);

AND2x2_ASAP7_75t_L g2613 ( 
.A(n_2390),
.B(n_1515),
.Y(n_2613)
);

INVx2_ASAP7_75t_L g2614 ( 
.A(n_2141),
.Y(n_2614)
);

INVx2_ASAP7_75t_L g2615 ( 
.A(n_2178),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2240),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2268),
.Y(n_2617)
);

AO21x2_ASAP7_75t_L g2618 ( 
.A1(n_2194),
.A2(n_1359),
.B(n_1356),
.Y(n_2618)
);

INVx2_ASAP7_75t_L g2619 ( 
.A(n_2279),
.Y(n_2619)
);

INVxp67_ASAP7_75t_L g2620 ( 
.A(n_2180),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_SL g2621 ( 
.A(n_2328),
.B(n_1251),
.Y(n_2621)
);

NOR2xp33_ASAP7_75t_L g2622 ( 
.A(n_2097),
.B(n_1516),
.Y(n_2622)
);

BUFx2_ASAP7_75t_L g2623 ( 
.A(n_2166),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_2279),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2278),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2168),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2257),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_L g2628 ( 
.A(n_2337),
.B(n_1256),
.Y(n_2628)
);

INVx3_ASAP7_75t_L g2629 ( 
.A(n_2340),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2314),
.Y(n_2630)
);

INVx2_ASAP7_75t_L g2631 ( 
.A(n_2315),
.Y(n_2631)
);

INVx2_ASAP7_75t_SL g2632 ( 
.A(n_2366),
.Y(n_2632)
);

BUFx2_ASAP7_75t_L g2633 ( 
.A(n_2166),
.Y(n_2633)
);

BUFx3_ASAP7_75t_L g2634 ( 
.A(n_2158),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2184),
.Y(n_2635)
);

INVx5_ASAP7_75t_L g2636 ( 
.A(n_2366),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2315),
.Y(n_2637)
);

AND2x2_ASAP7_75t_L g2638 ( 
.A(n_2393),
.B(n_1516),
.Y(n_2638)
);

BUFx6f_ASAP7_75t_L g2639 ( 
.A(n_2367),
.Y(n_2639)
);

INVx2_ASAP7_75t_SL g2640 ( 
.A(n_2367),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_SL g2641 ( 
.A(n_2326),
.B(n_1259),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2329),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_2149),
.Y(n_2643)
);

OR2x2_ASAP7_75t_L g2644 ( 
.A(n_2219),
.B(n_2255),
.Y(n_2644)
);

INVx2_ASAP7_75t_L g2645 ( 
.A(n_2205),
.Y(n_2645)
);

BUFx6f_ASAP7_75t_SL g2646 ( 
.A(n_2150),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2205),
.Y(n_2647)
);

NAND2xp5_ASAP7_75t_L g2648 ( 
.A(n_2252),
.B(n_1263),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2121),
.Y(n_2649)
);

CKINVDCx5p33_ASAP7_75t_R g2650 ( 
.A(n_2249),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2310),
.Y(n_2651)
);

INVx3_ASAP7_75t_L g2652 ( 
.A(n_2369),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_SL g2653 ( 
.A(n_2378),
.B(n_1264),
.Y(n_2653)
);

BUFx6f_ASAP7_75t_SL g2654 ( 
.A(n_2183),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2128),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2134),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_SL g2657 ( 
.A(n_2209),
.B(n_2221),
.Y(n_2657)
);

AND2x2_ASAP7_75t_L g2658 ( 
.A(n_2089),
.B(n_1519),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2215),
.B(n_1266),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2282),
.Y(n_2660)
);

INVxp67_ASAP7_75t_R g2661 ( 
.A(n_2197),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_SL g2662 ( 
.A(n_2284),
.B(n_2288),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2116),
.Y(n_2663)
);

BUFx10_ASAP7_75t_L g2664 ( 
.A(n_2286),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2254),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2283),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2287),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2295),
.Y(n_2668)
);

INVx2_ASAP7_75t_SL g2669 ( 
.A(n_2369),
.Y(n_2669)
);

NOR2xp33_ASAP7_75t_L g2670 ( 
.A(n_2199),
.B(n_1519),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2242),
.Y(n_2671)
);

INVx2_ASAP7_75t_L g2672 ( 
.A(n_2222),
.Y(n_2672)
);

NAND2xp33_ASAP7_75t_L g2673 ( 
.A(n_2384),
.B(n_1267),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_2135),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2237),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2331),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2387),
.Y(n_2677)
);

OR2x2_ASAP7_75t_L g2678 ( 
.A(n_2219),
.B(n_1213),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2226),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2384),
.Y(n_2680)
);

NOR2xp33_ASAP7_75t_L g2681 ( 
.A(n_2303),
.B(n_1523),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_2388),
.Y(n_2682)
);

AND3x2_ASAP7_75t_L g2683 ( 
.A(n_2292),
.B(n_1564),
.C(n_1523),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2262),
.B(n_2306),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2388),
.Y(n_2685)
);

NOR2xp33_ASAP7_75t_L g2686 ( 
.A(n_2304),
.B(n_1564),
.Y(n_2686)
);

AOI21x1_ASAP7_75t_L g2687 ( 
.A1(n_2260),
.A2(n_1367),
.B(n_1360),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2308),
.Y(n_2688)
);

INVx3_ASAP7_75t_L g2689 ( 
.A(n_2379),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2290),
.Y(n_2690)
);

NOR2xp33_ASAP7_75t_SL g2691 ( 
.A(n_2313),
.B(n_1571),
.Y(n_2691)
);

BUFx10_ASAP7_75t_L g2692 ( 
.A(n_2286),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2320),
.B(n_1268),
.Y(n_2693)
);

AND3x2_ASAP7_75t_L g2694 ( 
.A(n_2273),
.B(n_1584),
.C(n_1571),
.Y(n_2694)
);

INVx2_ASAP7_75t_L g2695 ( 
.A(n_2318),
.Y(n_2695)
);

INVx2_ASAP7_75t_L g2696 ( 
.A(n_2305),
.Y(n_2696)
);

INVx8_ASAP7_75t_L g2697 ( 
.A(n_2298),
.Y(n_2697)
);

AOI21x1_ASAP7_75t_L g2698 ( 
.A1(n_2311),
.A2(n_1386),
.B(n_1377),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_L g2699 ( 
.A(n_2289),
.B(n_1275),
.Y(n_2699)
);

INVx2_ASAP7_75t_L g2700 ( 
.A(n_2317),
.Y(n_2700)
);

NAND2xp33_ASAP7_75t_SL g2701 ( 
.A(n_2298),
.B(n_1584),
.Y(n_2701)
);

INVx3_ASAP7_75t_L g2702 ( 
.A(n_2183),
.Y(n_2702)
);

AND2x2_ASAP7_75t_SL g2703 ( 
.A(n_2153),
.B(n_1593),
.Y(n_2703)
);

AND2x2_ASAP7_75t_SL g2704 ( 
.A(n_2155),
.B(n_1593),
.Y(n_2704)
);

INVx2_ASAP7_75t_L g2705 ( 
.A(n_2291),
.Y(n_2705)
);

AND2x2_ASAP7_75t_L g2706 ( 
.A(n_2312),
.B(n_1596),
.Y(n_2706)
);

BUFx10_ASAP7_75t_L g2707 ( 
.A(n_2198),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_SL g2708 ( 
.A(n_2198),
.B(n_1276),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2189),
.Y(n_2709)
);

BUFx6f_ASAP7_75t_SL g2710 ( 
.A(n_2231),
.Y(n_2710)
);

BUFx3_ASAP7_75t_L g2711 ( 
.A(n_2322),
.Y(n_2711)
);

CKINVDCx16_ASAP7_75t_R g2712 ( 
.A(n_2123),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2203),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2206),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2214),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_SL g2716 ( 
.A(n_2231),
.B(n_1278),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2220),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2247),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2245),
.Y(n_2719)
);

INVx2_ASAP7_75t_L g2720 ( 
.A(n_2245),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_2248),
.Y(n_2721)
);

AO21x2_ASAP7_75t_L g2722 ( 
.A1(n_2316),
.A2(n_1407),
.B(n_1395),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2248),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2186),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2188),
.Y(n_2725)
);

INVx2_ASAP7_75t_SL g2726 ( 
.A(n_2112),
.Y(n_2726)
);

NOR2xp33_ASAP7_75t_L g2727 ( 
.A(n_2321),
.B(n_2196),
.Y(n_2727)
);

INVx2_ASAP7_75t_L g2728 ( 
.A(n_2148),
.Y(n_2728)
);

INVx5_ASAP7_75t_L g2729 ( 
.A(n_2300),
.Y(n_2729)
);

INVx3_ASAP7_75t_L g2730 ( 
.A(n_2202),
.Y(n_2730)
);

INVx8_ASAP7_75t_L g2731 ( 
.A(n_2132),
.Y(n_2731)
);

AND2x2_ASAP7_75t_L g2732 ( 
.A(n_2204),
.B(n_1596),
.Y(n_2732)
);

INVx2_ASAP7_75t_L g2733 ( 
.A(n_2136),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2223),
.Y(n_2734)
);

BUFx10_ASAP7_75t_L g2735 ( 
.A(n_2234),
.Y(n_2735)
);

BUFx10_ASAP7_75t_L g2736 ( 
.A(n_2256),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_SL g2737 ( 
.A(n_2265),
.B(n_1279),
.Y(n_2737)
);

INVx2_ASAP7_75t_L g2738 ( 
.A(n_2126),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2165),
.Y(n_2739)
);

AND2x2_ASAP7_75t_L g2740 ( 
.A(n_2110),
.B(n_1600),
.Y(n_2740)
);

CKINVDCx20_ASAP7_75t_R g2741 ( 
.A(n_2217),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_2218),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2271),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2092),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2251),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2092),
.Y(n_2746)
);

INVx3_ASAP7_75t_L g2747 ( 
.A(n_2347),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_2092),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2251),
.Y(n_2749)
);

NOR2xp33_ASAP7_75t_L g2750 ( 
.A(n_2364),
.B(n_1600),
.Y(n_2750)
);

INVx2_ASAP7_75t_L g2751 ( 
.A(n_2092),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2251),
.Y(n_2752)
);

INVx2_ASAP7_75t_SL g2753 ( 
.A(n_2391),
.Y(n_2753)
);

AND3x2_ASAP7_75t_L g2754 ( 
.A(n_2137),
.B(n_1689),
.C(n_1686),
.Y(n_2754)
);

INVx3_ASAP7_75t_L g2755 ( 
.A(n_2347),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_2092),
.Y(n_2756)
);

INVx2_ASAP7_75t_SL g2757 ( 
.A(n_2391),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_SL g2758 ( 
.A(n_2391),
.B(n_1280),
.Y(n_2758)
);

OR2x2_ASAP7_75t_L g2759 ( 
.A(n_2358),
.B(n_1214),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_SL g2760 ( 
.A(n_2391),
.B(n_1281),
.Y(n_2760)
);

NAND3xp33_ASAP7_75t_L g2761 ( 
.A(n_2365),
.B(n_1291),
.C(n_1288),
.Y(n_2761)
);

AOI21x1_ASAP7_75t_L g2762 ( 
.A1(n_2092),
.A2(n_1420),
.B(n_1419),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2251),
.Y(n_2763)
);

INVx4_ASAP7_75t_L g2764 ( 
.A(n_2133),
.Y(n_2764)
);

INVx2_ASAP7_75t_SL g2765 ( 
.A(n_2391),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2251),
.Y(n_2766)
);

INVx3_ASAP7_75t_L g2767 ( 
.A(n_2347),
.Y(n_2767)
);

INVx8_ASAP7_75t_L g2768 ( 
.A(n_2345),
.Y(n_2768)
);

INVx2_ASAP7_75t_L g2769 ( 
.A(n_2092),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2099),
.B(n_1292),
.Y(n_2770)
);

AND2x2_ASAP7_75t_L g2771 ( 
.A(n_2391),
.B(n_1686),
.Y(n_2771)
);

NOR2xp33_ASAP7_75t_L g2772 ( 
.A(n_2364),
.B(n_1689),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_SL g2773 ( 
.A(n_2391),
.B(n_1293),
.Y(n_2773)
);

OR2x2_ASAP7_75t_L g2774 ( 
.A(n_2358),
.B(n_1287),
.Y(n_2774)
);

NAND3xp33_ASAP7_75t_L g2775 ( 
.A(n_2365),
.B(n_1295),
.C(n_1294),
.Y(n_2775)
);

OR2x2_ASAP7_75t_L g2776 ( 
.A(n_2358),
.B(n_1321),
.Y(n_2776)
);

CKINVDCx6p67_ASAP7_75t_R g2777 ( 
.A(n_2391),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2092),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2251),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_2092),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2251),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2251),
.Y(n_2782)
);

INVx3_ASAP7_75t_L g2783 ( 
.A(n_2347),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2092),
.Y(n_2784)
);

BUFx4f_ASAP7_75t_L g2785 ( 
.A(n_2354),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2251),
.Y(n_2786)
);

NOR2x1p5_ASAP7_75t_L g2787 ( 
.A(n_2354),
.B(n_1296),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2251),
.Y(n_2788)
);

BUFx6f_ASAP7_75t_L g2789 ( 
.A(n_2092),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2092),
.Y(n_2790)
);

INVx3_ASAP7_75t_L g2791 ( 
.A(n_2347),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2092),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2251),
.Y(n_2793)
);

XNOR2x2_ASAP7_75t_SL g2794 ( 
.A(n_2417),
.B(n_1717),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2615),
.B(n_1297),
.Y(n_2795)
);

INVx3_ASAP7_75t_L g2796 ( 
.A(n_2639),
.Y(n_2796)
);

AND2x4_ASAP7_75t_L g2797 ( 
.A(n_2616),
.B(n_2617),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2443),
.Y(n_2798)
);

INVx2_ASAP7_75t_L g2799 ( 
.A(n_2418),
.Y(n_2799)
);

NOR2xp33_ASAP7_75t_L g2800 ( 
.A(n_2513),
.B(n_2507),
.Y(n_2800)
);

INVx4_ASAP7_75t_L g2801 ( 
.A(n_2697),
.Y(n_2801)
);

NAND2x1p5_ASAP7_75t_L g2802 ( 
.A(n_2785),
.B(n_2764),
.Y(n_2802)
);

CKINVDCx5p33_ASAP7_75t_R g2803 ( 
.A(n_2495),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2418),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2443),
.Y(n_2805)
);

AND2x4_ASAP7_75t_L g2806 ( 
.A(n_2616),
.B(n_1717),
.Y(n_2806)
);

CKINVDCx5p33_ASAP7_75t_R g2807 ( 
.A(n_2504),
.Y(n_2807)
);

INVx1_ASAP7_75t_SL g2808 ( 
.A(n_2416),
.Y(n_2808)
);

AOI22xp33_ASAP7_75t_L g2809 ( 
.A1(n_2676),
.A2(n_1319),
.B1(n_1442),
.B2(n_1290),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2444),
.Y(n_2810)
);

CKINVDCx20_ASAP7_75t_R g2811 ( 
.A(n_2421),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2444),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_2679),
.B(n_1298),
.Y(n_2813)
);

AND2x6_ASAP7_75t_L g2814 ( 
.A(n_2406),
.B(n_1527),
.Y(n_2814)
);

AND2x4_ASAP7_75t_L g2815 ( 
.A(n_2617),
.B(n_1527),
.Y(n_2815)
);

INVx2_ASAP7_75t_L g2816 ( 
.A(n_2418),
.Y(n_2816)
);

BUFx6f_ASAP7_75t_L g2817 ( 
.A(n_2571),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2679),
.B(n_1299),
.Y(n_2818)
);

BUFx3_ASAP7_75t_L g2819 ( 
.A(n_2697),
.Y(n_2819)
);

BUFx3_ASAP7_75t_L g2820 ( 
.A(n_2482),
.Y(n_2820)
);

NOR2xp33_ASAP7_75t_L g2821 ( 
.A(n_2538),
.B(n_1301),
.Y(n_2821)
);

NOR2x1p5_ASAP7_75t_L g2822 ( 
.A(n_2515),
.B(n_1305),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_SL g2823 ( 
.A(n_2593),
.B(n_1306),
.Y(n_2823)
);

HB1xp67_ASAP7_75t_L g2824 ( 
.A(n_2415),
.Y(n_2824)
);

AND2x4_ASAP7_75t_L g2825 ( 
.A(n_2663),
.B(n_1528),
.Y(n_2825)
);

AND2x2_ASAP7_75t_L g2826 ( 
.A(n_2414),
.B(n_1319),
.Y(n_2826)
);

INVx2_ASAP7_75t_L g2827 ( 
.A(n_2435),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2436),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2493),
.Y(n_2829)
);

BUFx2_ASAP7_75t_L g2830 ( 
.A(n_2403),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2493),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2501),
.Y(n_2832)
);

OA22x2_ASAP7_75t_L g2833 ( 
.A1(n_2544),
.A2(n_1308),
.B1(n_1312),
.B2(n_1307),
.Y(n_2833)
);

AND2x2_ASAP7_75t_L g2834 ( 
.A(n_2658),
.B(n_1319),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2452),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_L g2836 ( 
.A(n_2676),
.B(n_1313),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2462),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_L g2838 ( 
.A(n_2677),
.B(n_1315),
.Y(n_2838)
);

NOR2xp33_ASAP7_75t_L g2839 ( 
.A(n_2568),
.B(n_2430),
.Y(n_2839)
);

AND2x4_ASAP7_75t_L g2840 ( 
.A(n_2663),
.B(n_1528),
.Y(n_2840)
);

INVx2_ASAP7_75t_L g2841 ( 
.A(n_2438),
.Y(n_2841)
);

BUFx3_ASAP7_75t_L g2842 ( 
.A(n_2482),
.Y(n_2842)
);

INVx1_ASAP7_75t_SL g2843 ( 
.A(n_2777),
.Y(n_2843)
);

AOI22xp33_ASAP7_75t_L g2844 ( 
.A1(n_2677),
.A2(n_1568),
.B1(n_1591),
.B2(n_1442),
.Y(n_2844)
);

AOI22xp33_ASAP7_75t_L g2845 ( 
.A1(n_2688),
.A2(n_1568),
.B1(n_1591),
.B2(n_1442),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_2406),
.Y(n_2846)
);

BUFx2_ASAP7_75t_L g2847 ( 
.A(n_2421),
.Y(n_2847)
);

NAND2xp33_ASAP7_75t_L g2848 ( 
.A(n_2571),
.B(n_1316),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2466),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2467),
.Y(n_2850)
);

BUFx4f_ASAP7_75t_L g2851 ( 
.A(n_2768),
.Y(n_2851)
);

OA22x2_ASAP7_75t_L g2852 ( 
.A1(n_2575),
.A2(n_1320),
.B1(n_1322),
.B2(n_1317),
.Y(n_2852)
);

AND2x2_ASAP7_75t_L g2853 ( 
.A(n_2771),
.B(n_1568),
.Y(n_2853)
);

INVx2_ASAP7_75t_SL g2854 ( 
.A(n_2768),
.Y(n_2854)
);

OAI22xp5_ASAP7_75t_L g2855 ( 
.A1(n_2649),
.A2(n_1324),
.B1(n_1325),
.B2(n_1323),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2688),
.B(n_1327),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_SL g2857 ( 
.A(n_2405),
.B(n_2753),
.Y(n_2857)
);

INVx3_ASAP7_75t_L g2858 ( 
.A(n_2639),
.Y(n_2858)
);

INVx4_ASAP7_75t_L g2859 ( 
.A(n_2785),
.Y(n_2859)
);

OR2x2_ASAP7_75t_L g2860 ( 
.A(n_2413),
.B(n_1363),
.Y(n_2860)
);

BUFx3_ASAP7_75t_L g2861 ( 
.A(n_2527),
.Y(n_2861)
);

BUFx10_ASAP7_75t_L g2862 ( 
.A(n_2567),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2471),
.Y(n_2863)
);

AND2x2_ASAP7_75t_L g2864 ( 
.A(n_2579),
.B(n_1591),
.Y(n_2864)
);

INVx2_ASAP7_75t_L g2865 ( 
.A(n_2407),
.Y(n_2865)
);

INVx4_ASAP7_75t_L g2866 ( 
.A(n_2527),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2407),
.Y(n_2867)
);

INVx2_ASAP7_75t_L g2868 ( 
.A(n_2440),
.Y(n_2868)
);

BUFx8_ASAP7_75t_SL g2869 ( 
.A(n_2634),
.Y(n_2869)
);

NAND3x1_ASAP7_75t_L g2870 ( 
.A(n_2489),
.B(n_1434),
.C(n_1423),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2603),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2626),
.B(n_1329),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2626),
.B(n_1331),
.Y(n_2873)
);

INVx3_ASAP7_75t_L g2874 ( 
.A(n_2639),
.Y(n_2874)
);

AND2x2_ASAP7_75t_L g2875 ( 
.A(n_2759),
.B(n_1647),
.Y(n_2875)
);

INVx2_ASAP7_75t_L g2876 ( 
.A(n_2440),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2603),
.Y(n_2877)
);

AND2x4_ASAP7_75t_L g2878 ( 
.A(n_2625),
.B(n_2672),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2606),
.Y(n_2879)
);

INVxp67_ASAP7_75t_L g2880 ( 
.A(n_2455),
.Y(n_2880)
);

AND2x6_ASAP7_75t_L g2881 ( 
.A(n_2745),
.B(n_1531),
.Y(n_2881)
);

INVx5_ASAP7_75t_L g2882 ( 
.A(n_2564),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2606),
.Y(n_2883)
);

AND2x2_ASAP7_75t_L g2884 ( 
.A(n_2774),
.B(n_1647),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2478),
.Y(n_2885)
);

INVx2_ASAP7_75t_SL g2886 ( 
.A(n_2564),
.Y(n_2886)
);

OR2x2_ASAP7_75t_L g2887 ( 
.A(n_2776),
.B(n_1394),
.Y(n_2887)
);

BUFx6f_ASAP7_75t_L g2888 ( 
.A(n_2571),
.Y(n_2888)
);

INVx1_ASAP7_75t_SL g2889 ( 
.A(n_2439),
.Y(n_2889)
);

AND2x4_ASAP7_75t_L g2890 ( 
.A(n_2635),
.B(n_1531),
.Y(n_2890)
);

BUFx6f_ASAP7_75t_L g2891 ( 
.A(n_2789),
.Y(n_2891)
);

AOI22xp5_ASAP7_75t_L g2892 ( 
.A1(n_2454),
.A2(n_2750),
.B1(n_2772),
.B2(n_2425),
.Y(n_2892)
);

AND2x4_ASAP7_75t_L g2893 ( 
.A(n_2635),
.B(n_1567),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2483),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2486),
.Y(n_2895)
);

INVx4_ASAP7_75t_L g2896 ( 
.A(n_2528),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2487),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_SL g2898 ( 
.A(n_2757),
.B(n_1336),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_2655),
.B(n_1337),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2745),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_SL g2901 ( 
.A(n_2765),
.B(n_2437),
.Y(n_2901)
);

NOR2xp33_ASAP7_75t_L g2902 ( 
.A(n_2681),
.B(n_1340),
.Y(n_2902)
);

INVx2_ASAP7_75t_L g2903 ( 
.A(n_2749),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2655),
.B(n_1341),
.Y(n_2904)
);

INVx3_ASAP7_75t_L g2905 ( 
.A(n_2424),
.Y(n_2905)
);

BUFx6f_ASAP7_75t_L g2906 ( 
.A(n_2789),
.Y(n_2906)
);

NOR2xp33_ASAP7_75t_L g2907 ( 
.A(n_2686),
.B(n_1342),
.Y(n_2907)
);

CKINVDCx5p33_ASAP7_75t_R g2908 ( 
.A(n_2589),
.Y(n_2908)
);

BUFx2_ASAP7_75t_L g2909 ( 
.A(n_2408),
.Y(n_2909)
);

INVxp33_ASAP7_75t_SL g2910 ( 
.A(n_2691),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2453),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2456),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_2656),
.B(n_1344),
.Y(n_2913)
);

INVx4_ASAP7_75t_L g2914 ( 
.A(n_2528),
.Y(n_2914)
);

NOR2xp33_ASAP7_75t_L g2915 ( 
.A(n_2670),
.B(n_1345),
.Y(n_2915)
);

INVx2_ASAP7_75t_L g2916 ( 
.A(n_2749),
.Y(n_2916)
);

OAI22xp33_ASAP7_75t_L g2917 ( 
.A1(n_2661),
.A2(n_1349),
.B1(n_1351),
.B2(n_1347),
.Y(n_2917)
);

INVxp67_ASAP7_75t_L g2918 ( 
.A(n_2701),
.Y(n_2918)
);

INVx4_ASAP7_75t_L g2919 ( 
.A(n_2587),
.Y(n_2919)
);

INVx2_ASAP7_75t_SL g2920 ( 
.A(n_2596),
.Y(n_2920)
);

BUFx10_ASAP7_75t_L g2921 ( 
.A(n_2584),
.Y(n_2921)
);

BUFx4f_ASAP7_75t_L g2922 ( 
.A(n_2497),
.Y(n_2922)
);

AND2x2_ASAP7_75t_L g2923 ( 
.A(n_2554),
.B(n_1647),
.Y(n_2923)
);

INVx4_ASAP7_75t_L g2924 ( 
.A(n_2587),
.Y(n_2924)
);

NAND2xp5_ASAP7_75t_SL g2925 ( 
.A(n_2423),
.B(n_1354),
.Y(n_2925)
);

NAND2x1p5_ASAP7_75t_L g2926 ( 
.A(n_2764),
.B(n_1402),
.Y(n_2926)
);

CKINVDCx5p33_ASAP7_75t_R g2927 ( 
.A(n_2741),
.Y(n_2927)
);

INVx2_ASAP7_75t_L g2928 ( 
.A(n_2752),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2460),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2501),
.Y(n_2930)
);

INVx3_ASAP7_75t_L g2931 ( 
.A(n_2424),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2506),
.Y(n_2932)
);

NOR2xp33_ASAP7_75t_L g2933 ( 
.A(n_2600),
.B(n_1355),
.Y(n_2933)
);

INVx4_ASAP7_75t_L g2934 ( 
.A(n_2587),
.Y(n_2934)
);

BUFx2_ASAP7_75t_L g2935 ( 
.A(n_2584),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2506),
.Y(n_2936)
);

NAND2xp33_ASAP7_75t_L g2937 ( 
.A(n_2752),
.B(n_1357),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2520),
.Y(n_2938)
);

BUFx6f_ASAP7_75t_L g2939 ( 
.A(n_2789),
.Y(n_2939)
);

NOR2xp33_ASAP7_75t_L g2940 ( 
.A(n_2446),
.B(n_1361),
.Y(n_2940)
);

INVx2_ASAP7_75t_L g2941 ( 
.A(n_2763),
.Y(n_2941)
);

INVxp67_ASAP7_75t_SL g2942 ( 
.A(n_2763),
.Y(n_2942)
);

AND2x2_ASAP7_75t_L g2943 ( 
.A(n_2613),
.B(n_1688),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2520),
.Y(n_2944)
);

INVx2_ASAP7_75t_SL g2945 ( 
.A(n_2596),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2523),
.Y(n_2946)
);

BUFx4f_ASAP7_75t_L g2947 ( 
.A(n_2497),
.Y(n_2947)
);

CKINVDCx20_ASAP7_75t_R g2948 ( 
.A(n_2712),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2523),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2766),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_SL g2951 ( 
.A(n_2423),
.B(n_1362),
.Y(n_2951)
);

INVx2_ASAP7_75t_L g2952 ( 
.A(n_2766),
.Y(n_2952)
);

CKINVDCx5p33_ASAP7_75t_R g2953 ( 
.A(n_2511),
.Y(n_2953)
);

INVxp67_ASAP7_75t_SL g2954 ( 
.A(n_2779),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2525),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2525),
.Y(n_2956)
);

CKINVDCx5p33_ASAP7_75t_R g2957 ( 
.A(n_2650),
.Y(n_2957)
);

INVx1_ASAP7_75t_SL g2958 ( 
.A(n_2550),
.Y(n_2958)
);

AND2x6_ASAP7_75t_L g2959 ( 
.A(n_2779),
.B(n_1567),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_L g2960 ( 
.A(n_2656),
.B(n_1365),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2535),
.Y(n_2961)
);

AO22x2_ASAP7_75t_L g2962 ( 
.A1(n_2781),
.A2(n_1467),
.B1(n_1471),
.B2(n_1456),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2781),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_L g2964 ( 
.A(n_2667),
.B(n_1366),
.Y(n_2964)
);

INVx2_ASAP7_75t_SL g2965 ( 
.A(n_2664),
.Y(n_2965)
);

INVx2_ASAP7_75t_SL g2966 ( 
.A(n_2664),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2535),
.Y(n_2967)
);

OR2x6_ASAP7_75t_L g2968 ( 
.A(n_2731),
.B(n_1573),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2540),
.Y(n_2969)
);

BUFx8_ASAP7_75t_SL g2970 ( 
.A(n_2605),
.Y(n_2970)
);

INVx1_ASAP7_75t_SL g2971 ( 
.A(n_2623),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2540),
.Y(n_2972)
);

NAND2xp33_ASAP7_75t_L g2973 ( 
.A(n_2782),
.B(n_1368),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2549),
.Y(n_2974)
);

AND2x6_ASAP7_75t_L g2975 ( 
.A(n_2782),
.B(n_1573),
.Y(n_2975)
);

INVx4_ASAP7_75t_L g2976 ( 
.A(n_2636),
.Y(n_2976)
);

BUFx6f_ASAP7_75t_L g2977 ( 
.A(n_2451),
.Y(n_2977)
);

AND2x6_ASAP7_75t_L g2978 ( 
.A(n_2786),
.B(n_1577),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_L g2979 ( 
.A(n_2667),
.B(n_1369),
.Y(n_2979)
);

INVxp33_ASAP7_75t_SL g2980 ( 
.A(n_2732),
.Y(n_2980)
);

INVx5_ASAP7_75t_L g2981 ( 
.A(n_2692),
.Y(n_2981)
);

INVx3_ASAP7_75t_L g2982 ( 
.A(n_2441),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_L g2983 ( 
.A(n_2649),
.B(n_1370),
.Y(n_2983)
);

INVx4_ASAP7_75t_L g2984 ( 
.A(n_2636),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2668),
.B(n_1371),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2549),
.Y(n_2986)
);

AOI22xp5_ASAP7_75t_L g2987 ( 
.A1(n_2576),
.A2(n_1374),
.B1(n_1375),
.B2(n_1373),
.Y(n_2987)
);

NOR2xp33_ASAP7_75t_L g2988 ( 
.A(n_2684),
.B(n_1376),
.Y(n_2988)
);

INVx2_ASAP7_75t_L g2989 ( 
.A(n_2786),
.Y(n_2989)
);

AOI22xp33_ASAP7_75t_L g2990 ( 
.A1(n_2638),
.A2(n_1688),
.B1(n_1606),
.B2(n_1643),
.Y(n_2990)
);

INVxp33_ASAP7_75t_L g2991 ( 
.A(n_2706),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_SL g2992 ( 
.A(n_2636),
.B(n_1378),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2788),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2788),
.Y(n_2994)
);

HB1xp67_ASAP7_75t_L g2995 ( 
.A(n_2633),
.Y(n_2995)
);

NAND2x1p5_ASAP7_75t_L g2996 ( 
.A(n_2465),
.B(n_2702),
.Y(n_2996)
);

INVx2_ASAP7_75t_SL g2997 ( 
.A(n_2692),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2557),
.Y(n_2998)
);

BUFx6f_ASAP7_75t_L g2999 ( 
.A(n_2451),
.Y(n_2999)
);

BUFx3_ASAP7_75t_L g3000 ( 
.A(n_2707),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2557),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2793),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2668),
.B(n_1379),
.Y(n_3003)
);

BUFx3_ASAP7_75t_L g3004 ( 
.A(n_2707),
.Y(n_3004)
);

INVx2_ASAP7_75t_L g3005 ( 
.A(n_2793),
.Y(n_3005)
);

NOR2xp33_ASAP7_75t_L g3006 ( 
.A(n_2610),
.B(n_1382),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_SL g3007 ( 
.A(n_2470),
.B(n_1385),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2570),
.Y(n_3008)
);

CKINVDCx5p33_ASAP7_75t_R g3009 ( 
.A(n_2731),
.Y(n_3009)
);

INVx6_ASAP7_75t_L g3010 ( 
.A(n_2735),
.Y(n_3010)
);

AND2x4_ASAP7_75t_SL g3011 ( 
.A(n_2735),
.B(n_1688),
.Y(n_3011)
);

NOR2xp33_ASAP7_75t_L g3012 ( 
.A(n_2622),
.B(n_1388),
.Y(n_3012)
);

BUFx2_ASAP7_75t_L g3013 ( 
.A(n_2754),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2570),
.Y(n_3014)
);

AND2x2_ASAP7_75t_SL g3015 ( 
.A(n_2703),
.B(n_1148),
.Y(n_3015)
);

OR2x6_ASAP7_75t_L g3016 ( 
.A(n_2574),
.B(n_1577),
.Y(n_3016)
);

NOR2xp33_ASAP7_75t_L g3017 ( 
.A(n_2620),
.B(n_1389),
.Y(n_3017)
);

BUFx2_ASAP7_75t_L g3018 ( 
.A(n_2694),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_2572),
.B(n_1391),
.Y(n_3019)
);

BUFx2_ASAP7_75t_L g3020 ( 
.A(n_2683),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2572),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2573),
.Y(n_3022)
);

AND2x2_ASAP7_75t_L g3023 ( 
.A(n_2583),
.B(n_1392),
.Y(n_3023)
);

NAND2x1p5_ASAP7_75t_L g3024 ( 
.A(n_2702),
.B(n_1495),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2573),
.Y(n_3025)
);

NOR2xp33_ASAP7_75t_L g3026 ( 
.A(n_2484),
.B(n_1396),
.Y(n_3026)
);

INVx2_ASAP7_75t_L g3027 ( 
.A(n_2585),
.Y(n_3027)
);

BUFx6f_ASAP7_75t_L g3028 ( 
.A(n_2451),
.Y(n_3028)
);

INVx2_ASAP7_75t_SL g3029 ( 
.A(n_2562),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2585),
.Y(n_3030)
);

NOR2xp33_ASAP7_75t_L g3031 ( 
.A(n_2491),
.B(n_1397),
.Y(n_3031)
);

INVx2_ASAP7_75t_L g3032 ( 
.A(n_2577),
.Y(n_3032)
);

INVx2_ASAP7_75t_L g3033 ( 
.A(n_2578),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2502),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2627),
.B(n_1398),
.Y(n_3035)
);

AND2x4_ASAP7_75t_L g3036 ( 
.A(n_2696),
.B(n_1606),
.Y(n_3036)
);

NOR2xp33_ASAP7_75t_L g3037 ( 
.A(n_2598),
.B(n_1400),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2503),
.Y(n_3038)
);

NOR2xp33_ASAP7_75t_L g3039 ( 
.A(n_2643),
.B(n_1401),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2505),
.Y(n_3040)
);

NAND3xp33_ASAP7_75t_SL g3041 ( 
.A(n_2410),
.B(n_1406),
.C(n_1405),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_SL g3042 ( 
.A(n_2470),
.B(n_1408),
.Y(n_3042)
);

AND2x4_ASAP7_75t_L g3043 ( 
.A(n_2700),
.B(n_1643),
.Y(n_3043)
);

BUFx6f_ASAP7_75t_L g3044 ( 
.A(n_2565),
.Y(n_3044)
);

NOR2xp33_ASAP7_75t_L g3045 ( 
.A(n_2590),
.B(n_2724),
.Y(n_3045)
);

INVx3_ASAP7_75t_L g3046 ( 
.A(n_2441),
.Y(n_3046)
);

INVx3_ASAP7_75t_L g3047 ( 
.A(n_2473),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_SL g3048 ( 
.A(n_2468),
.B(n_1409),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2508),
.Y(n_3049)
);

BUFx2_ASAP7_75t_L g3050 ( 
.A(n_2704),
.Y(n_3050)
);

NOR2xp33_ASAP7_75t_SL g3051 ( 
.A(n_2605),
.B(n_2646),
.Y(n_3051)
);

AND2x2_ASAP7_75t_L g3052 ( 
.A(n_2492),
.B(n_1410),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_SL g3053 ( 
.A(n_2699),
.B(n_1411),
.Y(n_3053)
);

INVx3_ASAP7_75t_L g3054 ( 
.A(n_2473),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2509),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_2580),
.B(n_1413),
.Y(n_3056)
);

INVx3_ASAP7_75t_L g3057 ( 
.A(n_2747),
.Y(n_3057)
);

BUFx3_ASAP7_75t_L g3058 ( 
.A(n_2711),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_SL g3059 ( 
.A(n_2597),
.B(n_1414),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2581),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2582),
.Y(n_3061)
);

AOI22xp5_ASAP7_75t_L g3062 ( 
.A1(n_2727),
.A2(n_1416),
.B1(n_1417),
.B2(n_1415),
.Y(n_3062)
);

BUFx2_ASAP7_75t_L g3063 ( 
.A(n_2678),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2588),
.Y(n_3064)
);

BUFx2_ASAP7_75t_L g3065 ( 
.A(n_2644),
.Y(n_3065)
);

AND3x1_ASAP7_75t_L g3066 ( 
.A(n_2740),
.B(n_1711),
.C(n_1708),
.Y(n_3066)
);

OR2x6_ASAP7_75t_L g3067 ( 
.A(n_2787),
.B(n_1155),
.Y(n_3067)
);

OR2x6_ASAP7_75t_L g3068 ( 
.A(n_2726),
.B(n_1248),
.Y(n_3068)
);

CKINVDCx5p33_ASAP7_75t_R g3069 ( 
.A(n_2646),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2591),
.Y(n_3070)
);

BUFx6f_ASAP7_75t_L g3071 ( 
.A(n_2566),
.Y(n_3071)
);

INVx2_ASAP7_75t_L g3072 ( 
.A(n_2595),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2602),
.Y(n_3073)
);

HB1xp67_ASAP7_75t_L g3074 ( 
.A(n_2654),
.Y(n_3074)
);

INVx2_ASAP7_75t_L g3075 ( 
.A(n_2604),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2690),
.Y(n_3076)
);

AND2x6_ASAP7_75t_L g3077 ( 
.A(n_2592),
.B(n_1159),
.Y(n_3077)
);

OAI22xp33_ASAP7_75t_L g3078 ( 
.A1(n_2536),
.A2(n_1422),
.B1(n_1427),
.B2(n_1421),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2690),
.Y(n_3079)
);

INVx3_ASAP7_75t_L g3080 ( 
.A(n_2747),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2404),
.B(n_1428),
.Y(n_3081)
);

AOI22xp33_ASAP7_75t_L g3082 ( 
.A1(n_2725),
.A2(n_1430),
.B1(n_1433),
.B2(n_1429),
.Y(n_3082)
);

INVx3_ASAP7_75t_L g3083 ( 
.A(n_2755),
.Y(n_3083)
);

AND2x6_ASAP7_75t_L g3084 ( 
.A(n_2592),
.B(n_2599),
.Y(n_3084)
);

NOR2xp33_ASAP7_75t_L g3085 ( 
.A(n_2594),
.B(n_2738),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2510),
.Y(n_3086)
);

BUFx4f_ASAP7_75t_L g3087 ( 
.A(n_2730),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2512),
.Y(n_3088)
);

BUFx3_ASAP7_75t_L g3089 ( 
.A(n_2736),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2514),
.Y(n_3090)
);

BUFx6f_ASAP7_75t_L g3091 ( 
.A(n_2399),
.Y(n_3091)
);

AND2x2_ASAP7_75t_L g3092 ( 
.A(n_2518),
.B(n_1435),
.Y(n_3092)
);

BUFx6f_ASAP7_75t_L g3093 ( 
.A(n_2744),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_2770),
.B(n_2545),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2628),
.B(n_1436),
.Y(n_3095)
);

AND2x6_ASAP7_75t_L g3096 ( 
.A(n_2599),
.B(n_1164),
.Y(n_3096)
);

HB1xp67_ASAP7_75t_L g3097 ( 
.A(n_2654),
.Y(n_3097)
);

AND2x2_ASAP7_75t_L g3098 ( 
.A(n_2548),
.B(n_1437),
.Y(n_3098)
);

INVxp67_ASAP7_75t_L g3099 ( 
.A(n_2458),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2517),
.Y(n_3100)
);

AND2x4_ASAP7_75t_L g3101 ( 
.A(n_2660),
.B(n_1439),
.Y(n_3101)
);

AND2x6_ASAP7_75t_L g3102 ( 
.A(n_2666),
.B(n_1164),
.Y(n_3102)
);

OR2x6_ASAP7_75t_L g3103 ( 
.A(n_2730),
.B(n_2494),
.Y(n_3103)
);

BUFx8_ASAP7_75t_SL g3104 ( 
.A(n_2710),
.Y(n_3104)
);

NOR2xp33_ASAP7_75t_L g3105 ( 
.A(n_2742),
.B(n_1438),
.Y(n_3105)
);

NOR2xp33_ASAP7_75t_L g3106 ( 
.A(n_2743),
.B(n_1443),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_2521),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_L g3108 ( 
.A(n_2659),
.B(n_1448),
.Y(n_3108)
);

AND2x2_ASAP7_75t_L g3109 ( 
.A(n_2555),
.B(n_1450),
.Y(n_3109)
);

AOI22xp5_ASAP7_75t_L g3110 ( 
.A1(n_2531),
.A2(n_1452),
.B1(n_1455),
.B2(n_1451),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2524),
.Y(n_3111)
);

CKINVDCx5p33_ASAP7_75t_R g3112 ( 
.A(n_2710),
.Y(n_3112)
);

INVx3_ASAP7_75t_L g3113 ( 
.A(n_2755),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_2722),
.B(n_1458),
.Y(n_3114)
);

NOR2xp33_ASAP7_75t_L g3115 ( 
.A(n_2729),
.B(n_1459),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2526),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2539),
.Y(n_3117)
);

AND2x2_ASAP7_75t_L g3118 ( 
.A(n_2433),
.B(n_2464),
.Y(n_3118)
);

INVx2_ASAP7_75t_L g3119 ( 
.A(n_2541),
.Y(n_3119)
);

INVx2_ASAP7_75t_SL g3120 ( 
.A(n_2562),
.Y(n_3120)
);

INVx2_ASAP7_75t_L g3121 ( 
.A(n_2542),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2546),
.Y(n_3122)
);

BUFx3_ASAP7_75t_L g3123 ( 
.A(n_2736),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2601),
.B(n_1461),
.Y(n_3124)
);

INVxp67_ASAP7_75t_SL g3125 ( 
.A(n_2472),
.Y(n_3125)
);

INVx6_ASAP7_75t_L g3126 ( 
.A(n_2729),
.Y(n_3126)
);

BUFx3_ASAP7_75t_L g3127 ( 
.A(n_2629),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_SL g3128 ( 
.A(n_2556),
.B(n_1462),
.Y(n_3128)
);

AOI22xp33_ASAP7_75t_L g3129 ( 
.A1(n_2530),
.A2(n_1469),
.B1(n_1470),
.B2(n_1465),
.Y(n_3129)
);

AND2x4_ASAP7_75t_L g3130 ( 
.A(n_2695),
.B(n_1440),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_SL g3131 ( 
.A(n_2561),
.B(n_1472),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_SL g3132 ( 
.A(n_2561),
.B(n_1475),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2559),
.Y(n_3133)
);

INVx1_ASAP7_75t_SL g3134 ( 
.A(n_2729),
.Y(n_3134)
);

INVx2_ASAP7_75t_L g3135 ( 
.A(n_2447),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2560),
.Y(n_3136)
);

AND2x2_ASAP7_75t_L g3137 ( 
.A(n_2532),
.B(n_1476),
.Y(n_3137)
);

INVx2_ASAP7_75t_L g3138 ( 
.A(n_2448),
.Y(n_3138)
);

CKINVDCx5p33_ASAP7_75t_R g3139 ( 
.A(n_2519),
.Y(n_3139)
);

BUFx3_ASAP7_75t_L g3140 ( 
.A(n_2629),
.Y(n_3140)
);

NAND2xp33_ASAP7_75t_L g3141 ( 
.A(n_2746),
.B(n_1480),
.Y(n_3141)
);

AND2x4_ASAP7_75t_L g3142 ( 
.A(n_2657),
.B(n_1441),
.Y(n_3142)
);

BUFx6f_ASAP7_75t_L g3143 ( 
.A(n_2748),
.Y(n_3143)
);

OAI22xp5_ASAP7_75t_L g3144 ( 
.A1(n_2563),
.A2(n_1488),
.B1(n_1489),
.B2(n_1484),
.Y(n_3144)
);

INVx1_ASAP7_75t_SL g3145 ( 
.A(n_2422),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_SL g3146 ( 
.A(n_2551),
.B(n_1490),
.Y(n_3146)
);

INVx3_ASAP7_75t_L g3147 ( 
.A(n_2767),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2698),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_2705),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2450),
.Y(n_3150)
);

OAI22xp33_ASAP7_75t_L g3151 ( 
.A1(n_2537),
.A2(n_1493),
.B1(n_1494),
.B2(n_1492),
.Y(n_3151)
);

BUFx6f_ASAP7_75t_L g3152 ( 
.A(n_2751),
.Y(n_3152)
);

INVx4_ASAP7_75t_L g3153 ( 
.A(n_2689),
.Y(n_3153)
);

INVx3_ASAP7_75t_L g3154 ( 
.A(n_2767),
.Y(n_3154)
);

AND2x4_ASAP7_75t_L g3155 ( 
.A(n_2662),
.B(n_1447),
.Y(n_3155)
);

NAND2x1p5_ASAP7_75t_L g3156 ( 
.A(n_2652),
.B(n_1526),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2687),
.Y(n_3157)
);

BUFx10_ASAP7_75t_L g3158 ( 
.A(n_2739),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2618),
.B(n_1496),
.Y(n_3159)
);

AND2x6_ASAP7_75t_L g3160 ( 
.A(n_2457),
.B(n_2459),
.Y(n_3160)
);

NOR2xp33_ASAP7_75t_L g3161 ( 
.A(n_2739),
.B(n_1498),
.Y(n_3161)
);

INVx2_ASAP7_75t_SL g3162 ( 
.A(n_2652),
.Y(n_3162)
);

INVx3_ASAP7_75t_L g3163 ( 
.A(n_2783),
.Y(n_3163)
);

AND2x4_ASAP7_75t_L g3164 ( 
.A(n_2675),
.B(n_1454),
.Y(n_3164)
);

INVx1_ASAP7_75t_L g3165 ( 
.A(n_2461),
.Y(n_3165)
);

BUFx10_ASAP7_75t_L g3166 ( 
.A(n_2723),
.Y(n_3166)
);

INVx8_ASAP7_75t_L g3167 ( 
.A(n_2689),
.Y(n_3167)
);

NAND2xp33_ASAP7_75t_SL g3168 ( 
.A(n_2648),
.B(n_1701),
.Y(n_3168)
);

INVx3_ASAP7_75t_L g3169 ( 
.A(n_2783),
.Y(n_3169)
);

BUFx3_ASAP7_75t_L g3170 ( 
.A(n_2632),
.Y(n_3170)
);

INVx5_ASAP7_75t_L g3171 ( 
.A(n_2791),
.Y(n_3171)
);

BUFx10_ASAP7_75t_L g3172 ( 
.A(n_2709),
.Y(n_3172)
);

INVx5_ASAP7_75t_L g3173 ( 
.A(n_2791),
.Y(n_3173)
);

AND2x4_ASAP7_75t_L g3174 ( 
.A(n_2675),
.B(n_1457),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_L g3175 ( 
.A(n_2619),
.B(n_1500),
.Y(n_3175)
);

OR2x2_ASAP7_75t_L g3176 ( 
.A(n_2411),
.B(n_1691),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_2463),
.Y(n_3177)
);

NOR2xp33_ASAP7_75t_SL g3178 ( 
.A(n_2734),
.B(n_1503),
.Y(n_3178)
);

BUFx2_ASAP7_75t_L g3179 ( 
.A(n_2558),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2469),
.Y(n_3180)
);

AND2x2_ASAP7_75t_SL g3181 ( 
.A(n_2673),
.B(n_2609),
.Y(n_3181)
);

NOR2xp33_ASAP7_75t_L g3182 ( 
.A(n_2498),
.B(n_1504),
.Y(n_3182)
);

BUFx6f_ASAP7_75t_L g3183 ( 
.A(n_2756),
.Y(n_3183)
);

BUFx3_ASAP7_75t_L g3184 ( 
.A(n_2640),
.Y(n_3184)
);

INVx2_ASAP7_75t_L g3185 ( 
.A(n_2474),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2476),
.Y(n_3186)
);

BUFx6f_ASAP7_75t_L g3187 ( 
.A(n_2769),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2624),
.Y(n_3188)
);

AOI22xp5_ASAP7_75t_L g3189 ( 
.A1(n_2733),
.A2(n_1506),
.B1(n_1508),
.B2(n_1505),
.Y(n_3189)
);

AND2x6_ASAP7_75t_L g3190 ( 
.A(n_2479),
.B(n_1164),
.Y(n_3190)
);

INVx5_ASAP7_75t_L g3191 ( 
.A(n_2669),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_2480),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_SL g3193 ( 
.A(n_2761),
.B(n_1509),
.Y(n_3193)
);

INVx5_ASAP7_75t_L g3194 ( 
.A(n_2563),
.Y(n_3194)
);

INVx2_ASAP7_75t_L g3195 ( 
.A(n_2481),
.Y(n_3195)
);

INVx2_ASAP7_75t_L g3196 ( 
.A(n_2485),
.Y(n_3196)
);

NAND2xp33_ASAP7_75t_L g3197 ( 
.A(n_2778),
.B(n_1512),
.Y(n_3197)
);

AND2x4_ASAP7_75t_L g3198 ( 
.A(n_2674),
.B(n_1460),
.Y(n_3198)
);

AND2x2_ASAP7_75t_L g3199 ( 
.A(n_2645),
.B(n_1510),
.Y(n_3199)
);

INVx3_ASAP7_75t_L g3200 ( 
.A(n_2533),
.Y(n_3200)
);

NOR2xp33_ASAP7_75t_L g3201 ( 
.A(n_2516),
.B(n_1511),
.Y(n_3201)
);

INVx1_ASAP7_75t_SL g3202 ( 
.A(n_2522),
.Y(n_3202)
);

INVx4_ASAP7_75t_L g3203 ( 
.A(n_2534),
.Y(n_3203)
);

NOR3xp33_ASAP7_75t_SL g3204 ( 
.A(n_2737),
.B(n_2445),
.C(n_2428),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_2693),
.B(n_1514),
.Y(n_3205)
);

INVx2_ASAP7_75t_L g3206 ( 
.A(n_2488),
.Y(n_3206)
);

INVx3_ASAP7_75t_L g3207 ( 
.A(n_2533),
.Y(n_3207)
);

INVx4_ASAP7_75t_L g3208 ( 
.A(n_2534),
.Y(n_3208)
);

AND2x2_ASAP7_75t_L g3209 ( 
.A(n_2647),
.B(n_1517),
.Y(n_3209)
);

INVx1_ASAP7_75t_SL g3210 ( 
.A(n_2529),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_L g3211 ( 
.A(n_2621),
.B(n_1518),
.Y(n_3211)
);

AND2x2_ASAP7_75t_L g3212 ( 
.A(n_2494),
.B(n_1520),
.Y(n_3212)
);

INVx2_ASAP7_75t_L g3213 ( 
.A(n_2490),
.Y(n_3213)
);

BUFx6f_ASAP7_75t_SL g3214 ( 
.A(n_2713),
.Y(n_3214)
);

AOI22xp5_ASAP7_75t_L g3215 ( 
.A1(n_2775),
.A2(n_1524),
.B1(n_1529),
.B2(n_1522),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_2496),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_2499),
.Y(n_3217)
);

OR2x2_ASAP7_75t_L g3218 ( 
.A(n_2419),
.B(n_1551),
.Y(n_3218)
);

OR2x2_ASAP7_75t_L g3219 ( 
.A(n_2449),
.B(n_1556),
.Y(n_3219)
);

INVx2_ASAP7_75t_L g3220 ( 
.A(n_2500),
.Y(n_3220)
);

INVx1_ASAP7_75t_SL g3221 ( 
.A(n_2409),
.Y(n_3221)
);

NOR2xp33_ASAP7_75t_R g3222 ( 
.A(n_2728),
.B(n_1532),
.Y(n_3222)
);

AND2x4_ASAP7_75t_L g3223 ( 
.A(n_2614),
.B(n_1466),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_2552),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_SL g3225 ( 
.A(n_2714),
.B(n_2715),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_L g3226 ( 
.A(n_2641),
.B(n_1533),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_L g3227 ( 
.A(n_2653),
.B(n_1534),
.Y(n_3227)
);

AOI22xp5_ASAP7_75t_SL g3228 ( 
.A1(n_2718),
.A2(n_1720),
.B1(n_1718),
.B2(n_1539),
.Y(n_3228)
);

NOR2xp33_ASAP7_75t_L g3229 ( 
.A(n_2758),
.B(n_2760),
.Y(n_3229)
);

INVx3_ASAP7_75t_L g3230 ( 
.A(n_2547),
.Y(n_3230)
);

BUFx6f_ASAP7_75t_L g3231 ( 
.A(n_2780),
.Y(n_3231)
);

AND2x4_ASAP7_75t_L g3232 ( 
.A(n_2719),
.B(n_1468),
.Y(n_3232)
);

OAI22xp5_ASAP7_75t_L g3233 ( 
.A1(n_2784),
.A2(n_1542),
.B1(n_1543),
.B2(n_1537),
.Y(n_3233)
);

BUFx8_ASAP7_75t_SL g3234 ( 
.A(n_2720),
.Y(n_3234)
);

NOR2xp33_ASAP7_75t_L g3235 ( 
.A(n_2773),
.B(n_1544),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_L g3236 ( 
.A(n_2607),
.B(n_1545),
.Y(n_3236)
);

NOR2xp33_ASAP7_75t_L g3237 ( 
.A(n_2717),
.B(n_1548),
.Y(n_3237)
);

AND2x4_ASAP7_75t_L g3238 ( 
.A(n_2721),
.B(n_1477),
.Y(n_3238)
);

BUFx6f_ASAP7_75t_L g3239 ( 
.A(n_2790),
.Y(n_3239)
);

NOR2xp33_ASAP7_75t_L g3240 ( 
.A(n_2708),
.B(n_1550),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_2400),
.Y(n_3241)
);

INVx2_ASAP7_75t_L g3242 ( 
.A(n_2612),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_L g3243 ( 
.A(n_2553),
.B(n_1552),
.Y(n_3243)
);

NOR2xp33_ASAP7_75t_L g3244 ( 
.A(n_2716),
.B(n_1553),
.Y(n_3244)
);

INVx3_ASAP7_75t_L g3245 ( 
.A(n_2547),
.Y(n_3245)
);

CKINVDCx8_ASAP7_75t_R g3246 ( 
.A(n_2680),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_2611),
.B(n_1555),
.Y(n_3247)
);

AND2x6_ASAP7_75t_L g3248 ( 
.A(n_2792),
.B(n_1164),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_L g3249 ( 
.A(n_2682),
.B(n_1557),
.Y(n_3249)
);

AND2x6_ASAP7_75t_L g3250 ( 
.A(n_2665),
.B(n_1201),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_2401),
.Y(n_3251)
);

AND2x2_ASAP7_75t_L g3252 ( 
.A(n_2685),
.B(n_1558),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_2402),
.Y(n_3253)
);

INVx4_ASAP7_75t_L g3254 ( 
.A(n_2412),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_L g3255 ( 
.A(n_2642),
.B(n_1559),
.Y(n_3255)
);

INVxp33_ASAP7_75t_L g3256 ( 
.A(n_2420),
.Y(n_3256)
);

INVx2_ASAP7_75t_L g3257 ( 
.A(n_2762),
.Y(n_3257)
);

INVx3_ASAP7_75t_L g3258 ( 
.A(n_2426),
.Y(n_3258)
);

INVx3_ASAP7_75t_L g3259 ( 
.A(n_2427),
.Y(n_3259)
);

NOR2xp33_ASAP7_75t_L g3260 ( 
.A(n_2429),
.B(n_1560),
.Y(n_3260)
);

INVx3_ASAP7_75t_L g3261 ( 
.A(n_2432),
.Y(n_3261)
);

NOR2xp33_ASAP7_75t_L g3262 ( 
.A(n_2434),
.B(n_1565),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_2586),
.B(n_1569),
.Y(n_3263)
);

NOR2xp33_ASAP7_75t_L g3264 ( 
.A(n_2671),
.B(n_1570),
.Y(n_3264)
);

BUFx3_ASAP7_75t_L g3265 ( 
.A(n_2671),
.Y(n_3265)
);

HB1xp67_ASAP7_75t_L g3266 ( 
.A(n_2431),
.Y(n_3266)
);

CKINVDCx20_ASAP7_75t_R g3267 ( 
.A(n_2665),
.Y(n_3267)
);

NOR2x1p5_ASAP7_75t_L g3268 ( 
.A(n_2442),
.B(n_1572),
.Y(n_3268)
);

AOI22xp33_ASAP7_75t_L g3269 ( 
.A1(n_2651),
.A2(n_1576),
.B1(n_1579),
.B2(n_1575),
.Y(n_3269)
);

INVx2_ASAP7_75t_L g3270 ( 
.A(n_2608),
.Y(n_3270)
);

INVx3_ASAP7_75t_L g3271 ( 
.A(n_2637),
.Y(n_3271)
);

NOR2xp33_ASAP7_75t_L g3272 ( 
.A(n_2475),
.B(n_1582),
.Y(n_3272)
);

BUFx6f_ASAP7_75t_SL g3273 ( 
.A(n_2477),
.Y(n_3273)
);

INVx2_ASAP7_75t_L g3274 ( 
.A(n_2543),
.Y(n_3274)
);

INVx2_ASAP7_75t_SL g3275 ( 
.A(n_2630),
.Y(n_3275)
);

AND2x4_ASAP7_75t_L g3276 ( 
.A(n_2631),
.B(n_1478),
.Y(n_3276)
);

CKINVDCx16_ASAP7_75t_R g3277 ( 
.A(n_2569),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_2615),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_2615),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_2615),
.Y(n_3280)
);

INVxp67_ASAP7_75t_L g3281 ( 
.A(n_2416),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_2615),
.Y(n_3282)
);

INVx2_ASAP7_75t_L g3283 ( 
.A(n_2418),
.Y(n_3283)
);

INVxp67_ASAP7_75t_SL g3284 ( 
.A(n_2416),
.Y(n_3284)
);

INVx2_ASAP7_75t_L g3285 ( 
.A(n_2418),
.Y(n_3285)
);

CKINVDCx16_ASAP7_75t_R g3286 ( 
.A(n_2691),
.Y(n_3286)
);

AOI22xp33_ASAP7_75t_L g3287 ( 
.A1(n_2676),
.A2(n_1587),
.B1(n_1590),
.B2(n_1583),
.Y(n_3287)
);

INVx3_ASAP7_75t_L g3288 ( 
.A(n_2639),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_L g3289 ( 
.A(n_2615),
.B(n_1592),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_2615),
.Y(n_3290)
);

BUFx6f_ASAP7_75t_L g3291 ( 
.A(n_2571),
.Y(n_3291)
);

INVx2_ASAP7_75t_L g3292 ( 
.A(n_2418),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_2615),
.Y(n_3293)
);

NOR2xp33_ASAP7_75t_L g3294 ( 
.A(n_2513),
.B(n_1594),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_2615),
.Y(n_3295)
);

AND2x6_ASAP7_75t_L g3296 ( 
.A(n_2406),
.B(n_1201),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_SL g3297 ( 
.A(n_2593),
.B(n_1595),
.Y(n_3297)
);

AND2x4_ASAP7_75t_L g3298 ( 
.A(n_2615),
.B(n_1479),
.Y(n_3298)
);

INVx3_ASAP7_75t_L g3299 ( 
.A(n_2639),
.Y(n_3299)
);

INVx2_ASAP7_75t_L g3300 ( 
.A(n_2418),
.Y(n_3300)
);

INVx2_ASAP7_75t_L g3301 ( 
.A(n_2418),
.Y(n_3301)
);

NOR2xp33_ASAP7_75t_L g3302 ( 
.A(n_2513),
.B(n_1597),
.Y(n_3302)
);

INVx3_ASAP7_75t_L g3303 ( 
.A(n_2639),
.Y(n_3303)
);

INVx1_ASAP7_75t_SL g3304 ( 
.A(n_2416),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_2615),
.Y(n_3305)
);

OR2x6_ASAP7_75t_L g3306 ( 
.A(n_2421),
.B(n_1698),
.Y(n_3306)
);

AOI22xp5_ASAP7_75t_L g3307 ( 
.A1(n_2430),
.A2(n_1601),
.B1(n_1602),
.B2(n_1598),
.Y(n_3307)
);

INVx1_ASAP7_75t_L g3308 ( 
.A(n_2615),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_2615),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_2615),
.B(n_1603),
.Y(n_3310)
);

AND2x4_ASAP7_75t_L g3311 ( 
.A(n_2615),
.B(n_1482),
.Y(n_3311)
);

INVx3_ASAP7_75t_L g3312 ( 
.A(n_2639),
.Y(n_3312)
);

NOR2xp33_ASAP7_75t_L g3313 ( 
.A(n_2513),
.B(n_1604),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_2615),
.B(n_1605),
.Y(n_3314)
);

AND2x2_ASAP7_75t_L g3315 ( 
.A(n_2414),
.B(n_1607),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_2615),
.Y(n_3316)
);

INVx2_ASAP7_75t_L g3317 ( 
.A(n_2418),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_L g3318 ( 
.A(n_2615),
.B(n_1609),
.Y(n_3318)
);

INVx2_ASAP7_75t_SL g3319 ( 
.A(n_2482),
.Y(n_3319)
);

INVx4_ASAP7_75t_L g3320 ( 
.A(n_2697),
.Y(n_3320)
);

BUFx6f_ASAP7_75t_L g3321 ( 
.A(n_2571),
.Y(n_3321)
);

HB1xp67_ASAP7_75t_L g3322 ( 
.A(n_2416),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_2615),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_L g3324 ( 
.A(n_2615),
.B(n_1612),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_L g3325 ( 
.A(n_2615),
.B(n_1613),
.Y(n_3325)
);

INVxp67_ASAP7_75t_SL g3326 ( 
.A(n_2416),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_2615),
.Y(n_3327)
);

BUFx6f_ASAP7_75t_L g3328 ( 
.A(n_2571),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_2615),
.Y(n_3329)
);

INVx3_ASAP7_75t_L g3330 ( 
.A(n_2639),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_2615),
.B(n_1614),
.Y(n_3331)
);

BUFx3_ASAP7_75t_L g3332 ( 
.A(n_2697),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_SL g3333 ( 
.A(n_2593),
.B(n_1617),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_2615),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_L g3335 ( 
.A(n_2615),
.B(n_1619),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_2615),
.Y(n_3336)
);

INVx4_ASAP7_75t_SL g3337 ( 
.A(n_2515),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_SL g3338 ( 
.A(n_2593),
.B(n_1620),
.Y(n_3338)
);

OR2x2_ASAP7_75t_L g3339 ( 
.A(n_2417),
.B(n_1629),
.Y(n_3339)
);

CKINVDCx16_ASAP7_75t_R g3340 ( 
.A(n_2691),
.Y(n_3340)
);

INVx4_ASAP7_75t_L g3341 ( 
.A(n_2697),
.Y(n_3341)
);

NAND2xp33_ASAP7_75t_SL g3342 ( 
.A(n_2437),
.B(n_1697),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_2615),
.Y(n_3343)
);

INVx1_ASAP7_75t_SL g3344 ( 
.A(n_2416),
.Y(n_3344)
);

INVxp67_ASAP7_75t_SL g3345 ( 
.A(n_2416),
.Y(n_3345)
);

BUFx6f_ASAP7_75t_L g3346 ( 
.A(n_2571),
.Y(n_3346)
);

INVx3_ASAP7_75t_L g3347 ( 
.A(n_2639),
.Y(n_3347)
);

OR2x6_ASAP7_75t_L g3348 ( 
.A(n_2421),
.B(n_1698),
.Y(n_3348)
);

AND2x2_ASAP7_75t_SL g3349 ( 
.A(n_2691),
.B(n_1248),
.Y(n_3349)
);

INVx1_ASAP7_75t_SL g3350 ( 
.A(n_2416),
.Y(n_3350)
);

INVx4_ASAP7_75t_L g3351 ( 
.A(n_2697),
.Y(n_3351)
);

INVx2_ASAP7_75t_L g3352 ( 
.A(n_2418),
.Y(n_3352)
);

AND2x6_ASAP7_75t_L g3353 ( 
.A(n_2406),
.B(n_1201),
.Y(n_3353)
);

AND2x2_ASAP7_75t_L g3354 ( 
.A(n_2414),
.B(n_1621),
.Y(n_3354)
);

NOR2xp33_ASAP7_75t_L g3355 ( 
.A(n_2513),
.B(n_1622),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_2615),
.Y(n_3356)
);

INVx2_ASAP7_75t_L g3357 ( 
.A(n_2418),
.Y(n_3357)
);

AND2x2_ASAP7_75t_L g3358 ( 
.A(n_2414),
.B(n_1632),
.Y(n_3358)
);

INVx2_ASAP7_75t_SL g3359 ( 
.A(n_2482),
.Y(n_3359)
);

INVx4_ASAP7_75t_L g3360 ( 
.A(n_2697),
.Y(n_3360)
);

INVx2_ASAP7_75t_SL g3361 ( 
.A(n_2482),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_L g3362 ( 
.A(n_2615),
.B(n_1635),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_SL g3363 ( 
.A(n_2593),
.B(n_1639),
.Y(n_3363)
);

BUFx4f_ASAP7_75t_L g3364 ( 
.A(n_2777),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_2615),
.Y(n_3365)
);

AND2x6_ASAP7_75t_L g3366 ( 
.A(n_2406),
.B(n_1201),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_2615),
.Y(n_3367)
);

BUFx6f_ASAP7_75t_L g3368 ( 
.A(n_2571),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_2615),
.B(n_1646),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_L g3370 ( 
.A(n_2615),
.B(n_1648),
.Y(n_3370)
);

INVx3_ASAP7_75t_L g3371 ( 
.A(n_2639),
.Y(n_3371)
);

BUFx3_ASAP7_75t_L g3372 ( 
.A(n_2697),
.Y(n_3372)
);

INVx1_ASAP7_75t_L g3373 ( 
.A(n_2615),
.Y(n_3373)
);

INVx4_ASAP7_75t_L g3374 ( 
.A(n_2697),
.Y(n_3374)
);

INVx2_ASAP7_75t_L g3375 ( 
.A(n_2418),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_2615),
.Y(n_3376)
);

AND2x4_ASAP7_75t_L g3377 ( 
.A(n_2615),
.B(n_1483),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_L g3378 ( 
.A(n_2615),
.B(n_1650),
.Y(n_3378)
);

INVx2_ASAP7_75t_L g3379 ( 
.A(n_2418),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_2615),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_2615),
.Y(n_3381)
);

AND2x4_ASAP7_75t_L g3382 ( 
.A(n_2615),
.B(n_1486),
.Y(n_3382)
);

NOR2xp33_ASAP7_75t_L g3383 ( 
.A(n_2513),
.B(n_1651),
.Y(n_3383)
);

NOR2xp33_ASAP7_75t_L g3384 ( 
.A(n_2513),
.B(n_1652),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_2615),
.B(n_1653),
.Y(n_3385)
);

AND2x4_ASAP7_75t_L g3386 ( 
.A(n_2615),
.B(n_1487),
.Y(n_3386)
);

INVx1_ASAP7_75t_SL g3387 ( 
.A(n_2416),
.Y(n_3387)
);

OAI22xp33_ASAP7_75t_SL g3388 ( 
.A1(n_2455),
.A2(n_1656),
.B1(n_1657),
.B2(n_1654),
.Y(n_3388)
);

NOR2xp33_ASAP7_75t_L g3389 ( 
.A(n_2513),
.B(n_1659),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_2615),
.B(n_1660),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_2443),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_2443),
.Y(n_3392)
);

AOI22xp33_ASAP7_75t_L g3393 ( 
.A1(n_2676),
.A2(n_1667),
.B1(n_1669),
.B2(n_1665),
.Y(n_3393)
);

INVx2_ASAP7_75t_SL g3394 ( 
.A(n_2482),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_L g3395 ( 
.A(n_2615),
.B(n_1670),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_2443),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_2443),
.Y(n_3397)
);

INVxp67_ASAP7_75t_L g3398 ( 
.A(n_2416),
.Y(n_3398)
);

INVx1_ASAP7_75t_SL g3399 ( 
.A(n_2416),
.Y(n_3399)
);

NOR2xp33_ASAP7_75t_R g3400 ( 
.A(n_2495),
.B(n_1671),
.Y(n_3400)
);

BUFx3_ASAP7_75t_L g3401 ( 
.A(n_2697),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_2615),
.B(n_1672),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_2443),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_2443),
.Y(n_3404)
);

INVx2_ASAP7_75t_L g3405 ( 
.A(n_2418),
.Y(n_3405)
);

BUFx6f_ASAP7_75t_L g3406 ( 
.A(n_2571),
.Y(n_3406)
);

NOR2xp33_ASAP7_75t_L g3407 ( 
.A(n_2513),
.B(n_1673),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_2443),
.Y(n_3408)
);

INVx1_ASAP7_75t_L g3409 ( 
.A(n_2443),
.Y(n_3409)
);

AND2x2_ASAP7_75t_L g3410 ( 
.A(n_2414),
.B(n_1674),
.Y(n_3410)
);

AND2x6_ASAP7_75t_L g3411 ( 
.A(n_2406),
.B(n_1254),
.Y(n_3411)
);

INVx4_ASAP7_75t_L g3412 ( 
.A(n_2697),
.Y(n_3412)
);

INVxp67_ASAP7_75t_L g3413 ( 
.A(n_2416),
.Y(n_3413)
);

CKINVDCx5p33_ASAP7_75t_R g3414 ( 
.A(n_2495),
.Y(n_3414)
);

AND2x4_ASAP7_75t_L g3415 ( 
.A(n_2615),
.B(n_1491),
.Y(n_3415)
);

NOR2xp33_ASAP7_75t_L g3416 ( 
.A(n_2513),
.B(n_1675),
.Y(n_3416)
);

INVx2_ASAP7_75t_L g3417 ( 
.A(n_2418),
.Y(n_3417)
);

NAND3xp33_ASAP7_75t_L g3418 ( 
.A(n_2455),
.B(n_1703),
.C(n_1702),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_2615),
.B(n_1676),
.Y(n_3419)
);

INVx1_ASAP7_75t_L g3420 ( 
.A(n_2443),
.Y(n_3420)
);

INVx2_ASAP7_75t_SL g3421 ( 
.A(n_2482),
.Y(n_3421)
);

INVx4_ASAP7_75t_SL g3422 ( 
.A(n_2515),
.Y(n_3422)
);

AND2x2_ASAP7_75t_SL g3423 ( 
.A(n_2691),
.B(n_1271),
.Y(n_3423)
);

NOR2xp33_ASAP7_75t_L g3424 ( 
.A(n_2513),
.B(n_1677),
.Y(n_3424)
);

INVx2_ASAP7_75t_L g3425 ( 
.A(n_2418),
.Y(n_3425)
);

BUFx4_ASAP7_75t_L g3426 ( 
.A(n_2785),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_2443),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_2443),
.Y(n_3428)
);

INVx2_ASAP7_75t_L g3429 ( 
.A(n_2418),
.Y(n_3429)
);

INVx2_ASAP7_75t_L g3430 ( 
.A(n_2418),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_L g3431 ( 
.A(n_2615),
.B(n_1678),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_L g3432 ( 
.A(n_2615),
.B(n_1679),
.Y(n_3432)
);

CKINVDCx5p33_ASAP7_75t_R g3433 ( 
.A(n_2495),
.Y(n_3433)
);

NAND3xp33_ASAP7_75t_L g3434 ( 
.A(n_2455),
.B(n_1706),
.C(n_1704),
.Y(n_3434)
);

BUFx2_ASAP7_75t_L g3435 ( 
.A(n_2415),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_2443),
.Y(n_3436)
);

BUFx4f_ASAP7_75t_L g3437 ( 
.A(n_2777),
.Y(n_3437)
);

AND2x2_ASAP7_75t_L g3438 ( 
.A(n_2414),
.B(n_1680),
.Y(n_3438)
);

INVx2_ASAP7_75t_L g3439 ( 
.A(n_2418),
.Y(n_3439)
);

OAI22xp5_ASAP7_75t_L g3440 ( 
.A1(n_2615),
.A2(n_1682),
.B1(n_1685),
.B2(n_1681),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_SL g3441 ( 
.A(n_2593),
.B(n_1687),
.Y(n_3441)
);

INVx2_ASAP7_75t_L g3442 ( 
.A(n_2418),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_SL g3443 ( 
.A(n_2593),
.B(n_1690),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_2443),
.Y(n_3444)
);

BUFx3_ASAP7_75t_L g3445 ( 
.A(n_2697),
.Y(n_3445)
);

BUFx3_ASAP7_75t_L g3446 ( 
.A(n_2697),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_2443),
.Y(n_3447)
);

NOR2xp33_ASAP7_75t_L g3448 ( 
.A(n_2513),
.B(n_1692),
.Y(n_3448)
);

AND2x2_ASAP7_75t_L g3449 ( 
.A(n_2414),
.B(n_1710),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_SL g3450 ( 
.A(n_2593),
.B(n_1713),
.Y(n_3450)
);

OAI22xp5_ASAP7_75t_L g3451 ( 
.A1(n_2615),
.A2(n_1649),
.B1(n_1630),
.B2(n_1271),
.Y(n_3451)
);

NAND2xp33_ASAP7_75t_L g3452 ( 
.A(n_2571),
.B(n_1254),
.Y(n_3452)
);

INVx4_ASAP7_75t_L g3453 ( 
.A(n_2697),
.Y(n_3453)
);

CKINVDCx5p33_ASAP7_75t_R g3454 ( 
.A(n_2495),
.Y(n_3454)
);

INVx4_ASAP7_75t_L g3455 ( 
.A(n_2697),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_L g3456 ( 
.A(n_2797),
.B(n_3118),
.Y(n_3456)
);

NOR2xp33_ASAP7_75t_SL g3457 ( 
.A(n_2922),
.B(n_1114),
.Y(n_3457)
);

AO22x2_ASAP7_75t_L g3458 ( 
.A1(n_2942),
.A2(n_1339),
.B1(n_1346),
.B2(n_1338),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_L g3459 ( 
.A(n_2797),
.B(n_1497),
.Y(n_3459)
);

NOR2xp33_ASAP7_75t_L g3460 ( 
.A(n_2980),
.B(n_1499),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_L g3461 ( 
.A(n_3298),
.B(n_1501),
.Y(n_3461)
);

INVx2_ASAP7_75t_L g3462 ( 
.A(n_2846),
.Y(n_3462)
);

INVx2_ASAP7_75t_L g3463 ( 
.A(n_2865),
.Y(n_3463)
);

NOR2xp67_ASAP7_75t_L g3464 ( 
.A(n_2859),
.B(n_43),
.Y(n_3464)
);

OAI22xp5_ASAP7_75t_L g3465 ( 
.A1(n_2892),
.A2(n_1339),
.B1(n_1346),
.B2(n_1338),
.Y(n_3465)
);

O2A1O1Ixp5_ASAP7_75t_L g3466 ( 
.A1(n_3148),
.A2(n_3272),
.B(n_3157),
.C(n_3270),
.Y(n_3466)
);

INVx1_ASAP7_75t_L g3467 ( 
.A(n_3278),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_L g3468 ( 
.A(n_3298),
.B(n_3311),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_L g3469 ( 
.A(n_3311),
.B(n_1513),
.Y(n_3469)
);

NOR2xp33_ASAP7_75t_L g3470 ( 
.A(n_2839),
.B(n_1521),
.Y(n_3470)
);

INVx2_ASAP7_75t_L g3471 ( 
.A(n_2867),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_L g3472 ( 
.A(n_3377),
.B(n_1535),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_L g3473 ( 
.A(n_3377),
.B(n_1538),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_3382),
.B(n_1540),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_L g3475 ( 
.A(n_3382),
.B(n_1541),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3279),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3280),
.Y(n_3477)
);

NOR2xp33_ASAP7_75t_L g3478 ( 
.A(n_2800),
.B(n_2806),
.Y(n_3478)
);

NOR2xp33_ASAP7_75t_L g3479 ( 
.A(n_2806),
.B(n_1549),
.Y(n_3479)
);

INVx2_ASAP7_75t_L g3480 ( 
.A(n_2868),
.Y(n_3480)
);

INVx2_ASAP7_75t_L g3481 ( 
.A(n_2876),
.Y(n_3481)
);

CKINVDCx5p33_ASAP7_75t_R g3482 ( 
.A(n_2970),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_SL g3483 ( 
.A(n_3349),
.B(n_3423),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_3386),
.B(n_1562),
.Y(n_3484)
);

AOI221xp5_ASAP7_75t_L g3485 ( 
.A1(n_3066),
.A2(n_1580),
.B1(n_1581),
.B2(n_1574),
.C(n_1566),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_L g3486 ( 
.A(n_3386),
.B(n_1585),
.Y(n_3486)
);

OAI22xp5_ASAP7_75t_L g3487 ( 
.A1(n_2962),
.A2(n_1383),
.B1(n_1390),
.B2(n_1358),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3282),
.Y(n_3488)
);

NOR2xp33_ASAP7_75t_L g3489 ( 
.A(n_2991),
.B(n_1588),
.Y(n_3489)
);

NOR2xp33_ASAP7_75t_L g3490 ( 
.A(n_3050),
.B(n_1589),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_3290),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_SL g3492 ( 
.A(n_3286),
.B(n_1254),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_3293),
.Y(n_3493)
);

INVx2_ASAP7_75t_SL g3494 ( 
.A(n_3426),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_SL g3495 ( 
.A(n_3340),
.B(n_1254),
.Y(n_3495)
);

NOR2xp33_ASAP7_75t_L g3496 ( 
.A(n_3015),
.B(n_1608),
.Y(n_3496)
);

NAND3xp33_ASAP7_75t_L g3497 ( 
.A(n_2988),
.B(n_1372),
.C(n_1328),
.Y(n_3497)
);

NOR2xp33_ASAP7_75t_R g3498 ( 
.A(n_2922),
.B(n_1),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_SL g3499 ( 
.A(n_2910),
.B(n_1328),
.Y(n_3499)
);

OR2x2_ASAP7_75t_L g3500 ( 
.A(n_2860),
.B(n_1721),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_L g3501 ( 
.A(n_3415),
.B(n_1611),
.Y(n_3501)
);

NOR2xp33_ASAP7_75t_L g3502 ( 
.A(n_2834),
.B(n_1615),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_SL g3503 ( 
.A(n_3178),
.B(n_1328),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_3415),
.B(n_1616),
.Y(n_3504)
);

BUFx6f_ASAP7_75t_L g3505 ( 
.A(n_2817),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_SL g3506 ( 
.A(n_2947),
.B(n_1328),
.Y(n_3506)
);

NAND3xp33_ASAP7_75t_L g3507 ( 
.A(n_3026),
.B(n_1536),
.C(n_1372),
.Y(n_3507)
);

INVx2_ASAP7_75t_SL g3508 ( 
.A(n_3364),
.Y(n_3508)
);

INVx2_ASAP7_75t_L g3509 ( 
.A(n_2900),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_L g3510 ( 
.A(n_2878),
.B(n_1624),
.Y(n_3510)
);

INVx2_ASAP7_75t_L g3511 ( 
.A(n_2903),
.Y(n_3511)
);

A2O1A1Ixp33_ASAP7_75t_L g3512 ( 
.A1(n_3094),
.A2(n_2818),
.B(n_2813),
.C(n_2856),
.Y(n_3512)
);

O2A1O1Ixp33_ASAP7_75t_L g3513 ( 
.A1(n_2836),
.A2(n_1633),
.B(n_1636),
.C(n_1628),
.Y(n_3513)
);

HB1xp67_ASAP7_75t_L g3514 ( 
.A(n_2808),
.Y(n_3514)
);

NOR2xp33_ASAP7_75t_L g3515 ( 
.A(n_2909),
.B(n_1638),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3295),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_SL g3517 ( 
.A(n_2947),
.B(n_3222),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_L g3518 ( 
.A(n_2878),
.B(n_1641),
.Y(n_3518)
);

NAND3xp33_ASAP7_75t_L g3519 ( 
.A(n_3031),
.B(n_1536),
.C(n_1372),
.Y(n_3519)
);

AO221x1_ASAP7_75t_L g3520 ( 
.A1(n_2962),
.A2(n_1372),
.B1(n_1640),
.B2(n_1578),
.C(n_1536),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_3076),
.B(n_1642),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3305),
.Y(n_3522)
);

BUFx6f_ASAP7_75t_L g3523 ( 
.A(n_2817),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3308),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3309),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_3316),
.Y(n_3526)
);

NAND2xp33_ASAP7_75t_L g3527 ( 
.A(n_3084),
.B(n_1536),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_3323),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3327),
.Y(n_3529)
);

HB1xp67_ASAP7_75t_L g3530 ( 
.A(n_3304),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_3079),
.B(n_1644),
.Y(n_3531)
);

INVx3_ASAP7_75t_L g3532 ( 
.A(n_3084),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3329),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_L g3534 ( 
.A(n_3334),
.B(n_1645),
.Y(n_3534)
);

NAND2xp5_ASAP7_75t_L g3535 ( 
.A(n_3336),
.B(n_1655),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_SL g3536 ( 
.A(n_2926),
.B(n_1578),
.Y(n_3536)
);

AOI22xp5_ASAP7_75t_L g3537 ( 
.A1(n_2902),
.A2(n_1662),
.B1(n_1663),
.B2(n_1658),
.Y(n_3537)
);

OAI22xp33_ASAP7_75t_L g3538 ( 
.A1(n_2968),
.A2(n_1684),
.B1(n_1694),
.B2(n_1664),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_3343),
.Y(n_3539)
);

NOR2xp67_ASAP7_75t_SL g3540 ( 
.A(n_2953),
.B(n_1151),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3356),
.Y(n_3541)
);

AOI21xp5_ASAP7_75t_L g3542 ( 
.A1(n_2937),
.A2(n_1383),
.B(n_1358),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_3365),
.Y(n_3543)
);

OR2x2_ASAP7_75t_L g3544 ( 
.A(n_2887),
.B(n_1696),
.Y(n_3544)
);

NOR2xp67_ASAP7_75t_L g3545 ( 
.A(n_2859),
.B(n_43),
.Y(n_3545)
);

INVx2_ASAP7_75t_L g3546 ( 
.A(n_2916),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_3367),
.B(n_1699),
.Y(n_3547)
);

INVx1_ASAP7_75t_SL g3548 ( 
.A(n_2889),
.Y(n_3548)
);

INVxp67_ASAP7_75t_L g3549 ( 
.A(n_3284),
.Y(n_3549)
);

NOR2xp33_ASAP7_75t_L g3550 ( 
.A(n_3063),
.B(n_1700),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_SL g3551 ( 
.A(n_2880),
.B(n_1578),
.Y(n_3551)
);

INVx2_ASAP7_75t_SL g3552 ( 
.A(n_3364),
.Y(n_3552)
);

NOR2xp33_ASAP7_75t_L g3553 ( 
.A(n_2918),
.B(n_1715),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_3373),
.Y(n_3554)
);

NOR2xp67_ASAP7_75t_L g3555 ( 
.A(n_3171),
.B(n_43),
.Y(n_3555)
);

AOI22xp33_ASAP7_75t_L g3556 ( 
.A1(n_3103),
.A2(n_1640),
.B1(n_1668),
.B2(n_1578),
.Y(n_3556)
);

INVxp67_ASAP7_75t_L g3557 ( 
.A(n_3326),
.Y(n_3557)
);

NOR2xp33_ASAP7_75t_L g3558 ( 
.A(n_3339),
.B(n_1722),
.Y(n_3558)
);

AOI22xp33_ASAP7_75t_L g3559 ( 
.A1(n_3103),
.A2(n_1668),
.B1(n_1695),
.B2(n_1640),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3376),
.Y(n_3560)
);

INVxp67_ASAP7_75t_L g3561 ( 
.A(n_3345),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_SL g3562 ( 
.A(n_2882),
.B(n_1640),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_SL g3563 ( 
.A(n_2882),
.B(n_1668),
.Y(n_3563)
);

AND2x4_ASAP7_75t_L g3564 ( 
.A(n_3380),
.B(n_1390),
.Y(n_3564)
);

INVx2_ASAP7_75t_L g3565 ( 
.A(n_2928),
.Y(n_3565)
);

INVx2_ASAP7_75t_SL g3566 ( 
.A(n_3437),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3381),
.Y(n_3567)
);

AND2x2_ASAP7_75t_L g3568 ( 
.A(n_3315),
.B(n_1464),
.Y(n_3568)
);

NOR2xp33_ASAP7_75t_SL g3569 ( 
.A(n_3437),
.B(n_1233),
.Y(n_3569)
);

AOI22xp5_ASAP7_75t_L g3570 ( 
.A1(n_3451),
.A2(n_1485),
.B1(n_1507),
.B2(n_1464),
.Y(n_3570)
);

BUFx6f_ASAP7_75t_L g3571 ( 
.A(n_2817),
.Y(n_3571)
);

NOR2xp33_ASAP7_75t_L g3572 ( 
.A(n_2958),
.B(n_1485),
.Y(n_3572)
);

INVx3_ASAP7_75t_L g3573 ( 
.A(n_3084),
.Y(n_3573)
);

NOR3xp33_ASAP7_75t_L g3574 ( 
.A(n_3041),
.B(n_1554),
.C(n_1507),
.Y(n_3574)
);

BUFx3_ASAP7_75t_L g3575 ( 
.A(n_2819),
.Y(n_3575)
);

INVx2_ASAP7_75t_L g3576 ( 
.A(n_2941),
.Y(n_3576)
);

INVx2_ASAP7_75t_L g3577 ( 
.A(n_2950),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_SL g3578 ( 
.A(n_2882),
.B(n_1668),
.Y(n_3578)
);

INVx1_ASAP7_75t_L g3579 ( 
.A(n_2835),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_2798),
.B(n_1554),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_SL g3581 ( 
.A(n_2981),
.B(n_1695),
.Y(n_3581)
);

INVxp67_ASAP7_75t_L g3582 ( 
.A(n_3322),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_2798),
.B(n_1563),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_2837),
.Y(n_3584)
);

NAND2xp5_ASAP7_75t_SL g3585 ( 
.A(n_2981),
.B(n_1695),
.Y(n_3585)
);

INVx2_ASAP7_75t_L g3586 ( 
.A(n_2952),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_2805),
.B(n_1563),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_2849),
.Y(n_3588)
);

AOI21xp5_ASAP7_75t_L g3589 ( 
.A1(n_2973),
.A2(n_2954),
.B(n_3141),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_2805),
.B(n_1599),
.Y(n_3590)
);

INVx1_ASAP7_75t_L g3591 ( 
.A(n_2850),
.Y(n_3591)
);

NOR3xp33_ASAP7_75t_L g3592 ( 
.A(n_2821),
.B(n_1625),
.C(n_1599),
.Y(n_3592)
);

INVxp67_ASAP7_75t_L g3593 ( 
.A(n_3065),
.Y(n_3593)
);

OR2x6_ASAP7_75t_L g3594 ( 
.A(n_2968),
.B(n_3016),
.Y(n_3594)
);

INVx3_ASAP7_75t_L g3595 ( 
.A(n_3084),
.Y(n_3595)
);

INVx1_ASAP7_75t_L g3596 ( 
.A(n_2863),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_L g3597 ( 
.A(n_2810),
.B(n_2812),
.Y(n_3597)
);

INVx2_ASAP7_75t_SL g3598 ( 
.A(n_2981),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_SL g3599 ( 
.A(n_3344),
.B(n_1695),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_SL g3600 ( 
.A(n_3350),
.B(n_1625),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_L g3601 ( 
.A(n_2810),
.B(n_1627),
.Y(n_3601)
);

INVx2_ASAP7_75t_L g3602 ( 
.A(n_2963),
.Y(n_3602)
);

INVxp33_ASAP7_75t_L g3603 ( 
.A(n_3400),
.Y(n_3603)
);

AND2x2_ASAP7_75t_L g3604 ( 
.A(n_3354),
.B(n_1627),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_L g3605 ( 
.A(n_2812),
.B(n_44),
.Y(n_3605)
);

INVx2_ASAP7_75t_L g3606 ( 
.A(n_2989),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_SL g3607 ( 
.A(n_3387),
.B(n_44),
.Y(n_3607)
);

O2A1O1Ixp5_ASAP7_75t_L g3608 ( 
.A1(n_3243),
.A2(n_45),
.B(n_46),
.C(n_44),
.Y(n_3608)
);

AOI22xp33_ASAP7_75t_L g3609 ( 
.A1(n_3294),
.A2(n_47),
.B1(n_49),
.B2(n_46),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_2885),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_SL g3611 ( 
.A(n_3399),
.B(n_46),
.Y(n_3611)
);

BUFx2_ASAP7_75t_L g3612 ( 
.A(n_3306),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_2894),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_2895),
.Y(n_3614)
);

NOR2xp33_ASAP7_75t_L g3615 ( 
.A(n_2971),
.B(n_49),
.Y(n_3615)
);

AND2x2_ASAP7_75t_L g3616 ( 
.A(n_3358),
.B(n_49),
.Y(n_3616)
);

NAND2xp5_ASAP7_75t_L g3617 ( 
.A(n_2829),
.B(n_50),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_2897),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_SL g3619 ( 
.A(n_3078),
.B(n_50),
.Y(n_3619)
);

INVx1_ASAP7_75t_SL g3620 ( 
.A(n_2820),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_SL g3621 ( 
.A(n_3228),
.B(n_50),
.Y(n_3621)
);

NOR2xp67_ASAP7_75t_L g3622 ( 
.A(n_3171),
.B(n_51),
.Y(n_3622)
);

NAND2xp5_ASAP7_75t_SL g3623 ( 
.A(n_2921),
.B(n_51),
.Y(n_3623)
);

INVx4_ASAP7_75t_L g3624 ( 
.A(n_2801),
.Y(n_3624)
);

INVx1_ASAP7_75t_L g3625 ( 
.A(n_2911),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_SL g3626 ( 
.A(n_2921),
.B(n_3388),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_2912),
.Y(n_3627)
);

BUFx8_ASAP7_75t_L g3628 ( 
.A(n_2847),
.Y(n_3628)
);

AOI22xp5_ASAP7_75t_L g3629 ( 
.A1(n_2838),
.A2(n_1066),
.B1(n_1067),
.B2(n_1065),
.Y(n_3629)
);

BUFx3_ASAP7_75t_L g3630 ( 
.A(n_3332),
.Y(n_3630)
);

AOI22xp5_ASAP7_75t_L g3631 ( 
.A1(n_3045),
.A2(n_1066),
.B1(n_1067),
.B2(n_1065),
.Y(n_3631)
);

BUFx8_ASAP7_75t_L g3632 ( 
.A(n_3435),
.Y(n_3632)
);

INVx2_ASAP7_75t_L g3633 ( 
.A(n_2993),
.Y(n_3633)
);

AOI22xp33_ASAP7_75t_L g3634 ( 
.A1(n_3302),
.A2(n_53),
.B1(n_54),
.B2(n_52),
.Y(n_3634)
);

BUFx4f_ASAP7_75t_L g3635 ( 
.A(n_3016),
.Y(n_3635)
);

NOR2xp33_ASAP7_75t_L g3636 ( 
.A(n_3218),
.B(n_52),
.Y(n_3636)
);

INVxp67_ASAP7_75t_SL g3637 ( 
.A(n_3281),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_SL g3638 ( 
.A(n_3267),
.B(n_52),
.Y(n_3638)
);

NAND2xp5_ASAP7_75t_SL g3639 ( 
.A(n_2935),
.B(n_53),
.Y(n_3639)
);

NOR2xp67_ASAP7_75t_L g3640 ( 
.A(n_3171),
.B(n_54),
.Y(n_3640)
);

INVx2_ASAP7_75t_L g3641 ( 
.A(n_2994),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_SL g3642 ( 
.A(n_3024),
.B(n_54),
.Y(n_3642)
);

NAND2xp5_ASAP7_75t_L g3643 ( 
.A(n_2829),
.B(n_55),
.Y(n_3643)
);

AND2x6_ASAP7_75t_L g3644 ( 
.A(n_2831),
.B(n_55),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_L g3645 ( 
.A(n_2831),
.B(n_56),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_2929),
.Y(n_3646)
);

OR2x2_ASAP7_75t_SL g3647 ( 
.A(n_3010),
.B(n_56),
.Y(n_3647)
);

OR2x2_ASAP7_75t_L g3648 ( 
.A(n_3068),
.B(n_56),
.Y(n_3648)
);

INVx2_ASAP7_75t_L g3649 ( 
.A(n_3002),
.Y(n_3649)
);

INVx2_ASAP7_75t_SL g3650 ( 
.A(n_3010),
.Y(n_3650)
);

INVxp67_ASAP7_75t_L g3651 ( 
.A(n_3068),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_3061),
.Y(n_3652)
);

INVx1_ASAP7_75t_L g3653 ( 
.A(n_3064),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_SL g3654 ( 
.A(n_3342),
.B(n_3087),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3073),
.Y(n_3655)
);

NOR2xp33_ASAP7_75t_L g3656 ( 
.A(n_3313),
.B(n_3355),
.Y(n_3656)
);

INVx3_ASAP7_75t_L g3657 ( 
.A(n_3160),
.Y(n_3657)
);

INVx1_ASAP7_75t_L g3658 ( 
.A(n_3060),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_L g3659 ( 
.A(n_2832),
.B(n_57),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3060),
.Y(n_3660)
);

AO22x2_ASAP7_75t_L g3661 ( 
.A1(n_3005),
.A2(n_58),
.B1(n_59),
.B2(n_57),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_L g3662 ( 
.A(n_2832),
.B(n_57),
.Y(n_3662)
);

O2A1O1Ixp33_ASAP7_75t_L g3663 ( 
.A1(n_3059),
.A2(n_59),
.B(n_60),
.C(n_58),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3133),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_3136),
.Y(n_3665)
);

AOI221xp5_ASAP7_75t_L g3666 ( 
.A1(n_3037),
.A2(n_61),
.B1(n_62),
.B2(n_60),
.C(n_58),
.Y(n_3666)
);

AND2x4_ASAP7_75t_L g3667 ( 
.A(n_2944),
.B(n_61),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_2944),
.B(n_61),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_L g3669 ( 
.A(n_2946),
.B(n_63),
.Y(n_3669)
);

INVx8_ASAP7_75t_L g3670 ( 
.A(n_3167),
.Y(n_3670)
);

NAND3xp33_ASAP7_75t_L g3671 ( 
.A(n_3383),
.B(n_64),
.C(n_63),
.Y(n_3671)
);

NAND2xp33_ASAP7_75t_L g3672 ( 
.A(n_2814),
.B(n_2881),
.Y(n_3672)
);

AND2x2_ASAP7_75t_L g3673 ( 
.A(n_3410),
.B(n_63),
.Y(n_3673)
);

AND2x2_ASAP7_75t_L g3674 ( 
.A(n_3438),
.B(n_64),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_L g3675 ( 
.A(n_2946),
.B(n_2949),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_2949),
.B(n_65),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_L g3677 ( 
.A(n_2955),
.B(n_66),
.Y(n_3677)
);

NAND2xp5_ASAP7_75t_L g3678 ( 
.A(n_2955),
.B(n_66),
.Y(n_3678)
);

NAND2xp33_ASAP7_75t_L g3679 ( 
.A(n_2814),
.B(n_67),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3149),
.Y(n_3680)
);

AND2x4_ASAP7_75t_L g3681 ( 
.A(n_3014),
.B(n_67),
.Y(n_3681)
);

INVx2_ASAP7_75t_SL g3682 ( 
.A(n_3372),
.Y(n_3682)
);

NOR3xp33_ASAP7_75t_L g3683 ( 
.A(n_3384),
.B(n_68),
.C(n_67),
.Y(n_3683)
);

INVx3_ASAP7_75t_L g3684 ( 
.A(n_3160),
.Y(n_3684)
);

NOR2xp67_ASAP7_75t_L g3685 ( 
.A(n_3173),
.B(n_68),
.Y(n_3685)
);

NAND2xp33_ASAP7_75t_L g3686 ( 
.A(n_2814),
.B(n_68),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_3150),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_L g3688 ( 
.A(n_3014),
.B(n_69),
.Y(n_3688)
);

OAI22xp33_ASAP7_75t_SL g3689 ( 
.A1(n_3306),
.A2(n_70),
.B1(n_71),
.B2(n_69),
.Y(n_3689)
);

NAND2xp5_ASAP7_75t_SL g3690 ( 
.A(n_3087),
.B(n_69),
.Y(n_3690)
);

NAND2xp33_ASAP7_75t_L g3691 ( 
.A(n_2814),
.B(n_70),
.Y(n_3691)
);

INVx2_ASAP7_75t_L g3692 ( 
.A(n_3027),
.Y(n_3692)
);

INVx2_ASAP7_75t_L g3693 ( 
.A(n_3021),
.Y(n_3693)
);

AOI22xp33_ASAP7_75t_L g3694 ( 
.A1(n_3389),
.A2(n_72),
.B1(n_73),
.B2(n_71),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_L g3695 ( 
.A(n_3021),
.B(n_72),
.Y(n_3695)
);

NOR3xp33_ASAP7_75t_L g3696 ( 
.A(n_3407),
.B(n_74),
.C(n_73),
.Y(n_3696)
);

NAND2xp5_ASAP7_75t_L g3697 ( 
.A(n_3022),
.B(n_74),
.Y(n_3697)
);

INVxp33_ASAP7_75t_L g3698 ( 
.A(n_2995),
.Y(n_3698)
);

CKINVDCx20_ASAP7_75t_R g3699 ( 
.A(n_3104),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_L g3700 ( 
.A(n_3022),
.B(n_74),
.Y(n_3700)
);

AOI22xp5_ASAP7_75t_L g3701 ( 
.A1(n_3181),
.A2(n_1074),
.B1(n_1075),
.B2(n_1073),
.Y(n_3701)
);

INVx2_ASAP7_75t_SL g3702 ( 
.A(n_3401),
.Y(n_3702)
);

NOR2xp33_ASAP7_75t_L g3703 ( 
.A(n_3416),
.B(n_75),
.Y(n_3703)
);

INVx2_ASAP7_75t_L g3704 ( 
.A(n_3025),
.Y(n_3704)
);

NAND2xp5_ASAP7_75t_L g3705 ( 
.A(n_3025),
.B(n_75),
.Y(n_3705)
);

NOR2xp33_ASAP7_75t_L g3706 ( 
.A(n_3424),
.B(n_76),
.Y(n_3706)
);

INVx2_ASAP7_75t_SL g3707 ( 
.A(n_3445),
.Y(n_3707)
);

NOR2xp33_ASAP7_75t_L g3708 ( 
.A(n_3448),
.B(n_76),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_SL g3709 ( 
.A(n_3156),
.B(n_77),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3150),
.Y(n_3710)
);

NOR2xp33_ASAP7_75t_L g3711 ( 
.A(n_3151),
.B(n_77),
.Y(n_3711)
);

INVxp67_ASAP7_75t_L g3712 ( 
.A(n_3179),
.Y(n_3712)
);

NOR2xp33_ASAP7_75t_L g3713 ( 
.A(n_2830),
.B(n_2907),
.Y(n_3713)
);

OAI22xp33_ASAP7_75t_L g3714 ( 
.A1(n_3348),
.A2(n_78),
.B1(n_79),
.B2(n_77),
.Y(n_3714)
);

AND2x4_ASAP7_75t_L g3715 ( 
.A(n_3030),
.B(n_78),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_L g3716 ( 
.A(n_3030),
.B(n_78),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_L g3717 ( 
.A(n_3391),
.B(n_79),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3165),
.Y(n_3718)
);

NAND2xp5_ASAP7_75t_L g3719 ( 
.A(n_3391),
.B(n_79),
.Y(n_3719)
);

INVx1_ASAP7_75t_L g3720 ( 
.A(n_3165),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_3177),
.Y(n_3721)
);

NOR2xp33_ASAP7_75t_L g3722 ( 
.A(n_2915),
.B(n_80),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_SL g3723 ( 
.A(n_3194),
.B(n_80),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3177),
.Y(n_3724)
);

INVxp67_ASAP7_75t_L g3725 ( 
.A(n_2826),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3180),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_SL g3727 ( 
.A(n_3194),
.B(n_80),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_L g3728 ( 
.A(n_3392),
.B(n_81),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_L g3729 ( 
.A(n_3392),
.B(n_81),
.Y(n_3729)
);

INVx2_ASAP7_75t_L g3730 ( 
.A(n_3396),
.Y(n_3730)
);

INVx2_ASAP7_75t_L g3731 ( 
.A(n_3396),
.Y(n_3731)
);

NAND2xp5_ASAP7_75t_L g3732 ( 
.A(n_3397),
.B(n_82),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_3180),
.Y(n_3733)
);

BUFx3_ASAP7_75t_L g3734 ( 
.A(n_3446),
.Y(n_3734)
);

NAND2xp5_ASAP7_75t_L g3735 ( 
.A(n_3397),
.B(n_82),
.Y(n_3735)
);

INVx2_ASAP7_75t_SL g3736 ( 
.A(n_2842),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_3403),
.B(n_83),
.Y(n_3737)
);

AOI22xp5_ASAP7_75t_L g3738 ( 
.A1(n_3006),
.A2(n_84),
.B1(n_85),
.B2(n_83),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3186),
.Y(n_3739)
);

INVx2_ASAP7_75t_L g3740 ( 
.A(n_3403),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_3404),
.B(n_84),
.Y(n_3741)
);

AND2x6_ASAP7_75t_SL g3742 ( 
.A(n_3067),
.B(n_0),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_3404),
.B(n_84),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3186),
.Y(n_3744)
);

NAND2xp5_ASAP7_75t_L g3745 ( 
.A(n_3408),
.B(n_85),
.Y(n_3745)
);

CKINVDCx5p33_ASAP7_75t_R g3746 ( 
.A(n_2869),
.Y(n_3746)
);

INVxp67_ASAP7_75t_L g3747 ( 
.A(n_3449),
.Y(n_3747)
);

INVx3_ASAP7_75t_L g3748 ( 
.A(n_3160),
.Y(n_3748)
);

NAND2xp5_ASAP7_75t_L g3749 ( 
.A(n_3408),
.B(n_85),
.Y(n_3749)
);

INVx2_ASAP7_75t_L g3750 ( 
.A(n_3409),
.Y(n_3750)
);

NAND2xp33_ASAP7_75t_L g3751 ( 
.A(n_2881),
.B(n_86),
.Y(n_3751)
);

AND2x2_ASAP7_75t_SL g3752 ( 
.A(n_2851),
.B(n_86),
.Y(n_3752)
);

O2A1O1Ixp5_ASAP7_75t_L g3753 ( 
.A1(n_3159),
.A2(n_3114),
.B(n_3263),
.C(n_3274),
.Y(n_3753)
);

INVx2_ASAP7_75t_L g3754 ( 
.A(n_3409),
.Y(n_3754)
);

NAND2xp33_ASAP7_75t_SL g3755 ( 
.A(n_2919),
.B(n_86),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3032),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3033),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_SL g3758 ( 
.A(n_3194),
.B(n_87),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3070),
.Y(n_3759)
);

AND2x2_ASAP7_75t_L g3760 ( 
.A(n_2875),
.B(n_87),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3072),
.Y(n_3761)
);

INVx2_ASAP7_75t_SL g3762 ( 
.A(n_2862),
.Y(n_3762)
);

OR2x2_ASAP7_75t_L g3763 ( 
.A(n_3398),
.B(n_87),
.Y(n_3763)
);

NAND2xp5_ASAP7_75t_L g3764 ( 
.A(n_3420),
.B(n_88),
.Y(n_3764)
);

INVx2_ASAP7_75t_L g3765 ( 
.A(n_3420),
.Y(n_3765)
);

NOR2xp33_ASAP7_75t_L g3766 ( 
.A(n_3202),
.B(n_88),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_SL g3767 ( 
.A(n_3277),
.B(n_88),
.Y(n_3767)
);

INVxp67_ASAP7_75t_L g3768 ( 
.A(n_2884),
.Y(n_3768)
);

INVx4_ASAP7_75t_L g3769 ( 
.A(n_2801),
.Y(n_3769)
);

NAND2xp33_ASAP7_75t_L g3770 ( 
.A(n_2881),
.B(n_2959),
.Y(n_3770)
);

NAND2xp5_ASAP7_75t_L g3771 ( 
.A(n_3427),
.B(n_89),
.Y(n_3771)
);

AND2x2_ASAP7_75t_L g3772 ( 
.A(n_2923),
.B(n_2864),
.Y(n_3772)
);

NAND2xp5_ASAP7_75t_L g3773 ( 
.A(n_3427),
.B(n_3428),
.Y(n_3773)
);

AO22x2_ASAP7_75t_L g3774 ( 
.A1(n_2794),
.A2(n_90),
.B1(n_91),
.B2(n_89),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_3428),
.B(n_89),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_SL g3776 ( 
.A(n_3418),
.B(n_90),
.Y(n_3776)
);

INVx2_ASAP7_75t_L g3777 ( 
.A(n_3436),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3075),
.Y(n_3778)
);

INVx1_ASAP7_75t_L g3779 ( 
.A(n_3216),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_3436),
.B(n_90),
.Y(n_3780)
);

AOI22xp5_ASAP7_75t_L g3781 ( 
.A1(n_3012),
.A2(n_92),
.B1(n_93),
.B2(n_91),
.Y(n_3781)
);

INVx1_ASAP7_75t_L g3782 ( 
.A(n_3217),
.Y(n_3782)
);

AOI21xp5_ASAP7_75t_L g3783 ( 
.A1(n_3197),
.A2(n_93),
.B(n_92),
.Y(n_3783)
);

OAI221xp5_ASAP7_75t_L g3784 ( 
.A1(n_2990),
.A2(n_95),
.B1(n_96),
.B2(n_94),
.C(n_92),
.Y(n_3784)
);

INVx2_ASAP7_75t_L g3785 ( 
.A(n_3444),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_L g3786 ( 
.A(n_3444),
.B(n_95),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3034),
.Y(n_3787)
);

BUFx5_ASAP7_75t_L g3788 ( 
.A(n_3077),
.Y(n_3788)
);

NAND2xp5_ASAP7_75t_L g3789 ( 
.A(n_3447),
.B(n_95),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3034),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_L g3791 ( 
.A(n_3447),
.B(n_96),
.Y(n_3791)
);

NOR2xp67_ASAP7_75t_L g3792 ( 
.A(n_3173),
.B(n_96),
.Y(n_3792)
);

INVx2_ASAP7_75t_L g3793 ( 
.A(n_2871),
.Y(n_3793)
);

BUFx6f_ASAP7_75t_L g3794 ( 
.A(n_2888),
.Y(n_3794)
);

NAND2xp5_ASAP7_75t_L g3795 ( 
.A(n_2877),
.B(n_97),
.Y(n_3795)
);

AOI22xp5_ASAP7_75t_L g3796 ( 
.A1(n_3017),
.A2(n_98),
.B1(n_99),
.B2(n_97),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_SL g3797 ( 
.A(n_3434),
.B(n_3413),
.Y(n_3797)
);

NOR2xp33_ASAP7_75t_L g3798 ( 
.A(n_3210),
.B(n_3099),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_L g3799 ( 
.A(n_2879),
.B(n_97),
.Y(n_3799)
);

INVx3_ASAP7_75t_L g3800 ( 
.A(n_3160),
.Y(n_3800)
);

NAND2xp5_ASAP7_75t_L g3801 ( 
.A(n_2883),
.B(n_2930),
.Y(n_3801)
);

INVx4_ASAP7_75t_L g3802 ( 
.A(n_3320),
.Y(n_3802)
);

NAND2xp33_ASAP7_75t_SL g3803 ( 
.A(n_2919),
.B(n_98),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_2932),
.B(n_99),
.Y(n_3804)
);

NAND2xp5_ASAP7_75t_SL g3805 ( 
.A(n_3191),
.B(n_100),
.Y(n_3805)
);

BUFx6f_ASAP7_75t_SL g3806 ( 
.A(n_2862),
.Y(n_3806)
);

OR2x6_ASAP7_75t_L g3807 ( 
.A(n_3348),
.B(n_100),
.Y(n_3807)
);

INVx2_ASAP7_75t_L g3808 ( 
.A(n_2936),
.Y(n_3808)
);

NAND2xp5_ASAP7_75t_SL g3809 ( 
.A(n_3191),
.B(n_100),
.Y(n_3809)
);

NOR2xp33_ASAP7_75t_L g3810 ( 
.A(n_2917),
.B(n_102),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_SL g3811 ( 
.A(n_3191),
.B(n_102),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_SL g3812 ( 
.A(n_3018),
.B(n_103),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3038),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_L g3814 ( 
.A(n_2938),
.B(n_103),
.Y(n_3814)
);

NAND2xp5_ASAP7_75t_L g3815 ( 
.A(n_2956),
.B(n_103),
.Y(n_3815)
);

NAND2xp5_ASAP7_75t_L g3816 ( 
.A(n_2961),
.B(n_104),
.Y(n_3816)
);

NOR2xp33_ASAP7_75t_L g3817 ( 
.A(n_3176),
.B(n_104),
.Y(n_3817)
);

NAND2xp5_ASAP7_75t_L g3818 ( 
.A(n_2967),
.B(n_105),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_SL g3819 ( 
.A(n_2825),
.B(n_105),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_2969),
.B(n_106),
.Y(n_3820)
);

HB1xp67_ASAP7_75t_L g3821 ( 
.A(n_3000),
.Y(n_3821)
);

NAND2xp5_ASAP7_75t_L g3822 ( 
.A(n_2972),
.B(n_2974),
.Y(n_3822)
);

INVx2_ASAP7_75t_L g3823 ( 
.A(n_2986),
.Y(n_3823)
);

BUFx6f_ASAP7_75t_L g3824 ( 
.A(n_2888),
.Y(n_3824)
);

CKINVDCx5p33_ASAP7_75t_R g3825 ( 
.A(n_2803),
.Y(n_3825)
);

NAND2xp5_ASAP7_75t_L g3826 ( 
.A(n_2998),
.B(n_3001),
.Y(n_3826)
);

INVx2_ASAP7_75t_L g3827 ( 
.A(n_3008),
.Y(n_3827)
);

NAND2xp5_ASAP7_75t_SL g3828 ( 
.A(n_2825),
.B(n_106),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_3092),
.B(n_107),
.Y(n_3829)
);

NAND2xp33_ASAP7_75t_L g3830 ( 
.A(n_2881),
.B(n_107),
.Y(n_3830)
);

NOR2xp33_ASAP7_75t_L g3831 ( 
.A(n_2943),
.B(n_108),
.Y(n_3831)
);

INVx2_ASAP7_75t_L g3832 ( 
.A(n_3038),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_SL g3833 ( 
.A(n_2840),
.B(n_108),
.Y(n_3833)
);

NOR2xp33_ASAP7_75t_L g3834 ( 
.A(n_3007),
.B(n_108),
.Y(n_3834)
);

NAND2xp5_ASAP7_75t_L g3835 ( 
.A(n_2840),
.B(n_109),
.Y(n_3835)
);

INVx2_ASAP7_75t_L g3836 ( 
.A(n_3040),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_2815),
.B(n_109),
.Y(n_3837)
);

INVx2_ASAP7_75t_L g3838 ( 
.A(n_3040),
.Y(n_3838)
);

O2A1O1Ixp5_ASAP7_75t_L g3839 ( 
.A1(n_2992),
.A2(n_111),
.B(n_112),
.C(n_110),
.Y(n_3839)
);

BUFx6f_ASAP7_75t_L g3840 ( 
.A(n_2888),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_2815),
.B(n_2890),
.Y(n_3841)
);

NOR2xp33_ASAP7_75t_L g3842 ( 
.A(n_3042),
.B(n_110),
.Y(n_3842)
);

AOI22xp33_ASAP7_75t_L g3843 ( 
.A1(n_3212),
.A2(n_111),
.B1(n_112),
.B2(n_110),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3049),
.Y(n_3844)
);

INVx2_ASAP7_75t_SL g3845 ( 
.A(n_3320),
.Y(n_3845)
);

NAND2xp5_ASAP7_75t_L g3846 ( 
.A(n_2890),
.B(n_111),
.Y(n_3846)
);

OAI22xp5_ASAP7_75t_SL g3847 ( 
.A1(n_3067),
.A2(n_2948),
.B1(n_3013),
.B2(n_2811),
.Y(n_3847)
);

INVx1_ASAP7_75t_L g3848 ( 
.A(n_3049),
.Y(n_3848)
);

NAND2xp5_ASAP7_75t_SL g3849 ( 
.A(n_2851),
.B(n_112),
.Y(n_3849)
);

INVx1_ASAP7_75t_L g3850 ( 
.A(n_3055),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_L g3851 ( 
.A(n_2893),
.B(n_113),
.Y(n_3851)
);

INVx2_ASAP7_75t_SL g3852 ( 
.A(n_3341),
.Y(n_3852)
);

NOR2xp33_ASAP7_75t_L g3853 ( 
.A(n_2823),
.B(n_113),
.Y(n_3853)
);

NAND2xp5_ASAP7_75t_SL g3854 ( 
.A(n_3173),
.B(n_113),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_L g3855 ( 
.A(n_2893),
.B(n_114),
.Y(n_3855)
);

INVx2_ASAP7_75t_L g3856 ( 
.A(n_3055),
.Y(n_3856)
);

INVx2_ASAP7_75t_L g3857 ( 
.A(n_3135),
.Y(n_3857)
);

AOI22xp5_ASAP7_75t_L g3858 ( 
.A1(n_2855),
.A2(n_115),
.B1(n_116),
.B2(n_114),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_3086),
.Y(n_3859)
);

HB1xp67_ASAP7_75t_L g3860 ( 
.A(n_3004),
.Y(n_3860)
);

INVx2_ASAP7_75t_L g3861 ( 
.A(n_3138),
.Y(n_3861)
);

OAI22xp5_ASAP7_75t_L g3862 ( 
.A1(n_2899),
.A2(n_116),
.B1(n_117),
.B2(n_115),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_L g3863 ( 
.A(n_3098),
.B(n_3109),
.Y(n_3863)
);

INVx2_ASAP7_75t_L g3864 ( 
.A(n_3185),
.Y(n_3864)
);

INVx2_ASAP7_75t_SL g3865 ( 
.A(n_3341),
.Y(n_3865)
);

AOI21xp5_ASAP7_75t_L g3866 ( 
.A1(n_3257),
.A2(n_117),
.B(n_115),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3088),
.Y(n_3867)
);

AOI22xp33_ASAP7_75t_L g3868 ( 
.A1(n_3023),
.A2(n_2833),
.B1(n_2852),
.B2(n_3052),
.Y(n_3868)
);

NAND2xp33_ASAP7_75t_L g3869 ( 
.A(n_2959),
.B(n_118),
.Y(n_3869)
);

INVx1_ASAP7_75t_L g3870 ( 
.A(n_3090),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_3100),
.Y(n_3871)
);

INVxp67_ASAP7_75t_L g3872 ( 
.A(n_2853),
.Y(n_3872)
);

INVx2_ASAP7_75t_L g3873 ( 
.A(n_3192),
.Y(n_3873)
);

NAND2xp5_ASAP7_75t_SL g3874 ( 
.A(n_3254),
.B(n_118),
.Y(n_3874)
);

INVx8_ASAP7_75t_L g3875 ( 
.A(n_3167),
.Y(n_3875)
);

INVx1_ASAP7_75t_L g3876 ( 
.A(n_3111),
.Y(n_3876)
);

INVx2_ASAP7_75t_L g3877 ( 
.A(n_3195),
.Y(n_3877)
);

NAND2xp5_ASAP7_75t_L g3878 ( 
.A(n_3198),
.B(n_119),
.Y(n_3878)
);

INVx2_ASAP7_75t_L g3879 ( 
.A(n_3196),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_L g3880 ( 
.A(n_3198),
.B(n_119),
.Y(n_3880)
);

NAND2xp5_ASAP7_75t_L g3881 ( 
.A(n_2985),
.B(n_119),
.Y(n_3881)
);

OAI221xp5_ASAP7_75t_L g3882 ( 
.A1(n_2809),
.A2(n_122),
.B1(n_123),
.B2(n_121),
.C(n_120),
.Y(n_3882)
);

AOI21xp5_ASAP7_75t_L g3883 ( 
.A1(n_3266),
.A2(n_122),
.B(n_121),
.Y(n_3883)
);

CKINVDCx5p33_ASAP7_75t_R g3884 ( 
.A(n_2807),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_SL g3885 ( 
.A(n_3254),
.B(n_121),
.Y(n_3885)
);

O2A1O1Ixp5_ASAP7_75t_L g3886 ( 
.A1(n_3125),
.A2(n_125),
.B(n_126),
.C(n_124),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3116),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_L g3888 ( 
.A(n_3003),
.B(n_124),
.Y(n_3888)
);

NOR3xp33_ASAP7_75t_L g3889 ( 
.A(n_3168),
.B(n_126),
.C(n_124),
.Y(n_3889)
);

NAND2xp5_ASAP7_75t_SL g3890 ( 
.A(n_3153),
.B(n_126),
.Y(n_3890)
);

NAND2xp5_ASAP7_75t_L g3891 ( 
.A(n_2904),
.B(n_127),
.Y(n_3891)
);

NAND3xp33_ASAP7_75t_L g3892 ( 
.A(n_3115),
.B(n_129),
.C(n_128),
.Y(n_3892)
);

INVxp67_ASAP7_75t_L g3893 ( 
.A(n_2933),
.Y(n_3893)
);

NAND2xp5_ASAP7_75t_SL g3894 ( 
.A(n_3153),
.B(n_128),
.Y(n_3894)
);

INVx1_ASAP7_75t_L g3895 ( 
.A(n_3117),
.Y(n_3895)
);

NAND2xp5_ASAP7_75t_SL g3896 ( 
.A(n_3020),
.B(n_128),
.Y(n_3896)
);

NOR2xp33_ASAP7_75t_L g3897 ( 
.A(n_3297),
.B(n_129),
.Y(n_3897)
);

AOI22xp33_ASAP7_75t_L g3898 ( 
.A1(n_3161),
.A2(n_130),
.B1(n_131),
.B2(n_129),
.Y(n_3898)
);

INVx3_ASAP7_75t_L g3899 ( 
.A(n_2924),
.Y(n_3899)
);

INVxp67_ASAP7_75t_L g3900 ( 
.A(n_2940),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_3122),
.Y(n_3901)
);

INVx2_ASAP7_75t_L g3902 ( 
.A(n_3206),
.Y(n_3902)
);

INVx2_ASAP7_75t_L g3903 ( 
.A(n_3213),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_SL g3904 ( 
.A(n_3291),
.B(n_130),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3220),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_2913),
.B(n_130),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_L g3907 ( 
.A(n_2960),
.B(n_131),
.Y(n_3907)
);

AOI22xp33_ASAP7_75t_L g3908 ( 
.A1(n_3085),
.A2(n_132),
.B1(n_133),
.B2(n_131),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3101),
.Y(n_3909)
);

NAND2xp5_ASAP7_75t_L g3910 ( 
.A(n_2983),
.B(n_132),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_SL g3911 ( 
.A(n_3291),
.B(n_132),
.Y(n_3911)
);

BUFx6f_ASAP7_75t_L g3912 ( 
.A(n_3291),
.Y(n_3912)
);

A2O1A1Ixp33_ASAP7_75t_L g3913 ( 
.A1(n_3264),
.A2(n_3268),
.B(n_2979),
.C(n_2964),
.Y(n_3913)
);

BUFx3_ASAP7_75t_L g3914 ( 
.A(n_2861),
.Y(n_3914)
);

NOR2xp67_ASAP7_75t_L g3915 ( 
.A(n_3203),
.B(n_133),
.Y(n_3915)
);

INVx2_ASAP7_75t_L g3916 ( 
.A(n_2827),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_SL g3917 ( 
.A(n_3321),
.B(n_134),
.Y(n_3917)
);

AOI221xp5_ASAP7_75t_L g3918 ( 
.A1(n_3039),
.A2(n_136),
.B1(n_137),
.B2(n_135),
.C(n_134),
.Y(n_3918)
);

NOR2xp33_ASAP7_75t_R g3919 ( 
.A(n_3414),
.B(n_3433),
.Y(n_3919)
);

INVx2_ASAP7_75t_L g3920 ( 
.A(n_2828),
.Y(n_3920)
);

AND2x4_ASAP7_75t_L g3921 ( 
.A(n_2924),
.B(n_135),
.Y(n_3921)
);

OR2x2_ASAP7_75t_L g3922 ( 
.A(n_3219),
.B(n_135),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3101),
.Y(n_3923)
);

NOR2xp33_ASAP7_75t_L g3924 ( 
.A(n_3333),
.B(n_136),
.Y(n_3924)
);

INVxp67_ASAP7_75t_L g3925 ( 
.A(n_2927),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_L g3926 ( 
.A(n_3130),
.B(n_136),
.Y(n_3926)
);

OR2x2_ASAP7_75t_L g3927 ( 
.A(n_3440),
.B(n_138),
.Y(n_3927)
);

CKINVDCx5p33_ASAP7_75t_R g3928 ( 
.A(n_3454),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_L g3929 ( 
.A(n_3130),
.B(n_138),
.Y(n_3929)
);

NOR2xp33_ASAP7_75t_L g3930 ( 
.A(n_3338),
.B(n_138),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3224),
.Y(n_3931)
);

NAND2xp5_ASAP7_75t_SL g3932 ( 
.A(n_3321),
.B(n_139),
.Y(n_3932)
);

BUFx8_ASAP7_75t_L g3933 ( 
.A(n_3214),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_2872),
.B(n_139),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3036),
.Y(n_3935)
);

INVx2_ASAP7_75t_SL g3936 ( 
.A(n_3351),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3036),
.Y(n_3937)
);

NAND2xp5_ASAP7_75t_SL g3938 ( 
.A(n_3321),
.B(n_139),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3043),
.Y(n_3939)
);

BUFx3_ASAP7_75t_L g3940 ( 
.A(n_3351),
.Y(n_3940)
);

INVx1_ASAP7_75t_L g3941 ( 
.A(n_3043),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_SL g3942 ( 
.A(n_3328),
.B(n_140),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3241),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3251),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3253),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3188),
.Y(n_3946)
);

INVxp33_ASAP7_75t_L g3947 ( 
.A(n_2824),
.Y(n_3947)
);

BUFx6f_ASAP7_75t_SL g3948 ( 
.A(n_3089),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_SL g3949 ( 
.A(n_3328),
.B(n_140),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_L g3950 ( 
.A(n_2873),
.B(n_140),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_SL g3951 ( 
.A(n_3328),
.B(n_141),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_L g3952 ( 
.A(n_3142),
.B(n_141),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_L g3953 ( 
.A(n_3142),
.B(n_141),
.Y(n_3953)
);

BUFx6f_ASAP7_75t_L g3954 ( 
.A(n_3346),
.Y(n_3954)
);

NAND2xp5_ASAP7_75t_L g3955 ( 
.A(n_3155),
.B(n_3164),
.Y(n_3955)
);

NOR2xp33_ASAP7_75t_L g3956 ( 
.A(n_3363),
.B(n_142),
.Y(n_3956)
);

INVxp33_ASAP7_75t_L g3957 ( 
.A(n_2857),
.Y(n_3957)
);

INVx2_ASAP7_75t_L g3958 ( 
.A(n_2841),
.Y(n_3958)
);

INVx1_ASAP7_75t_L g3959 ( 
.A(n_3223),
.Y(n_3959)
);

INVx2_ASAP7_75t_SL g3960 ( 
.A(n_3360),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_SL g3961 ( 
.A(n_3346),
.B(n_142),
.Y(n_3961)
);

INVx2_ASAP7_75t_SL g3962 ( 
.A(n_3360),
.Y(n_3962)
);

AND2x6_ASAP7_75t_SL g3963 ( 
.A(n_3337),
.B(n_0),
.Y(n_3963)
);

AND2x2_ASAP7_75t_SL g3964 ( 
.A(n_3051),
.B(n_143),
.Y(n_3964)
);

A2O1A1Ixp33_ASAP7_75t_L g3965 ( 
.A1(n_3229),
.A2(n_3),
.B(n_1),
.C(n_2),
.Y(n_3965)
);

NOR2xp33_ASAP7_75t_L g3966 ( 
.A(n_3441),
.B(n_143),
.Y(n_3966)
);

NAND2xp5_ASAP7_75t_SL g3967 ( 
.A(n_3346),
.B(n_143),
.Y(n_3967)
);

OAI22xp5_ASAP7_75t_L g3968 ( 
.A1(n_3307),
.A2(n_145),
.B1(n_146),
.B2(n_144),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_SL g3969 ( 
.A(n_3368),
.B(n_144),
.Y(n_3969)
);

NAND2xp5_ASAP7_75t_SL g3970 ( 
.A(n_3368),
.B(n_144),
.Y(n_3970)
);

INVx1_ASAP7_75t_L g3971 ( 
.A(n_3223),
.Y(n_3971)
);

INVx8_ASAP7_75t_L g3972 ( 
.A(n_3077),
.Y(n_3972)
);

INVxp67_ASAP7_75t_L g3973 ( 
.A(n_3237),
.Y(n_3973)
);

BUFx6f_ASAP7_75t_L g3974 ( 
.A(n_3368),
.Y(n_3974)
);

NOR3xp33_ASAP7_75t_L g3975 ( 
.A(n_3443),
.B(n_146),
.C(n_145),
.Y(n_3975)
);

NOR3xp33_ASAP7_75t_L g3976 ( 
.A(n_3450),
.B(n_148),
.C(n_147),
.Y(n_3976)
);

INVx2_ASAP7_75t_SL g3977 ( 
.A(n_3374),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_SL g3978 ( 
.A(n_3406),
.B(n_147),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_L g3979 ( 
.A(n_3155),
.B(n_147),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_SL g3980 ( 
.A(n_3406),
.B(n_148),
.Y(n_3980)
);

INVx1_ASAP7_75t_L g3981 ( 
.A(n_3107),
.Y(n_3981)
);

AND2x2_ASAP7_75t_L g3982 ( 
.A(n_3199),
.B(n_148),
.Y(n_3982)
);

NOR2xp67_ASAP7_75t_L g3983 ( 
.A(n_3203),
.B(n_149),
.Y(n_3983)
);

NAND2xp5_ASAP7_75t_SL g3984 ( 
.A(n_3406),
.B(n_149),
.Y(n_3984)
);

NAND2xp5_ASAP7_75t_L g3985 ( 
.A(n_3164),
.B(n_149),
.Y(n_3985)
);

OAI22xp5_ASAP7_75t_L g3986 ( 
.A1(n_2987),
.A2(n_151),
.B1(n_152),
.B2(n_150),
.Y(n_3986)
);

OAI22xp5_ASAP7_75t_L g3987 ( 
.A1(n_3287),
.A2(n_151),
.B1(n_152),
.B2(n_150),
.Y(n_3987)
);

INVx2_ASAP7_75t_SL g3988 ( 
.A(n_3374),
.Y(n_3988)
);

INVx1_ASAP7_75t_L g3989 ( 
.A(n_3119),
.Y(n_3989)
);

INVx1_ASAP7_75t_L g3990 ( 
.A(n_3121),
.Y(n_3990)
);

INVx2_ASAP7_75t_SL g3991 ( 
.A(n_3412),
.Y(n_3991)
);

NAND2xp5_ASAP7_75t_SL g3992 ( 
.A(n_3233),
.B(n_152),
.Y(n_3992)
);

INVx1_ASAP7_75t_L g3993 ( 
.A(n_3242),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_L g3994 ( 
.A(n_3174),
.B(n_153),
.Y(n_3994)
);

OR2x2_ASAP7_75t_L g3995 ( 
.A(n_3144),
.B(n_154),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_L g3996 ( 
.A(n_3174),
.B(n_154),
.Y(n_3996)
);

INVxp67_ASAP7_75t_L g3997 ( 
.A(n_3137),
.Y(n_3997)
);

BUFx6f_ASAP7_75t_SL g3998 ( 
.A(n_3123),
.Y(n_3998)
);

OR2x2_ASAP7_75t_L g3999 ( 
.A(n_2795),
.B(n_154),
.Y(n_3999)
);

INVx1_ASAP7_75t_SL g4000 ( 
.A(n_3234),
.Y(n_4000)
);

BUFx2_ASAP7_75t_L g4001 ( 
.A(n_3412),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_3209),
.B(n_155),
.Y(n_4002)
);

INVx2_ASAP7_75t_L g4003 ( 
.A(n_3044),
.Y(n_4003)
);

INVx1_ASAP7_75t_L g4004 ( 
.A(n_3232),
.Y(n_4004)
);

INVxp67_ASAP7_75t_SL g4005 ( 
.A(n_3044),
.Y(n_4005)
);

O2A1O1Ixp33_ASAP7_75t_L g4006 ( 
.A1(n_3108),
.A2(n_157),
.B(n_158),
.C(n_156),
.Y(n_4006)
);

AOI22xp5_ASAP7_75t_L g4007 ( 
.A1(n_3110),
.A2(n_157),
.B1(n_158),
.B2(n_156),
.Y(n_4007)
);

BUFx3_ASAP7_75t_L g4008 ( 
.A(n_3453),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_L g4009 ( 
.A(n_3393),
.B(n_157),
.Y(n_4009)
);

NOR2xp33_ASAP7_75t_L g4010 ( 
.A(n_3221),
.B(n_159),
.Y(n_4010)
);

NOR2xp33_ASAP7_75t_L g4011 ( 
.A(n_2925),
.B(n_159),
.Y(n_4011)
);

INVxp33_ASAP7_75t_L g4012 ( 
.A(n_3453),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_L g4013 ( 
.A(n_3289),
.B(n_3310),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_L g4014 ( 
.A(n_3314),
.B(n_160),
.Y(n_4014)
);

AOI22xp5_ASAP7_75t_SL g4015 ( 
.A1(n_2908),
.A2(n_161),
.B1(n_162),
.B2(n_160),
.Y(n_4015)
);

NAND2xp5_ASAP7_75t_SL g4016 ( 
.A(n_2934),
.B(n_160),
.Y(n_4016)
);

NAND2xp5_ASAP7_75t_L g4017 ( 
.A(n_3318),
.B(n_161),
.Y(n_4017)
);

INVx2_ASAP7_75t_L g4018 ( 
.A(n_3044),
.Y(n_4018)
);

INVx1_ASAP7_75t_L g4019 ( 
.A(n_3232),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_3238),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3238),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_3324),
.B(n_163),
.Y(n_4022)
);

OR2x2_ASAP7_75t_L g4023 ( 
.A(n_3325),
.B(n_163),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_L g4024 ( 
.A(n_3331),
.B(n_163),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3276),
.Y(n_4025)
);

INVxp67_ASAP7_75t_L g4026 ( 
.A(n_3319),
.Y(n_4026)
);

AOI22x1_ASAP7_75t_L g4027 ( 
.A1(n_2796),
.A2(n_165),
.B1(n_166),
.B2(n_164),
.Y(n_4027)
);

NAND2xp5_ASAP7_75t_SL g4028 ( 
.A(n_2934),
.B(n_164),
.Y(n_4028)
);

NAND2xp5_ASAP7_75t_L g4029 ( 
.A(n_3335),
.B(n_3362),
.Y(n_4029)
);

AND2x2_ASAP7_75t_L g4030 ( 
.A(n_3062),
.B(n_164),
.Y(n_4030)
);

OAI22x1_ASAP7_75t_SL g4031 ( 
.A1(n_3139),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_3579),
.Y(n_4032)
);

INVx2_ASAP7_75t_L g4033 ( 
.A(n_3832),
.Y(n_4033)
);

AOI22xp5_ASAP7_75t_L g4034 ( 
.A1(n_3478),
.A2(n_2870),
.B1(n_3106),
.B2(n_3105),
.Y(n_4034)
);

AND2x6_ASAP7_75t_SL g4035 ( 
.A(n_3594),
.B(n_2957),
.Y(n_4035)
);

NOR2xp33_ASAP7_75t_L g4036 ( 
.A(n_3957),
.B(n_2854),
.Y(n_4036)
);

INVx2_ASAP7_75t_L g4037 ( 
.A(n_3836),
.Y(n_4037)
);

INVx1_ASAP7_75t_L g4038 ( 
.A(n_3584),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_SL g4039 ( 
.A(n_3635),
.B(n_3071),
.Y(n_4039)
);

AOI22xp5_ASAP7_75t_L g4040 ( 
.A1(n_3656),
.A2(n_3182),
.B1(n_3201),
.B2(n_3235),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_SL g4041 ( 
.A(n_3635),
.B(n_3071),
.Y(n_4041)
);

O2A1O1Ixp5_ASAP7_75t_L g4042 ( 
.A1(n_3483),
.A2(n_2984),
.B(n_2976),
.C(n_2858),
.Y(n_4042)
);

AOI22xp33_ASAP7_75t_L g4043 ( 
.A1(n_3683),
.A2(n_2959),
.B1(n_2978),
.B2(n_2975),
.Y(n_4043)
);

AND2x4_ASAP7_75t_L g4044 ( 
.A(n_3532),
.B(n_2905),
.Y(n_4044)
);

INVx1_ASAP7_75t_L g4045 ( 
.A(n_3588),
.Y(n_4045)
);

AND2x4_ASAP7_75t_L g4046 ( 
.A(n_3532),
.B(n_2905),
.Y(n_4046)
);

INVx1_ASAP7_75t_SL g4047 ( 
.A(n_3620),
.Y(n_4047)
);

INVx1_ASAP7_75t_L g4048 ( 
.A(n_3591),
.Y(n_4048)
);

INVx1_ASAP7_75t_L g4049 ( 
.A(n_3596),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_3610),
.Y(n_4050)
);

INVxp67_ASAP7_75t_L g4051 ( 
.A(n_3514),
.Y(n_4051)
);

BUFx3_ASAP7_75t_L g4052 ( 
.A(n_3670),
.Y(n_4052)
);

OR2x2_ASAP7_75t_L g4053 ( 
.A(n_3456),
.B(n_3359),
.Y(n_4053)
);

NAND2xp33_ASAP7_75t_SL g4054 ( 
.A(n_3498),
.B(n_2822),
.Y(n_4054)
);

INVx2_ASAP7_75t_L g4055 ( 
.A(n_3838),
.Y(n_4055)
);

INVx2_ASAP7_75t_L g4056 ( 
.A(n_3856),
.Y(n_4056)
);

NOR2xp33_ASAP7_75t_R g4057 ( 
.A(n_3699),
.B(n_3009),
.Y(n_4057)
);

NOR3xp33_ASAP7_75t_SL g4058 ( 
.A(n_3482),
.B(n_3112),
.C(n_3069),
.Y(n_4058)
);

INVx2_ASAP7_75t_SL g4059 ( 
.A(n_3670),
.Y(n_4059)
);

INVx1_ASAP7_75t_SL g4060 ( 
.A(n_4001),
.Y(n_4060)
);

INVx5_ASAP7_75t_L g4061 ( 
.A(n_3670),
.Y(n_4061)
);

INVx2_ASAP7_75t_L g4062 ( 
.A(n_3692),
.Y(n_4062)
);

HB1xp67_ASAP7_75t_L g4063 ( 
.A(n_3530),
.Y(n_4063)
);

AOI22xp5_ASAP7_75t_L g4064 ( 
.A1(n_3807),
.A2(n_3538),
.B1(n_3713),
.B2(n_3460),
.Y(n_4064)
);

BUFx12f_ASAP7_75t_L g4065 ( 
.A(n_3746),
.Y(n_4065)
);

BUFx3_ASAP7_75t_L g4066 ( 
.A(n_3875),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_3558),
.B(n_3369),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_3613),
.Y(n_4068)
);

NAND2xp5_ASAP7_75t_L g4069 ( 
.A(n_3772),
.B(n_3370),
.Y(n_4069)
);

NOR2xp33_ASAP7_75t_L g4070 ( 
.A(n_3863),
.B(n_2951),
.Y(n_4070)
);

INVx2_ASAP7_75t_L g4071 ( 
.A(n_3693),
.Y(n_4071)
);

BUFx2_ASAP7_75t_L g4072 ( 
.A(n_3594),
.Y(n_4072)
);

INVx4_ASAP7_75t_L g4073 ( 
.A(n_3875),
.Y(n_4073)
);

INVx2_ASAP7_75t_SL g4074 ( 
.A(n_3875),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_L g4075 ( 
.A(n_3479),
.B(n_3378),
.Y(n_4075)
);

OAI21xp5_ASAP7_75t_L g4076 ( 
.A1(n_3512),
.A2(n_3095),
.B(n_3081),
.Y(n_4076)
);

BUFx3_ASAP7_75t_L g4077 ( 
.A(n_3940),
.Y(n_4077)
);

AOI22xp33_ASAP7_75t_L g4078 ( 
.A1(n_3696),
.A2(n_2959),
.B1(n_2978),
.B2(n_2975),
.Y(n_4078)
);

NAND2xp5_ASAP7_75t_L g4079 ( 
.A(n_3470),
.B(n_3385),
.Y(n_4079)
);

INVx4_ASAP7_75t_L g4080 ( 
.A(n_3624),
.Y(n_4080)
);

BUFx6f_ASAP7_75t_L g4081 ( 
.A(n_3972),
.Y(n_4081)
);

CKINVDCx6p67_ASAP7_75t_R g4082 ( 
.A(n_3806),
.Y(n_4082)
);

INVx2_ASAP7_75t_SL g4083 ( 
.A(n_4008),
.Y(n_4083)
);

NAND2xp5_ASAP7_75t_L g4084 ( 
.A(n_3747),
.B(n_3390),
.Y(n_4084)
);

INVxp67_ASAP7_75t_SL g4085 ( 
.A(n_3527),
.Y(n_4085)
);

INVx2_ASAP7_75t_L g4086 ( 
.A(n_3704),
.Y(n_4086)
);

BUFx2_ASAP7_75t_L g4087 ( 
.A(n_3594),
.Y(n_4087)
);

NAND2xp5_ASAP7_75t_L g4088 ( 
.A(n_3502),
.B(n_3395),
.Y(n_4088)
);

AOI22xp33_ASAP7_75t_L g4089 ( 
.A1(n_3807),
.A2(n_2975),
.B1(n_2978),
.B2(n_3265),
.Y(n_4089)
);

HB1xp67_ASAP7_75t_L g4090 ( 
.A(n_3549),
.Y(n_4090)
);

AOI22xp5_ASAP7_75t_L g4091 ( 
.A1(n_3807),
.A2(n_3240),
.B1(n_3244),
.B2(n_3011),
.Y(n_4091)
);

INVxp67_ASAP7_75t_L g4092 ( 
.A(n_3637),
.Y(n_4092)
);

INVx1_ASAP7_75t_L g4093 ( 
.A(n_3614),
.Y(n_4093)
);

INVxp67_ASAP7_75t_L g4094 ( 
.A(n_3821),
.Y(n_4094)
);

AO22x1_ASAP7_75t_L g4095 ( 
.A1(n_3933),
.A2(n_2978),
.B1(n_2975),
.B2(n_3190),
.Y(n_4095)
);

NAND2xp5_ASAP7_75t_SL g4096 ( 
.A(n_3788),
.B(n_3071),
.Y(n_4096)
);

INVx2_ASAP7_75t_L g4097 ( 
.A(n_3730),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_L g4098 ( 
.A(n_3500),
.B(n_3402),
.Y(n_4098)
);

NAND2xp5_ASAP7_75t_L g4099 ( 
.A(n_3544),
.B(n_3419),
.Y(n_4099)
);

AOI22xp5_ASAP7_75t_L g4100 ( 
.A1(n_3752),
.A2(n_2844),
.B1(n_2845),
.B2(n_3048),
.Y(n_4100)
);

AND2x4_ASAP7_75t_L g4101 ( 
.A(n_3573),
.B(n_2931),
.Y(n_4101)
);

BUFx2_ASAP7_75t_L g4102 ( 
.A(n_3632),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_3618),
.Y(n_4103)
);

NAND2xp5_ASAP7_75t_L g4104 ( 
.A(n_3872),
.B(n_3431),
.Y(n_4104)
);

NAND3xp33_ASAP7_75t_SL g4105 ( 
.A(n_3457),
.B(n_3701),
.C(n_3569),
.Y(n_4105)
);

AND2x2_ASAP7_75t_L g4106 ( 
.A(n_3774),
.B(n_3252),
.Y(n_4106)
);

INVx1_ASAP7_75t_L g4107 ( 
.A(n_3625),
.Y(n_4107)
);

INVx2_ASAP7_75t_L g4108 ( 
.A(n_3731),
.Y(n_4108)
);

AOI22xp5_ASAP7_75t_L g4109 ( 
.A1(n_3893),
.A2(n_3128),
.B1(n_3053),
.B2(n_3205),
.Y(n_4109)
);

BUFx3_ASAP7_75t_L g4110 ( 
.A(n_3575),
.Y(n_4110)
);

BUFx3_ASAP7_75t_L g4111 ( 
.A(n_3630),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_3725),
.B(n_3432),
.Y(n_4112)
);

AOI22xp33_ASAP7_75t_L g4113 ( 
.A1(n_3889),
.A2(n_3158),
.B1(n_3214),
.B2(n_3276),
.Y(n_4113)
);

AND2x2_ASAP7_75t_L g4114 ( 
.A(n_3774),
.B(n_3256),
.Y(n_4114)
);

INVx3_ASAP7_75t_L g4115 ( 
.A(n_3624),
.Y(n_4115)
);

INVx2_ASAP7_75t_L g4116 ( 
.A(n_3740),
.Y(n_4116)
);

NOR2xp33_ASAP7_75t_L g4117 ( 
.A(n_3900),
.B(n_2898),
.Y(n_4117)
);

NAND2xp5_ASAP7_75t_L g4118 ( 
.A(n_3568),
.B(n_3604),
.Y(n_4118)
);

NOR2xp33_ASAP7_75t_L g4119 ( 
.A(n_3973),
.B(n_2901),
.Y(n_4119)
);

INVx1_ASAP7_75t_L g4120 ( 
.A(n_3627),
.Y(n_4120)
);

AND2x4_ASAP7_75t_L g4121 ( 
.A(n_3573),
.B(n_2931),
.Y(n_4121)
);

INVx5_ASAP7_75t_L g4122 ( 
.A(n_3972),
.Y(n_4122)
);

AOI22xp33_ASAP7_75t_L g4123 ( 
.A1(n_3722),
.A2(n_3158),
.B1(n_3190),
.B2(n_3273),
.Y(n_4123)
);

NAND2xp5_ASAP7_75t_SL g4124 ( 
.A(n_3788),
.B(n_2976),
.Y(n_4124)
);

NAND2xp5_ASAP7_75t_L g4125 ( 
.A(n_3768),
.B(n_3019),
.Y(n_4125)
);

AOI22xp5_ASAP7_75t_L g4126 ( 
.A1(n_3636),
.A2(n_3124),
.B1(n_3262),
.B2(n_3260),
.Y(n_4126)
);

NOR2xp33_ASAP7_75t_L g4127 ( 
.A(n_3997),
.B(n_3134),
.Y(n_4127)
);

OR2x6_ASAP7_75t_L g4128 ( 
.A(n_3494),
.B(n_3455),
.Y(n_4128)
);

NAND2xp5_ASAP7_75t_L g4129 ( 
.A(n_3646),
.B(n_3204),
.Y(n_4129)
);

INVx3_ASAP7_75t_L g4130 ( 
.A(n_3769),
.Y(n_4130)
);

INVx2_ASAP7_75t_SL g4131 ( 
.A(n_3769),
.Y(n_4131)
);

AOI22xp33_ASAP7_75t_L g4132 ( 
.A1(n_3703),
.A2(n_3190),
.B1(n_3273),
.B2(n_3096),
.Y(n_4132)
);

AOI22xp33_ASAP7_75t_L g4133 ( 
.A1(n_3706),
.A2(n_3190),
.B1(n_3096),
.B2(n_3077),
.Y(n_4133)
);

AO22x1_ASAP7_75t_L g4134 ( 
.A1(n_3933),
.A2(n_3353),
.B1(n_3366),
.B2(n_3296),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_L g4135 ( 
.A(n_3468),
.B(n_3056),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_L g4136 ( 
.A(n_3550),
.B(n_3035),
.Y(n_4136)
);

NOR2xp33_ASAP7_75t_L g4137 ( 
.A(n_3651),
.B(n_3455),
.Y(n_4137)
);

NOR2xp33_ASAP7_75t_L g4138 ( 
.A(n_3612),
.B(n_2843),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_3489),
.B(n_3082),
.Y(n_4139)
);

AND2x6_ASAP7_75t_L g4140 ( 
.A(n_3595),
.B(n_3657),
.Y(n_4140)
);

NAND2xp5_ASAP7_75t_L g4141 ( 
.A(n_3537),
.B(n_3189),
.Y(n_4141)
);

INVx2_ASAP7_75t_L g4142 ( 
.A(n_3750),
.Y(n_4142)
);

INVx2_ASAP7_75t_L g4143 ( 
.A(n_3754),
.Y(n_4143)
);

NAND2xp5_ASAP7_75t_L g4144 ( 
.A(n_3708),
.B(n_3129),
.Y(n_4144)
);

HB1xp67_ASAP7_75t_L g4145 ( 
.A(n_3557),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_3652),
.Y(n_4146)
);

A2O1A1Ixp33_ASAP7_75t_L g4147 ( 
.A1(n_3755),
.A2(n_3803),
.B(n_3679),
.C(n_3691),
.Y(n_4147)
);

NAND2xp5_ASAP7_75t_L g4148 ( 
.A(n_3955),
.B(n_3269),
.Y(n_4148)
);

INVx2_ASAP7_75t_SL g4149 ( 
.A(n_3802),
.Y(n_4149)
);

INVx3_ASAP7_75t_L g4150 ( 
.A(n_3802),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_SL g4151 ( 
.A(n_3788),
.B(n_2984),
.Y(n_4151)
);

BUFx2_ASAP7_75t_L g4152 ( 
.A(n_3632),
.Y(n_4152)
);

NAND2xp5_ASAP7_75t_L g4153 ( 
.A(n_3570),
.B(n_3175),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_L g4154 ( 
.A(n_3570),
.B(n_3361),
.Y(n_4154)
);

AND2x4_ASAP7_75t_L g4155 ( 
.A(n_3595),
.B(n_2982),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_3653),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_3655),
.Y(n_4157)
);

AND2x2_ASAP7_75t_L g4158 ( 
.A(n_3616),
.B(n_3394),
.Y(n_4158)
);

NAND2xp5_ASAP7_75t_L g4159 ( 
.A(n_4030),
.B(n_3421),
.Y(n_4159)
);

INVx1_ASAP7_75t_L g4160 ( 
.A(n_3664),
.Y(n_4160)
);

HB1xp67_ASAP7_75t_L g4161 ( 
.A(n_3561),
.Y(n_4161)
);

INVx1_ASAP7_75t_SL g4162 ( 
.A(n_3734),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_3665),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_L g4164 ( 
.A(n_4013),
.B(n_2886),
.Y(n_4164)
);

AOI21xp5_ASAP7_75t_L g4165 ( 
.A1(n_3672),
.A2(n_2999),
.B(n_2977),
.Y(n_4165)
);

BUFx6f_ASAP7_75t_L g4166 ( 
.A(n_3972),
.Y(n_4166)
);

INVx2_ASAP7_75t_L g4167 ( 
.A(n_3765),
.Y(n_4167)
);

INVx2_ASAP7_75t_L g4168 ( 
.A(n_3777),
.Y(n_4168)
);

AOI21xp5_ASAP7_75t_L g4169 ( 
.A1(n_3770),
.A2(n_2999),
.B(n_2977),
.Y(n_4169)
);

BUFx8_ASAP7_75t_L g4170 ( 
.A(n_3806),
.Y(n_4170)
);

NAND2xp5_ASAP7_75t_L g4171 ( 
.A(n_4029),
.B(n_2920),
.Y(n_4171)
);

NOR3xp33_ASAP7_75t_L g4172 ( 
.A(n_3487),
.B(n_3193),
.C(n_3146),
.Y(n_4172)
);

CKINVDCx5p33_ASAP7_75t_R g4173 ( 
.A(n_3919),
.Y(n_4173)
);

BUFx3_ASAP7_75t_L g4174 ( 
.A(n_3914),
.Y(n_4174)
);

INVx5_ASAP7_75t_L g4175 ( 
.A(n_3644),
.Y(n_4175)
);

CKINVDCx5p33_ASAP7_75t_R g4176 ( 
.A(n_3825),
.Y(n_4176)
);

NOR2xp33_ASAP7_75t_L g4177 ( 
.A(n_3925),
.B(n_3074),
.Y(n_4177)
);

NAND3xp33_ASAP7_75t_SL g4178 ( 
.A(n_3701),
.B(n_2802),
.C(n_3215),
.Y(n_4178)
);

INVx2_ASAP7_75t_L g4179 ( 
.A(n_3785),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_L g4180 ( 
.A(n_3817),
.B(n_2945),
.Y(n_4180)
);

INVx2_ASAP7_75t_L g4181 ( 
.A(n_3462),
.Y(n_4181)
);

AOI21x1_ASAP7_75t_L g4182 ( 
.A1(n_3589),
.A2(n_2804),
.B(n_2799),
.Y(n_4182)
);

NAND2xp5_ASAP7_75t_L g4183 ( 
.A(n_3793),
.B(n_3808),
.Y(n_4183)
);

BUFx6f_ASAP7_75t_L g4184 ( 
.A(n_3505),
.Y(n_4184)
);

INVx1_ASAP7_75t_L g4185 ( 
.A(n_3680),
.Y(n_4185)
);

NAND2xp5_ASAP7_75t_L g4186 ( 
.A(n_3823),
.B(n_2965),
.Y(n_4186)
);

OAI21xp5_ASAP7_75t_L g4187 ( 
.A1(n_3513),
.A2(n_3227),
.B(n_3226),
.Y(n_4187)
);

AOI22x1_ASAP7_75t_L g4188 ( 
.A1(n_3458),
.A2(n_3097),
.B1(n_2996),
.B2(n_2997),
.Y(n_4188)
);

NAND2x1p5_ASAP7_75t_L g4189 ( 
.A(n_3508),
.B(n_2866),
.Y(n_4189)
);

CKINVDCx5p33_ASAP7_75t_R g4190 ( 
.A(n_3884),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_SL g4191 ( 
.A(n_3788),
.B(n_2796),
.Y(n_4191)
);

BUFx3_ASAP7_75t_L g4192 ( 
.A(n_3628),
.Y(n_4192)
);

NAND2xp5_ASAP7_75t_L g4193 ( 
.A(n_3827),
.B(n_3496),
.Y(n_4193)
);

INVx2_ASAP7_75t_L g4194 ( 
.A(n_3463),
.Y(n_4194)
);

INVx2_ASAP7_75t_L g4195 ( 
.A(n_3471),
.Y(n_4195)
);

BUFx6f_ASAP7_75t_L g4196 ( 
.A(n_3505),
.Y(n_4196)
);

BUFx2_ASAP7_75t_L g4197 ( 
.A(n_3628),
.Y(n_4197)
);

NAND2xp5_ASAP7_75t_L g4198 ( 
.A(n_3673),
.B(n_3674),
.Y(n_4198)
);

INVx1_ASAP7_75t_SL g4199 ( 
.A(n_3548),
.Y(n_4199)
);

AOI22xp33_ASAP7_75t_L g4200 ( 
.A1(n_3619),
.A2(n_3077),
.B1(n_3096),
.B2(n_3126),
.Y(n_4200)
);

AOI22xp5_ASAP7_75t_L g4201 ( 
.A1(n_3711),
.A2(n_3810),
.B1(n_3831),
.B2(n_3638),
.Y(n_4201)
);

INVxp67_ASAP7_75t_L g4202 ( 
.A(n_3860),
.Y(n_4202)
);

AOI22xp5_ASAP7_75t_L g4203 ( 
.A1(n_3964),
.A2(n_3975),
.B1(n_3976),
.B2(n_3644),
.Y(n_4203)
);

HB1xp67_ASAP7_75t_L g4204 ( 
.A(n_3712),
.Y(n_4204)
);

AOI22xp33_ASAP7_75t_L g4205 ( 
.A1(n_3458),
.A2(n_3096),
.B1(n_3126),
.B2(n_3258),
.Y(n_4205)
);

INVx2_ASAP7_75t_L g4206 ( 
.A(n_3480),
.Y(n_4206)
);

NAND2xp5_ASAP7_75t_L g4207 ( 
.A(n_3868),
.B(n_2966),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_L g4208 ( 
.A(n_3801),
.B(n_3029),
.Y(n_4208)
);

NOR2x2_ASAP7_75t_L g4209 ( 
.A(n_3742),
.B(n_3337),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_L g4210 ( 
.A(n_3822),
.B(n_3120),
.Y(n_4210)
);

INVx2_ASAP7_75t_SL g4211 ( 
.A(n_3845),
.Y(n_4211)
);

INVx1_ASAP7_75t_L g4212 ( 
.A(n_3779),
.Y(n_4212)
);

INVx4_ASAP7_75t_L g4213 ( 
.A(n_3948),
.Y(n_4213)
);

NOR2x1p5_ASAP7_75t_L g4214 ( 
.A(n_3648),
.B(n_2866),
.Y(n_4214)
);

INVx3_ASAP7_75t_L g4215 ( 
.A(n_3852),
.Y(n_4215)
);

BUFx2_ASAP7_75t_L g4216 ( 
.A(n_3598),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_3782),
.Y(n_4217)
);

NAND2xp5_ASAP7_75t_SL g4218 ( 
.A(n_3788),
.B(n_2858),
.Y(n_4218)
);

BUFx3_ASAP7_75t_L g4219 ( 
.A(n_3865),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_SL g4220 ( 
.A(n_3915),
.B(n_2874),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_3467),
.Y(n_4221)
);

AND2x4_ASAP7_75t_L g4222 ( 
.A(n_3899),
.B(n_2982),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_SL g4223 ( 
.A(n_3915),
.B(n_2874),
.Y(n_4223)
);

AOI22xp5_ASAP7_75t_L g4224 ( 
.A1(n_3644),
.A2(n_3211),
.B1(n_3145),
.B2(n_3255),
.Y(n_4224)
);

NOR2x2_ASAP7_75t_L g4225 ( 
.A(n_3603),
.B(n_3422),
.Y(n_4225)
);

AND2x2_ASAP7_75t_L g4226 ( 
.A(n_3982),
.B(n_3170),
.Y(n_4226)
);

INVx1_ASAP7_75t_L g4227 ( 
.A(n_3476),
.Y(n_4227)
);

AOI22xp33_ASAP7_75t_L g4228 ( 
.A1(n_3644),
.A2(n_3258),
.B1(n_3261),
.B2(n_3259),
.Y(n_4228)
);

INVx4_ASAP7_75t_L g4229 ( 
.A(n_3948),
.Y(n_4229)
);

AOI22xp33_ASAP7_75t_L g4230 ( 
.A1(n_3767),
.A2(n_3259),
.B1(n_3261),
.B2(n_3296),
.Y(n_4230)
);

BUFx3_ASAP7_75t_L g4231 ( 
.A(n_3936),
.Y(n_4231)
);

NOR3xp33_ASAP7_75t_SL g4232 ( 
.A(n_3928),
.B(n_3132),
.C(n_3131),
.Y(n_4232)
);

CKINVDCx5p33_ASAP7_75t_R g4233 ( 
.A(n_3998),
.Y(n_4233)
);

CKINVDCx5p33_ASAP7_75t_R g4234 ( 
.A(n_3998),
.Y(n_4234)
);

OR2x6_ASAP7_75t_L g4235 ( 
.A(n_3517),
.B(n_2914),
.Y(n_4235)
);

NAND2xp5_ASAP7_75t_SL g4236 ( 
.A(n_3983),
.B(n_3288),
.Y(n_4236)
);

NAND2xp5_ASAP7_75t_L g4237 ( 
.A(n_3826),
.B(n_3236),
.Y(n_4237)
);

AND2x2_ASAP7_75t_L g4238 ( 
.A(n_3760),
.B(n_3184),
.Y(n_4238)
);

NOR2xp33_ASAP7_75t_L g4239 ( 
.A(n_3698),
.B(n_3947),
.Y(n_4239)
);

NAND2xp5_ASAP7_75t_SL g4240 ( 
.A(n_3983),
.B(n_3288),
.Y(n_4240)
);

AOI22xp5_ASAP7_75t_L g4241 ( 
.A1(n_3686),
.A2(n_3247),
.B1(n_2848),
.B2(n_3102),
.Y(n_4241)
);

INVx2_ASAP7_75t_SL g4242 ( 
.A(n_3960),
.Y(n_4242)
);

NAND2xp5_ASAP7_75t_SL g4243 ( 
.A(n_3555),
.B(n_3299),
.Y(n_4243)
);

AO22x1_ASAP7_75t_L g4244 ( 
.A1(n_4000),
.A2(n_3296),
.B1(n_3366),
.B2(n_3353),
.Y(n_4244)
);

INVx5_ASAP7_75t_L g4245 ( 
.A(n_3505),
.Y(n_4245)
);

BUFx3_ASAP7_75t_L g4246 ( 
.A(n_3962),
.Y(n_4246)
);

INVx3_ASAP7_75t_L g4247 ( 
.A(n_3977),
.Y(n_4247)
);

AOI22xp5_ASAP7_75t_L g4248 ( 
.A1(n_3751),
.A2(n_3102),
.B1(n_3353),
.B2(n_3296),
.Y(n_4248)
);

INVx1_ASAP7_75t_L g4249 ( 
.A(n_3477),
.Y(n_4249)
);

BUFx3_ASAP7_75t_L g4250 ( 
.A(n_3988),
.Y(n_4250)
);

INVx2_ASAP7_75t_L g4251 ( 
.A(n_3481),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_SL g4252 ( 
.A(n_3555),
.B(n_3299),
.Y(n_4252)
);

BUFx4f_ASAP7_75t_L g4253 ( 
.A(n_3552),
.Y(n_4253)
);

INVx2_ASAP7_75t_L g4254 ( 
.A(n_3509),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_3488),
.Y(n_4255)
);

NAND2x1p5_ASAP7_75t_L g4256 ( 
.A(n_3566),
.B(n_2896),
.Y(n_4256)
);

AOI22xp33_ASAP7_75t_L g4257 ( 
.A1(n_3592),
.A2(n_3353),
.B1(n_3411),
.B2(n_3366),
.Y(n_4257)
);

BUFx12f_ASAP7_75t_L g4258 ( 
.A(n_3963),
.Y(n_4258)
);

INVx5_ASAP7_75t_L g4259 ( 
.A(n_3523),
.Y(n_4259)
);

AOI21xp5_ASAP7_75t_L g4260 ( 
.A1(n_3830),
.A2(n_2999),
.B(n_2977),
.Y(n_4260)
);

BUFx6f_ASAP7_75t_L g4261 ( 
.A(n_3523),
.Y(n_4261)
);

BUFx12f_ASAP7_75t_L g4262 ( 
.A(n_3762),
.Y(n_4262)
);

OAI22xp5_ASAP7_75t_L g4263 ( 
.A1(n_3647),
.A2(n_3246),
.B1(n_3046),
.B2(n_3054),
.Y(n_4263)
);

AND3x1_ASAP7_75t_L g4264 ( 
.A(n_3615),
.B(n_3422),
.C(n_3047),
.Y(n_4264)
);

NAND2xp5_ASAP7_75t_SL g4265 ( 
.A(n_3622),
.B(n_3640),
.Y(n_4265)
);

BUFx6f_ASAP7_75t_L g4266 ( 
.A(n_3523),
.Y(n_4266)
);

AND2x4_ASAP7_75t_L g4267 ( 
.A(n_3899),
.B(n_3046),
.Y(n_4267)
);

INVx2_ASAP7_75t_L g4268 ( 
.A(n_3511),
.Y(n_4268)
);

INVx2_ASAP7_75t_L g4269 ( 
.A(n_3546),
.Y(n_4269)
);

INVx1_ASAP7_75t_L g4270 ( 
.A(n_3491),
.Y(n_4270)
);

INVx3_ASAP7_75t_L g4271 ( 
.A(n_3991),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_SL g4272 ( 
.A(n_3622),
.B(n_3371),
.Y(n_4272)
);

NOR2xp33_ASAP7_75t_L g4273 ( 
.A(n_3593),
.B(n_3058),
.Y(n_4273)
);

AO21x1_ASAP7_75t_L g4274 ( 
.A1(n_3869),
.A2(n_3208),
.B(n_3357),
.Y(n_4274)
);

NAND2xp5_ASAP7_75t_L g4275 ( 
.A(n_3658),
.B(n_3249),
.Y(n_4275)
);

NAND2xp5_ASAP7_75t_SL g4276 ( 
.A(n_3640),
.B(n_3371),
.Y(n_4276)
);

BUFx3_ASAP7_75t_L g4277 ( 
.A(n_3736),
.Y(n_4277)
);

INVx1_ASAP7_75t_L g4278 ( 
.A(n_3493),
.Y(n_4278)
);

CKINVDCx5p33_ASAP7_75t_R g4279 ( 
.A(n_3847),
.Y(n_4279)
);

INVx1_ASAP7_75t_L g4280 ( 
.A(n_3516),
.Y(n_4280)
);

OR2x6_ASAP7_75t_L g4281 ( 
.A(n_3654),
.B(n_2896),
.Y(n_4281)
);

AOI22xp5_ASAP7_75t_L g4282 ( 
.A1(n_3834),
.A2(n_3102),
.B1(n_3411),
.B2(n_3366),
.Y(n_4282)
);

BUFx6f_ASAP7_75t_L g4283 ( 
.A(n_3571),
.Y(n_4283)
);

NAND2xp5_ASAP7_75t_L g4284 ( 
.A(n_3660),
.B(n_3687),
.Y(n_4284)
);

INVx2_ASAP7_75t_L g4285 ( 
.A(n_3565),
.Y(n_4285)
);

CKINVDCx5p33_ASAP7_75t_R g4286 ( 
.A(n_4031),
.Y(n_4286)
);

INVx3_ASAP7_75t_L g4287 ( 
.A(n_3682),
.Y(n_4287)
);

INVx2_ASAP7_75t_L g4288 ( 
.A(n_3576),
.Y(n_4288)
);

HB1xp67_ASAP7_75t_L g4289 ( 
.A(n_3582),
.Y(n_4289)
);

NAND2xp5_ASAP7_75t_SL g4290 ( 
.A(n_3685),
.B(n_3303),
.Y(n_4290)
);

BUFx6f_ASAP7_75t_L g4291 ( 
.A(n_3571),
.Y(n_4291)
);

NAND2xp5_ASAP7_75t_SL g4292 ( 
.A(n_3685),
.B(n_3303),
.Y(n_4292)
);

CKINVDCx5p33_ASAP7_75t_R g4293 ( 
.A(n_3702),
.Y(n_4293)
);

INVx4_ASAP7_75t_L g4294 ( 
.A(n_3657),
.Y(n_4294)
);

CKINVDCx5p33_ASAP7_75t_R g4295 ( 
.A(n_3707),
.Y(n_4295)
);

AND2x4_ASAP7_75t_L g4296 ( 
.A(n_3684),
.B(n_3047),
.Y(n_4296)
);

AND2x4_ASAP7_75t_L g4297 ( 
.A(n_3684),
.B(n_3054),
.Y(n_4297)
);

AOI22xp33_ASAP7_75t_L g4298 ( 
.A1(n_3671),
.A2(n_3411),
.B1(n_3102),
.B2(n_3250),
.Y(n_4298)
);

BUFx3_ASAP7_75t_L g4299 ( 
.A(n_3650),
.Y(n_4299)
);

NOR2xp33_ASAP7_75t_L g4300 ( 
.A(n_3626),
.B(n_2914),
.Y(n_4300)
);

NAND2xp5_ASAP7_75t_L g4301 ( 
.A(n_3710),
.B(n_3127),
.Y(n_4301)
);

CKINVDCx5p33_ASAP7_75t_R g4302 ( 
.A(n_4015),
.Y(n_4302)
);

BUFx6f_ASAP7_75t_L g4303 ( 
.A(n_3571),
.Y(n_4303)
);

NOR2xp33_ASAP7_75t_L g4304 ( 
.A(n_3621),
.B(n_3172),
.Y(n_4304)
);

INVx3_ASAP7_75t_L g4305 ( 
.A(n_3921),
.Y(n_4305)
);

BUFx6f_ASAP7_75t_L g4306 ( 
.A(n_3794),
.Y(n_4306)
);

OR2x2_ASAP7_75t_SL g4307 ( 
.A(n_3995),
.B(n_165),
.Y(n_4307)
);

INVx2_ASAP7_75t_L g4308 ( 
.A(n_3577),
.Y(n_4308)
);

HB1xp67_ASAP7_75t_L g4309 ( 
.A(n_3667),
.Y(n_4309)
);

OR2x6_ASAP7_75t_L g4310 ( 
.A(n_3667),
.B(n_3208),
.Y(n_4310)
);

INVx1_ASAP7_75t_L g4311 ( 
.A(n_3522),
.Y(n_4311)
);

NAND2xp5_ASAP7_75t_L g4312 ( 
.A(n_3718),
.B(n_3140),
.Y(n_4312)
);

AND2x4_ASAP7_75t_SL g4313 ( 
.A(n_3921),
.B(n_3172),
.Y(n_4313)
);

AOI22xp5_ASAP7_75t_L g4314 ( 
.A1(n_3842),
.A2(n_3411),
.B1(n_3225),
.B2(n_3207),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_3524),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_3525),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_3526),
.Y(n_4317)
);

AOI22xp33_ASAP7_75t_SL g4318 ( 
.A1(n_3520),
.A2(n_3715),
.B1(n_3681),
.B2(n_3689),
.Y(n_4318)
);

OR2x6_ASAP7_75t_L g4319 ( 
.A(n_3681),
.B(n_3715),
.Y(n_4319)
);

INVx1_ASAP7_75t_L g4320 ( 
.A(n_3528),
.Y(n_4320)
);

NAND2xp5_ASAP7_75t_L g4321 ( 
.A(n_3720),
.B(n_3057),
.Y(n_4321)
);

INVx5_ASAP7_75t_L g4322 ( 
.A(n_3794),
.Y(n_4322)
);

AND2x4_ASAP7_75t_L g4323 ( 
.A(n_3748),
.B(n_3057),
.Y(n_4323)
);

AO22x1_ASAP7_75t_L g4324 ( 
.A1(n_4012),
.A2(n_3248),
.B1(n_3250),
.B2(n_3083),
.Y(n_4324)
);

AOI22xp5_ASAP7_75t_L g4325 ( 
.A1(n_3853),
.A2(n_3207),
.B1(n_3200),
.B2(n_3250),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_3529),
.Y(n_4326)
);

BUFx3_ASAP7_75t_L g4327 ( 
.A(n_3564),
.Y(n_4327)
);

NAND2xp5_ASAP7_75t_SL g4328 ( 
.A(n_3792),
.B(n_3312),
.Y(n_4328)
);

NOR2xp67_ASAP7_75t_L g4329 ( 
.A(n_4026),
.B(n_3312),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_3533),
.Y(n_4330)
);

AOI22xp33_ASAP7_75t_L g4331 ( 
.A1(n_3882),
.A2(n_3250),
.B1(n_3200),
.B2(n_3080),
.Y(n_4331)
);

AOI22xp5_ASAP7_75t_L g4332 ( 
.A1(n_3897),
.A2(n_3080),
.B1(n_3113),
.B2(n_3083),
.Y(n_4332)
);

AND2x4_ASAP7_75t_L g4333 ( 
.A(n_3748),
.B(n_3113),
.Y(n_4333)
);

AND2x2_ASAP7_75t_L g4334 ( 
.A(n_3564),
.B(n_3166),
.Y(n_4334)
);

INVx2_ASAP7_75t_L g4335 ( 
.A(n_3586),
.Y(n_4335)
);

NAND2xp5_ASAP7_75t_L g4336 ( 
.A(n_3721),
.B(n_3147),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_3539),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_3541),
.Y(n_4338)
);

AND2x2_ASAP7_75t_L g4339 ( 
.A(n_3922),
.B(n_3166),
.Y(n_4339)
);

INVx2_ASAP7_75t_L g4340 ( 
.A(n_3602),
.Y(n_4340)
);

AND2x4_ASAP7_75t_L g4341 ( 
.A(n_3800),
.B(n_3147),
.Y(n_4341)
);

NOR3xp33_ASAP7_75t_SL g4342 ( 
.A(n_3714),
.B(n_167),
.C(n_166),
.Y(n_4342)
);

NAND2xp5_ASAP7_75t_L g4343 ( 
.A(n_3724),
.B(n_3154),
.Y(n_4343)
);

INVx2_ASAP7_75t_L g4344 ( 
.A(n_3606),
.Y(n_4344)
);

NOR3xp33_ASAP7_75t_SL g4345 ( 
.A(n_3812),
.B(n_167),
.C(n_166),
.Y(n_4345)
);

INVx2_ASAP7_75t_SL g4346 ( 
.A(n_3536),
.Y(n_4346)
);

INVx2_ASAP7_75t_L g4347 ( 
.A(n_3633),
.Y(n_4347)
);

NAND2xp5_ASAP7_75t_L g4348 ( 
.A(n_3726),
.B(n_3154),
.Y(n_4348)
);

INVx1_ASAP7_75t_L g4349 ( 
.A(n_3543),
.Y(n_4349)
);

BUFx6f_ASAP7_75t_L g4350 ( 
.A(n_3794),
.Y(n_4350)
);

NOR2xp33_ASAP7_75t_L g4351 ( 
.A(n_3841),
.B(n_3230),
.Y(n_4351)
);

INVx1_ASAP7_75t_L g4352 ( 
.A(n_3554),
.Y(n_4352)
);

AND2x6_ASAP7_75t_SL g4353 ( 
.A(n_3798),
.B(n_1),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_3560),
.Y(n_4354)
);

INVx2_ASAP7_75t_SL g4355 ( 
.A(n_3567),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_3859),
.Y(n_4356)
);

NAND2xp5_ASAP7_75t_L g4357 ( 
.A(n_3733),
.B(n_3163),
.Y(n_4357)
);

INVx2_ASAP7_75t_L g4358 ( 
.A(n_3641),
.Y(n_4358)
);

NAND2xp5_ASAP7_75t_L g4359 ( 
.A(n_3739),
.B(n_3163),
.Y(n_4359)
);

AND2x4_ASAP7_75t_L g4360 ( 
.A(n_3800),
.B(n_3169),
.Y(n_4360)
);

AOI21xp5_ASAP7_75t_L g4361 ( 
.A1(n_3466),
.A2(n_3028),
.B(n_3301),
.Y(n_4361)
);

NOR2xp33_ASAP7_75t_L g4362 ( 
.A(n_3642),
.B(n_3230),
.Y(n_4362)
);

AOI21xp5_ASAP7_75t_L g4363 ( 
.A1(n_3753),
.A2(n_3028),
.B(n_3352),
.Y(n_4363)
);

INVx4_ASAP7_75t_L g4364 ( 
.A(n_3824),
.Y(n_4364)
);

AOI22xp5_ASAP7_75t_L g4365 ( 
.A1(n_3924),
.A2(n_3169),
.B1(n_3162),
.B2(n_3245),
.Y(n_4365)
);

NAND2xp5_ASAP7_75t_SL g4366 ( 
.A(n_3792),
.B(n_3330),
.Y(n_4366)
);

INVx1_ASAP7_75t_L g4367 ( 
.A(n_3867),
.Y(n_4367)
);

BUFx8_ASAP7_75t_L g4368 ( 
.A(n_3763),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_3870),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_3871),
.Y(n_4370)
);

NAND2xp5_ASAP7_75t_L g4371 ( 
.A(n_3744),
.B(n_3245),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_3876),
.Y(n_4372)
);

NOR2xp33_ASAP7_75t_L g4373 ( 
.A(n_3709),
.B(n_3330),
.Y(n_4373)
);

CKINVDCx5p33_ASAP7_75t_R g4374 ( 
.A(n_3572),
.Y(n_4374)
);

BUFx6f_ASAP7_75t_L g4375 ( 
.A(n_3824),
.Y(n_4375)
);

AND2x2_ASAP7_75t_L g4376 ( 
.A(n_3756),
.B(n_167),
.Y(n_4376)
);

AND2x2_ASAP7_75t_L g4377 ( 
.A(n_3757),
.B(n_168),
.Y(n_4377)
);

INVx2_ASAP7_75t_L g4378 ( 
.A(n_3649),
.Y(n_4378)
);

NAND2xp5_ASAP7_75t_SL g4379 ( 
.A(n_3464),
.B(n_3347),
.Y(n_4379)
);

INVx2_ASAP7_75t_L g4380 ( 
.A(n_3857),
.Y(n_4380)
);

INVx1_ASAP7_75t_L g4381 ( 
.A(n_3887),
.Y(n_4381)
);

AND2x2_ASAP7_75t_L g4382 ( 
.A(n_3759),
.B(n_168),
.Y(n_4382)
);

NOR2xp33_ASAP7_75t_L g4383 ( 
.A(n_3797),
.B(n_3347),
.Y(n_4383)
);

BUFx2_ASAP7_75t_L g4384 ( 
.A(n_3861),
.Y(n_4384)
);

AND2x6_ASAP7_75t_L g4385 ( 
.A(n_3824),
.B(n_3028),
.Y(n_4385)
);

NAND2xp5_ASAP7_75t_SL g4386 ( 
.A(n_3464),
.B(n_3091),
.Y(n_4386)
);

INVx1_ASAP7_75t_SL g4387 ( 
.A(n_3600),
.Y(n_4387)
);

BUFx2_ASAP7_75t_L g4388 ( 
.A(n_3864),
.Y(n_4388)
);

BUFx4f_ASAP7_75t_SL g4389 ( 
.A(n_3623),
.Y(n_4389)
);

CKINVDCx5p33_ASAP7_75t_R g4390 ( 
.A(n_3930),
.Y(n_4390)
);

NAND2xp5_ASAP7_75t_L g4391 ( 
.A(n_3461),
.B(n_3275),
.Y(n_4391)
);

OAI22xp5_ASAP7_75t_L g4392 ( 
.A1(n_3631),
.A2(n_3283),
.B1(n_3285),
.B2(n_2816),
.Y(n_4392)
);

NAND2xp5_ASAP7_75t_L g4393 ( 
.A(n_3469),
.B(n_3271),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_3895),
.Y(n_4394)
);

BUFx3_ASAP7_75t_L g4395 ( 
.A(n_3761),
.Y(n_4395)
);

INVx3_ASAP7_75t_L g4396 ( 
.A(n_3873),
.Y(n_4396)
);

CKINVDCx5p33_ASAP7_75t_R g4397 ( 
.A(n_3956),
.Y(n_4397)
);

INVx1_ASAP7_75t_SL g4398 ( 
.A(n_3835),
.Y(n_4398)
);

INVx2_ASAP7_75t_SL g4399 ( 
.A(n_3877),
.Y(n_4399)
);

NAND2xp5_ASAP7_75t_L g4400 ( 
.A(n_3472),
.B(n_3271),
.Y(n_4400)
);

INVx1_ASAP7_75t_L g4401 ( 
.A(n_3901),
.Y(n_4401)
);

INVx4_ASAP7_75t_L g4402 ( 
.A(n_3840),
.Y(n_4402)
);

NAND2xp5_ASAP7_75t_SL g4403 ( 
.A(n_3545),
.B(n_3091),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_3931),
.Y(n_4404)
);

INVx2_ASAP7_75t_L g4405 ( 
.A(n_3879),
.Y(n_4405)
);

INVx1_ASAP7_75t_L g4406 ( 
.A(n_3943),
.Y(n_4406)
);

AOI22xp5_ASAP7_75t_L g4407 ( 
.A1(n_3966),
.A2(n_3248),
.B1(n_3300),
.B2(n_3292),
.Y(n_4407)
);

AOI22xp33_ASAP7_75t_L g4408 ( 
.A1(n_3992),
.A2(n_3248),
.B1(n_3375),
.B2(n_3317),
.Y(n_4408)
);

INVx1_ASAP7_75t_L g4409 ( 
.A(n_3944),
.Y(n_4409)
);

AND2x2_ASAP7_75t_SL g4410 ( 
.A(n_3631),
.B(n_3439),
.Y(n_4410)
);

AOI21xp5_ASAP7_75t_L g4411 ( 
.A1(n_3597),
.A2(n_3405),
.B(n_3379),
.Y(n_4411)
);

NAND2xp5_ASAP7_75t_L g4412 ( 
.A(n_3473),
.B(n_169),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_3945),
.Y(n_4413)
);

BUFx3_ASAP7_75t_L g4414 ( 
.A(n_3778),
.Y(n_4414)
);

OR2x6_ASAP7_75t_L g4415 ( 
.A(n_3545),
.B(n_3417),
.Y(n_4415)
);

NOR2xp33_ASAP7_75t_L g4416 ( 
.A(n_3639),
.B(n_169),
.Y(n_4416)
);

AOI21xp5_ASAP7_75t_L g4417 ( 
.A1(n_3675),
.A2(n_3429),
.B(n_3425),
.Y(n_4417)
);

AND2x2_ASAP7_75t_L g4418 ( 
.A(n_3905),
.B(n_169),
.Y(n_4418)
);

INVx1_ASAP7_75t_L g4419 ( 
.A(n_3946),
.Y(n_4419)
);

NAND2xp5_ASAP7_75t_L g4420 ( 
.A(n_3474),
.B(n_170),
.Y(n_4420)
);

AND2x4_ASAP7_75t_L g4421 ( 
.A(n_3787),
.B(n_3248),
.Y(n_4421)
);

BUFx2_ASAP7_75t_L g4422 ( 
.A(n_3902),
.Y(n_4422)
);

OR2x6_ASAP7_75t_L g4423 ( 
.A(n_3506),
.B(n_3442),
.Y(n_4423)
);

NOR2xp33_ASAP7_75t_L g4424 ( 
.A(n_3829),
.B(n_170),
.Y(n_4424)
);

NAND2xp5_ASAP7_75t_L g4425 ( 
.A(n_3475),
.B(n_170),
.Y(n_4425)
);

AND2x6_ASAP7_75t_SL g4426 ( 
.A(n_4010),
.B(n_2),
.Y(n_4426)
);

O2A1O1Ixp33_ASAP7_75t_L g4427 ( 
.A1(n_3913),
.A2(n_3896),
.B(n_3611),
.C(n_3607),
.Y(n_4427)
);

INVx1_ASAP7_75t_L g4428 ( 
.A(n_3661),
.Y(n_4428)
);

INVx3_ASAP7_75t_SL g4429 ( 
.A(n_3849),
.Y(n_4429)
);

NAND2xp5_ASAP7_75t_SL g4430 ( 
.A(n_3783),
.B(n_3091),
.Y(n_4430)
);

NOR2xp33_ASAP7_75t_L g4431 ( 
.A(n_4011),
.B(n_172),
.Y(n_4431)
);

AOI22xp33_ASAP7_75t_L g4432 ( 
.A1(n_3574),
.A2(n_3666),
.B1(n_3828),
.B2(n_3819),
.Y(n_4432)
);

NAND2xp5_ASAP7_75t_L g4433 ( 
.A(n_3484),
.B(n_172),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_L g4434 ( 
.A(n_3486),
.B(n_173),
.Y(n_4434)
);

INVx1_ASAP7_75t_L g4435 ( 
.A(n_3661),
.Y(n_4435)
);

INVx1_ASAP7_75t_L g4436 ( 
.A(n_3790),
.Y(n_4436)
);

NAND2xp5_ASAP7_75t_L g4437 ( 
.A(n_3501),
.B(n_173),
.Y(n_4437)
);

INVx2_ASAP7_75t_L g4438 ( 
.A(n_3903),
.Y(n_4438)
);

INVx1_ASAP7_75t_SL g4439 ( 
.A(n_3837),
.Y(n_4439)
);

INVx1_ASAP7_75t_L g4440 ( 
.A(n_3813),
.Y(n_4440)
);

NOR2xp33_ASAP7_75t_L g4441 ( 
.A(n_3999),
.B(n_173),
.Y(n_4441)
);

INVx2_ASAP7_75t_L g4442 ( 
.A(n_3916),
.Y(n_4442)
);

AOI22xp5_ASAP7_75t_L g4443 ( 
.A1(n_3490),
.A2(n_3430),
.B1(n_3452),
.B2(n_3143),
.Y(n_4443)
);

NAND2xp5_ASAP7_75t_L g4444 ( 
.A(n_3504),
.B(n_3844),
.Y(n_4444)
);

INVx4_ASAP7_75t_L g4445 ( 
.A(n_3840),
.Y(n_4445)
);

BUFx2_ASAP7_75t_L g4446 ( 
.A(n_3920),
.Y(n_4446)
);

INVx1_ASAP7_75t_L g4447 ( 
.A(n_3848),
.Y(n_4447)
);

BUFx8_ASAP7_75t_L g4448 ( 
.A(n_3959),
.Y(n_4448)
);

BUFx6f_ASAP7_75t_L g4449 ( 
.A(n_3840),
.Y(n_4449)
);

NAND2xp5_ASAP7_75t_SL g4450 ( 
.A(n_3556),
.B(n_3093),
.Y(n_4450)
);

INVx1_ASAP7_75t_L g4451 ( 
.A(n_3850),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_L g4452 ( 
.A(n_3909),
.B(n_174),
.Y(n_4452)
);

OR2x6_ASAP7_75t_L g4453 ( 
.A(n_3492),
.B(n_2891),
.Y(n_4453)
);

CKINVDCx5p33_ASAP7_75t_R g4454 ( 
.A(n_3766),
.Y(n_4454)
);

INVxp33_ASAP7_75t_SL g4455 ( 
.A(n_3540),
.Y(n_4455)
);

INVx2_ASAP7_75t_SL g4456 ( 
.A(n_3981),
.Y(n_4456)
);

NAND2xp5_ASAP7_75t_L g4457 ( 
.A(n_3923),
.B(n_174),
.Y(n_4457)
);

INVx2_ASAP7_75t_L g4458 ( 
.A(n_3958),
.Y(n_4458)
);

BUFx6f_ASAP7_75t_L g4459 ( 
.A(n_3912),
.Y(n_4459)
);

BUFx6f_ASAP7_75t_L g4460 ( 
.A(n_3912),
.Y(n_4460)
);

NAND2xp5_ASAP7_75t_L g4461 ( 
.A(n_3459),
.B(n_175),
.Y(n_4461)
);

NOR2xp33_ASAP7_75t_L g4462 ( 
.A(n_4023),
.B(n_4002),
.Y(n_4462)
);

AND2x4_ASAP7_75t_L g4463 ( 
.A(n_3773),
.B(n_2891),
.Y(n_4463)
);

OR2x6_ASAP7_75t_L g4464 ( 
.A(n_3495),
.B(n_2891),
.Y(n_4464)
);

INVx1_ASAP7_75t_L g4465 ( 
.A(n_3989),
.Y(n_4465)
);

NAND2xp5_ASAP7_75t_L g4466 ( 
.A(n_4009),
.B(n_175),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_L g4467 ( 
.A(n_3881),
.B(n_175),
.Y(n_4467)
);

BUFx6f_ASAP7_75t_L g4468 ( 
.A(n_3912),
.Y(n_4468)
);

AND2x2_ASAP7_75t_L g4469 ( 
.A(n_3990),
.B(n_176),
.Y(n_4469)
);

NAND2xp5_ASAP7_75t_L g4470 ( 
.A(n_3888),
.B(n_176),
.Y(n_4470)
);

BUFx6f_ASAP7_75t_L g4471 ( 
.A(n_3954),
.Y(n_4471)
);

AOI221xp5_ASAP7_75t_L g4472 ( 
.A1(n_3485),
.A2(n_3239),
.B1(n_3093),
.B2(n_3183),
.C(n_3152),
.Y(n_4472)
);

AOI22xp5_ASAP7_75t_L g4473 ( 
.A1(n_3833),
.A2(n_3143),
.B1(n_3152),
.B2(n_3093),
.Y(n_4473)
);

NOR2xp33_ASAP7_75t_L g4474 ( 
.A(n_3846),
.B(n_176),
.Y(n_4474)
);

NAND2xp5_ASAP7_75t_L g4475 ( 
.A(n_3891),
.B(n_177),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_3993),
.Y(n_4476)
);

OR2x6_ASAP7_75t_L g4477 ( 
.A(n_3690),
.B(n_2906),
.Y(n_4477)
);

AND2x2_ASAP7_75t_L g4478 ( 
.A(n_3971),
.B(n_3927),
.Y(n_4478)
);

NOR2xp33_ASAP7_75t_L g4479 ( 
.A(n_3851),
.B(n_177),
.Y(n_4479)
);

NAND2xp5_ASAP7_75t_L g4480 ( 
.A(n_3906),
.B(n_178),
.Y(n_4480)
);

OR2x2_ASAP7_75t_L g4481 ( 
.A(n_3926),
.B(n_178),
.Y(n_4481)
);

NAND2xp5_ASAP7_75t_L g4482 ( 
.A(n_3907),
.B(n_179),
.Y(n_4482)
);

INVx2_ASAP7_75t_L g4483 ( 
.A(n_4027),
.Y(n_4483)
);

INVx2_ASAP7_75t_L g4484 ( 
.A(n_3605),
.Y(n_4484)
);

INVx1_ASAP7_75t_L g4485 ( 
.A(n_3510),
.Y(n_4485)
);

NAND2xp5_ASAP7_75t_L g4486 ( 
.A(n_3910),
.B(n_179),
.Y(n_4486)
);

OAI22xp5_ASAP7_75t_L g4487 ( 
.A1(n_3629),
.A2(n_3143),
.B1(n_3183),
.B2(n_3152),
.Y(n_4487)
);

NAND2xp5_ASAP7_75t_L g4488 ( 
.A(n_3934),
.B(n_179),
.Y(n_4488)
);

NAND2xp5_ASAP7_75t_SL g4489 ( 
.A(n_3559),
.B(n_3183),
.Y(n_4489)
);

BUFx4f_ASAP7_75t_L g4490 ( 
.A(n_3935),
.Y(n_4490)
);

INVxp67_ASAP7_75t_SL g4491 ( 
.A(n_4005),
.Y(n_4491)
);

NAND2xp5_ASAP7_75t_L g4492 ( 
.A(n_3950),
.B(n_180),
.Y(n_4492)
);

OAI21xp33_ASAP7_75t_L g4493 ( 
.A1(n_3515),
.A2(n_3231),
.B(n_3187),
.Y(n_4493)
);

AND2x4_ASAP7_75t_L g4494 ( 
.A(n_4004),
.B(n_2906),
.Y(n_4494)
);

AND2x2_ASAP7_75t_L g4495 ( 
.A(n_3843),
.B(n_180),
.Y(n_4495)
);

HB1xp67_ASAP7_75t_L g4496 ( 
.A(n_3855),
.Y(n_4496)
);

INVx1_ASAP7_75t_L g4497 ( 
.A(n_3518),
.Y(n_4497)
);

INVxp67_ASAP7_75t_L g4498 ( 
.A(n_3952),
.Y(n_4498)
);

INVx1_ASAP7_75t_L g4499 ( 
.A(n_3795),
.Y(n_4499)
);

AOI22xp5_ASAP7_75t_L g4500 ( 
.A1(n_3968),
.A2(n_3231),
.B1(n_3239),
.B2(n_3187),
.Y(n_4500)
);

NOR2xp33_ASAP7_75t_L g4501 ( 
.A(n_3985),
.B(n_180),
.Y(n_4501)
);

AO22x1_ASAP7_75t_L g4502 ( 
.A1(n_3986),
.A2(n_2939),
.B1(n_2906),
.B2(n_3187),
.Y(n_4502)
);

AOI22xp5_ASAP7_75t_L g4503 ( 
.A1(n_3987),
.A2(n_3231),
.B1(n_3239),
.B2(n_2939),
.Y(n_4503)
);

INVx3_ASAP7_75t_L g4504 ( 
.A(n_3954),
.Y(n_4504)
);

INVx2_ASAP7_75t_SL g4505 ( 
.A(n_3937),
.Y(n_4505)
);

INVx2_ASAP7_75t_L g4506 ( 
.A(n_3617),
.Y(n_4506)
);

NAND2xp5_ASAP7_75t_L g4507 ( 
.A(n_3553),
.B(n_181),
.Y(n_4507)
);

NAND2xp5_ASAP7_75t_L g4508 ( 
.A(n_4019),
.B(n_181),
.Y(n_4508)
);

AND2x4_ASAP7_75t_L g4509 ( 
.A(n_4020),
.B(n_2939),
.Y(n_4509)
);

INVx2_ASAP7_75t_L g4510 ( 
.A(n_3643),
.Y(n_4510)
);

INVx1_ASAP7_75t_L g4511 ( 
.A(n_3799),
.Y(n_4511)
);

BUFx4f_ASAP7_75t_L g4512 ( 
.A(n_3939),
.Y(n_4512)
);

NAND2xp5_ASAP7_75t_SL g4513 ( 
.A(n_3954),
.B(n_181),
.Y(n_4513)
);

AOI22xp5_ASAP7_75t_L g4514 ( 
.A1(n_3629),
.A2(n_183),
.B1(n_184),
.B2(n_182),
.Y(n_4514)
);

BUFx6f_ASAP7_75t_L g4515 ( 
.A(n_3974),
.Y(n_4515)
);

BUFx6f_ASAP7_75t_SL g4516 ( 
.A(n_3941),
.Y(n_4516)
);

NAND2xp5_ASAP7_75t_L g4517 ( 
.A(n_4021),
.B(n_182),
.Y(n_4517)
);

NOR2xp33_ASAP7_75t_L g4518 ( 
.A(n_3994),
.B(n_184),
.Y(n_4518)
);

INVx1_ASAP7_75t_SL g4519 ( 
.A(n_3503),
.Y(n_4519)
);

INVx1_ASAP7_75t_L g4520 ( 
.A(n_3804),
.Y(n_4520)
);

HB1xp67_ASAP7_75t_L g4521 ( 
.A(n_3953),
.Y(n_4521)
);

INVx2_ASAP7_75t_L g4522 ( 
.A(n_3645),
.Y(n_4522)
);

NOR2xp33_ASAP7_75t_L g4523 ( 
.A(n_3996),
.B(n_3979),
.Y(n_4523)
);

NOR2xp33_ASAP7_75t_L g4524 ( 
.A(n_3929),
.B(n_3878),
.Y(n_4524)
);

INVx1_ASAP7_75t_L g4525 ( 
.A(n_3814),
.Y(n_4525)
);

INVx1_ASAP7_75t_L g4526 ( 
.A(n_3815),
.Y(n_4526)
);

INVx2_ASAP7_75t_L g4527 ( 
.A(n_3659),
.Y(n_4527)
);

INVx1_ASAP7_75t_L g4528 ( 
.A(n_3816),
.Y(n_4528)
);

NAND2xp5_ASAP7_75t_L g4529 ( 
.A(n_4025),
.B(n_184),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_L g4530 ( 
.A(n_4014),
.B(n_185),
.Y(n_4530)
);

INVx2_ASAP7_75t_L g4531 ( 
.A(n_3662),
.Y(n_4531)
);

AOI21xp5_ASAP7_75t_L g4532 ( 
.A1(n_4003),
.A2(n_186),
.B(n_185),
.Y(n_4532)
);

BUFx6f_ASAP7_75t_L g4533 ( 
.A(n_3974),
.Y(n_4533)
);

AOI22xp5_ASAP7_75t_L g4534 ( 
.A1(n_3862),
.A2(n_186),
.B1(n_187),
.B2(n_185),
.Y(n_4534)
);

INVx1_ASAP7_75t_L g4535 ( 
.A(n_3818),
.Y(n_4535)
);

NAND2xp5_ASAP7_75t_SL g4536 ( 
.A(n_3974),
.B(n_186),
.Y(n_4536)
);

NAND2xp5_ASAP7_75t_L g4537 ( 
.A(n_4017),
.B(n_187),
.Y(n_4537)
);

INVx2_ASAP7_75t_SL g4538 ( 
.A(n_3805),
.Y(n_4538)
);

OAI221xp5_ASAP7_75t_L g4539 ( 
.A1(n_3796),
.A2(n_189),
.B1(n_190),
.B2(n_188),
.C(n_187),
.Y(n_4539)
);

O2A1O1Ixp5_ASAP7_75t_L g4540 ( 
.A1(n_3599),
.A2(n_189),
.B(n_190),
.C(n_188),
.Y(n_4540)
);

INVx1_ASAP7_75t_L g4541 ( 
.A(n_3820),
.Y(n_4541)
);

NAND2xp5_ASAP7_75t_L g4542 ( 
.A(n_4022),
.B(n_188),
.Y(n_4542)
);

INVx2_ASAP7_75t_L g4543 ( 
.A(n_3668),
.Y(n_4543)
);

INVx5_ASAP7_75t_L g4544 ( 
.A(n_4018),
.Y(n_4544)
);

NAND2xp5_ASAP7_75t_SL g4545 ( 
.A(n_3499),
.B(n_191),
.Y(n_4545)
);

NAND2xp5_ASAP7_75t_L g4546 ( 
.A(n_4024),
.B(n_191),
.Y(n_4546)
);

AND2x2_ASAP7_75t_L g4547 ( 
.A(n_3880),
.B(n_1077),
.Y(n_4547)
);

NAND2xp5_ASAP7_75t_L g4548 ( 
.A(n_3465),
.B(n_191),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_3534),
.Y(n_4549)
);

INVx1_ASAP7_75t_L g4550 ( 
.A(n_3535),
.Y(n_4550)
);

BUFx3_ASAP7_75t_L g4551 ( 
.A(n_3547),
.Y(n_4551)
);

BUFx2_ASAP7_75t_L g4552 ( 
.A(n_3669),
.Y(n_4552)
);

BUFx3_ASAP7_75t_L g4553 ( 
.A(n_3676),
.Y(n_4553)
);

INVx1_ASAP7_75t_L g4554 ( 
.A(n_3677),
.Y(n_4554)
);

NAND2xp5_ASAP7_75t_L g4555 ( 
.A(n_3678),
.B(n_192),
.Y(n_4555)
);

AOI22xp5_ASAP7_75t_L g4556 ( 
.A1(n_3738),
.A2(n_193),
.B1(n_194),
.B2(n_192),
.Y(n_4556)
);

INVx2_ASAP7_75t_L g4557 ( 
.A(n_3688),
.Y(n_4557)
);

INVx2_ASAP7_75t_L g4558 ( 
.A(n_3695),
.Y(n_4558)
);

INVx3_ASAP7_75t_L g4559 ( 
.A(n_3697),
.Y(n_4559)
);

NAND2x1p5_ASAP7_75t_L g4560 ( 
.A(n_3809),
.B(n_200),
.Y(n_4560)
);

INVx1_ASAP7_75t_L g4561 ( 
.A(n_3700),
.Y(n_4561)
);

HB1xp67_ASAP7_75t_L g4562 ( 
.A(n_3874),
.Y(n_4562)
);

INVx1_ASAP7_75t_L g4563 ( 
.A(n_3705),
.Y(n_4563)
);

NAND3xp33_ASAP7_75t_SL g4564 ( 
.A(n_3918),
.B(n_2),
.C(n_3),
.Y(n_4564)
);

INVx2_ASAP7_75t_SL g4565 ( 
.A(n_3811),
.Y(n_4565)
);

INVx1_ASAP7_75t_L g4566 ( 
.A(n_3716),
.Y(n_4566)
);

NAND2xp5_ASAP7_75t_L g4567 ( 
.A(n_3717),
.B(n_193),
.Y(n_4567)
);

OAI22xp5_ASAP7_75t_L g4568 ( 
.A1(n_3781),
.A2(n_195),
.B1(n_196),
.B2(n_194),
.Y(n_4568)
);

INVx4_ASAP7_75t_L g4569 ( 
.A(n_3562),
.Y(n_4569)
);

NAND2xp5_ASAP7_75t_L g4570 ( 
.A(n_3719),
.B(n_195),
.Y(n_4570)
);

NAND2xp5_ASAP7_75t_L g4571 ( 
.A(n_3728),
.B(n_3729),
.Y(n_4571)
);

INVxp67_ASAP7_75t_L g4572 ( 
.A(n_3890),
.Y(n_4572)
);

INVx1_ASAP7_75t_L g4573 ( 
.A(n_3732),
.Y(n_4573)
);

CKINVDCx5p33_ASAP7_75t_R g4574 ( 
.A(n_3858),
.Y(n_4574)
);

NAND2xp5_ASAP7_75t_SL g4575 ( 
.A(n_3507),
.B(n_195),
.Y(n_4575)
);

BUFx3_ASAP7_75t_L g4576 ( 
.A(n_3735),
.Y(n_4576)
);

NOR2xp33_ASAP7_75t_L g4577 ( 
.A(n_3521),
.B(n_196),
.Y(n_4577)
);

OR2x6_ASAP7_75t_L g4578 ( 
.A(n_4016),
.B(n_4028),
.Y(n_4578)
);

CKINVDCx5p33_ASAP7_75t_R g4579 ( 
.A(n_4007),
.Y(n_4579)
);

NAND2xp5_ASAP7_75t_SL g4580 ( 
.A(n_3519),
.B(n_196),
.Y(n_4580)
);

NOR2xp33_ASAP7_75t_L g4581 ( 
.A(n_3531),
.B(n_3776),
.Y(n_4581)
);

INVx5_ASAP7_75t_L g4582 ( 
.A(n_3563),
.Y(n_4582)
);

NAND2xp5_ASAP7_75t_SL g4583 ( 
.A(n_3885),
.B(n_3894),
.Y(n_4583)
);

BUFx2_ASAP7_75t_L g4584 ( 
.A(n_3737),
.Y(n_4584)
);

NAND2x1p5_ASAP7_75t_L g4585 ( 
.A(n_3854),
.B(n_197),
.Y(n_4585)
);

INVx1_ASAP7_75t_L g4586 ( 
.A(n_3741),
.Y(n_4586)
);

NAND2xp5_ASAP7_75t_SL g4587 ( 
.A(n_3578),
.B(n_197),
.Y(n_4587)
);

INVx1_ASAP7_75t_L g4588 ( 
.A(n_3743),
.Y(n_4588)
);

INVx1_ASAP7_75t_L g4589 ( 
.A(n_3745),
.Y(n_4589)
);

NAND2xp5_ASAP7_75t_L g4590 ( 
.A(n_3749),
.B(n_198),
.Y(n_4590)
);

NAND2xp5_ASAP7_75t_L g4591 ( 
.A(n_3764),
.B(n_198),
.Y(n_4591)
);

NAND2xp5_ASAP7_75t_SL g4592 ( 
.A(n_3581),
.B(n_198),
.Y(n_4592)
);

NOR2xp33_ASAP7_75t_L g4593 ( 
.A(n_3723),
.B(n_199),
.Y(n_4593)
);

BUFx2_ASAP7_75t_L g4594 ( 
.A(n_3771),
.Y(n_4594)
);

INVx2_ASAP7_75t_SL g4595 ( 
.A(n_3585),
.Y(n_4595)
);

NAND2xp5_ASAP7_75t_SL g4596 ( 
.A(n_3497),
.B(n_199),
.Y(n_4596)
);

INVx2_ASAP7_75t_L g4597 ( 
.A(n_3775),
.Y(n_4597)
);

NOR2xp33_ASAP7_75t_L g4598 ( 
.A(n_3727),
.B(n_199),
.Y(n_4598)
);

OAI21x1_ASAP7_75t_L g4599 ( 
.A1(n_3551),
.A2(n_202),
.B(n_201),
.Y(n_4599)
);

INVx2_ASAP7_75t_L g4600 ( 
.A(n_4033),
.Y(n_4600)
);

NAND2x1p5_ASAP7_75t_L g4601 ( 
.A(n_4061),
.B(n_3758),
.Y(n_4601)
);

NAND2xp5_ASAP7_75t_L g4602 ( 
.A(n_4485),
.B(n_3780),
.Y(n_4602)
);

AOI22xp5_ASAP7_75t_L g4603 ( 
.A1(n_4054),
.A2(n_3784),
.B1(n_3898),
.B2(n_3694),
.Y(n_4603)
);

AOI22xp5_ASAP7_75t_L g4604 ( 
.A1(n_4574),
.A2(n_3634),
.B1(n_3609),
.B2(n_3892),
.Y(n_4604)
);

AOI21xp5_ASAP7_75t_L g4605 ( 
.A1(n_4085),
.A2(n_3969),
.B(n_3967),
.Y(n_4605)
);

OAI21xp5_ASAP7_75t_L g4606 ( 
.A1(n_4076),
.A2(n_3608),
.B(n_3886),
.Y(n_4606)
);

NAND2xp5_ASAP7_75t_L g4607 ( 
.A(n_4497),
.B(n_3786),
.Y(n_4607)
);

AOI22xp33_ASAP7_75t_L g4608 ( 
.A1(n_4410),
.A2(n_3908),
.B1(n_3911),
.B2(n_3904),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_4032),
.Y(n_4609)
);

AND2x2_ASAP7_75t_L g4610 ( 
.A(n_4198),
.B(n_200),
.Y(n_4610)
);

INVx1_ASAP7_75t_L g4611 ( 
.A(n_4038),
.Y(n_4611)
);

AOI21x1_ASAP7_75t_L g4612 ( 
.A1(n_4095),
.A2(n_3932),
.B(n_3917),
.Y(n_4612)
);

INVx4_ASAP7_75t_L g4613 ( 
.A(n_4061),
.Y(n_4613)
);

NAND2xp5_ASAP7_75t_SL g4614 ( 
.A(n_4175),
.B(n_4006),
.Y(n_4614)
);

NAND3xp33_ASAP7_75t_L g4615 ( 
.A(n_4431),
.B(n_3965),
.C(n_3839),
.Y(n_4615)
);

NAND2xp5_ASAP7_75t_SL g4616 ( 
.A(n_4175),
.B(n_3883),
.Y(n_4616)
);

HB1xp67_ASAP7_75t_L g4617 ( 
.A(n_4090),
.Y(n_4617)
);

OAI22xp5_ASAP7_75t_L g4618 ( 
.A1(n_4319),
.A2(n_3791),
.B1(n_3789),
.B2(n_3938),
.Y(n_4618)
);

AOI21xp5_ASAP7_75t_L g4619 ( 
.A1(n_4134),
.A2(n_3970),
.B(n_3961),
.Y(n_4619)
);

NOR2x1_ASAP7_75t_L g4620 ( 
.A(n_4080),
.B(n_4115),
.Y(n_4620)
);

AO31x2_ASAP7_75t_L g4621 ( 
.A1(n_4487),
.A2(n_4274),
.A3(n_4483),
.B(n_4392),
.Y(n_4621)
);

O2A1O1Ixp33_ASAP7_75t_L g4622 ( 
.A1(n_4079),
.A2(n_3663),
.B(n_3949),
.C(n_3942),
.Y(n_4622)
);

NOR2xp33_ASAP7_75t_L g4623 ( 
.A(n_4374),
.B(n_202),
.Y(n_4623)
);

NAND2xp5_ASAP7_75t_L g4624 ( 
.A(n_4478),
.B(n_3580),
.Y(n_4624)
);

INVx2_ASAP7_75t_L g4625 ( 
.A(n_4037),
.Y(n_4625)
);

BUFx6f_ASAP7_75t_L g4626 ( 
.A(n_4061),
.Y(n_4626)
);

NAND2xp5_ASAP7_75t_L g4627 ( 
.A(n_4045),
.B(n_3583),
.Y(n_4627)
);

BUFx8_ASAP7_75t_L g4628 ( 
.A(n_4197),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_4048),
.Y(n_4629)
);

NOR2xp33_ASAP7_75t_SL g4630 ( 
.A(n_4080),
.B(n_4073),
.Y(n_4630)
);

NAND2xp5_ASAP7_75t_L g4631 ( 
.A(n_4049),
.B(n_3587),
.Y(n_4631)
);

NAND2xp5_ASAP7_75t_L g4632 ( 
.A(n_4050),
.B(n_3590),
.Y(n_4632)
);

AOI21xp5_ASAP7_75t_L g4633 ( 
.A1(n_4244),
.A2(n_3978),
.B(n_3951),
.Y(n_4633)
);

NOR2xp33_ASAP7_75t_L g4634 ( 
.A(n_4073),
.B(n_202),
.Y(n_4634)
);

NOR2x1_ASAP7_75t_L g4635 ( 
.A(n_4130),
.B(n_4150),
.Y(n_4635)
);

AND2x2_ASAP7_75t_L g4636 ( 
.A(n_4158),
.B(n_203),
.Y(n_4636)
);

NAND2xp5_ASAP7_75t_L g4637 ( 
.A(n_4068),
.B(n_3601),
.Y(n_4637)
);

AND2x2_ASAP7_75t_L g4638 ( 
.A(n_4395),
.B(n_4414),
.Y(n_4638)
);

AOI21xp5_ASAP7_75t_L g4639 ( 
.A1(n_4248),
.A2(n_3984),
.B(n_3980),
.Y(n_4639)
);

O2A1O1Ixp5_ASAP7_75t_L g4640 ( 
.A1(n_4324),
.A2(n_3866),
.B(n_3542),
.C(n_204),
.Y(n_4640)
);

AOI21xp5_ASAP7_75t_L g4641 ( 
.A1(n_4147),
.A2(n_204),
.B(n_203),
.Y(n_4641)
);

AOI21xp5_ASAP7_75t_L g4642 ( 
.A1(n_4260),
.A2(n_205),
.B(n_204),
.Y(n_4642)
);

AOI21xp5_ASAP7_75t_L g4643 ( 
.A1(n_4386),
.A2(n_4403),
.B(n_4502),
.Y(n_4643)
);

AOI21xp5_ASAP7_75t_L g4644 ( 
.A1(n_4430),
.A2(n_206),
.B(n_205),
.Y(n_4644)
);

INVx2_ASAP7_75t_L g4645 ( 
.A(n_4055),
.Y(n_4645)
);

NAND2xp5_ASAP7_75t_L g4646 ( 
.A(n_4093),
.B(n_4103),
.Y(n_4646)
);

NAND2xp5_ASAP7_75t_L g4647 ( 
.A(n_4107),
.B(n_205),
.Y(n_4647)
);

NOR2xp33_ASAP7_75t_SL g4648 ( 
.A(n_4170),
.B(n_206),
.Y(n_4648)
);

O2A1O1Ixp33_ASAP7_75t_L g4649 ( 
.A1(n_4427),
.A2(n_207),
.B(n_208),
.C(n_206),
.Y(n_4649)
);

O2A1O1Ixp5_ASAP7_75t_L g4650 ( 
.A1(n_4265),
.A2(n_208),
.B(n_209),
.C(n_207),
.Y(n_4650)
);

OAI22xp5_ASAP7_75t_SL g4651 ( 
.A1(n_4302),
.A2(n_210),
.B1(n_211),
.B2(n_209),
.Y(n_4651)
);

A2O1A1Ixp33_ASAP7_75t_L g4652 ( 
.A1(n_4203),
.A2(n_211),
.B(n_212),
.C(n_210),
.Y(n_4652)
);

INVx1_ASAP7_75t_L g4653 ( 
.A(n_4120),
.Y(n_4653)
);

AOI21xp5_ASAP7_75t_L g4654 ( 
.A1(n_4257),
.A2(n_211),
.B(n_210),
.Y(n_4654)
);

AOI21xp5_ASAP7_75t_L g4655 ( 
.A1(n_4089),
.A2(n_213),
.B(n_212),
.Y(n_4655)
);

OAI21x1_ASAP7_75t_L g4656 ( 
.A1(n_4182),
.A2(n_213),
.B(n_212),
.Y(n_4656)
);

O2A1O1Ixp33_ASAP7_75t_L g4657 ( 
.A1(n_4067),
.A2(n_215),
.B(n_216),
.C(n_214),
.Y(n_4657)
);

AND2x2_ASAP7_75t_L g4658 ( 
.A(n_4226),
.B(n_4384),
.Y(n_4658)
);

HB1xp67_ASAP7_75t_L g4659 ( 
.A(n_4145),
.Y(n_4659)
);

AO22x1_ASAP7_75t_L g4660 ( 
.A1(n_4170),
.A2(n_215),
.B1(n_216),
.B2(n_214),
.Y(n_4660)
);

OAI21x1_ASAP7_75t_L g4661 ( 
.A1(n_4363),
.A2(n_216),
.B(n_215),
.Y(n_4661)
);

NAND2xp5_ASAP7_75t_L g4662 ( 
.A(n_4146),
.B(n_217),
.Y(n_4662)
);

OAI22xp5_ASAP7_75t_L g4663 ( 
.A1(n_4319),
.A2(n_4307),
.B1(n_4064),
.B2(n_4175),
.Y(n_4663)
);

AOI21xp5_ASAP7_75t_L g4664 ( 
.A1(n_4421),
.A2(n_219),
.B(n_218),
.Y(n_4664)
);

AND2x2_ASAP7_75t_SL g4665 ( 
.A(n_4313),
.B(n_218),
.Y(n_4665)
);

AOI22xp5_ASAP7_75t_L g4666 ( 
.A1(n_4579),
.A2(n_1075),
.B1(n_1076),
.B2(n_1074),
.Y(n_4666)
);

A2O1A1Ixp33_ASAP7_75t_L g4667 ( 
.A1(n_4342),
.A2(n_220),
.B(n_221),
.C(n_219),
.Y(n_4667)
);

NAND2xp5_ASAP7_75t_L g4668 ( 
.A(n_4156),
.B(n_220),
.Y(n_4668)
);

INVx1_ASAP7_75t_L g4669 ( 
.A(n_4157),
.Y(n_4669)
);

AOI21xp5_ASAP7_75t_L g4670 ( 
.A1(n_4421),
.A2(n_221),
.B(n_220),
.Y(n_4670)
);

OAI22xp5_ASAP7_75t_L g4671 ( 
.A1(n_4310),
.A2(n_222),
.B1(n_223),
.B2(n_221),
.Y(n_4671)
);

INVx2_ASAP7_75t_L g4672 ( 
.A(n_4056),
.Y(n_4672)
);

NOR2xp33_ASAP7_75t_L g4673 ( 
.A(n_4390),
.B(n_223),
.Y(n_4673)
);

INVx2_ASAP7_75t_L g4674 ( 
.A(n_4062),
.Y(n_4674)
);

NOR2xp33_ASAP7_75t_L g4675 ( 
.A(n_4397),
.B(n_223),
.Y(n_4675)
);

NAND2xp5_ASAP7_75t_L g4676 ( 
.A(n_4160),
.B(n_224),
.Y(n_4676)
);

NAND2xp5_ASAP7_75t_SL g4677 ( 
.A(n_4318),
.B(n_4263),
.Y(n_4677)
);

INVx4_ASAP7_75t_L g4678 ( 
.A(n_4122),
.Y(n_4678)
);

INVx2_ASAP7_75t_L g4679 ( 
.A(n_4181),
.Y(n_4679)
);

OAI21xp5_ASAP7_75t_L g4680 ( 
.A1(n_4540),
.A2(n_226),
.B(n_225),
.Y(n_4680)
);

AOI21xp5_ASAP7_75t_L g4681 ( 
.A1(n_4165),
.A2(n_226),
.B(n_225),
.Y(n_4681)
);

BUFx3_ASAP7_75t_L g4682 ( 
.A(n_4052),
.Y(n_4682)
);

NAND2xp5_ASAP7_75t_L g4683 ( 
.A(n_4163),
.B(n_4185),
.Y(n_4683)
);

AOI21xp5_ASAP7_75t_L g4684 ( 
.A1(n_4169),
.A2(n_227),
.B(n_225),
.Y(n_4684)
);

INVx2_ASAP7_75t_L g4685 ( 
.A(n_4194),
.Y(n_4685)
);

OAI21x1_ASAP7_75t_L g4686 ( 
.A1(n_4361),
.A2(n_228),
.B(n_227),
.Y(n_4686)
);

A2O1A1Ixp33_ASAP7_75t_L g4687 ( 
.A1(n_4345),
.A2(n_229),
.B(n_230),
.C(n_227),
.Y(n_4687)
);

INVx3_ASAP7_75t_L g4688 ( 
.A(n_4122),
.Y(n_4688)
);

A2O1A1Ixp33_ASAP7_75t_L g4689 ( 
.A1(n_4105),
.A2(n_230),
.B(n_231),
.C(n_229),
.Y(n_4689)
);

INVx2_ASAP7_75t_SL g4690 ( 
.A(n_4066),
.Y(n_4690)
);

AND2x2_ASAP7_75t_L g4691 ( 
.A(n_4388),
.B(n_229),
.Y(n_4691)
);

AO32x2_ASAP7_75t_L g4692 ( 
.A1(n_4355),
.A2(n_246),
.A3(n_254),
.B1(n_238),
.B2(n_230),
.Y(n_4692)
);

NAND2xp5_ASAP7_75t_L g4693 ( 
.A(n_4212),
.B(n_231),
.Y(n_4693)
);

NAND2xp5_ASAP7_75t_SL g4694 ( 
.A(n_4188),
.B(n_231),
.Y(n_4694)
);

CKINVDCx20_ASAP7_75t_R g4695 ( 
.A(n_4057),
.Y(n_4695)
);

AOI21xp5_ASAP7_75t_L g4696 ( 
.A1(n_4096),
.A2(n_233),
.B(n_232),
.Y(n_4696)
);

AOI21xp5_ASAP7_75t_L g4697 ( 
.A1(n_4310),
.A2(n_233),
.B(n_232),
.Y(n_4697)
);

AND2x4_ASAP7_75t_L g4698 ( 
.A(n_4122),
.B(n_232),
.Y(n_4698)
);

AOI22xp5_ASAP7_75t_L g4699 ( 
.A1(n_4034),
.A2(n_1076),
.B1(n_1077),
.B2(n_1073),
.Y(n_4699)
);

OAI22xp5_ASAP7_75t_L g4700 ( 
.A1(n_4043),
.A2(n_235),
.B1(n_236),
.B2(n_234),
.Y(n_4700)
);

AOI21xp5_ASAP7_75t_L g4701 ( 
.A1(n_4282),
.A2(n_235),
.B(n_234),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4217),
.Y(n_4702)
);

NAND2xp5_ASAP7_75t_L g4703 ( 
.A(n_4221),
.B(n_234),
.Y(n_4703)
);

HB1xp67_ASAP7_75t_L g4704 ( 
.A(n_4161),
.Y(n_4704)
);

AOI21x1_ASAP7_75t_L g4705 ( 
.A1(n_4415),
.A2(n_4151),
.B(n_4124),
.Y(n_4705)
);

AND2x2_ASAP7_75t_L g4706 ( 
.A(n_4422),
.B(n_235),
.Y(n_4706)
);

NAND2xp5_ASAP7_75t_SL g4707 ( 
.A(n_4131),
.B(n_236),
.Y(n_4707)
);

NOR2xp33_ASAP7_75t_L g4708 ( 
.A(n_4389),
.B(n_236),
.Y(n_4708)
);

NAND2xp5_ASAP7_75t_L g4709 ( 
.A(n_4227),
.B(n_237),
.Y(n_4709)
);

NAND2xp5_ASAP7_75t_L g4710 ( 
.A(n_4249),
.B(n_237),
.Y(n_4710)
);

INVx2_ASAP7_75t_L g4711 ( 
.A(n_4195),
.Y(n_4711)
);

AOI21xp5_ASAP7_75t_L g4712 ( 
.A1(n_4220),
.A2(n_238),
.B(n_237),
.Y(n_4712)
);

AOI21x1_ASAP7_75t_L g4713 ( 
.A1(n_4415),
.A2(n_240),
.B(n_239),
.Y(n_4713)
);

BUFx4f_ASAP7_75t_L g4714 ( 
.A(n_4082),
.Y(n_4714)
);

NOR2xp33_ASAP7_75t_L g4715 ( 
.A(n_4162),
.B(n_4429),
.Y(n_4715)
);

NAND2x1p5_ASAP7_75t_L g4716 ( 
.A(n_4192),
.B(n_239),
.Y(n_4716)
);

NAND2xp5_ASAP7_75t_L g4717 ( 
.A(n_4255),
.B(n_241),
.Y(n_4717)
);

OAI21xp5_ASAP7_75t_L g4718 ( 
.A1(n_4126),
.A2(n_242),
.B(n_241),
.Y(n_4718)
);

AND2x2_ASAP7_75t_L g4719 ( 
.A(n_4446),
.B(n_241),
.Y(n_4719)
);

AOI22xp5_ASAP7_75t_L g4720 ( 
.A1(n_4201),
.A2(n_1065),
.B1(n_1066),
.B2(n_1064),
.Y(n_4720)
);

BUFx6f_ASAP7_75t_L g4721 ( 
.A(n_4081),
.Y(n_4721)
);

AOI21xp33_ASAP7_75t_L g4722 ( 
.A1(n_4581),
.A2(n_243),
.B(n_242),
.Y(n_4722)
);

OAI22xp5_ASAP7_75t_L g4723 ( 
.A1(n_4078),
.A2(n_243),
.B1(n_244),
.B2(n_242),
.Y(n_4723)
);

INVx1_ASAP7_75t_L g4724 ( 
.A(n_4270),
.Y(n_4724)
);

NAND2xp5_ASAP7_75t_L g4725 ( 
.A(n_4278),
.B(n_245),
.Y(n_4725)
);

NAND2xp5_ASAP7_75t_L g4726 ( 
.A(n_4280),
.B(n_245),
.Y(n_4726)
);

AOI21xp5_ASAP7_75t_L g4727 ( 
.A1(n_4223),
.A2(n_246),
.B(n_245),
.Y(n_4727)
);

NAND2xp5_ASAP7_75t_L g4728 ( 
.A(n_4311),
.B(n_247),
.Y(n_4728)
);

CKINVDCx20_ASAP7_75t_R g4729 ( 
.A(n_4173),
.Y(n_4729)
);

AOI21xp5_ASAP7_75t_L g4730 ( 
.A1(n_4236),
.A2(n_248),
.B(n_247),
.Y(n_4730)
);

BUFx6f_ASAP7_75t_L g4731 ( 
.A(n_4081),
.Y(n_4731)
);

NAND2xp5_ASAP7_75t_L g4732 ( 
.A(n_4315),
.B(n_247),
.Y(n_4732)
);

INVx1_ASAP7_75t_L g4733 ( 
.A(n_4316),
.Y(n_4733)
);

AOI21xp5_ASAP7_75t_L g4734 ( 
.A1(n_4240),
.A2(n_249),
.B(n_248),
.Y(n_4734)
);

BUFx2_ASAP7_75t_L g4735 ( 
.A(n_4077),
.Y(n_4735)
);

AOI21xp5_ASAP7_75t_L g4736 ( 
.A1(n_4472),
.A2(n_249),
.B(n_248),
.Y(n_4736)
);

INVx2_ASAP7_75t_L g4737 ( 
.A(n_4206),
.Y(n_4737)
);

NOR2x1_ASAP7_75t_L g4738 ( 
.A(n_4213),
.B(n_249),
.Y(n_4738)
);

AO21x1_ASAP7_75t_L g4739 ( 
.A1(n_4428),
.A2(n_251),
.B(n_250),
.Y(n_4739)
);

NAND2xp5_ASAP7_75t_L g4740 ( 
.A(n_4317),
.B(n_250),
.Y(n_4740)
);

NAND2xp5_ASAP7_75t_SL g4741 ( 
.A(n_4149),
.B(n_250),
.Y(n_4741)
);

AOI21xp5_ASAP7_75t_L g4742 ( 
.A1(n_4450),
.A2(n_252),
.B(n_251),
.Y(n_4742)
);

INVx1_ASAP7_75t_L g4743 ( 
.A(n_4320),
.Y(n_4743)
);

A2O1A1Ixp33_ASAP7_75t_L g4744 ( 
.A1(n_4304),
.A2(n_252),
.B(n_253),
.C(n_251),
.Y(n_4744)
);

NAND2xp5_ASAP7_75t_L g4745 ( 
.A(n_4326),
.B(n_253),
.Y(n_4745)
);

AOI21xp5_ASAP7_75t_L g4746 ( 
.A1(n_4489),
.A2(n_254),
.B(n_253),
.Y(n_4746)
);

AOI21x1_ASAP7_75t_L g4747 ( 
.A1(n_4435),
.A2(n_255),
.B(n_254),
.Y(n_4747)
);

INVx2_ASAP7_75t_L g4748 ( 
.A(n_4251),
.Y(n_4748)
);

NAND2xp5_ASAP7_75t_L g4749 ( 
.A(n_4330),
.B(n_255),
.Y(n_4749)
);

O2A1O1Ixp33_ASAP7_75t_SL g4750 ( 
.A1(n_4178),
.A2(n_257),
.B(n_258),
.C(n_256),
.Y(n_4750)
);

AND2x2_ASAP7_75t_L g4751 ( 
.A(n_4238),
.B(n_257),
.Y(n_4751)
);

AOI21xp5_ASAP7_75t_L g4752 ( 
.A1(n_4493),
.A2(n_258),
.B(n_257),
.Y(n_4752)
);

NOR2x1_ASAP7_75t_L g4753 ( 
.A(n_4213),
.B(n_258),
.Y(n_4753)
);

BUFx3_ASAP7_75t_L g4754 ( 
.A(n_4110),
.Y(n_4754)
);

A2O1A1Ixp33_ASAP7_75t_L g4755 ( 
.A1(n_4241),
.A2(n_260),
.B(n_261),
.C(n_259),
.Y(n_4755)
);

INVx1_ASAP7_75t_L g4756 ( 
.A(n_4337),
.Y(n_4756)
);

NAND2xp5_ASAP7_75t_L g4757 ( 
.A(n_4338),
.B(n_4349),
.Y(n_4757)
);

OAI21x1_ASAP7_75t_L g4758 ( 
.A1(n_4411),
.A2(n_261),
.B(n_260),
.Y(n_4758)
);

INVx3_ASAP7_75t_L g4759 ( 
.A(n_4189),
.Y(n_4759)
);

NAND2xp5_ASAP7_75t_L g4760 ( 
.A(n_4352),
.B(n_260),
.Y(n_4760)
);

OAI21xp5_ASAP7_75t_L g4761 ( 
.A1(n_4187),
.A2(n_4564),
.B(n_4432),
.Y(n_4761)
);

INVx1_ASAP7_75t_L g4762 ( 
.A(n_4354),
.Y(n_4762)
);

INVx2_ASAP7_75t_L g4763 ( 
.A(n_4254),
.Y(n_4763)
);

AOI22xp5_ASAP7_75t_L g4764 ( 
.A1(n_4551),
.A2(n_1072),
.B1(n_1073),
.B2(n_1071),
.Y(n_4764)
);

AOI21xp5_ASAP7_75t_L g4765 ( 
.A1(n_4379),
.A2(n_263),
.B(n_262),
.Y(n_4765)
);

INVx3_ASAP7_75t_L g4766 ( 
.A(n_4081),
.Y(n_4766)
);

INVx2_ASAP7_75t_L g4767 ( 
.A(n_4268),
.Y(n_4767)
);

INVx1_ASAP7_75t_L g4768 ( 
.A(n_4356),
.Y(n_4768)
);

AO21x1_ASAP7_75t_L g4769 ( 
.A1(n_4106),
.A2(n_263),
.B(n_262),
.Y(n_4769)
);

AOI21xp5_ASAP7_75t_L g4770 ( 
.A1(n_4243),
.A2(n_264),
.B(n_263),
.Y(n_4770)
);

AND2x4_ASAP7_75t_L g4771 ( 
.A(n_4166),
.B(n_265),
.Y(n_4771)
);

NAND2xp5_ASAP7_75t_L g4772 ( 
.A(n_4367),
.B(n_265),
.Y(n_4772)
);

INVx2_ASAP7_75t_L g4773 ( 
.A(n_4269),
.Y(n_4773)
);

INVx1_ASAP7_75t_SL g4774 ( 
.A(n_4111),
.Y(n_4774)
);

OR2x6_ASAP7_75t_SL g4775 ( 
.A(n_4279),
.B(n_1055),
.Y(n_4775)
);

NAND3xp33_ASAP7_75t_L g4776 ( 
.A(n_4424),
.B(n_267),
.C(n_266),
.Y(n_4776)
);

AOI21xp5_ASAP7_75t_L g4777 ( 
.A1(n_4252),
.A2(n_267),
.B(n_266),
.Y(n_4777)
);

OAI21xp5_ASAP7_75t_L g4778 ( 
.A1(n_4144),
.A2(n_267),
.B(n_266),
.Y(n_4778)
);

OAI21xp5_ASAP7_75t_L g4779 ( 
.A1(n_4224),
.A2(n_269),
.B(n_268),
.Y(n_4779)
);

INVx2_ASAP7_75t_L g4780 ( 
.A(n_4285),
.Y(n_4780)
);

NAND2xp5_ASAP7_75t_L g4781 ( 
.A(n_4369),
.B(n_268),
.Y(n_4781)
);

NAND2xp5_ASAP7_75t_L g4782 ( 
.A(n_4370),
.B(n_268),
.Y(n_4782)
);

AOI221xp5_ASAP7_75t_L g4783 ( 
.A1(n_4577),
.A2(n_4441),
.B1(n_4088),
.B2(n_4518),
.C(n_4501),
.Y(n_4783)
);

NOR3xp33_ASAP7_75t_L g4784 ( 
.A(n_4129),
.B(n_277),
.C(n_269),
.Y(n_4784)
);

HB1xp67_ASAP7_75t_L g4785 ( 
.A(n_4092),
.Y(n_4785)
);

NAND2xp5_ASAP7_75t_L g4786 ( 
.A(n_4372),
.B(n_270),
.Y(n_4786)
);

NAND2xp5_ASAP7_75t_L g4787 ( 
.A(n_4381),
.B(n_270),
.Y(n_4787)
);

NOR2xp33_ASAP7_75t_L g4788 ( 
.A(n_4177),
.B(n_270),
.Y(n_4788)
);

NAND2xp5_ASAP7_75t_L g4789 ( 
.A(n_4394),
.B(n_271),
.Y(n_4789)
);

INVx4_ASAP7_75t_L g4790 ( 
.A(n_4128),
.Y(n_4790)
);

A2O1A1Ixp33_ASAP7_75t_L g4791 ( 
.A1(n_4514),
.A2(n_272),
.B(n_273),
.C(n_271),
.Y(n_4791)
);

NAND2xp5_ASAP7_75t_L g4792 ( 
.A(n_4401),
.B(n_271),
.Y(n_4792)
);

O2A1O1Ixp33_ASAP7_75t_L g4793 ( 
.A1(n_4075),
.A2(n_274),
.B(n_275),
.C(n_272),
.Y(n_4793)
);

AOI21xp5_ASAP7_75t_L g4794 ( 
.A1(n_4272),
.A2(n_274),
.B(n_272),
.Y(n_4794)
);

A2O1A1Ixp33_ASAP7_75t_L g4795 ( 
.A1(n_4205),
.A2(n_275),
.B(n_276),
.C(n_274),
.Y(n_4795)
);

NOR3xp33_ASAP7_75t_L g4796 ( 
.A(n_4207),
.B(n_285),
.C(n_275),
.Y(n_4796)
);

NAND2xp5_ASAP7_75t_L g4797 ( 
.A(n_4404),
.B(n_276),
.Y(n_4797)
);

AOI21xp5_ASAP7_75t_L g4798 ( 
.A1(n_4276),
.A2(n_277),
.B(n_276),
.Y(n_4798)
);

NAND2xp5_ASAP7_75t_L g4799 ( 
.A(n_4406),
.B(n_4409),
.Y(n_4799)
);

INVx2_ASAP7_75t_L g4800 ( 
.A(n_4288),
.Y(n_4800)
);

BUFx4_ASAP7_75t_SL g4801 ( 
.A(n_4035),
.Y(n_4801)
);

NAND2xp5_ASAP7_75t_SL g4802 ( 
.A(n_4060),
.B(n_4582),
.Y(n_4802)
);

NOR2xp33_ASAP7_75t_L g4803 ( 
.A(n_4047),
.B(n_277),
.Y(n_4803)
);

AOI21xp5_ASAP7_75t_L g4804 ( 
.A1(n_4290),
.A2(n_281),
.B(n_278),
.Y(n_4804)
);

AOI21xp5_ASAP7_75t_L g4805 ( 
.A1(n_4292),
.A2(n_281),
.B(n_278),
.Y(n_4805)
);

O2A1O1Ixp33_ASAP7_75t_SL g4806 ( 
.A1(n_4039),
.A2(n_281),
.B(n_282),
.C(n_278),
.Y(n_4806)
);

INVx1_ASAP7_75t_L g4807 ( 
.A(n_4413),
.Y(n_4807)
);

AOI21xp5_ASAP7_75t_L g4808 ( 
.A1(n_4328),
.A2(n_283),
.B(n_282),
.Y(n_4808)
);

AOI21xp5_ASAP7_75t_L g4809 ( 
.A1(n_4366),
.A2(n_283),
.B(n_282),
.Y(n_4809)
);

OAI22xp5_ASAP7_75t_L g4810 ( 
.A1(n_4331),
.A2(n_284),
.B1(n_285),
.B2(n_283),
.Y(n_4810)
);

NAND2xp5_ASAP7_75t_L g4811 ( 
.A(n_4419),
.B(n_284),
.Y(n_4811)
);

NAND2xp5_ASAP7_75t_SL g4812 ( 
.A(n_4582),
.B(n_284),
.Y(n_4812)
);

INVx1_ASAP7_75t_SL g4813 ( 
.A(n_4174),
.Y(n_4813)
);

NAND2xp5_ASAP7_75t_L g4814 ( 
.A(n_4549),
.B(n_286),
.Y(n_4814)
);

NAND2xp5_ASAP7_75t_L g4815 ( 
.A(n_4550),
.B(n_286),
.Y(n_4815)
);

NAND2xp5_ASAP7_75t_L g4816 ( 
.A(n_4444),
.B(n_287),
.Y(n_4816)
);

O2A1O1Ixp33_ASAP7_75t_L g4817 ( 
.A1(n_4136),
.A2(n_288),
.B(n_289),
.C(n_287),
.Y(n_4817)
);

NAND2xp5_ASAP7_75t_L g4818 ( 
.A(n_4436),
.B(n_287),
.Y(n_4818)
);

AOI21xp5_ASAP7_75t_L g4819 ( 
.A1(n_4228),
.A2(n_289),
.B(n_288),
.Y(n_4819)
);

INVx1_ASAP7_75t_L g4820 ( 
.A(n_4465),
.Y(n_4820)
);

OAI22xp5_ASAP7_75t_L g4821 ( 
.A1(n_4309),
.A2(n_291),
.B1(n_292),
.B2(n_290),
.Y(n_4821)
);

HB1xp67_ASAP7_75t_L g4822 ( 
.A(n_4063),
.Y(n_4822)
);

AOI21xp5_ASAP7_75t_L g4823 ( 
.A1(n_4133),
.A2(n_291),
.B(n_290),
.Y(n_4823)
);

AOI21xp5_ASAP7_75t_L g4824 ( 
.A1(n_4191),
.A2(n_291),
.B(n_290),
.Y(n_4824)
);

NAND2xp5_ASAP7_75t_L g4825 ( 
.A(n_4440),
.B(n_292),
.Y(n_4825)
);

AOI21xp5_ASAP7_75t_L g4826 ( 
.A1(n_4218),
.A2(n_293),
.B(n_292),
.Y(n_4826)
);

NAND2xp5_ASAP7_75t_L g4827 ( 
.A(n_4447),
.B(n_293),
.Y(n_4827)
);

AND2x4_ASAP7_75t_L g4828 ( 
.A(n_4166),
.B(n_293),
.Y(n_4828)
);

OAI21xp5_ASAP7_75t_L g4829 ( 
.A1(n_4572),
.A2(n_295),
.B(n_294),
.Y(n_4829)
);

BUFx6f_ASAP7_75t_L g4830 ( 
.A(n_4166),
.Y(n_4830)
);

INVx2_ASAP7_75t_SL g4831 ( 
.A(n_4059),
.Y(n_4831)
);

INVx1_ASAP7_75t_L g4832 ( 
.A(n_4476),
.Y(n_4832)
);

A2O1A1Ixp33_ASAP7_75t_L g4833 ( 
.A1(n_4091),
.A2(n_296),
.B(n_297),
.C(n_294),
.Y(n_4833)
);

AOI21x1_ASAP7_75t_L g4834 ( 
.A1(n_4583),
.A2(n_297),
.B(n_296),
.Y(n_4834)
);

AND2x2_ASAP7_75t_L g4835 ( 
.A(n_4118),
.B(n_296),
.Y(n_4835)
);

BUFx6f_ASAP7_75t_L g4836 ( 
.A(n_4184),
.Y(n_4836)
);

A2O1A1Ixp33_ASAP7_75t_L g4837 ( 
.A1(n_4539),
.A2(n_298),
.B(n_300),
.C(n_297),
.Y(n_4837)
);

NOR2x1_ASAP7_75t_L g4838 ( 
.A(n_4229),
.B(n_298),
.Y(n_4838)
);

AOI21xp33_ASAP7_75t_L g4839 ( 
.A1(n_4562),
.A2(n_300),
.B(n_298),
.Y(n_4839)
);

INVx4_ASAP7_75t_L g4840 ( 
.A(n_4128),
.Y(n_4840)
);

INVx2_ASAP7_75t_SL g4841 ( 
.A(n_4074),
.Y(n_4841)
);

AOI21xp5_ASAP7_75t_L g4842 ( 
.A1(n_4463),
.A2(n_302),
.B(n_301),
.Y(n_4842)
);

AOI21xp5_ASAP7_75t_L g4843 ( 
.A1(n_4463),
.A2(n_302),
.B(n_301),
.Y(n_4843)
);

AOI21xp5_ASAP7_75t_L g4844 ( 
.A1(n_4417),
.A2(n_302),
.B(n_301),
.Y(n_4844)
);

A2O1A1Ixp33_ASAP7_75t_L g4845 ( 
.A1(n_4534),
.A2(n_4598),
.B(n_4593),
.C(n_4556),
.Y(n_4845)
);

O2A1O1Ixp33_ASAP7_75t_L g4846 ( 
.A1(n_4141),
.A2(n_304),
.B(n_305),
.C(n_303),
.Y(n_4846)
);

NAND2x1_ASAP7_75t_L g4847 ( 
.A(n_4294),
.B(n_303),
.Y(n_4847)
);

O2A1O1Ixp33_ASAP7_75t_SL g4848 ( 
.A1(n_4041),
.A2(n_304),
.B(n_305),
.C(n_303),
.Y(n_4848)
);

INVx1_ASAP7_75t_L g4849 ( 
.A(n_4451),
.Y(n_4849)
);

NAND3xp33_ASAP7_75t_L g4850 ( 
.A(n_4416),
.B(n_306),
.C(n_304),
.Y(n_4850)
);

AND2x2_ASAP7_75t_L g4851 ( 
.A(n_4456),
.B(n_307),
.Y(n_4851)
);

INVx2_ASAP7_75t_L g4852 ( 
.A(n_4308),
.Y(n_4852)
);

INVx1_ASAP7_75t_L g4853 ( 
.A(n_4183),
.Y(n_4853)
);

NAND2xp5_ASAP7_75t_L g4854 ( 
.A(n_4521),
.B(n_307),
.Y(n_4854)
);

AOI22xp5_ASAP7_75t_L g4855 ( 
.A1(n_4040),
.A2(n_1064),
.B1(n_1068),
.B2(n_1063),
.Y(n_4855)
);

OAI22xp5_ASAP7_75t_L g4856 ( 
.A1(n_4230),
.A2(n_4123),
.B1(n_4132),
.B2(n_4578),
.Y(n_4856)
);

INVx1_ASAP7_75t_L g4857 ( 
.A(n_4284),
.Y(n_4857)
);

OAI21x1_ASAP7_75t_L g4858 ( 
.A1(n_4503),
.A2(n_309),
.B(n_308),
.Y(n_4858)
);

NOR3xp33_ASAP7_75t_L g4859 ( 
.A(n_4180),
.B(n_316),
.C(n_308),
.Y(n_4859)
);

AOI21xp5_ASAP7_75t_L g4860 ( 
.A1(n_4298),
.A2(n_309),
.B(n_308),
.Y(n_4860)
);

INVx2_ASAP7_75t_L g4861 ( 
.A(n_4335),
.Y(n_4861)
);

NAND2xp5_ASAP7_75t_L g4862 ( 
.A(n_4499),
.B(n_309),
.Y(n_4862)
);

NAND2xp5_ASAP7_75t_L g4863 ( 
.A(n_4511),
.B(n_310),
.Y(n_4863)
);

AOI21xp5_ASAP7_75t_L g4864 ( 
.A1(n_4408),
.A2(n_311),
.B(n_310),
.Y(n_4864)
);

INVx2_ASAP7_75t_L g4865 ( 
.A(n_4340),
.Y(n_4865)
);

NAND2xp5_ASAP7_75t_L g4866 ( 
.A(n_4520),
.B(n_310),
.Y(n_4866)
);

BUFx2_ASAP7_75t_L g4867 ( 
.A(n_4219),
.Y(n_4867)
);

AOI22xp33_ASAP7_75t_L g4868 ( 
.A1(n_4553),
.A2(n_312),
.B1(n_313),
.B2(n_311),
.Y(n_4868)
);

NAND3xp33_ASAP7_75t_L g4869 ( 
.A(n_4474),
.B(n_312),
.C(n_311),
.Y(n_4869)
);

OAI21xp5_ASAP7_75t_L g4870 ( 
.A1(n_4599),
.A2(n_313),
.B(n_312),
.Y(n_4870)
);

NAND3xp33_ASAP7_75t_SL g4871 ( 
.A(n_4286),
.B(n_3),
.C(n_4),
.Y(n_4871)
);

AOI21xp5_ASAP7_75t_L g4872 ( 
.A1(n_4571),
.A2(n_314),
.B(n_313),
.Y(n_4872)
);

NOR2xp33_ASAP7_75t_L g4873 ( 
.A(n_4454),
.B(n_314),
.Y(n_4873)
);

AOI22xp5_ASAP7_75t_L g4874 ( 
.A1(n_4462),
.A2(n_4070),
.B1(n_4100),
.B2(n_4523),
.Y(n_4874)
);

AOI22xp5_ASAP7_75t_L g4875 ( 
.A1(n_4524),
.A2(n_1055),
.B1(n_1056),
.B2(n_1054),
.Y(n_4875)
);

CKINVDCx10_ASAP7_75t_R g4876 ( 
.A(n_4235),
.Y(n_4876)
);

AOI21xp5_ASAP7_75t_L g4877 ( 
.A1(n_4407),
.A2(n_4519),
.B(n_4491),
.Y(n_4877)
);

AOI21xp5_ASAP7_75t_L g4878 ( 
.A1(n_4153),
.A2(n_316),
.B(n_315),
.Y(n_4878)
);

AOI22xp5_ASAP7_75t_L g4879 ( 
.A1(n_4139),
.A2(n_1056),
.B1(n_1057),
.B2(n_1055),
.Y(n_4879)
);

NOR2xp33_ASAP7_75t_L g4880 ( 
.A(n_4119),
.B(n_315),
.Y(n_4880)
);

INVx11_ASAP7_75t_L g4881 ( 
.A(n_4065),
.Y(n_4881)
);

AOI21xp5_ASAP7_75t_L g4882 ( 
.A1(n_4500),
.A2(n_317),
.B(n_316),
.Y(n_4882)
);

O2A1O1Ixp5_ASAP7_75t_L g4883 ( 
.A1(n_4596),
.A2(n_318),
.B(n_319),
.C(n_317),
.Y(n_4883)
);

INVx2_ASAP7_75t_L g4884 ( 
.A(n_4344),
.Y(n_4884)
);

NAND2xp5_ASAP7_75t_SL g4885 ( 
.A(n_4582),
.B(n_317),
.Y(n_4885)
);

NOR2xp33_ASAP7_75t_L g4886 ( 
.A(n_4159),
.B(n_318),
.Y(n_4886)
);

NOR2xp33_ASAP7_75t_L g4887 ( 
.A(n_4072),
.B(n_318),
.Y(n_4887)
);

NOR2xp33_ASAP7_75t_L g4888 ( 
.A(n_4087),
.B(n_319),
.Y(n_4888)
);

INVx2_ASAP7_75t_L g4889 ( 
.A(n_4347),
.Y(n_4889)
);

AOI21xp5_ASAP7_75t_L g4890 ( 
.A1(n_4071),
.A2(n_320),
.B(n_319),
.Y(n_4890)
);

INVx4_ASAP7_75t_L g4891 ( 
.A(n_4231),
.Y(n_4891)
);

AOI21xp5_ASAP7_75t_L g4892 ( 
.A1(n_4086),
.A2(n_321),
.B(n_320),
.Y(n_4892)
);

AOI21xp5_ASAP7_75t_L g4893 ( 
.A1(n_4097),
.A2(n_322),
.B(n_320),
.Y(n_4893)
);

NAND2x1p5_ASAP7_75t_L g4894 ( 
.A(n_4102),
.B(n_322),
.Y(n_4894)
);

NAND2xp5_ASAP7_75t_L g4895 ( 
.A(n_4525),
.B(n_322),
.Y(n_4895)
);

NAND2xp5_ASAP7_75t_L g4896 ( 
.A(n_4526),
.B(n_323),
.Y(n_4896)
);

AOI22xp33_ASAP7_75t_L g4897 ( 
.A1(n_4576),
.A2(n_324),
.B1(n_325),
.B2(n_323),
.Y(n_4897)
);

O2A1O1Ixp33_ASAP7_75t_L g4898 ( 
.A1(n_4098),
.A2(n_324),
.B(n_325),
.C(n_323),
.Y(n_4898)
);

INVx1_ASAP7_75t_L g4899 ( 
.A(n_4358),
.Y(n_4899)
);

NOR2xp33_ASAP7_75t_SL g4900 ( 
.A(n_4152),
.B(n_4258),
.Y(n_4900)
);

NAND2xp5_ASAP7_75t_L g4901 ( 
.A(n_4528),
.B(n_324),
.Y(n_4901)
);

AOI21xp5_ASAP7_75t_L g4902 ( 
.A1(n_4108),
.A2(n_4142),
.B(n_4116),
.Y(n_4902)
);

AOI21xp5_ASAP7_75t_L g4903 ( 
.A1(n_4143),
.A2(n_326),
.B(n_325),
.Y(n_4903)
);

A2O1A1Ixp33_ASAP7_75t_L g4904 ( 
.A1(n_4200),
.A2(n_327),
.B(n_329),
.C(n_326),
.Y(n_4904)
);

NOR3xp33_ASAP7_75t_L g4905 ( 
.A(n_4300),
.B(n_338),
.C(n_330),
.Y(n_4905)
);

AO21x1_ASAP7_75t_L g4906 ( 
.A1(n_4513),
.A2(n_331),
.B(n_327),
.Y(n_4906)
);

NOR2xp33_ASAP7_75t_L g4907 ( 
.A(n_4138),
.B(n_331),
.Y(n_4907)
);

AOI221xp5_ASAP7_75t_L g4908 ( 
.A1(n_4568),
.A2(n_333),
.B1(n_334),
.B2(n_332),
.C(n_331),
.Y(n_4908)
);

INVx1_ASAP7_75t_L g4909 ( 
.A(n_4378),
.Y(n_4909)
);

BUFx3_ASAP7_75t_L g4910 ( 
.A(n_4293),
.Y(n_4910)
);

NAND2xp5_ASAP7_75t_L g4911 ( 
.A(n_4535),
.B(n_332),
.Y(n_4911)
);

O2A1O1Ixp5_ASAP7_75t_L g4912 ( 
.A1(n_4575),
.A2(n_333),
.B(n_334),
.C(n_332),
.Y(n_4912)
);

NAND2x1p5_ASAP7_75t_L g4913 ( 
.A(n_4229),
.B(n_335),
.Y(n_4913)
);

OR2x6_ASAP7_75t_L g4914 ( 
.A(n_4214),
.B(n_335),
.Y(n_4914)
);

NOR2xp33_ASAP7_75t_L g4915 ( 
.A(n_4036),
.B(n_335),
.Y(n_4915)
);

HB1xp67_ASAP7_75t_L g4916 ( 
.A(n_4289),
.Y(n_4916)
);

NOR2xp33_ASAP7_75t_L g4917 ( 
.A(n_4069),
.B(n_336),
.Y(n_4917)
);

BUFx2_ASAP7_75t_SL g4918 ( 
.A(n_4083),
.Y(n_4918)
);

BUFx12f_ASAP7_75t_L g4919 ( 
.A(n_4176),
.Y(n_4919)
);

NOR2xp33_ASAP7_75t_L g4920 ( 
.A(n_4117),
.B(n_336),
.Y(n_4920)
);

NAND2xp5_ASAP7_75t_L g4921 ( 
.A(n_4541),
.B(n_337),
.Y(n_4921)
);

OAI22xp5_ASAP7_75t_L g4922 ( 
.A1(n_4578),
.A2(n_338),
.B1(n_339),
.B2(n_337),
.Y(n_4922)
);

AOI22xp5_ASAP7_75t_L g4923 ( 
.A1(n_4114),
.A2(n_1068),
.B1(n_1069),
.B2(n_1064),
.Y(n_4923)
);

NOR2xp67_ASAP7_75t_L g4924 ( 
.A(n_4211),
.B(n_4242),
.Y(n_4924)
);

BUFx4f_ASAP7_75t_L g4925 ( 
.A(n_4256),
.Y(n_4925)
);

NAND2xp5_ASAP7_75t_L g4926 ( 
.A(n_4193),
.B(n_337),
.Y(n_4926)
);

AOI21xp5_ASAP7_75t_L g4927 ( 
.A1(n_4167),
.A2(n_340),
.B(n_339),
.Y(n_4927)
);

AOI21xp5_ASAP7_75t_L g4928 ( 
.A1(n_4168),
.A2(n_340),
.B(n_339),
.Y(n_4928)
);

AOI22xp5_ASAP7_75t_L g4929 ( 
.A1(n_4172),
.A2(n_1072),
.B1(n_1071),
.B2(n_342),
.Y(n_4929)
);

NAND2xp5_ASAP7_75t_L g4930 ( 
.A(n_4498),
.B(n_341),
.Y(n_4930)
);

INVx3_ASAP7_75t_L g4931 ( 
.A(n_4245),
.Y(n_4931)
);

INVx1_ASAP7_75t_L g4932 ( 
.A(n_4380),
.Y(n_4932)
);

OAI22xp5_ASAP7_75t_L g4933 ( 
.A1(n_4113),
.A2(n_342),
.B1(n_343),
.B2(n_341),
.Y(n_4933)
);

AND2x2_ASAP7_75t_L g4934 ( 
.A(n_4053),
.B(n_341),
.Y(n_4934)
);

NAND2xp5_ASAP7_75t_L g4935 ( 
.A(n_4554),
.B(n_343),
.Y(n_4935)
);

AOI21xp33_ASAP7_75t_L g4936 ( 
.A1(n_4346),
.A2(n_4373),
.B(n_4538),
.Y(n_4936)
);

OAI22xp5_ASAP7_75t_L g4937 ( 
.A1(n_4585),
.A2(n_345),
.B1(n_346),
.B2(n_343),
.Y(n_4937)
);

AOI22xp33_ASAP7_75t_L g4938 ( 
.A1(n_4552),
.A2(n_346),
.B1(n_347),
.B2(n_345),
.Y(n_4938)
);

INVx2_ASAP7_75t_L g4939 ( 
.A(n_4405),
.Y(n_4939)
);

INVx2_ASAP7_75t_L g4940 ( 
.A(n_4438),
.Y(n_4940)
);

OAI21xp5_ASAP7_75t_L g4941 ( 
.A1(n_4580),
.A2(n_346),
.B(n_345),
.Y(n_4941)
);

OAI22xp5_ASAP7_75t_L g4942 ( 
.A1(n_4560),
.A2(n_348),
.B1(n_349),
.B2(n_347),
.Y(n_4942)
);

NAND2xp5_ASAP7_75t_L g4943 ( 
.A(n_4561),
.B(n_347),
.Y(n_4943)
);

BUFx6f_ASAP7_75t_L g4944 ( 
.A(n_4184),
.Y(n_4944)
);

NAND2xp5_ASAP7_75t_L g4945 ( 
.A(n_4563),
.B(n_348),
.Y(n_4945)
);

BUFx6f_ASAP7_75t_L g4946 ( 
.A(n_4184),
.Y(n_4946)
);

AND2x4_ASAP7_75t_L g4947 ( 
.A(n_4294),
.B(n_348),
.Y(n_4947)
);

NAND3xp33_ASAP7_75t_SL g4948 ( 
.A(n_4295),
.B(n_4),
.C(n_5),
.Y(n_4948)
);

INVx2_ASAP7_75t_L g4949 ( 
.A(n_4442),
.Y(n_4949)
);

INVx1_ASAP7_75t_L g4950 ( 
.A(n_4458),
.Y(n_4950)
);

OAI21xp5_ASAP7_75t_L g4951 ( 
.A1(n_4532),
.A2(n_350),
.B(n_349),
.Y(n_4951)
);

NAND2xp5_ASAP7_75t_SL g4952 ( 
.A(n_4245),
.B(n_349),
.Y(n_4952)
);

OAI22xp5_ASAP7_75t_L g4953 ( 
.A1(n_4154),
.A2(n_352),
.B1(n_353),
.B2(n_351),
.Y(n_4953)
);

AOI22xp5_ASAP7_75t_L g4954 ( 
.A1(n_4479),
.A2(n_1062),
.B1(n_1063),
.B2(n_1061),
.Y(n_4954)
);

NAND2xp5_ASAP7_75t_L g4955 ( 
.A(n_4566),
.B(n_351),
.Y(n_4955)
);

NAND2xp5_ASAP7_75t_SL g4956 ( 
.A(n_4245),
.B(n_351),
.Y(n_4956)
);

AOI21xp5_ASAP7_75t_L g4957 ( 
.A1(n_4179),
.A2(n_354),
.B(n_352),
.Y(n_4957)
);

INVx1_ASAP7_75t_L g4958 ( 
.A(n_4186),
.Y(n_4958)
);

O2A1O1Ixp33_ASAP7_75t_L g4959 ( 
.A1(n_4099),
.A2(n_354),
.B(n_355),
.C(n_352),
.Y(n_4959)
);

NAND2xp5_ASAP7_75t_SL g4960 ( 
.A(n_4259),
.B(n_355),
.Y(n_4960)
);

NAND2xp5_ASAP7_75t_SL g4961 ( 
.A(n_4259),
.B(n_355),
.Y(n_4961)
);

NOR2xp33_ASAP7_75t_L g4962 ( 
.A(n_4164),
.B(n_356),
.Y(n_4962)
);

AOI21xp5_ASAP7_75t_L g4963 ( 
.A1(n_4423),
.A2(n_357),
.B(n_356),
.Y(n_4963)
);

NAND2xp5_ASAP7_75t_L g4964 ( 
.A(n_4573),
.B(n_356),
.Y(n_4964)
);

BUFx6f_ASAP7_75t_L g4965 ( 
.A(n_4196),
.Y(n_4965)
);

AOI21xp5_ASAP7_75t_L g4966 ( 
.A1(n_4423),
.A2(n_358),
.B(n_357),
.Y(n_4966)
);

NOR2xp33_ASAP7_75t_L g4967 ( 
.A(n_4171),
.B(n_357),
.Y(n_4967)
);

AOI21xp5_ASAP7_75t_L g4968 ( 
.A1(n_4399),
.A2(n_359),
.B(n_358),
.Y(n_4968)
);

NAND2xp5_ASAP7_75t_SL g4969 ( 
.A(n_4259),
.B(n_359),
.Y(n_4969)
);

O2A1O1Ixp33_ASAP7_75t_SL g4970 ( 
.A1(n_4545),
.A2(n_4536),
.B(n_4592),
.C(n_4587),
.Y(n_4970)
);

AOI21xp5_ASAP7_75t_L g4971 ( 
.A1(n_4595),
.A2(n_360),
.B(n_359),
.Y(n_4971)
);

AND2x2_ASAP7_75t_L g4972 ( 
.A(n_4208),
.B(n_360),
.Y(n_4972)
);

NAND2xp5_ASAP7_75t_SL g4973 ( 
.A(n_4322),
.B(n_360),
.Y(n_4973)
);

NOR2xp33_ASAP7_75t_L g4974 ( 
.A(n_4273),
.B(n_361),
.Y(n_4974)
);

O2A1O1Ixp33_ASAP7_75t_L g4975 ( 
.A1(n_4507),
.A2(n_362),
.B(n_363),
.C(n_361),
.Y(n_4975)
);

CKINVDCx8_ASAP7_75t_R g4976 ( 
.A(n_4190),
.Y(n_4976)
);

NAND2xp5_ASAP7_75t_L g4977 ( 
.A(n_4586),
.B(n_361),
.Y(n_4977)
);

AOI21xp5_ASAP7_75t_L g4978 ( 
.A1(n_4473),
.A2(n_363),
.B(n_362),
.Y(n_4978)
);

INVx1_ASAP7_75t_L g4979 ( 
.A(n_4210),
.Y(n_4979)
);

INVx3_ASAP7_75t_L g4980 ( 
.A(n_4322),
.Y(n_4980)
);

NAND2xp5_ASAP7_75t_L g4981 ( 
.A(n_4588),
.B(n_363),
.Y(n_4981)
);

NAND2xp5_ASAP7_75t_SL g4982 ( 
.A(n_4322),
.B(n_364),
.Y(n_4982)
);

NOR2xp33_ASAP7_75t_SL g4983 ( 
.A(n_4233),
.B(n_1057),
.Y(n_4983)
);

NAND2xp5_ASAP7_75t_L g4984 ( 
.A(n_4589),
.B(n_364),
.Y(n_4984)
);

INVxp67_ASAP7_75t_L g4985 ( 
.A(n_4246),
.Y(n_4985)
);

NAND2xp5_ASAP7_75t_L g4986 ( 
.A(n_4584),
.B(n_4594),
.Y(n_4986)
);

AOI21xp5_ASAP7_75t_L g4987 ( 
.A1(n_4477),
.A2(n_365),
.B(n_364),
.Y(n_4987)
);

AOI22xp5_ASAP7_75t_L g4988 ( 
.A1(n_4495),
.A2(n_1058),
.B1(n_1060),
.B2(n_1057),
.Y(n_4988)
);

AOI21xp5_ASAP7_75t_L g4989 ( 
.A1(n_4477),
.A2(n_366),
.B(n_365),
.Y(n_4989)
);

OR2x2_ASAP7_75t_L g4990 ( 
.A(n_4199),
.B(n_365),
.Y(n_4990)
);

AOI21xp5_ASAP7_75t_L g4991 ( 
.A1(n_4494),
.A2(n_367),
.B(n_366),
.Y(n_4991)
);

NAND2xp5_ASAP7_75t_L g4992 ( 
.A(n_4496),
.B(n_367),
.Y(n_4992)
);

OR2x2_ASAP7_75t_L g4993 ( 
.A(n_4204),
.B(n_367),
.Y(n_4993)
);

INVx5_ASAP7_75t_L g4994 ( 
.A(n_4385),
.Y(n_4994)
);

NAND2x1p5_ASAP7_75t_L g4995 ( 
.A(n_4253),
.B(n_368),
.Y(n_4995)
);

NOR2xp33_ASAP7_75t_L g4996 ( 
.A(n_4368),
.B(n_368),
.Y(n_4996)
);

BUFx2_ASAP7_75t_L g4997 ( 
.A(n_4250),
.Y(n_4997)
);

NAND2xp5_ASAP7_75t_L g4998 ( 
.A(n_4398),
.B(n_368),
.Y(n_4998)
);

INVx3_ASAP7_75t_L g4999 ( 
.A(n_4364),
.Y(n_4999)
);

NAND2xp5_ASAP7_75t_SL g5000 ( 
.A(n_4569),
.B(n_369),
.Y(n_5000)
);

OAI21xp33_ASAP7_75t_SL g5001 ( 
.A1(n_4329),
.A2(n_371),
.B(n_369),
.Y(n_5001)
);

AOI21xp5_ASAP7_75t_L g5002 ( 
.A1(n_4494),
.A2(n_370),
.B(n_369),
.Y(n_5002)
);

AOI21xp5_ASAP7_75t_L g5003 ( 
.A1(n_4509),
.A2(n_371),
.B(n_370),
.Y(n_5003)
);

INVx1_ASAP7_75t_SL g5004 ( 
.A(n_4277),
.Y(n_5004)
);

AO21x1_ASAP7_75t_L g5005 ( 
.A1(n_4569),
.A2(n_372),
.B(n_371),
.Y(n_5005)
);

A2O1A1Ixp33_ASAP7_75t_L g5006 ( 
.A1(n_4305),
.A2(n_373),
.B(n_374),
.C(n_372),
.Y(n_5006)
);

AOI21x1_ASAP7_75t_L g5007 ( 
.A1(n_4453),
.A2(n_374),
.B(n_373),
.Y(n_5007)
);

NOR3xp33_ASAP7_75t_L g5008 ( 
.A(n_4084),
.B(n_383),
.C(n_375),
.Y(n_5008)
);

OAI22xp5_ASAP7_75t_L g5009 ( 
.A1(n_4327),
.A2(n_375),
.B1(n_376),
.B2(n_374),
.Y(n_5009)
);

OAI22xp5_ASAP7_75t_L g5010 ( 
.A1(n_4387),
.A2(n_376),
.B1(n_377),
.B2(n_375),
.Y(n_5010)
);

NAND2xp5_ASAP7_75t_L g5011 ( 
.A(n_4439),
.B(n_377),
.Y(n_5011)
);

NAND2xp5_ASAP7_75t_L g5012 ( 
.A(n_4484),
.B(n_377),
.Y(n_5012)
);

OAI22xp5_ASAP7_75t_L g5013 ( 
.A1(n_4559),
.A2(n_379),
.B1(n_380),
.B2(n_378),
.Y(n_5013)
);

HB1xp67_ASAP7_75t_L g5014 ( 
.A(n_4051),
.Y(n_5014)
);

NAND2xp5_ASAP7_75t_SL g5015 ( 
.A(n_4264),
.B(n_378),
.Y(n_5015)
);

NAND2xp5_ASAP7_75t_L g5016 ( 
.A(n_4506),
.B(n_379),
.Y(n_5016)
);

BUFx3_ASAP7_75t_L g5017 ( 
.A(n_4262),
.Y(n_5017)
);

OAI21xp5_ASAP7_75t_L g5018 ( 
.A1(n_4548),
.A2(n_380),
.B(n_379),
.Y(n_5018)
);

INVx1_ASAP7_75t_SL g5019 ( 
.A(n_4209),
.Y(n_5019)
);

AO32x2_ASAP7_75t_L g5020 ( 
.A1(n_4505),
.A2(n_398),
.A3(n_406),
.B1(n_390),
.B2(n_382),
.Y(n_5020)
);

NAND2xp5_ASAP7_75t_SL g5021 ( 
.A(n_4216),
.B(n_381),
.Y(n_5021)
);

NAND2xp5_ASAP7_75t_L g5022 ( 
.A(n_4510),
.B(n_381),
.Y(n_5022)
);

BUFx2_ASAP7_75t_L g5023 ( 
.A(n_4094),
.Y(n_5023)
);

AOI21xp5_ASAP7_75t_L g5024 ( 
.A1(n_4509),
.A2(n_382),
.B(n_381),
.Y(n_5024)
);

INVx1_ASAP7_75t_L g5025 ( 
.A(n_4376),
.Y(n_5025)
);

OAI21x1_ASAP7_75t_L g5026 ( 
.A1(n_4504),
.A2(n_383),
.B(n_382),
.Y(n_5026)
);

OAI21xp5_ASAP7_75t_L g5027 ( 
.A1(n_4109),
.A2(n_384),
.B(n_383),
.Y(n_5027)
);

INVx5_ASAP7_75t_L g5028 ( 
.A(n_4385),
.Y(n_5028)
);

AOI21x1_ASAP7_75t_L g5029 ( 
.A1(n_4453),
.A2(n_385),
.B(n_384),
.Y(n_5029)
);

AND2x2_ASAP7_75t_L g5030 ( 
.A(n_4339),
.B(n_385),
.Y(n_5030)
);

OAI22xp5_ASAP7_75t_L g5031 ( 
.A1(n_4202),
.A2(n_386),
.B1(n_387),
.B2(n_385),
.Y(n_5031)
);

O2A1O1Ixp33_ASAP7_75t_L g5032 ( 
.A1(n_4237),
.A2(n_387),
.B(n_388),
.C(n_386),
.Y(n_5032)
);

NOR2xp33_ASAP7_75t_SL g5033 ( 
.A(n_4234),
.B(n_1069),
.Y(n_5033)
);

AND2x2_ASAP7_75t_L g5034 ( 
.A(n_4334),
.B(n_386),
.Y(n_5034)
);

A2O1A1Ixp33_ASAP7_75t_L g5035 ( 
.A1(n_4565),
.A2(n_388),
.B(n_389),
.C(n_387),
.Y(n_5035)
);

NAND2xp5_ASAP7_75t_L g5036 ( 
.A(n_4522),
.B(n_389),
.Y(n_5036)
);

AOI21xp5_ASAP7_75t_L g5037 ( 
.A1(n_4527),
.A2(n_4543),
.B(n_4531),
.Y(n_5037)
);

AOI21xp5_ASAP7_75t_L g5038 ( 
.A1(n_4557),
.A2(n_4597),
.B(n_4558),
.Y(n_5038)
);

NOR2xp33_ASAP7_75t_L g5039 ( 
.A(n_4368),
.B(n_4455),
.Y(n_5039)
);

AOI22xp33_ASAP7_75t_L g5040 ( 
.A1(n_4547),
.A2(n_390),
.B1(n_391),
.B2(n_389),
.Y(n_5040)
);

NOR2xp33_ASAP7_75t_L g5041 ( 
.A(n_4137),
.B(n_391),
.Y(n_5041)
);

OAI22xp5_ASAP7_75t_L g5042 ( 
.A1(n_4325),
.A2(n_392),
.B1(n_393),
.B2(n_391),
.Y(n_5042)
);

INVx2_ASAP7_75t_L g5043 ( 
.A(n_4396),
.Y(n_5043)
);

NAND2xp5_ASAP7_75t_L g5044 ( 
.A(n_4377),
.B(n_393),
.Y(n_5044)
);

AND2x2_ASAP7_75t_L g5045 ( 
.A(n_4382),
.B(n_4418),
.Y(n_5045)
);

OA22x2_ASAP7_75t_L g5046 ( 
.A1(n_4281),
.A2(n_395),
.B1(n_396),
.B2(n_394),
.Y(n_5046)
);

NAND3x1_ASAP7_75t_L g5047 ( 
.A(n_4225),
.B(n_397),
.C(n_396),
.Y(n_5047)
);

NOR2xp33_ASAP7_75t_L g5048 ( 
.A(n_4287),
.B(n_397),
.Y(n_5048)
);

NAND2xp5_ASAP7_75t_L g5049 ( 
.A(n_4469),
.B(n_397),
.Y(n_5049)
);

NOR2xp33_ASAP7_75t_L g5050 ( 
.A(n_4239),
.B(n_398),
.Y(n_5050)
);

AOI21xp5_ASAP7_75t_L g5051 ( 
.A1(n_4314),
.A2(n_400),
.B(n_399),
.Y(n_5051)
);

NAND2xp5_ASAP7_75t_L g5052 ( 
.A(n_4135),
.B(n_400),
.Y(n_5052)
);

AOI21xp5_ASAP7_75t_L g5053 ( 
.A1(n_4464),
.A2(n_401),
.B(n_400),
.Y(n_5053)
);

NOR2xp33_ASAP7_75t_L g5054 ( 
.A(n_4426),
.B(n_4127),
.Y(n_5054)
);

NOR2xp33_ASAP7_75t_L g5055 ( 
.A(n_4299),
.B(n_401),
.Y(n_5055)
);

OAI22xp5_ASAP7_75t_L g5056 ( 
.A1(n_4464),
.A2(n_402),
.B1(n_403),
.B2(n_401),
.Y(n_5056)
);

AO21x1_ASAP7_75t_L g5057 ( 
.A1(n_4383),
.A2(n_403),
.B(n_402),
.Y(n_5057)
);

AOI21xp5_ASAP7_75t_L g5058 ( 
.A1(n_4321),
.A2(n_404),
.B(n_402),
.Y(n_5058)
);

NAND2xp5_ASAP7_75t_L g5059 ( 
.A(n_4125),
.B(n_404),
.Y(n_5059)
);

NAND2xp5_ASAP7_75t_L g5060 ( 
.A(n_4104),
.B(n_405),
.Y(n_5060)
);

BUFx6f_ASAP7_75t_L g5061 ( 
.A(n_4196),
.Y(n_5061)
);

AOI21xp5_ASAP7_75t_L g5062 ( 
.A1(n_4336),
.A2(n_406),
.B(n_405),
.Y(n_5062)
);

INVx2_ASAP7_75t_L g5063 ( 
.A(n_4371),
.Y(n_5063)
);

INVx2_ASAP7_75t_SL g5064 ( 
.A(n_4235),
.Y(n_5064)
);

AOI21xp5_ASAP7_75t_L g5065 ( 
.A1(n_4343),
.A2(n_407),
.B(n_406),
.Y(n_5065)
);

NAND2xp5_ASAP7_75t_L g5066 ( 
.A(n_4112),
.B(n_407),
.Y(n_5066)
);

NAND2xp5_ASAP7_75t_SL g5067 ( 
.A(n_4402),
.B(n_408),
.Y(n_5067)
);

INVx1_ASAP7_75t_SL g5068 ( 
.A(n_4215),
.Y(n_5068)
);

AOI22xp33_ASAP7_75t_SL g5069 ( 
.A1(n_4140),
.A2(n_409),
.B1(n_410),
.B2(n_408),
.Y(n_5069)
);

INVx2_ASAP7_75t_L g5070 ( 
.A(n_4348),
.Y(n_5070)
);

INVx3_ASAP7_75t_L g5071 ( 
.A(n_4281),
.Y(n_5071)
);

NAND2xp5_ASAP7_75t_SL g5072 ( 
.A(n_4445),
.B(n_409),
.Y(n_5072)
);

A2O1A1Ixp33_ASAP7_75t_L g5073 ( 
.A1(n_4490),
.A2(n_410),
.B(n_411),
.C(n_409),
.Y(n_5073)
);

NAND2xp5_ASAP7_75t_L g5074 ( 
.A(n_4275),
.B(n_411),
.Y(n_5074)
);

O2A1O1Ixp33_ASAP7_75t_L g5075 ( 
.A1(n_4467),
.A2(n_4475),
.B(n_4480),
.C(n_4470),
.Y(n_5075)
);

INVx3_ASAP7_75t_L g5076 ( 
.A(n_4247),
.Y(n_5076)
);

OAI21x1_ASAP7_75t_L g5077 ( 
.A1(n_4643),
.A2(n_4042),
.B(n_4357),
.Y(n_5077)
);

NAND2xp5_ASAP7_75t_L g5078 ( 
.A(n_4857),
.B(n_4481),
.Y(n_5078)
);

NAND2xp5_ASAP7_75t_SL g5079 ( 
.A(n_4630),
.B(n_4271),
.Y(n_5079)
);

AND2x2_ASAP7_75t_L g5080 ( 
.A(n_4658),
.B(n_4638),
.Y(n_5080)
);

INVx2_ASAP7_75t_L g5081 ( 
.A(n_4600),
.Y(n_5081)
);

A2O1A1Ixp33_ASAP7_75t_L g5082 ( 
.A1(n_4687),
.A2(n_4512),
.B(n_4362),
.C(n_4232),
.Y(n_5082)
);

OAI22xp5_ASAP7_75t_L g5083 ( 
.A1(n_4914),
.A2(n_4663),
.B1(n_4677),
.B2(n_5069),
.Y(n_5083)
);

AOI21xp5_ASAP7_75t_L g5084 ( 
.A1(n_4616),
.A2(n_4614),
.B(n_4633),
.Y(n_5084)
);

OAI21xp5_ASAP7_75t_L g5085 ( 
.A1(n_5001),
.A2(n_4486),
.B(n_4482),
.Y(n_5085)
);

NOR2x1_ASAP7_75t_L g5086 ( 
.A(n_4891),
.B(n_4364),
.Y(n_5086)
);

INVx1_ASAP7_75t_L g5087 ( 
.A(n_4609),
.Y(n_5087)
);

NOR2x1_ASAP7_75t_L g5088 ( 
.A(n_4891),
.B(n_4790),
.Y(n_5088)
);

AOI21xp5_ASAP7_75t_L g5089 ( 
.A1(n_4619),
.A2(n_4267),
.B(n_4222),
.Y(n_5089)
);

BUFx12f_ASAP7_75t_L g5090 ( 
.A(n_4628),
.Y(n_5090)
);

AOI21xp5_ASAP7_75t_L g5091 ( 
.A1(n_4605),
.A2(n_4267),
.B(n_4222),
.Y(n_5091)
);

AND2x2_ASAP7_75t_L g5092 ( 
.A(n_5045),
.B(n_4351),
.Y(n_5092)
);

OAI21xp5_ASAP7_75t_L g5093 ( 
.A1(n_4859),
.A2(n_4492),
.B(n_4488),
.Y(n_5093)
);

INVxp67_ASAP7_75t_L g5094 ( 
.A(n_4918),
.Y(n_5094)
);

AOI21xp5_ASAP7_75t_L g5095 ( 
.A1(n_4639),
.A2(n_4359),
.B(n_4261),
.Y(n_5095)
);

AOI21xp5_ASAP7_75t_L g5096 ( 
.A1(n_4877),
.A2(n_4261),
.B(n_4196),
.Y(n_5096)
);

OAI21xp5_ASAP7_75t_L g5097 ( 
.A1(n_5008),
.A2(n_4537),
.B(n_4530),
.Y(n_5097)
);

INVx5_ASAP7_75t_L g5098 ( 
.A(n_4613),
.Y(n_5098)
);

AOI21xp5_ASAP7_75t_L g5099 ( 
.A1(n_4618),
.A2(n_4266),
.B(n_4261),
.Y(n_5099)
);

NAND2xp5_ASAP7_75t_SL g5100 ( 
.A(n_4790),
.B(n_4266),
.Y(n_5100)
);

AND2x2_ASAP7_75t_L g5101 ( 
.A(n_4979),
.B(n_4301),
.Y(n_5101)
);

INVx3_ASAP7_75t_L g5102 ( 
.A(n_4925),
.Y(n_5102)
);

BUFx6f_ASAP7_75t_L g5103 ( 
.A(n_4626),
.Y(n_5103)
);

OAI21x1_ASAP7_75t_L g5104 ( 
.A1(n_4705),
.A2(n_4443),
.B(n_4400),
.Y(n_5104)
);

INVx3_ASAP7_75t_L g5105 ( 
.A(n_4682),
.Y(n_5105)
);

OAI21x1_ASAP7_75t_L g5106 ( 
.A1(n_4656),
.A2(n_4393),
.B(n_4332),
.Y(n_5106)
);

NAND2xp5_ASAP7_75t_L g5107 ( 
.A(n_4853),
.B(n_4412),
.Y(n_5107)
);

AOI221x1_ASAP7_75t_L g5108 ( 
.A1(n_4651),
.A2(n_4546),
.B1(n_4542),
.B2(n_4567),
.C(n_4555),
.Y(n_5108)
);

INVx2_ASAP7_75t_L g5109 ( 
.A(n_4625),
.Y(n_5109)
);

AND2x6_ASAP7_75t_SL g5110 ( 
.A(n_5039),
.B(n_4058),
.Y(n_5110)
);

NAND2xp5_ASAP7_75t_L g5111 ( 
.A(n_5025),
.B(n_4420),
.Y(n_5111)
);

INVxp67_ASAP7_75t_SL g5112 ( 
.A(n_4617),
.Y(n_5112)
);

INVx1_ASAP7_75t_L g5113 ( 
.A(n_4611),
.Y(n_5113)
);

AOI221x1_ASAP7_75t_L g5114 ( 
.A1(n_4796),
.A2(n_4591),
.B1(n_4590),
.B2(n_4570),
.C(n_4457),
.Y(n_5114)
);

AOI22xp33_ASAP7_75t_L g5115 ( 
.A1(n_4905),
.A2(n_4148),
.B1(n_4448),
.B2(n_4516),
.Y(n_5115)
);

OAI21x1_ASAP7_75t_L g5116 ( 
.A1(n_4620),
.A2(n_4365),
.B(n_4312),
.Y(n_5116)
);

INVxp67_ASAP7_75t_SL g5117 ( 
.A(n_4659),
.Y(n_5117)
);

AOI21xp5_ASAP7_75t_SL g5118 ( 
.A1(n_4914),
.A2(n_4297),
.B(n_4296),
.Y(n_5118)
);

NOR2x1_ASAP7_75t_R g5119 ( 
.A(n_5017),
.B(n_4353),
.Y(n_5119)
);

CKINVDCx5p33_ASAP7_75t_R g5120 ( 
.A(n_4801),
.Y(n_5120)
);

OA22x2_ASAP7_75t_L g5121 ( 
.A1(n_4840),
.A2(n_4297),
.B1(n_4323),
.B2(n_4296),
.Y(n_5121)
);

BUFx5_ASAP7_75t_L g5122 ( 
.A(n_4947),
.Y(n_5122)
);

BUFx8_ASAP7_75t_L g5123 ( 
.A(n_4919),
.Y(n_5123)
);

OAI21xp5_ASAP7_75t_L g5124 ( 
.A1(n_4776),
.A2(n_4433),
.B(n_4425),
.Y(n_5124)
);

AND2x2_ASAP7_75t_L g5125 ( 
.A(n_4751),
.B(n_4544),
.Y(n_5125)
);

OAI21xp5_ASAP7_75t_L g5126 ( 
.A1(n_4784),
.A2(n_4437),
.B(n_4434),
.Y(n_5126)
);

AND2x2_ASAP7_75t_L g5127 ( 
.A(n_4785),
.B(n_4544),
.Y(n_5127)
);

AO31x2_ASAP7_75t_L g5128 ( 
.A1(n_4856),
.A2(n_4466),
.A3(n_4517),
.B(n_4508),
.Y(n_5128)
);

NOR2xp33_ASAP7_75t_L g5129 ( 
.A(n_4774),
.B(n_4448),
.Y(n_5129)
);

AOI21x1_ASAP7_75t_SL g5130 ( 
.A1(n_4698),
.A2(n_4461),
.B(n_4529),
.Y(n_5130)
);

AOI21xp5_ASAP7_75t_L g5131 ( 
.A1(n_4606),
.A2(n_4283),
.B(n_4266),
.Y(n_5131)
);

AND2x2_ASAP7_75t_L g5132 ( 
.A(n_4958),
.B(n_4544),
.Y(n_5132)
);

OAI21x1_ASAP7_75t_L g5133 ( 
.A1(n_4661),
.A2(n_4452),
.B(n_4391),
.Y(n_5133)
);

AND2x2_ASAP7_75t_L g5134 ( 
.A(n_4636),
.B(n_4323),
.Y(n_5134)
);

AO21x2_ASAP7_75t_L g5135 ( 
.A1(n_4694),
.A2(n_4341),
.B(n_4333),
.Y(n_5135)
);

NAND2xp5_ASAP7_75t_L g5136 ( 
.A(n_4820),
.B(n_4333),
.Y(n_5136)
);

OAI21x1_ASAP7_75t_L g5137 ( 
.A1(n_4686),
.A2(n_4385),
.B(n_4140),
.Y(n_5137)
);

OAI21x1_ASAP7_75t_L g5138 ( 
.A1(n_4612),
.A2(n_4385),
.B(n_4140),
.Y(n_5138)
);

NAND2xp5_ASAP7_75t_L g5139 ( 
.A(n_4832),
.B(n_4341),
.Y(n_5139)
);

OAI21xp5_ASAP7_75t_L g5140 ( 
.A1(n_4869),
.A2(n_4046),
.B(n_4044),
.Y(n_5140)
);

AOI21xp5_ASAP7_75t_L g5141 ( 
.A1(n_4970),
.A2(n_4761),
.B(n_4640),
.Y(n_5141)
);

OAI21x1_ASAP7_75t_L g5142 ( 
.A1(n_4999),
.A2(n_4140),
.B(n_4283),
.Y(n_5142)
);

OAI21x1_ASAP7_75t_L g5143 ( 
.A1(n_4999),
.A2(n_4291),
.B(n_4283),
.Y(n_5143)
);

INVx5_ASAP7_75t_L g5144 ( 
.A(n_4613),
.Y(n_5144)
);

AOI21xp33_ASAP7_75t_L g5145 ( 
.A1(n_5075),
.A2(n_4360),
.B(n_4046),
.Y(n_5145)
);

AO21x2_ASAP7_75t_L g5146 ( 
.A1(n_4747),
.A2(n_4360),
.B(n_4101),
.Y(n_5146)
);

OAI21x1_ASAP7_75t_L g5147 ( 
.A1(n_4635),
.A2(n_4303),
.B(n_4291),
.Y(n_5147)
);

CKINVDCx5p33_ASAP7_75t_R g5148 ( 
.A(n_4628),
.Y(n_5148)
);

NOR2x1_ASAP7_75t_SL g5149 ( 
.A(n_4840),
.B(n_4994),
.Y(n_5149)
);

NOR2x1_ASAP7_75t_SL g5150 ( 
.A(n_4994),
.B(n_4291),
.Y(n_5150)
);

CKINVDCx5p33_ASAP7_75t_R g5151 ( 
.A(n_4714),
.Y(n_5151)
);

A2O1A1Ixp33_ASAP7_75t_L g5152 ( 
.A1(n_4665),
.A2(n_4101),
.B(n_4121),
.C(n_4044),
.Y(n_5152)
);

AND2x2_ASAP7_75t_SL g5153 ( 
.A(n_4678),
.B(n_4121),
.Y(n_5153)
);

NAND2xp5_ASAP7_75t_L g5154 ( 
.A(n_4629),
.B(n_4155),
.Y(n_5154)
);

INVx3_ASAP7_75t_L g5155 ( 
.A(n_4759),
.Y(n_5155)
);

INVx1_ASAP7_75t_L g5156 ( 
.A(n_4653),
.Y(n_5156)
);

INVx1_ASAP7_75t_L g5157 ( 
.A(n_4669),
.Y(n_5157)
);

INVx2_ASAP7_75t_L g5158 ( 
.A(n_4645),
.Y(n_5158)
);

OAI21x1_ASAP7_75t_L g5159 ( 
.A1(n_4858),
.A2(n_4306),
.B(n_4303),
.Y(n_5159)
);

AOI21xp5_ASAP7_75t_L g5160 ( 
.A1(n_4902),
.A2(n_4306),
.B(n_4303),
.Y(n_5160)
);

NAND2xp5_ASAP7_75t_L g5161 ( 
.A(n_4702),
.B(n_4155),
.Y(n_5161)
);

AOI21xp5_ASAP7_75t_L g5162 ( 
.A1(n_4750),
.A2(n_4350),
.B(n_4306),
.Y(n_5162)
);

NAND2xp5_ASAP7_75t_SL g5163 ( 
.A(n_4924),
.B(n_4350),
.Y(n_5163)
);

NAND2xp5_ASAP7_75t_L g5164 ( 
.A(n_4724),
.B(n_411),
.Y(n_5164)
);

NAND2xp5_ASAP7_75t_L g5165 ( 
.A(n_4733),
.B(n_412),
.Y(n_5165)
);

OAI21x1_ASAP7_75t_L g5166 ( 
.A1(n_4802),
.A2(n_4375),
.B(n_4350),
.Y(n_5166)
);

BUFx2_ASAP7_75t_L g5167 ( 
.A(n_4867),
.Y(n_5167)
);

OAI21xp5_ASAP7_75t_SL g5168 ( 
.A1(n_5019),
.A2(n_4449),
.B(n_4375),
.Y(n_5168)
);

AOI221xp5_ASAP7_75t_L g5169 ( 
.A1(n_4948),
.A2(n_4459),
.B1(n_4460),
.B2(n_4449),
.C(n_4375),
.Y(n_5169)
);

NAND2xp33_ASAP7_75t_L g5170 ( 
.A(n_4626),
.B(n_4449),
.Y(n_5170)
);

OAI21xp5_ASAP7_75t_L g5171 ( 
.A1(n_4689),
.A2(n_413),
.B(n_412),
.Y(n_5171)
);

AOI21xp5_ASAP7_75t_L g5172 ( 
.A1(n_5037),
.A2(n_4460),
.B(n_4459),
.Y(n_5172)
);

OAI21x1_ASAP7_75t_L g5173 ( 
.A1(n_5038),
.A2(n_4460),
.B(n_4459),
.Y(n_5173)
);

AOI21xp5_ASAP7_75t_L g5174 ( 
.A1(n_4622),
.A2(n_4847),
.B(n_4779),
.Y(n_5174)
);

AOI21xp33_ASAP7_75t_L g5175 ( 
.A1(n_4846),
.A2(n_4471),
.B(n_4468),
.Y(n_5175)
);

AOI21xp33_ASAP7_75t_L g5176 ( 
.A1(n_4649),
.A2(n_4817),
.B(n_4793),
.Y(n_5176)
);

INVx2_ASAP7_75t_L g5177 ( 
.A(n_4672),
.Y(n_5177)
);

NAND2xp5_ASAP7_75t_SL g5178 ( 
.A(n_4994),
.B(n_4468),
.Y(n_5178)
);

AND2x2_ASAP7_75t_SL g5179 ( 
.A(n_4678),
.B(n_4648),
.Y(n_5179)
);

AND2x2_ASAP7_75t_L g5180 ( 
.A(n_4704),
.B(n_4916),
.Y(n_5180)
);

OAI21x1_ASAP7_75t_L g5181 ( 
.A1(n_5007),
.A2(n_4471),
.B(n_4468),
.Y(n_5181)
);

CKINVDCx16_ASAP7_75t_R g5182 ( 
.A(n_4695),
.Y(n_5182)
);

OAI21x1_ASAP7_75t_SL g5183 ( 
.A1(n_4769),
.A2(n_413),
.B(n_412),
.Y(n_5183)
);

AOI21xp5_ASAP7_75t_L g5184 ( 
.A1(n_4755),
.A2(n_4515),
.B(n_4471),
.Y(n_5184)
);

BUFx2_ASAP7_75t_L g5185 ( 
.A(n_4836),
.Y(n_5185)
);

A2O1A1Ixp33_ASAP7_75t_L g5186 ( 
.A1(n_4634),
.A2(n_4533),
.B(n_4515),
.C(n_415),
.Y(n_5186)
);

OA21x2_ASAP7_75t_L g5187 ( 
.A1(n_4752),
.A2(n_4533),
.B(n_4515),
.Y(n_5187)
);

AOI21xp5_ASAP7_75t_L g5188 ( 
.A1(n_4627),
.A2(n_4533),
.B(n_415),
.Y(n_5188)
);

BUFx12f_ASAP7_75t_L g5189 ( 
.A(n_4735),
.Y(n_5189)
);

AND2x4_ASAP7_75t_L g5190 ( 
.A(n_5028),
.B(n_414),
.Y(n_5190)
);

NAND2xp5_ASAP7_75t_L g5191 ( 
.A(n_4743),
.B(n_414),
.Y(n_5191)
);

NAND2xp5_ASAP7_75t_L g5192 ( 
.A(n_4756),
.B(n_4762),
.Y(n_5192)
);

NAND2xp5_ASAP7_75t_L g5193 ( 
.A(n_4768),
.B(n_414),
.Y(n_5193)
);

NAND2xp5_ASAP7_75t_L g5194 ( 
.A(n_4807),
.B(n_416),
.Y(n_5194)
);

NAND2xp5_ASAP7_75t_L g5195 ( 
.A(n_4849),
.B(n_416),
.Y(n_5195)
);

INVx1_ASAP7_75t_L g5196 ( 
.A(n_4646),
.Y(n_5196)
);

AOI21xp5_ASAP7_75t_L g5197 ( 
.A1(n_4631),
.A2(n_417),
.B(n_416),
.Y(n_5197)
);

NAND2xp5_ASAP7_75t_L g5198 ( 
.A(n_5063),
.B(n_417),
.Y(n_5198)
);

OAI21x1_ASAP7_75t_L g5199 ( 
.A1(n_5029),
.A2(n_418),
.B(n_417),
.Y(n_5199)
);

OAI21xp5_ASAP7_75t_L g5200 ( 
.A1(n_4850),
.A2(n_419),
.B(n_418),
.Y(n_5200)
);

AOI21xp5_ASAP7_75t_SL g5201 ( 
.A1(n_4698),
.A2(n_419),
.B(n_418),
.Y(n_5201)
);

AO31x2_ASAP7_75t_L g5202 ( 
.A1(n_5005),
.A2(n_420),
.A3(n_421),
.B(n_419),
.Y(n_5202)
);

OAI21x1_ASAP7_75t_L g5203 ( 
.A1(n_4758),
.A2(n_421),
.B(n_420),
.Y(n_5203)
);

NAND2xp5_ASAP7_75t_L g5204 ( 
.A(n_5070),
.B(n_420),
.Y(n_5204)
);

OAI21xp5_ASAP7_75t_L g5205 ( 
.A1(n_5073),
.A2(n_423),
.B(n_422),
.Y(n_5205)
);

INVxp67_ASAP7_75t_L g5206 ( 
.A(n_4997),
.Y(n_5206)
);

AOI21xp33_ASAP7_75t_L g5207 ( 
.A1(n_4657),
.A2(n_4975),
.B(n_4959),
.Y(n_5207)
);

HB1xp67_ASAP7_75t_L g5208 ( 
.A(n_4822),
.Y(n_5208)
);

NAND2xp5_ASAP7_75t_L g5209 ( 
.A(n_4899),
.B(n_422),
.Y(n_5209)
);

NOR2xp33_ASAP7_75t_L g5210 ( 
.A(n_4813),
.B(n_4),
.Y(n_5210)
);

AOI21xp5_ASAP7_75t_L g5211 ( 
.A1(n_4632),
.A2(n_424),
.B(n_423),
.Y(n_5211)
);

INVx3_ASAP7_75t_L g5212 ( 
.A(n_4626),
.Y(n_5212)
);

OAI21x1_ASAP7_75t_L g5213 ( 
.A1(n_4713),
.A2(n_424),
.B(n_423),
.Y(n_5213)
);

INVx1_ASAP7_75t_L g5214 ( 
.A(n_4683),
.Y(n_5214)
);

INVx2_ASAP7_75t_L g5215 ( 
.A(n_4674),
.Y(n_5215)
);

OAI21x1_ASAP7_75t_L g5216 ( 
.A1(n_4688),
.A2(n_425),
.B(n_424),
.Y(n_5216)
);

AOI21xp5_ASAP7_75t_L g5217 ( 
.A1(n_4637),
.A2(n_4624),
.B(n_4736),
.Y(n_5217)
);

OAI21x1_ASAP7_75t_L g5218 ( 
.A1(n_4688),
.A2(n_426),
.B(n_425),
.Y(n_5218)
);

AOI21xp5_ASAP7_75t_L g5219 ( 
.A1(n_4806),
.A2(n_426),
.B(n_425),
.Y(n_5219)
);

NOR2x1_ASAP7_75t_SL g5220 ( 
.A(n_5028),
.B(n_426),
.Y(n_5220)
);

NAND2xp5_ASAP7_75t_L g5221 ( 
.A(n_4909),
.B(n_427),
.Y(n_5221)
);

INVx4_ASAP7_75t_L g5222 ( 
.A(n_4754),
.Y(n_5222)
);

BUFx2_ASAP7_75t_L g5223 ( 
.A(n_4931),
.Y(n_5223)
);

BUFx10_ASAP7_75t_L g5224 ( 
.A(n_4690),
.Y(n_5224)
);

NAND2xp33_ASAP7_75t_L g5225 ( 
.A(n_5047),
.B(n_427),
.Y(n_5225)
);

AO31x2_ASAP7_75t_L g5226 ( 
.A1(n_4739),
.A2(n_428),
.A3(n_429),
.B(n_427),
.Y(n_5226)
);

OAI21x1_ASAP7_75t_L g5227 ( 
.A1(n_4931),
.A2(n_430),
.B(n_429),
.Y(n_5227)
);

AO21x2_ASAP7_75t_L g5228 ( 
.A1(n_5015),
.A2(n_430),
.B(n_429),
.Y(n_5228)
);

AOI21x1_ASAP7_75t_L g5229 ( 
.A1(n_5000),
.A2(n_431),
.B(n_430),
.Y(n_5229)
);

NAND2xp5_ASAP7_75t_L g5230 ( 
.A(n_4932),
.B(n_431),
.Y(n_5230)
);

OAI21x1_ASAP7_75t_L g5231 ( 
.A1(n_4980),
.A2(n_433),
.B(n_432),
.Y(n_5231)
);

INVx3_ASAP7_75t_L g5232 ( 
.A(n_4976),
.Y(n_5232)
);

OAI21x1_ASAP7_75t_L g5233 ( 
.A1(n_4980),
.A2(n_433),
.B(n_432),
.Y(n_5233)
);

INVxp67_ASAP7_75t_L g5234 ( 
.A(n_4986),
.Y(n_5234)
);

INVx1_ASAP7_75t_L g5235 ( 
.A(n_4757),
.Y(n_5235)
);

AOI21xp5_ASAP7_75t_L g5236 ( 
.A1(n_4848),
.A2(n_434),
.B(n_432),
.Y(n_5236)
);

OAI21xp5_ASAP7_75t_L g5237 ( 
.A1(n_4641),
.A2(n_435),
.B(n_434),
.Y(n_5237)
);

OAI21xp5_ASAP7_75t_L g5238 ( 
.A1(n_4652),
.A2(n_436),
.B(n_435),
.Y(n_5238)
);

NOR2x1_ASAP7_75t_L g5239 ( 
.A(n_4910),
.B(n_436),
.Y(n_5239)
);

INVx1_ASAP7_75t_SL g5240 ( 
.A(n_5004),
.Y(n_5240)
);

AOI21xp5_ASAP7_75t_L g5241 ( 
.A1(n_4812),
.A2(n_437),
.B(n_436),
.Y(n_5241)
);

INVx1_ASAP7_75t_L g5242 ( 
.A(n_4799),
.Y(n_5242)
);

OAI22x1_ASAP7_75t_L g5243 ( 
.A1(n_5023),
.A2(n_438),
.B1(n_439),
.B2(n_437),
.Y(n_5243)
);

INVx3_ASAP7_75t_L g5244 ( 
.A(n_4721),
.Y(n_5244)
);

AOI21xp33_ASAP7_75t_L g5245 ( 
.A1(n_4898),
.A2(n_438),
.B(n_437),
.Y(n_5245)
);

INVx3_ASAP7_75t_L g5246 ( 
.A(n_4721),
.Y(n_5246)
);

NAND2xp5_ASAP7_75t_L g5247 ( 
.A(n_4950),
.B(n_439),
.Y(n_5247)
);

AND2x6_ASAP7_75t_L g5248 ( 
.A(n_4947),
.B(n_439),
.Y(n_5248)
);

OAI21xp5_ASAP7_75t_L g5249 ( 
.A1(n_5046),
.A2(n_442),
.B(n_440),
.Y(n_5249)
);

NAND2xp5_ASAP7_75t_L g5250 ( 
.A(n_5014),
.B(n_440),
.Y(n_5250)
);

INVx2_ASAP7_75t_L g5251 ( 
.A(n_4679),
.Y(n_5251)
);

AOI21xp5_ASAP7_75t_L g5252 ( 
.A1(n_4885),
.A2(n_443),
.B(n_440),
.Y(n_5252)
);

NAND2xp5_ASAP7_75t_L g5253 ( 
.A(n_4874),
.B(n_443),
.Y(n_5253)
);

INVx1_ASAP7_75t_L g5254 ( 
.A(n_4685),
.Y(n_5254)
);

AOI21xp5_ASAP7_75t_L g5255 ( 
.A1(n_4882),
.A2(n_444),
.B(n_443),
.Y(n_5255)
);

NAND2xp5_ASAP7_75t_L g5256 ( 
.A(n_4711),
.B(n_444),
.Y(n_5256)
);

NAND2xp5_ASAP7_75t_L g5257 ( 
.A(n_4737),
.B(n_445),
.Y(n_5257)
);

BUFx10_ASAP7_75t_L g5258 ( 
.A(n_4715),
.Y(n_5258)
);

OA22x2_ASAP7_75t_L g5259 ( 
.A1(n_5064),
.A2(n_5071),
.B1(n_4923),
.B2(n_4985),
.Y(n_5259)
);

INVx3_ASAP7_75t_L g5260 ( 
.A(n_4721),
.Y(n_5260)
);

OAI22x1_ASAP7_75t_L g5261 ( 
.A1(n_4894),
.A2(n_446),
.B1(n_447),
.B2(n_445),
.Y(n_5261)
);

OAI21x1_ASAP7_75t_L g5262 ( 
.A1(n_4644),
.A2(n_446),
.B(n_445),
.Y(n_5262)
);

OAI21xp5_ASAP7_75t_SL g5263 ( 
.A1(n_4913),
.A2(n_447),
.B(n_446),
.Y(n_5263)
);

INVx5_ASAP7_75t_L g5264 ( 
.A(n_5028),
.Y(n_5264)
);

INVx4_ASAP7_75t_L g5265 ( 
.A(n_4881),
.Y(n_5265)
);

OR2x2_ASAP7_75t_L g5266 ( 
.A(n_4993),
.B(n_447),
.Y(n_5266)
);

INVx3_ASAP7_75t_SL g5267 ( 
.A(n_4729),
.Y(n_5267)
);

OAI21x1_ASAP7_75t_L g5268 ( 
.A1(n_5026),
.A2(n_449),
.B(n_448),
.Y(n_5268)
);

NAND2xp5_ASAP7_75t_L g5269 ( 
.A(n_4748),
.B(n_4763),
.Y(n_5269)
);

AND2x4_ASAP7_75t_L g5270 ( 
.A(n_4771),
.B(n_4828),
.Y(n_5270)
);

OAI21x1_ASAP7_75t_L g5271 ( 
.A1(n_4834),
.A2(n_4601),
.B(n_4642),
.Y(n_5271)
);

AOI21xp33_ASAP7_75t_L g5272 ( 
.A1(n_5032),
.A2(n_450),
.B(n_448),
.Y(n_5272)
);

CKINVDCx16_ASAP7_75t_R g5273 ( 
.A(n_4900),
.Y(n_5273)
);

AOI21xp33_ASAP7_75t_L g5274 ( 
.A1(n_4615),
.A2(n_5042),
.B(n_4718),
.Y(n_5274)
);

AOI21xp33_ASAP7_75t_L g5275 ( 
.A1(n_4953),
.A2(n_450),
.B(n_448),
.Y(n_5275)
);

AOI221x1_ASAP7_75t_L g5276 ( 
.A1(n_4871),
.A2(n_453),
.B1(n_454),
.B2(n_452),
.C(n_451),
.Y(n_5276)
);

AND2x4_ASAP7_75t_L g5277 ( 
.A(n_4771),
.B(n_451),
.Y(n_5277)
);

NAND2xp5_ASAP7_75t_L g5278 ( 
.A(n_4767),
.B(n_451),
.Y(n_5278)
);

NAND2xp5_ASAP7_75t_L g5279 ( 
.A(n_4773),
.B(n_452),
.Y(n_5279)
);

CKINVDCx16_ASAP7_75t_R g5280 ( 
.A(n_4775),
.Y(n_5280)
);

NAND2x1_ASAP7_75t_L g5281 ( 
.A(n_4828),
.B(n_452),
.Y(n_5281)
);

AND2x2_ASAP7_75t_L g5282 ( 
.A(n_5034),
.B(n_4),
.Y(n_5282)
);

AOI21xp33_ASAP7_75t_L g5283 ( 
.A1(n_5056),
.A2(n_454),
.B(n_453),
.Y(n_5283)
);

AND2x2_ASAP7_75t_L g5284 ( 
.A(n_5030),
.B(n_5),
.Y(n_5284)
);

OAI21x1_ASAP7_75t_SL g5285 ( 
.A1(n_5057),
.A2(n_454),
.B(n_453),
.Y(n_5285)
);

NAND2xp5_ASAP7_75t_L g5286 ( 
.A(n_4780),
.B(n_455),
.Y(n_5286)
);

INVx2_ASAP7_75t_L g5287 ( 
.A(n_4800),
.Y(n_5287)
);

AOI21xp5_ASAP7_75t_L g5288 ( 
.A1(n_4602),
.A2(n_457),
.B(n_456),
.Y(n_5288)
);

INVx4_ASAP7_75t_L g5289 ( 
.A(n_4731),
.Y(n_5289)
);

HB1xp67_ASAP7_75t_L g5290 ( 
.A(n_4852),
.Y(n_5290)
);

AND2x2_ASAP7_75t_L g5291 ( 
.A(n_5043),
.B(n_4691),
.Y(n_5291)
);

OAI21xp5_ASAP7_75t_L g5292 ( 
.A1(n_4650),
.A2(n_4833),
.B(n_4744),
.Y(n_5292)
);

INVx1_ASAP7_75t_L g5293 ( 
.A(n_4861),
.Y(n_5293)
);

OAI21x1_ASAP7_75t_L g5294 ( 
.A1(n_4742),
.A2(n_458),
.B(n_457),
.Y(n_5294)
);

NAND2xp5_ASAP7_75t_L g5295 ( 
.A(n_4865),
.B(n_457),
.Y(n_5295)
);

OAI21xp33_ASAP7_75t_L g5296 ( 
.A1(n_4983),
.A2(n_459),
.B(n_458),
.Y(n_5296)
);

O2A1O1Ixp5_ASAP7_75t_L g5297 ( 
.A1(n_4660),
.A2(n_461),
.B(n_462),
.C(n_460),
.Y(n_5297)
);

OAI21x1_ASAP7_75t_L g5298 ( 
.A1(n_4746),
.A2(n_4701),
.B(n_4870),
.Y(n_5298)
);

NAND2xp5_ASAP7_75t_L g5299 ( 
.A(n_4884),
.B(n_460),
.Y(n_5299)
);

AO21x1_ASAP7_75t_L g5300 ( 
.A1(n_5033),
.A2(n_461),
.B(n_460),
.Y(n_5300)
);

NAND2xp5_ASAP7_75t_SL g5301 ( 
.A(n_4731),
.B(n_461),
.Y(n_5301)
);

INVx2_ASAP7_75t_SL g5302 ( 
.A(n_4876),
.Y(n_5302)
);

HB1xp67_ASAP7_75t_L g5303 ( 
.A(n_4889),
.Y(n_5303)
);

NOR2xp67_ASAP7_75t_L g5304 ( 
.A(n_5076),
.B(n_465),
.Y(n_5304)
);

NAND2xp5_ASAP7_75t_L g5305 ( 
.A(n_4939),
.B(n_463),
.Y(n_5305)
);

AND2x2_ASAP7_75t_L g5306 ( 
.A(n_4706),
.B(n_5),
.Y(n_5306)
);

AOI21xp5_ASAP7_75t_L g5307 ( 
.A1(n_4607),
.A2(n_464),
.B(n_463),
.Y(n_5307)
);

NAND2xp5_ASAP7_75t_L g5308 ( 
.A(n_4940),
.B(n_464),
.Y(n_5308)
);

NAND2xp5_ASAP7_75t_L g5309 ( 
.A(n_4949),
.B(n_465),
.Y(n_5309)
);

OAI21x1_ASAP7_75t_L g5310 ( 
.A1(n_4681),
.A2(n_467),
.B(n_466),
.Y(n_5310)
);

AOI21xp5_ASAP7_75t_L g5311 ( 
.A1(n_4667),
.A2(n_468),
.B(n_466),
.Y(n_5311)
);

HB1xp67_ASAP7_75t_L g5312 ( 
.A(n_5068),
.Y(n_5312)
);

NAND2xp5_ASAP7_75t_SL g5313 ( 
.A(n_4731),
.B(n_4830),
.Y(n_5313)
);

OAI21xp5_ASAP7_75t_L g5314 ( 
.A1(n_5027),
.A2(n_469),
.B(n_468),
.Y(n_5314)
);

INVxp67_ASAP7_75t_L g5315 ( 
.A(n_4930),
.Y(n_5315)
);

NAND2xp5_ASAP7_75t_L g5316 ( 
.A(n_4719),
.B(n_469),
.Y(n_5316)
);

OAI21x1_ASAP7_75t_L g5317 ( 
.A1(n_4684),
.A2(n_5051),
.B(n_4978),
.Y(n_5317)
);

NOR2x1_ASAP7_75t_L g5318 ( 
.A(n_4738),
.B(n_469),
.Y(n_5318)
);

OA22x2_ASAP7_75t_L g5319 ( 
.A1(n_4666),
.A2(n_471),
.B1(n_472),
.B2(n_470),
.Y(n_5319)
);

AO21x1_ASAP7_75t_L g5320 ( 
.A1(n_4716),
.A2(n_4996),
.B(n_5021),
.Y(n_5320)
);

AOI21x1_ASAP7_75t_SL g5321 ( 
.A1(n_4854),
.A2(n_471),
.B(n_470),
.Y(n_5321)
);

AND2x2_ASAP7_75t_L g5322 ( 
.A(n_4934),
.B(n_6),
.Y(n_5322)
);

AOI21x1_ASAP7_75t_L g5323 ( 
.A1(n_5067),
.A2(n_471),
.B(n_470),
.Y(n_5323)
);

BUFx12f_ASAP7_75t_L g5324 ( 
.A(n_4995),
.Y(n_5324)
);

AOI21xp5_ASAP7_75t_L g5325 ( 
.A1(n_4680),
.A2(n_473),
.B(n_472),
.Y(n_5325)
);

AOI21x1_ASAP7_75t_L g5326 ( 
.A1(n_5072),
.A2(n_474),
.B(n_473),
.Y(n_5326)
);

A2O1A1Ixp33_ASAP7_75t_L g5327 ( 
.A1(n_4697),
.A2(n_475),
.B(n_476),
.C(n_474),
.Y(n_5327)
);

OAI21x1_ASAP7_75t_L g5328 ( 
.A1(n_4864),
.A2(n_4823),
.B(n_4844),
.Y(n_5328)
);

OAI21x1_ASAP7_75t_L g5329 ( 
.A1(n_4860),
.A2(n_476),
.B(n_475),
.Y(n_5329)
);

OAI22x1_ASAP7_75t_L g5330 ( 
.A1(n_5054),
.A2(n_477),
.B1(n_478),
.B2(n_476),
.Y(n_5330)
);

AND2x4_ASAP7_75t_L g5331 ( 
.A(n_4830),
.B(n_477),
.Y(n_5331)
);

BUFx6f_ASAP7_75t_L g5332 ( 
.A(n_4830),
.Y(n_5332)
);

CKINVDCx5p33_ASAP7_75t_R g5333 ( 
.A(n_4673),
.Y(n_5333)
);

NAND2xp5_ASAP7_75t_L g5334 ( 
.A(n_4835),
.B(n_478),
.Y(n_5334)
);

A2O1A1Ixp33_ASAP7_75t_L g5335 ( 
.A1(n_4778),
.A2(n_479),
.B(n_480),
.C(n_478),
.Y(n_5335)
);

INVx5_ASAP7_75t_L g5336 ( 
.A(n_4836),
.Y(n_5336)
);

AOI21xp33_ASAP7_75t_L g5337 ( 
.A1(n_5052),
.A2(n_480),
.B(n_479),
.Y(n_5337)
);

NOR2x1_ASAP7_75t_SL g5338 ( 
.A(n_4952),
.B(n_479),
.Y(n_5338)
);

INVx2_ASAP7_75t_SL g5339 ( 
.A(n_4831),
.Y(n_5339)
);

OAI21x1_ASAP7_75t_L g5340 ( 
.A1(n_4766),
.A2(n_481),
.B(n_480),
.Y(n_5340)
);

NOR2xp67_ASAP7_75t_L g5341 ( 
.A(n_4841),
.B(n_484),
.Y(n_5341)
);

A2O1A1Ixp33_ASAP7_75t_L g5342 ( 
.A1(n_4987),
.A2(n_482),
.B(n_483),
.C(n_481),
.Y(n_5342)
);

AOI21x1_ASAP7_75t_L g5343 ( 
.A1(n_4906),
.A2(n_482),
.B(n_481),
.Y(n_5343)
);

INVx1_ASAP7_75t_L g5344 ( 
.A(n_4992),
.Y(n_5344)
);

OAI21x1_ASAP7_75t_SL g5345 ( 
.A1(n_4829),
.A2(n_483),
.B(n_482),
.Y(n_5345)
);

OAI21x1_ASAP7_75t_L g5346 ( 
.A1(n_4766),
.A2(n_4912),
.B(n_4883),
.Y(n_5346)
);

AOI21xp5_ASAP7_75t_L g5347 ( 
.A1(n_4608),
.A2(n_484),
.B(n_483),
.Y(n_5347)
);

AO21x1_ASAP7_75t_L g5348 ( 
.A1(n_4922),
.A2(n_4671),
.B(n_4707),
.Y(n_5348)
);

OAI21x1_ASAP7_75t_L g5349 ( 
.A1(n_5053),
.A2(n_485),
.B(n_484),
.Y(n_5349)
);

CKINVDCx5p33_ASAP7_75t_R g5350 ( 
.A(n_4675),
.Y(n_5350)
);

NAND2xp5_ASAP7_75t_L g5351 ( 
.A(n_4610),
.B(n_485),
.Y(n_5351)
);

NAND2xp5_ASAP7_75t_SL g5352 ( 
.A(n_4753),
.B(n_485),
.Y(n_5352)
);

AND2x2_ASAP7_75t_L g5353 ( 
.A(n_4972),
.B(n_6),
.Y(n_5353)
);

AO21x2_ASAP7_75t_L g5354 ( 
.A1(n_4839),
.A2(n_487),
.B(n_486),
.Y(n_5354)
);

CKINVDCx5p33_ASAP7_75t_R g5355 ( 
.A(n_4873),
.Y(n_5355)
);

OAI21x1_ASAP7_75t_L g5356 ( 
.A1(n_4951),
.A2(n_487),
.B(n_486),
.Y(n_5356)
);

OAI21x1_ASAP7_75t_L g5357 ( 
.A1(n_4819),
.A2(n_488),
.B(n_486),
.Y(n_5357)
);

CKINVDCx11_ASAP7_75t_R g5358 ( 
.A(n_4836),
.Y(n_5358)
);

AOI21xp5_ASAP7_75t_L g5359 ( 
.A1(n_4845),
.A2(n_489),
.B(n_488),
.Y(n_5359)
);

AND2x2_ASAP7_75t_L g5360 ( 
.A(n_4851),
.B(n_6),
.Y(n_5360)
);

INVx1_ASAP7_75t_SL g5361 ( 
.A(n_4990),
.Y(n_5361)
);

AND2x2_ASAP7_75t_L g5362 ( 
.A(n_4803),
.B(n_4886),
.Y(n_5362)
);

OAI21x1_ASAP7_75t_L g5363 ( 
.A1(n_4696),
.A2(n_489),
.B(n_488),
.Y(n_5363)
);

INVx2_ASAP7_75t_L g5364 ( 
.A(n_4944),
.Y(n_5364)
);

OAI21x1_ASAP7_75t_L g5365 ( 
.A1(n_4989),
.A2(n_490),
.B(n_489),
.Y(n_5365)
);

AO21x1_ASAP7_75t_L g5366 ( 
.A1(n_4741),
.A2(n_492),
.B(n_491),
.Y(n_5366)
);

AOI22xp33_ASAP7_75t_L g5367 ( 
.A1(n_4783),
.A2(n_492),
.B1(n_493),
.B2(n_491),
.Y(n_5367)
);

INVx2_ASAP7_75t_SL g5368 ( 
.A(n_4944),
.Y(n_5368)
);

NAND2xp5_ASAP7_75t_L g5369 ( 
.A(n_4917),
.B(n_491),
.Y(n_5369)
);

AOI21x1_ASAP7_75t_L g5370 ( 
.A1(n_4956),
.A2(n_494),
.B(n_493),
.Y(n_5370)
);

OAI21x1_ASAP7_75t_L g5371 ( 
.A1(n_4654),
.A2(n_494),
.B(n_493),
.Y(n_5371)
);

AOI21x1_ASAP7_75t_L g5372 ( 
.A1(n_4960),
.A2(n_495),
.B(n_494),
.Y(n_5372)
);

BUFx3_ASAP7_75t_L g5373 ( 
.A(n_4944),
.Y(n_5373)
);

AOI21x1_ASAP7_75t_L g5374 ( 
.A1(n_4961),
.A2(n_497),
.B(n_496),
.Y(n_5374)
);

AOI22xp33_ASAP7_75t_SL g5375 ( 
.A1(n_4708),
.A2(n_1068),
.B1(n_1070),
.B2(n_1063),
.Y(n_5375)
);

NAND2xp5_ASAP7_75t_L g5376 ( 
.A(n_4816),
.B(n_496),
.Y(n_5376)
);

A2O1A1Ixp33_ASAP7_75t_L g5377 ( 
.A1(n_4838),
.A2(n_498),
.B(n_499),
.C(n_497),
.Y(n_5377)
);

OAI21x1_ASAP7_75t_L g5378 ( 
.A1(n_4655),
.A2(n_4670),
.B(n_4664),
.Y(n_5378)
);

INVx3_ASAP7_75t_SL g5379 ( 
.A(n_4946),
.Y(n_5379)
);

AO31x2_ASAP7_75t_L g5380 ( 
.A1(n_4795),
.A2(n_499),
.A3(n_500),
.B(n_498),
.Y(n_5380)
);

INVx3_ASAP7_75t_L g5381 ( 
.A(n_4946),
.Y(n_5381)
);

AOI21xp5_ASAP7_75t_L g5382 ( 
.A1(n_4936),
.A2(n_500),
.B(n_498),
.Y(n_5382)
);

AOI21xp5_ASAP7_75t_L g5383 ( 
.A1(n_4969),
.A2(n_501),
.B(n_500),
.Y(n_5383)
);

OAI21x1_ASAP7_75t_L g5384 ( 
.A1(n_4712),
.A2(n_4730),
.B(n_4727),
.Y(n_5384)
);

INVx6_ASAP7_75t_SL g5385 ( 
.A(n_5055),
.Y(n_5385)
);

INVx2_ASAP7_75t_L g5386 ( 
.A(n_4946),
.Y(n_5386)
);

INVxp67_ASAP7_75t_SL g5387 ( 
.A(n_4965),
.Y(n_5387)
);

OAI21x1_ASAP7_75t_L g5388 ( 
.A1(n_4734),
.A2(n_502),
.B(n_501),
.Y(n_5388)
);

OAI22xp5_ASAP7_75t_L g5389 ( 
.A1(n_4699),
.A2(n_503),
.B1(n_504),
.B2(n_502),
.Y(n_5389)
);

NAND2xp5_ASAP7_75t_L g5390 ( 
.A(n_4962),
.B(n_502),
.Y(n_5390)
);

NAND2xp5_ASAP7_75t_L g5391 ( 
.A(n_4967),
.B(n_504),
.Y(n_5391)
);

AOI21x1_ASAP7_75t_L g5392 ( 
.A1(n_4973),
.A2(n_4982),
.B(n_4966),
.Y(n_5392)
);

AOI21xp5_ASAP7_75t_L g5393 ( 
.A1(n_4837),
.A2(n_4963),
.B(n_4878),
.Y(n_5393)
);

NAND2xp5_ASAP7_75t_SL g5394 ( 
.A(n_4965),
.B(n_505),
.Y(n_5394)
);

OAI21x1_ASAP7_75t_L g5395 ( 
.A1(n_4765),
.A2(n_506),
.B(n_505),
.Y(n_5395)
);

OAI21xp5_ASAP7_75t_L g5396 ( 
.A1(n_4872),
.A2(n_507),
.B(n_505),
.Y(n_5396)
);

BUFx12f_ASAP7_75t_L g5397 ( 
.A(n_5090),
.Y(n_5397)
);

BUFx3_ASAP7_75t_L g5398 ( 
.A(n_5105),
.Y(n_5398)
);

INVx1_ASAP7_75t_SL g5399 ( 
.A(n_5222),
.Y(n_5399)
);

INVx3_ASAP7_75t_L g5400 ( 
.A(n_5224),
.Y(n_5400)
);

INVx11_ASAP7_75t_L g5401 ( 
.A(n_5123),
.Y(n_5401)
);

AOI21xp5_ASAP7_75t_L g5402 ( 
.A1(n_5118),
.A2(n_5079),
.B(n_5162),
.Y(n_5402)
);

AO21x2_ASAP7_75t_L g5403 ( 
.A1(n_5084),
.A2(n_5011),
.B(n_4998),
.Y(n_5403)
);

INVx1_ASAP7_75t_SL g5404 ( 
.A(n_5189),
.Y(n_5404)
);

INVx1_ASAP7_75t_L g5405 ( 
.A(n_5087),
.Y(n_5405)
);

AND2x2_ASAP7_75t_L g5406 ( 
.A(n_5080),
.B(n_4621),
.Y(n_5406)
);

BUFx2_ASAP7_75t_SL g5407 ( 
.A(n_5102),
.Y(n_5407)
);

INVx1_ASAP7_75t_L g5408 ( 
.A(n_5113),
.Y(n_5408)
);

INVx1_ASAP7_75t_L g5409 ( 
.A(n_5156),
.Y(n_5409)
);

INVx2_ASAP7_75t_L g5410 ( 
.A(n_5290),
.Y(n_5410)
);

NAND2xp5_ASAP7_75t_L g5411 ( 
.A(n_5196),
.B(n_5059),
.Y(n_5411)
);

INVx1_ASAP7_75t_L g5412 ( 
.A(n_5157),
.Y(n_5412)
);

NAND2xp5_ASAP7_75t_L g5413 ( 
.A(n_5214),
.B(n_5060),
.Y(n_5413)
);

INVxp67_ASAP7_75t_SL g5414 ( 
.A(n_5303),
.Y(n_5414)
);

INVx1_ASAP7_75t_L g5415 ( 
.A(n_5192),
.Y(n_5415)
);

INVx3_ASAP7_75t_L g5416 ( 
.A(n_5265),
.Y(n_5416)
);

INVx4_ASAP7_75t_L g5417 ( 
.A(n_5148),
.Y(n_5417)
);

INVx1_ASAP7_75t_L g5418 ( 
.A(n_5208),
.Y(n_5418)
);

BUFx3_ASAP7_75t_L g5419 ( 
.A(n_5167),
.Y(n_5419)
);

BUFx12f_ASAP7_75t_L g5420 ( 
.A(n_5151),
.Y(n_5420)
);

BUFx6f_ASAP7_75t_L g5421 ( 
.A(n_5358),
.Y(n_5421)
);

BUFx3_ASAP7_75t_L g5422 ( 
.A(n_5339),
.Y(n_5422)
);

BUFx2_ASAP7_75t_R g5423 ( 
.A(n_5120),
.Y(n_5423)
);

BUFx6f_ASAP7_75t_L g5424 ( 
.A(n_5103),
.Y(n_5424)
);

BUFx3_ASAP7_75t_L g5425 ( 
.A(n_5267),
.Y(n_5425)
);

BUFx2_ASAP7_75t_L g5426 ( 
.A(n_5088),
.Y(n_5426)
);

BUFx3_ASAP7_75t_L g5427 ( 
.A(n_5302),
.Y(n_5427)
);

BUFx3_ASAP7_75t_L g5428 ( 
.A(n_5324),
.Y(n_5428)
);

INVx1_ASAP7_75t_SL g5429 ( 
.A(n_5240),
.Y(n_5429)
);

BUFx12f_ASAP7_75t_L g5430 ( 
.A(n_5110),
.Y(n_5430)
);

BUFx12f_ASAP7_75t_L g5431 ( 
.A(n_5258),
.Y(n_5431)
);

INVxp67_ASAP7_75t_SL g5432 ( 
.A(n_5112),
.Y(n_5432)
);

BUFx6f_ASAP7_75t_L g5433 ( 
.A(n_5103),
.Y(n_5433)
);

NOR2xp33_ASAP7_75t_L g5434 ( 
.A(n_5119),
.B(n_4623),
.Y(n_5434)
);

AOI22xp33_ASAP7_75t_L g5435 ( 
.A1(n_5083),
.A2(n_4880),
.B1(n_4700),
.B2(n_4723),
.Y(n_5435)
);

INVx6_ASAP7_75t_L g5436 ( 
.A(n_5182),
.Y(n_5436)
);

INVx2_ASAP7_75t_SL g5437 ( 
.A(n_5086),
.Y(n_5437)
);

INVxp67_ASAP7_75t_SL g5438 ( 
.A(n_5117),
.Y(n_5438)
);

INVx1_ASAP7_75t_L g5439 ( 
.A(n_5235),
.Y(n_5439)
);

OR2x2_ASAP7_75t_L g5440 ( 
.A(n_5180),
.B(n_5012),
.Y(n_5440)
);

BUFx6f_ASAP7_75t_L g5441 ( 
.A(n_5332),
.Y(n_5441)
);

INVx3_ASAP7_75t_L g5442 ( 
.A(n_5098),
.Y(n_5442)
);

CKINVDCx11_ASAP7_75t_R g5443 ( 
.A(n_5273),
.Y(n_5443)
);

INVx1_ASAP7_75t_L g5444 ( 
.A(n_5242),
.Y(n_5444)
);

CKINVDCx11_ASAP7_75t_R g5445 ( 
.A(n_5280),
.Y(n_5445)
);

INVx1_ASAP7_75t_L g5446 ( 
.A(n_5254),
.Y(n_5446)
);

BUFx5_ASAP7_75t_L g5447 ( 
.A(n_5248),
.Y(n_5447)
);

CKINVDCx20_ASAP7_75t_R g5448 ( 
.A(n_5232),
.Y(n_5448)
);

INVx2_ASAP7_75t_SL g5449 ( 
.A(n_5127),
.Y(n_5449)
);

NOR2xp33_ASAP7_75t_L g5450 ( 
.A(n_5094),
.B(n_4920),
.Y(n_5450)
);

INVx1_ASAP7_75t_SL g5451 ( 
.A(n_5125),
.Y(n_5451)
);

INVx1_ASAP7_75t_L g5452 ( 
.A(n_5293),
.Y(n_5452)
);

INVx2_ASAP7_75t_L g5453 ( 
.A(n_5081),
.Y(n_5453)
);

BUFx2_ASAP7_75t_L g5454 ( 
.A(n_5223),
.Y(n_5454)
);

BUFx4_ASAP7_75t_R g5455 ( 
.A(n_5149),
.Y(n_5455)
);

INVx1_ASAP7_75t_SL g5456 ( 
.A(n_5312),
.Y(n_5456)
);

INVxp67_ASAP7_75t_SL g5457 ( 
.A(n_5269),
.Y(n_5457)
);

INVx2_ASAP7_75t_L g5458 ( 
.A(n_5109),
.Y(n_5458)
);

INVxp67_ASAP7_75t_SL g5459 ( 
.A(n_5158),
.Y(n_5459)
);

NAND2x1p5_ASAP7_75t_L g5460 ( 
.A(n_5098),
.B(n_5048),
.Y(n_5460)
);

NAND2xp5_ASAP7_75t_L g5461 ( 
.A(n_5344),
.B(n_5066),
.Y(n_5461)
);

INVx3_ASAP7_75t_L g5462 ( 
.A(n_5098),
.Y(n_5462)
);

BUFx3_ASAP7_75t_L g5463 ( 
.A(n_5129),
.Y(n_5463)
);

BUFx12f_ASAP7_75t_L g5464 ( 
.A(n_5179),
.Y(n_5464)
);

BUFx12f_ASAP7_75t_L g5465 ( 
.A(n_5248),
.Y(n_5465)
);

BUFx2_ASAP7_75t_L g5466 ( 
.A(n_5153),
.Y(n_5466)
);

INVx1_ASAP7_75t_SL g5467 ( 
.A(n_5379),
.Y(n_5467)
);

INVx6_ASAP7_75t_L g5468 ( 
.A(n_5144),
.Y(n_5468)
);

INVx1_ASAP7_75t_L g5469 ( 
.A(n_5177),
.Y(n_5469)
);

CKINVDCx20_ASAP7_75t_R g5470 ( 
.A(n_5333),
.Y(n_5470)
);

BUFx2_ASAP7_75t_L g5471 ( 
.A(n_5144),
.Y(n_5471)
);

BUFx6f_ASAP7_75t_L g5472 ( 
.A(n_5332),
.Y(n_5472)
);

AND2x2_ASAP7_75t_L g5473 ( 
.A(n_5092),
.B(n_4621),
.Y(n_5473)
);

BUFx2_ASAP7_75t_SL g5474 ( 
.A(n_5341),
.Y(n_5474)
);

NAND2xp5_ASAP7_75t_L g5475 ( 
.A(n_5234),
.B(n_4926),
.Y(n_5475)
);

INVx6_ASAP7_75t_L g5476 ( 
.A(n_5144),
.Y(n_5476)
);

INVx1_ASAP7_75t_L g5477 ( 
.A(n_5215),
.Y(n_5477)
);

BUFx12f_ASAP7_75t_L g5478 ( 
.A(n_5248),
.Y(n_5478)
);

NOR2xp33_ASAP7_75t_L g5479 ( 
.A(n_5350),
.B(n_5050),
.Y(n_5479)
);

CKINVDCx5p33_ASAP7_75t_R g5480 ( 
.A(n_5355),
.Y(n_5480)
);

BUFx6f_ASAP7_75t_L g5481 ( 
.A(n_5373),
.Y(n_5481)
);

INVx2_ASAP7_75t_SL g5482 ( 
.A(n_5155),
.Y(n_5482)
);

INVx2_ASAP7_75t_L g5483 ( 
.A(n_5251),
.Y(n_5483)
);

NOR2xp33_ASAP7_75t_L g5484 ( 
.A(n_5206),
.B(n_4788),
.Y(n_5484)
);

BUFx3_ASAP7_75t_L g5485 ( 
.A(n_5132),
.Y(n_5485)
);

BUFx2_ASAP7_75t_L g5486 ( 
.A(n_5289),
.Y(n_5486)
);

NAND2x1p5_ASAP7_75t_L g5487 ( 
.A(n_5190),
.B(n_4887),
.Y(n_5487)
);

BUFx4f_ASAP7_75t_SL g5488 ( 
.A(n_5385),
.Y(n_5488)
);

BUFx12f_ASAP7_75t_L g5489 ( 
.A(n_5190),
.Y(n_5489)
);

AOI22xp5_ASAP7_75t_L g5490 ( 
.A1(n_5263),
.A2(n_5348),
.B1(n_5225),
.B2(n_5259),
.Y(n_5490)
);

INVx2_ASAP7_75t_L g5491 ( 
.A(n_5287),
.Y(n_5491)
);

BUFx12f_ASAP7_75t_L g5492 ( 
.A(n_5277),
.Y(n_5492)
);

CKINVDCx5p33_ASAP7_75t_R g5493 ( 
.A(n_5385),
.Y(n_5493)
);

BUFx12f_ASAP7_75t_L g5494 ( 
.A(n_5277),
.Y(n_5494)
);

CKINVDCx16_ASAP7_75t_R g5495 ( 
.A(n_5282),
.Y(n_5495)
);

INVx1_ASAP7_75t_L g5496 ( 
.A(n_5101),
.Y(n_5496)
);

BUFx4f_ASAP7_75t_SL g5497 ( 
.A(n_5361),
.Y(n_5497)
);

INVx5_ASAP7_75t_L g5498 ( 
.A(n_5264),
.Y(n_5498)
);

INVx1_ASAP7_75t_L g5499 ( 
.A(n_5136),
.Y(n_5499)
);

BUFx12f_ASAP7_75t_L g5500 ( 
.A(n_5284),
.Y(n_5500)
);

BUFx2_ASAP7_75t_SL g5501 ( 
.A(n_5264),
.Y(n_5501)
);

BUFx3_ASAP7_75t_L g5502 ( 
.A(n_5212),
.Y(n_5502)
);

INVx8_ASAP7_75t_L g5503 ( 
.A(n_5264),
.Y(n_5503)
);

INVx2_ASAP7_75t_SL g5504 ( 
.A(n_5134),
.Y(n_5504)
);

INVx2_ASAP7_75t_SL g5505 ( 
.A(n_5244),
.Y(n_5505)
);

CKINVDCx5p33_ASAP7_75t_R g5506 ( 
.A(n_5210),
.Y(n_5506)
);

BUFx4_ASAP7_75t_SL g5507 ( 
.A(n_5266),
.Y(n_5507)
);

CKINVDCx5p33_ASAP7_75t_R g5508 ( 
.A(n_5322),
.Y(n_5508)
);

CKINVDCx20_ASAP7_75t_R g5509 ( 
.A(n_5291),
.Y(n_5509)
);

BUFx8_ASAP7_75t_SL g5510 ( 
.A(n_5306),
.Y(n_5510)
);

INVx3_ASAP7_75t_SL g5511 ( 
.A(n_5122),
.Y(n_5511)
);

BUFx3_ASAP7_75t_L g5512 ( 
.A(n_5246),
.Y(n_5512)
);

INVx3_ASAP7_75t_SL g5513 ( 
.A(n_5122),
.Y(n_5513)
);

NAND2x1p5_ASAP7_75t_L g5514 ( 
.A(n_5304),
.B(n_4888),
.Y(n_5514)
);

CKINVDCx20_ASAP7_75t_R g5515 ( 
.A(n_5360),
.Y(n_5515)
);

BUFx3_ASAP7_75t_L g5516 ( 
.A(n_5260),
.Y(n_5516)
);

NAND2x1p5_ASAP7_75t_L g5517 ( 
.A(n_5239),
.B(n_5041),
.Y(n_5517)
);

NAND2xp5_ASAP7_75t_L g5518 ( 
.A(n_5315),
.B(n_4862),
.Y(n_5518)
);

AND2x4_ASAP7_75t_L g5519 ( 
.A(n_5270),
.B(n_4965),
.Y(n_5519)
);

BUFx12f_ASAP7_75t_L g5520 ( 
.A(n_5331),
.Y(n_5520)
);

INVx1_ASAP7_75t_SL g5521 ( 
.A(n_5170),
.Y(n_5521)
);

INVx2_ASAP7_75t_SL g5522 ( 
.A(n_5336),
.Y(n_5522)
);

BUFx12f_ASAP7_75t_L g5523 ( 
.A(n_5331),
.Y(n_5523)
);

CKINVDCx14_ASAP7_75t_R g5524 ( 
.A(n_5353),
.Y(n_5524)
);

BUFx6f_ASAP7_75t_L g5525 ( 
.A(n_5336),
.Y(n_5525)
);

INVx2_ASAP7_75t_L g5526 ( 
.A(n_5122),
.Y(n_5526)
);

CKINVDCx5p33_ASAP7_75t_R g5527 ( 
.A(n_5261),
.Y(n_5527)
);

INVx1_ASAP7_75t_SL g5528 ( 
.A(n_5163),
.Y(n_5528)
);

INVx3_ASAP7_75t_L g5529 ( 
.A(n_5121),
.Y(n_5529)
);

INVx1_ASAP7_75t_SL g5530 ( 
.A(n_5313),
.Y(n_5530)
);

INVx1_ASAP7_75t_L g5531 ( 
.A(n_5139),
.Y(n_5531)
);

AND2x2_ASAP7_75t_L g5532 ( 
.A(n_5270),
.B(n_4621),
.Y(n_5532)
);

BUFx3_ASAP7_75t_L g5533 ( 
.A(n_5122),
.Y(n_5533)
);

BUFx12f_ASAP7_75t_L g5534 ( 
.A(n_5336),
.Y(n_5534)
);

CKINVDCx5p33_ASAP7_75t_R g5535 ( 
.A(n_5201),
.Y(n_5535)
);

NAND2xp5_ASAP7_75t_L g5536 ( 
.A(n_5078),
.B(n_4863),
.Y(n_5536)
);

INVx3_ASAP7_75t_L g5537 ( 
.A(n_5281),
.Y(n_5537)
);

INVx2_ASAP7_75t_SL g5538 ( 
.A(n_5381),
.Y(n_5538)
);

BUFx6f_ASAP7_75t_L g5539 ( 
.A(n_5185),
.Y(n_5539)
);

NAND2x1p5_ASAP7_75t_L g5540 ( 
.A(n_5318),
.B(n_4764),
.Y(n_5540)
);

BUFx6f_ASAP7_75t_L g5541 ( 
.A(n_5185),
.Y(n_5541)
);

NAND2xp5_ASAP7_75t_L g5542 ( 
.A(n_5111),
.B(n_4866),
.Y(n_5542)
);

INVx2_ASAP7_75t_SL g5543 ( 
.A(n_5368),
.Y(n_5543)
);

BUFx3_ASAP7_75t_L g5544 ( 
.A(n_5143),
.Y(n_5544)
);

NOR2xp33_ASAP7_75t_L g5545 ( 
.A(n_5362),
.B(n_4907),
.Y(n_5545)
);

BUFx4_ASAP7_75t_SL g5546 ( 
.A(n_5220),
.Y(n_5546)
);

BUFx12f_ASAP7_75t_L g5547 ( 
.A(n_5320),
.Y(n_5547)
);

INVx3_ASAP7_75t_L g5548 ( 
.A(n_5142),
.Y(n_5548)
);

INVx6_ASAP7_75t_L g5549 ( 
.A(n_5152),
.Y(n_5549)
);

INVx1_ASAP7_75t_SL g5550 ( 
.A(n_5250),
.Y(n_5550)
);

BUFx3_ASAP7_75t_L g5551 ( 
.A(n_5147),
.Y(n_5551)
);

INVx1_ASAP7_75t_L g5552 ( 
.A(n_5154),
.Y(n_5552)
);

BUFx2_ASAP7_75t_L g5553 ( 
.A(n_5387),
.Y(n_5553)
);

INVx1_ASAP7_75t_L g5554 ( 
.A(n_5161),
.Y(n_5554)
);

BUFx2_ASAP7_75t_SL g5555 ( 
.A(n_5300),
.Y(n_5555)
);

AOI22xp33_ASAP7_75t_SL g5556 ( 
.A1(n_5338),
.A2(n_4974),
.B1(n_4937),
.B2(n_4942),
.Y(n_5556)
);

BUFx8_ASAP7_75t_L g5557 ( 
.A(n_5364),
.Y(n_5557)
);

BUFx6f_ASAP7_75t_L g5558 ( 
.A(n_5386),
.Y(n_5558)
);

INVx4_ASAP7_75t_L g5559 ( 
.A(n_5228),
.Y(n_5559)
);

AND2x2_ASAP7_75t_L g5560 ( 
.A(n_5107),
.B(n_4915),
.Y(n_5560)
);

INVx1_ASAP7_75t_SL g5561 ( 
.A(n_5334),
.Y(n_5561)
);

AND2x2_ASAP7_75t_L g5562 ( 
.A(n_5145),
.B(n_5061),
.Y(n_5562)
);

CKINVDCx5p33_ASAP7_75t_R g5563 ( 
.A(n_5316),
.Y(n_5563)
);

INVx1_ASAP7_75t_L g5564 ( 
.A(n_5164),
.Y(n_5564)
);

INVx2_ASAP7_75t_SL g5565 ( 
.A(n_5100),
.Y(n_5565)
);

CKINVDCx5p33_ASAP7_75t_R g5566 ( 
.A(n_5351),
.Y(n_5566)
);

INVx1_ASAP7_75t_L g5567 ( 
.A(n_5165),
.Y(n_5567)
);

INVx4_ASAP7_75t_L g5568 ( 
.A(n_5135),
.Y(n_5568)
);

AND2x2_ASAP7_75t_L g5569 ( 
.A(n_5128),
.B(n_5061),
.Y(n_5569)
);

BUFx3_ASAP7_75t_L g5570 ( 
.A(n_5166),
.Y(n_5570)
);

INVxp67_ASAP7_75t_SL g5571 ( 
.A(n_5096),
.Y(n_5571)
);

INVx3_ASAP7_75t_SL g5572 ( 
.A(n_5178),
.Y(n_5572)
);

CKINVDCx20_ASAP7_75t_R g5573 ( 
.A(n_5390),
.Y(n_5573)
);

HB1xp67_ASAP7_75t_L g5574 ( 
.A(n_5128),
.Y(n_5574)
);

BUFx3_ASAP7_75t_L g5575 ( 
.A(n_5173),
.Y(n_5575)
);

BUFx6f_ASAP7_75t_L g5576 ( 
.A(n_5116),
.Y(n_5576)
);

INVx5_ASAP7_75t_L g5577 ( 
.A(n_5150),
.Y(n_5577)
);

NOR2x1_ASAP7_75t_L g5578 ( 
.A(n_5168),
.B(n_4647),
.Y(n_5578)
);

NAND2x1p5_ASAP7_75t_L g5579 ( 
.A(n_5227),
.B(n_4988),
.Y(n_5579)
);

BUFx3_ASAP7_75t_L g5580 ( 
.A(n_5231),
.Y(n_5580)
);

BUFx2_ASAP7_75t_SL g5581 ( 
.A(n_5366),
.Y(n_5581)
);

BUFx6f_ASAP7_75t_L g5582 ( 
.A(n_5233),
.Y(n_5582)
);

CKINVDCx16_ASAP7_75t_R g5583 ( 
.A(n_5249),
.Y(n_5583)
);

BUFx6f_ASAP7_75t_L g5584 ( 
.A(n_5216),
.Y(n_5584)
);

INVx1_ASAP7_75t_L g5585 ( 
.A(n_5191),
.Y(n_5585)
);

INVx1_ASAP7_75t_SL g5586 ( 
.A(n_5198),
.Y(n_5586)
);

INVx8_ASAP7_75t_L g5587 ( 
.A(n_5296),
.Y(n_5587)
);

CKINVDCx5p33_ASAP7_75t_R g5588 ( 
.A(n_5330),
.Y(n_5588)
);

HB1xp67_ASAP7_75t_L g5589 ( 
.A(n_5172),
.Y(n_5589)
);

OAI21x1_ASAP7_75t_L g5590 ( 
.A1(n_5402),
.A2(n_5138),
.B(n_5077),
.Y(n_5590)
);

AOI22xp33_ASAP7_75t_L g5591 ( 
.A1(n_5587),
.A2(n_5274),
.B1(n_5176),
.B2(n_5207),
.Y(n_5591)
);

NAND2xp5_ASAP7_75t_L g5592 ( 
.A(n_5457),
.B(n_5217),
.Y(n_5592)
);

AOI221xp5_ASAP7_75t_L g5593 ( 
.A1(n_5490),
.A2(n_5243),
.B1(n_5253),
.B2(n_5337),
.C(n_5391),
.Y(n_5593)
);

BUFx12f_ASAP7_75t_L g5594 ( 
.A(n_5397),
.Y(n_5594)
);

INVx2_ASAP7_75t_L g5595 ( 
.A(n_5553),
.Y(n_5595)
);

AND2x2_ASAP7_75t_L g5596 ( 
.A(n_5451),
.B(n_5104),
.Y(n_5596)
);

INVx3_ASAP7_75t_L g5597 ( 
.A(n_5399),
.Y(n_5597)
);

INVx1_ASAP7_75t_L g5598 ( 
.A(n_5414),
.Y(n_5598)
);

HB1xp67_ASAP7_75t_L g5599 ( 
.A(n_5410),
.Y(n_5599)
);

AND2x2_ASAP7_75t_L g5600 ( 
.A(n_5449),
.B(n_5485),
.Y(n_5600)
);

OAI21x1_ASAP7_75t_L g5601 ( 
.A1(n_5548),
.A2(n_5181),
.B(n_5089),
.Y(n_5601)
);

INVx2_ASAP7_75t_L g5602 ( 
.A(n_5454),
.Y(n_5602)
);

INVx1_ASAP7_75t_L g5603 ( 
.A(n_5405),
.Y(n_5603)
);

NOR2x1_ASAP7_75t_SL g5604 ( 
.A(n_5465),
.B(n_5146),
.Y(n_5604)
);

INVx1_ASAP7_75t_L g5605 ( 
.A(n_5408),
.Y(n_5605)
);

INVx1_ASAP7_75t_L g5606 ( 
.A(n_5409),
.Y(n_5606)
);

OAI21x1_ASAP7_75t_L g5607 ( 
.A1(n_5442),
.A2(n_5130),
.B(n_5099),
.Y(n_5607)
);

CKINVDCx11_ASAP7_75t_R g5608 ( 
.A(n_5445),
.Y(n_5608)
);

OAI22xp5_ASAP7_75t_L g5609 ( 
.A1(n_5478),
.A2(n_5115),
.B1(n_5186),
.B2(n_5174),
.Y(n_5609)
);

NOR4xp25_ASAP7_75t_L g5610 ( 
.A(n_5550),
.B(n_5352),
.C(n_5194),
.D(n_5195),
.Y(n_5610)
);

INVx1_ASAP7_75t_SL g5611 ( 
.A(n_5497),
.Y(n_5611)
);

AOI21xp5_ASAP7_75t_L g5612 ( 
.A1(n_5587),
.A2(n_5141),
.B(n_5184),
.Y(n_5612)
);

OAI22xp5_ASAP7_75t_L g5613 ( 
.A1(n_5524),
.A2(n_5169),
.B1(n_5082),
.B2(n_5091),
.Y(n_5613)
);

AOI22xp33_ASAP7_75t_L g5614 ( 
.A1(n_5549),
.A2(n_5319),
.B1(n_5175),
.B2(n_5285),
.Y(n_5614)
);

INVx2_ASAP7_75t_L g5615 ( 
.A(n_5453),
.Y(n_5615)
);

BUFx2_ASAP7_75t_SL g5616 ( 
.A(n_5577),
.Y(n_5616)
);

AO21x2_ASAP7_75t_L g5617 ( 
.A1(n_5574),
.A2(n_5193),
.B(n_5200),
.Y(n_5617)
);

OA21x2_ASAP7_75t_L g5618 ( 
.A1(n_5571),
.A2(n_5131),
.B(n_5160),
.Y(n_5618)
);

OAI21x1_ASAP7_75t_L g5619 ( 
.A1(n_5462),
.A2(n_5137),
.B(n_5271),
.Y(n_5619)
);

OAI21xp5_ASAP7_75t_L g5620 ( 
.A1(n_5517),
.A2(n_5297),
.B(n_5377),
.Y(n_5620)
);

OA21x2_ASAP7_75t_L g5621 ( 
.A1(n_5589),
.A2(n_5095),
.B(n_5106),
.Y(n_5621)
);

BUFx2_ASAP7_75t_L g5622 ( 
.A(n_5471),
.Y(n_5622)
);

HB1xp67_ASAP7_75t_L g5623 ( 
.A(n_5432),
.Y(n_5623)
);

BUFx12f_ASAP7_75t_L g5624 ( 
.A(n_5428),
.Y(n_5624)
);

AND2x4_ASAP7_75t_L g5625 ( 
.A(n_5419),
.B(n_5140),
.Y(n_5625)
);

OAI21xp5_ASAP7_75t_L g5626 ( 
.A1(n_5556),
.A2(n_5276),
.B(n_5335),
.Y(n_5626)
);

AND2x2_ASAP7_75t_L g5627 ( 
.A(n_5504),
.B(n_5187),
.Y(n_5627)
);

INVx2_ASAP7_75t_L g5628 ( 
.A(n_5458),
.Y(n_5628)
);

OAI21x1_ASAP7_75t_L g5629 ( 
.A1(n_5537),
.A2(n_5321),
.B(n_5343),
.Y(n_5629)
);

AND2x4_ASAP7_75t_L g5630 ( 
.A(n_5569),
.B(n_5159),
.Y(n_5630)
);

O2A1O1Ixp33_ASAP7_75t_SL g5631 ( 
.A1(n_5455),
.A2(n_5301),
.B(n_5327),
.C(n_5394),
.Y(n_5631)
);

INVx1_ASAP7_75t_L g5632 ( 
.A(n_5412),
.Y(n_5632)
);

OR2x6_ASAP7_75t_L g5633 ( 
.A(n_5464),
.B(n_5474),
.Y(n_5633)
);

INVx3_ASAP7_75t_L g5634 ( 
.A(n_5488),
.Y(n_5634)
);

AOI211xp5_ASAP7_75t_L g5635 ( 
.A1(n_5529),
.A2(n_5359),
.B(n_5245),
.C(n_5272),
.Y(n_5635)
);

AO21x2_ASAP7_75t_L g5636 ( 
.A1(n_5403),
.A2(n_5438),
.B(n_5418),
.Y(n_5636)
);

NAND2xp5_ASAP7_75t_L g5637 ( 
.A(n_5473),
.B(n_5204),
.Y(n_5637)
);

OAI221xp5_ASAP7_75t_L g5638 ( 
.A1(n_5435),
.A2(n_5375),
.B1(n_5097),
.B2(n_5093),
.C(n_5126),
.Y(n_5638)
);

INVx3_ASAP7_75t_L g5639 ( 
.A(n_5398),
.Y(n_5639)
);

OAI21x1_ASAP7_75t_L g5640 ( 
.A1(n_5578),
.A2(n_5460),
.B(n_5526),
.Y(n_5640)
);

OAI21x1_ASAP7_75t_L g5641 ( 
.A1(n_5532),
.A2(n_5229),
.B(n_5392),
.Y(n_5641)
);

AO31x2_ASAP7_75t_L g5642 ( 
.A1(n_5568),
.A2(n_5108),
.A3(n_5114),
.B(n_5209),
.Y(n_5642)
);

AOI21xp33_ASAP7_75t_L g5643 ( 
.A1(n_5547),
.A2(n_5376),
.B(n_5369),
.Y(n_5643)
);

NAND2xp5_ASAP7_75t_L g5644 ( 
.A(n_5406),
.B(n_5221),
.Y(n_5644)
);

INVx1_ASAP7_75t_L g5645 ( 
.A(n_5439),
.Y(n_5645)
);

OA21x2_ASAP7_75t_L g5646 ( 
.A1(n_5426),
.A2(n_5247),
.B(n_5230),
.Y(n_5646)
);

NAND2xp5_ASAP7_75t_L g5647 ( 
.A(n_5415),
.B(n_5256),
.Y(n_5647)
);

AO21x2_ASAP7_75t_L g5648 ( 
.A1(n_5518),
.A2(n_5183),
.B(n_5345),
.Y(n_5648)
);

OR2x6_ASAP7_75t_L g5649 ( 
.A(n_5503),
.B(n_5213),
.Y(n_5649)
);

OR2x2_ASAP7_75t_L g5650 ( 
.A(n_5459),
.B(n_5257),
.Y(n_5650)
);

AOI22xp33_ASAP7_75t_L g5651 ( 
.A1(n_5555),
.A2(n_5393),
.B1(n_5292),
.B2(n_5283),
.Y(n_5651)
);

INVx2_ASAP7_75t_L g5652 ( 
.A(n_5483),
.Y(n_5652)
);

INVx1_ASAP7_75t_L g5653 ( 
.A(n_5444),
.Y(n_5653)
);

OAI21x1_ASAP7_75t_L g5654 ( 
.A1(n_5487),
.A2(n_5326),
.B(n_5323),
.Y(n_5654)
);

NAND2xp5_ASAP7_75t_L g5655 ( 
.A(n_5496),
.B(n_5278),
.Y(n_5655)
);

INVx1_ASAP7_75t_L g5656 ( 
.A(n_5446),
.Y(n_5656)
);

AOI21x1_ASAP7_75t_L g5657 ( 
.A1(n_5486),
.A2(n_5372),
.B(n_5370),
.Y(n_5657)
);

AND2x2_ASAP7_75t_SL g5658 ( 
.A(n_5466),
.B(n_5187),
.Y(n_5658)
);

NOR2xp33_ASAP7_75t_L g5659 ( 
.A(n_5427),
.B(n_5074),
.Y(n_5659)
);

OAI21x1_ASAP7_75t_L g5660 ( 
.A1(n_5514),
.A2(n_5374),
.B(n_5199),
.Y(n_5660)
);

INVx1_ASAP7_75t_SL g5661 ( 
.A(n_5467),
.Y(n_5661)
);

AO21x2_ASAP7_75t_L g5662 ( 
.A1(n_5461),
.A2(n_5286),
.B(n_5279),
.Y(n_5662)
);

INVx4_ASAP7_75t_L g5663 ( 
.A(n_5401),
.Y(n_5663)
);

BUFx6f_ASAP7_75t_L g5664 ( 
.A(n_5534),
.Y(n_5664)
);

AOI22xp33_ASAP7_75t_L g5665 ( 
.A1(n_5581),
.A2(n_5314),
.B1(n_5298),
.B2(n_5205),
.Y(n_5665)
);

O2A1O1Ixp33_ASAP7_75t_SL g5666 ( 
.A1(n_5404),
.A2(n_5342),
.B(n_5035),
.C(n_5006),
.Y(n_5666)
);

AOI21xp5_ASAP7_75t_L g5667 ( 
.A1(n_5437),
.A2(n_5325),
.B(n_5085),
.Y(n_5667)
);

AO21x1_ASAP7_75t_L g5668 ( 
.A1(n_5559),
.A2(n_5236),
.B(n_5219),
.Y(n_5668)
);

AND2x2_ASAP7_75t_L g5669 ( 
.A(n_5456),
.B(n_5061),
.Y(n_5669)
);

OAI21x1_ASAP7_75t_L g5670 ( 
.A1(n_5400),
.A2(n_5346),
.B(n_5218),
.Y(n_5670)
);

BUFx3_ASAP7_75t_L g5671 ( 
.A(n_5416),
.Y(n_5671)
);

A2O1A1Ixp33_ASAP7_75t_L g5672 ( 
.A1(n_5535),
.A2(n_5307),
.B(n_5288),
.C(n_5211),
.Y(n_5672)
);

NAND2x1p5_ASAP7_75t_L g5673 ( 
.A(n_5577),
.B(n_5340),
.Y(n_5673)
);

INVx2_ASAP7_75t_L g5674 ( 
.A(n_5491),
.Y(n_5674)
);

OAI21x1_ASAP7_75t_L g5675 ( 
.A1(n_5562),
.A2(n_5133),
.B(n_5317),
.Y(n_5675)
);

AND2x2_ASAP7_75t_L g5676 ( 
.A(n_5495),
.B(n_5295),
.Y(n_5676)
);

OAI22xp33_ASAP7_75t_L g5677 ( 
.A1(n_5583),
.A2(n_4929),
.B1(n_4954),
.B2(n_4875),
.Y(n_5677)
);

AO21x2_ASAP7_75t_L g5678 ( 
.A1(n_5475),
.A2(n_5567),
.B(n_5564),
.Y(n_5678)
);

INVx1_ASAP7_75t_L g5679 ( 
.A(n_5452),
.Y(n_5679)
);

OA21x2_ASAP7_75t_L g5680 ( 
.A1(n_5411),
.A2(n_5305),
.B(n_5299),
.Y(n_5680)
);

BUFx3_ASAP7_75t_L g5681 ( 
.A(n_5421),
.Y(n_5681)
);

BUFx4f_ASAP7_75t_SL g5682 ( 
.A(n_5420),
.Y(n_5682)
);

OAI21x1_ASAP7_75t_L g5683 ( 
.A1(n_5579),
.A2(n_5378),
.B(n_5309),
.Y(n_5683)
);

CKINVDCx16_ASAP7_75t_R g5684 ( 
.A(n_5431),
.Y(n_5684)
);

OAI21xp5_ASAP7_75t_L g5685 ( 
.A1(n_5527),
.A2(n_5197),
.B(n_5382),
.Y(n_5685)
);

OAI21x1_ASAP7_75t_L g5686 ( 
.A1(n_5540),
.A2(n_5308),
.B(n_5268),
.Y(n_5686)
);

NOR2xp33_ASAP7_75t_L g5687 ( 
.A(n_5425),
.B(n_4895),
.Y(n_5687)
);

OR2x2_ASAP7_75t_L g5688 ( 
.A(n_5499),
.B(n_5016),
.Y(n_5688)
);

CKINVDCx16_ASAP7_75t_R g5689 ( 
.A(n_5421),
.Y(n_5689)
);

OAI21x1_ASAP7_75t_L g5690 ( 
.A1(n_5469),
.A2(n_5384),
.B(n_5356),
.Y(n_5690)
);

AO21x2_ASAP7_75t_L g5691 ( 
.A1(n_5585),
.A2(n_5124),
.B(n_4668),
.Y(n_5691)
);

O2A1O1Ixp33_ASAP7_75t_L g5692 ( 
.A1(n_5586),
.A2(n_5561),
.B(n_5413),
.C(n_5434),
.Y(n_5692)
);

A2O1A1Ixp33_ASAP7_75t_SL g5693 ( 
.A1(n_5450),
.A2(n_5396),
.B(n_5018),
.C(n_5367),
.Y(n_5693)
);

BUFx2_ASAP7_75t_L g5694 ( 
.A(n_5557),
.Y(n_5694)
);

CKINVDCx5p33_ASAP7_75t_R g5695 ( 
.A(n_5443),
.Y(n_5695)
);

A2O1A1Ixp33_ASAP7_75t_L g5696 ( 
.A1(n_5588),
.A2(n_5422),
.B(n_5407),
.C(n_5463),
.Y(n_5696)
);

OAI21x1_ASAP7_75t_L g5697 ( 
.A1(n_5477),
.A2(n_5203),
.B(n_5328),
.Y(n_5697)
);

OAI22xp33_ASAP7_75t_L g5698 ( 
.A1(n_5489),
.A2(n_5171),
.B1(n_5238),
.B2(n_4720),
.Y(n_5698)
);

OAI21x1_ASAP7_75t_SL g5699 ( 
.A1(n_5482),
.A2(n_5347),
.B(n_5252),
.Y(n_5699)
);

BUFx3_ASAP7_75t_L g5700 ( 
.A(n_5448),
.Y(n_5700)
);

AOI22xp33_ASAP7_75t_SL g5701 ( 
.A1(n_5447),
.A2(n_5237),
.B1(n_5354),
.B2(n_4821),
.Y(n_5701)
);

INVx1_ASAP7_75t_L g5702 ( 
.A(n_5531),
.Y(n_5702)
);

NAND2x1p5_ASAP7_75t_L g5703 ( 
.A(n_5498),
.B(n_5525),
.Y(n_5703)
);

OAI21x1_ASAP7_75t_L g5704 ( 
.A1(n_5546),
.A2(n_5440),
.B(n_5552),
.Y(n_5704)
);

AND2x4_ASAP7_75t_L g5705 ( 
.A(n_5519),
.B(n_5188),
.Y(n_5705)
);

OR2x6_ASAP7_75t_L g5706 ( 
.A(n_5503),
.B(n_5501),
.Y(n_5706)
);

BUFx3_ASAP7_75t_L g5707 ( 
.A(n_5493),
.Y(n_5707)
);

AND2x4_ASAP7_75t_L g5708 ( 
.A(n_5502),
.B(n_5512),
.Y(n_5708)
);

NAND2xp5_ASAP7_75t_L g5709 ( 
.A(n_5554),
.B(n_5542),
.Y(n_5709)
);

OAI21xp5_ASAP7_75t_L g5710 ( 
.A1(n_5515),
.A2(n_5484),
.B(n_5545),
.Y(n_5710)
);

INVx1_ASAP7_75t_L g5711 ( 
.A(n_5429),
.Y(n_5711)
);

INVx2_ASAP7_75t_L g5712 ( 
.A(n_5539),
.Y(n_5712)
);

INVx1_ASAP7_75t_SL g5713 ( 
.A(n_5509),
.Y(n_5713)
);

OAI21x1_ASAP7_75t_L g5714 ( 
.A1(n_5536),
.A2(n_5241),
.B(n_5349),
.Y(n_5714)
);

OAI21x1_ASAP7_75t_L g5715 ( 
.A1(n_5570),
.A2(n_5365),
.B(n_4676),
.Y(n_5715)
);

OAI211xp5_ASAP7_75t_SL g5716 ( 
.A1(n_5479),
.A2(n_5040),
.B(n_4879),
.C(n_4855),
.Y(n_5716)
);

OAI21x1_ASAP7_75t_L g5717 ( 
.A1(n_5551),
.A2(n_4693),
.B(n_4662),
.Y(n_5717)
);

OAI21x1_ASAP7_75t_L g5718 ( 
.A1(n_5447),
.A2(n_4709),
.B(n_4703),
.Y(n_5718)
);

BUFx3_ASAP7_75t_L g5719 ( 
.A(n_5470),
.Y(n_5719)
);

OAI21xp5_ASAP7_75t_L g5720 ( 
.A1(n_5573),
.A2(n_5383),
.B(n_5311),
.Y(n_5720)
);

OAI21x1_ASAP7_75t_L g5721 ( 
.A1(n_5447),
.A2(n_4717),
.B(n_4710),
.Y(n_5721)
);

AOI21xp5_ASAP7_75t_L g5722 ( 
.A1(n_5521),
.A2(n_5275),
.B(n_4843),
.Y(n_5722)
);

NOR2xp33_ASAP7_75t_L g5723 ( 
.A(n_5436),
.B(n_4896),
.Y(n_5723)
);

NAND2x1p5_ASAP7_75t_L g5724 ( 
.A(n_5498),
.B(n_5363),
.Y(n_5724)
);

INVx6_ASAP7_75t_L g5725 ( 
.A(n_5706),
.Y(n_5725)
);

BUFx3_ASAP7_75t_L g5726 ( 
.A(n_5694),
.Y(n_5726)
);

INVx2_ASAP7_75t_L g5727 ( 
.A(n_5623),
.Y(n_5727)
);

INVx1_ASAP7_75t_L g5728 ( 
.A(n_5599),
.Y(n_5728)
);

INVxp67_ASAP7_75t_L g5729 ( 
.A(n_5694),
.Y(n_5729)
);

AOI22xp33_ASAP7_75t_L g5730 ( 
.A1(n_5591),
.A2(n_5613),
.B1(n_5609),
.B2(n_5638),
.Y(n_5730)
);

INVx2_ASAP7_75t_L g5731 ( 
.A(n_5622),
.Y(n_5731)
);

INVx2_ASAP7_75t_L g5732 ( 
.A(n_5622),
.Y(n_5732)
);

AOI22xp33_ASAP7_75t_SL g5733 ( 
.A1(n_5616),
.A2(n_5447),
.B1(n_5494),
.B2(n_5492),
.Y(n_5733)
);

BUFx8_ASAP7_75t_L g5734 ( 
.A(n_5594),
.Y(n_5734)
);

INVx4_ASAP7_75t_L g5735 ( 
.A(n_5624),
.Y(n_5735)
);

INVx1_ASAP7_75t_L g5736 ( 
.A(n_5603),
.Y(n_5736)
);

INVx4_ASAP7_75t_L g5737 ( 
.A(n_5663),
.Y(n_5737)
);

INVx1_ASAP7_75t_L g5738 ( 
.A(n_5605),
.Y(n_5738)
);

AND2x2_ASAP7_75t_L g5739 ( 
.A(n_5600),
.B(n_5539),
.Y(n_5739)
);

AO21x2_ASAP7_75t_L g5740 ( 
.A1(n_5636),
.A2(n_4726),
.B(n_4725),
.Y(n_5740)
);

AOI21x1_ASAP7_75t_L g5741 ( 
.A1(n_5706),
.A2(n_5522),
.B(n_5560),
.Y(n_5741)
);

INVx2_ASAP7_75t_L g5742 ( 
.A(n_5595),
.Y(n_5742)
);

INVx4_ASAP7_75t_L g5743 ( 
.A(n_5682),
.Y(n_5743)
);

INVx6_ASAP7_75t_L g5744 ( 
.A(n_5684),
.Y(n_5744)
);

INVx1_ASAP7_75t_L g5745 ( 
.A(n_5606),
.Y(n_5745)
);

AND2x2_ASAP7_75t_L g5746 ( 
.A(n_5669),
.B(n_5541),
.Y(n_5746)
);

OAI22xp5_ASAP7_75t_L g5747 ( 
.A1(n_5616),
.A2(n_5572),
.B1(n_5508),
.B2(n_5476),
.Y(n_5747)
);

INVx1_ASAP7_75t_L g5748 ( 
.A(n_5632),
.Y(n_5748)
);

INVx3_ASAP7_75t_L g5749 ( 
.A(n_5671),
.Y(n_5749)
);

NOR2xp33_ASAP7_75t_L g5750 ( 
.A(n_5608),
.B(n_5430),
.Y(n_5750)
);

OAI21x1_ASAP7_75t_L g5751 ( 
.A1(n_5640),
.A2(n_5476),
.B(n_5423),
.Y(n_5751)
);

BUFx2_ASAP7_75t_R g5752 ( 
.A(n_5695),
.Y(n_5752)
);

INVx3_ASAP7_75t_L g5753 ( 
.A(n_5597),
.Y(n_5753)
);

INVx2_ASAP7_75t_L g5754 ( 
.A(n_5615),
.Y(n_5754)
);

AND2x4_ASAP7_75t_L g5755 ( 
.A(n_5708),
.B(n_5481),
.Y(n_5755)
);

INVx3_ASAP7_75t_L g5756 ( 
.A(n_5633),
.Y(n_5756)
);

INVx1_ASAP7_75t_L g5757 ( 
.A(n_5656),
.Y(n_5757)
);

OAI21xp5_ASAP7_75t_L g5758 ( 
.A1(n_5667),
.A2(n_5566),
.B(n_5506),
.Y(n_5758)
);

NOR2xp33_ASAP7_75t_L g5759 ( 
.A(n_5689),
.B(n_5417),
.Y(n_5759)
);

INVx6_ASAP7_75t_L g5760 ( 
.A(n_5664),
.Y(n_5760)
);

BUFx4_ASAP7_75t_R g5761 ( 
.A(n_5604),
.Y(n_5761)
);

NAND2xp5_ASAP7_75t_L g5762 ( 
.A(n_5592),
.B(n_5678),
.Y(n_5762)
);

INVx1_ASAP7_75t_L g5763 ( 
.A(n_5679),
.Y(n_5763)
);

BUFx2_ASAP7_75t_L g5764 ( 
.A(n_5639),
.Y(n_5764)
);

INVx3_ASAP7_75t_L g5765 ( 
.A(n_5633),
.Y(n_5765)
);

NAND2x1_ASAP7_75t_L g5766 ( 
.A(n_5625),
.B(n_5634),
.Y(n_5766)
);

INVx1_ASAP7_75t_L g5767 ( 
.A(n_5645),
.Y(n_5767)
);

INVx2_ASAP7_75t_SL g5768 ( 
.A(n_5664),
.Y(n_5768)
);

OAI22xp5_ASAP7_75t_L g5769 ( 
.A1(n_5713),
.A2(n_5513),
.B1(n_5511),
.B2(n_5520),
.Y(n_5769)
);

INVx2_ASAP7_75t_SL g5770 ( 
.A(n_5681),
.Y(n_5770)
);

INVx1_ASAP7_75t_L g5771 ( 
.A(n_5653),
.Y(n_5771)
);

INVx1_ASAP7_75t_L g5772 ( 
.A(n_5702),
.Y(n_5772)
);

INVx1_ASAP7_75t_L g5773 ( 
.A(n_5598),
.Y(n_5773)
);

BUFx2_ASAP7_75t_L g5774 ( 
.A(n_5703),
.Y(n_5774)
);

BUFx3_ASAP7_75t_L g5775 ( 
.A(n_5700),
.Y(n_5775)
);

OAI21xp5_ASAP7_75t_L g5776 ( 
.A1(n_5626),
.A2(n_5563),
.B(n_5565),
.Y(n_5776)
);

CKINVDCx5p33_ASAP7_75t_R g5777 ( 
.A(n_5719),
.Y(n_5777)
);

AOI22xp33_ASAP7_75t_L g5778 ( 
.A1(n_5701),
.A2(n_5523),
.B1(n_5580),
.B2(n_5582),
.Y(n_5778)
);

BUFx3_ASAP7_75t_L g5779 ( 
.A(n_5707),
.Y(n_5779)
);

INVx3_ASAP7_75t_L g5780 ( 
.A(n_5611),
.Y(n_5780)
);

BUFx6f_ASAP7_75t_L g5781 ( 
.A(n_5712),
.Y(n_5781)
);

CKINVDCx5p33_ASAP7_75t_R g5782 ( 
.A(n_5661),
.Y(n_5782)
);

AND2x2_ASAP7_75t_L g5783 ( 
.A(n_5602),
.B(n_5541),
.Y(n_5783)
);

INVx3_ASAP7_75t_L g5784 ( 
.A(n_5704),
.Y(n_5784)
);

OAI21x1_ASAP7_75t_L g5785 ( 
.A1(n_5601),
.A2(n_4732),
.B(n_4728),
.Y(n_5785)
);

INVx1_ASAP7_75t_L g5786 ( 
.A(n_5709),
.Y(n_5786)
);

OAI21x1_ASAP7_75t_L g5787 ( 
.A1(n_5590),
.A2(n_4745),
.B(n_4740),
.Y(n_5787)
);

INVx1_ASAP7_75t_L g5788 ( 
.A(n_5628),
.Y(n_5788)
);

INVx2_ASAP7_75t_L g5789 ( 
.A(n_5652),
.Y(n_5789)
);

HB1xp67_ASAP7_75t_SL g5790 ( 
.A(n_5659),
.Y(n_5790)
);

INVx6_ASAP7_75t_L g5791 ( 
.A(n_5649),
.Y(n_5791)
);

AOI22xp33_ASAP7_75t_L g5792 ( 
.A1(n_5685),
.A2(n_5584),
.B1(n_5582),
.B2(n_5500),
.Y(n_5792)
);

INVx1_ASAP7_75t_L g5793 ( 
.A(n_5674),
.Y(n_5793)
);

BUFx6f_ASAP7_75t_L g5794 ( 
.A(n_5670),
.Y(n_5794)
);

OAI21x1_ASAP7_75t_L g5795 ( 
.A1(n_5619),
.A2(n_4760),
.B(n_4749),
.Y(n_5795)
);

INVx1_ASAP7_75t_L g5796 ( 
.A(n_5650),
.Y(n_5796)
);

NAND2x1p5_ASAP7_75t_L g5797 ( 
.A(n_5654),
.B(n_5525),
.Y(n_5797)
);

INVx1_ASAP7_75t_L g5798 ( 
.A(n_5647),
.Y(n_5798)
);

INVx2_ASAP7_75t_L g5799 ( 
.A(n_5627),
.Y(n_5799)
);

INVx1_ASAP7_75t_L g5800 ( 
.A(n_5655),
.Y(n_5800)
);

AND2x2_ASAP7_75t_L g5801 ( 
.A(n_5711),
.B(n_5543),
.Y(n_5801)
);

INVx1_ASAP7_75t_L g5802 ( 
.A(n_5688),
.Y(n_5802)
);

INVx1_ASAP7_75t_L g5803 ( 
.A(n_5644),
.Y(n_5803)
);

INVx1_ASAP7_75t_L g5804 ( 
.A(n_5637),
.Y(n_5804)
);

BUFx2_ASAP7_75t_L g5805 ( 
.A(n_5696),
.Y(n_5805)
);

OAI22xp5_ASAP7_75t_L g5806 ( 
.A1(n_5649),
.A2(n_5468),
.B1(n_5528),
.B2(n_5481),
.Y(n_5806)
);

INVx2_ASAP7_75t_L g5807 ( 
.A(n_5697),
.Y(n_5807)
);

HB1xp67_ASAP7_75t_L g5808 ( 
.A(n_5596),
.Y(n_5808)
);

INVx2_ASAP7_75t_L g5809 ( 
.A(n_5618),
.Y(n_5809)
);

AOI22xp33_ASAP7_75t_SL g5810 ( 
.A1(n_5658),
.A2(n_5516),
.B1(n_5576),
.B2(n_5533),
.Y(n_5810)
);

AND2x4_ASAP7_75t_L g5811 ( 
.A(n_5705),
.B(n_5505),
.Y(n_5811)
);

AO21x1_ASAP7_75t_SL g5812 ( 
.A1(n_5651),
.A2(n_5507),
.B(n_5530),
.Y(n_5812)
);

AOI22xp33_ASAP7_75t_L g5813 ( 
.A1(n_5698),
.A2(n_5584),
.B1(n_5576),
.B2(n_5538),
.Y(n_5813)
);

OAI21xp5_ASAP7_75t_L g5814 ( 
.A1(n_5612),
.A2(n_4904),
.B(n_5262),
.Y(n_5814)
);

BUFx2_ASAP7_75t_L g5815 ( 
.A(n_5618),
.Y(n_5815)
);

INVx1_ASAP7_75t_L g5816 ( 
.A(n_5680),
.Y(n_5816)
);

INVx1_ASAP7_75t_L g5817 ( 
.A(n_5680),
.Y(n_5817)
);

AND2x2_ASAP7_75t_L g5818 ( 
.A(n_5676),
.B(n_5544),
.Y(n_5818)
);

AO21x1_ASAP7_75t_SL g5819 ( 
.A1(n_5665),
.A2(n_5510),
.B(n_5433),
.Y(n_5819)
);

INVx2_ASAP7_75t_L g5820 ( 
.A(n_5630),
.Y(n_5820)
);

HB1xp67_ASAP7_75t_SL g5821 ( 
.A(n_5687),
.Y(n_5821)
);

AND2x2_ASAP7_75t_L g5822 ( 
.A(n_5630),
.B(n_5558),
.Y(n_5822)
);

OR2x6_ASAP7_75t_L g5823 ( 
.A(n_5673),
.B(n_5424),
.Y(n_5823)
);

INVx1_ASAP7_75t_L g5824 ( 
.A(n_5662),
.Y(n_5824)
);

BUFx2_ASAP7_75t_L g5825 ( 
.A(n_5607),
.Y(n_5825)
);

AND2x2_ASAP7_75t_L g5826 ( 
.A(n_5675),
.B(n_5558),
.Y(n_5826)
);

INVx1_ASAP7_75t_L g5827 ( 
.A(n_5691),
.Y(n_5827)
);

INVx6_ASAP7_75t_L g5828 ( 
.A(n_5631),
.Y(n_5828)
);

BUFx2_ASAP7_75t_L g5829 ( 
.A(n_5710),
.Y(n_5829)
);

BUFx3_ASAP7_75t_L g5830 ( 
.A(n_5723),
.Y(n_5830)
);

OAI21xp5_ASAP7_75t_L g5831 ( 
.A1(n_5692),
.A2(n_5395),
.B(n_5388),
.Y(n_5831)
);

INVx1_ASAP7_75t_L g5832 ( 
.A(n_5646),
.Y(n_5832)
);

INVx1_ASAP7_75t_L g5833 ( 
.A(n_5646),
.Y(n_5833)
);

BUFx6f_ASAP7_75t_L g5834 ( 
.A(n_5660),
.Y(n_5834)
);

INVx1_ASAP7_75t_L g5835 ( 
.A(n_5690),
.Y(n_5835)
);

INVx1_ASAP7_75t_L g5836 ( 
.A(n_5617),
.Y(n_5836)
);

INVx1_ASAP7_75t_L g5837 ( 
.A(n_5683),
.Y(n_5837)
);

INVx1_ASAP7_75t_L g5838 ( 
.A(n_5642),
.Y(n_5838)
);

INVx3_ASAP7_75t_L g5839 ( 
.A(n_5724),
.Y(n_5839)
);

INVx3_ASAP7_75t_L g5840 ( 
.A(n_5657),
.Y(n_5840)
);

AOI22xp33_ASAP7_75t_L g5841 ( 
.A1(n_5668),
.A2(n_4722),
.B1(n_5389),
.B2(n_5575),
.Y(n_5841)
);

INVx1_ASAP7_75t_L g5842 ( 
.A(n_5642),
.Y(n_5842)
);

OAI21xp33_ASAP7_75t_L g5843 ( 
.A1(n_5614),
.A2(n_5480),
.B(n_4938),
.Y(n_5843)
);

AOI22xp33_ASAP7_75t_SL g5844 ( 
.A1(n_5699),
.A2(n_5424),
.B1(n_5433),
.B2(n_5441),
.Y(n_5844)
);

AOI21x1_ASAP7_75t_L g5845 ( 
.A1(n_5657),
.A2(n_4781),
.B(n_4772),
.Y(n_5845)
);

INVx2_ASAP7_75t_L g5846 ( 
.A(n_5621),
.Y(n_5846)
);

BUFx2_ASAP7_75t_L g5847 ( 
.A(n_5621),
.Y(n_5847)
);

INVx1_ASAP7_75t_L g5848 ( 
.A(n_5717),
.Y(n_5848)
);

INVx1_ASAP7_75t_L g5849 ( 
.A(n_5641),
.Y(n_5849)
);

INVx8_ASAP7_75t_L g5850 ( 
.A(n_5610),
.Y(n_5850)
);

CKINVDCx20_ASAP7_75t_R g5851 ( 
.A(n_5643),
.Y(n_5851)
);

HB1xp67_ASAP7_75t_L g5852 ( 
.A(n_5648),
.Y(n_5852)
);

INVx1_ASAP7_75t_L g5853 ( 
.A(n_5715),
.Y(n_5853)
);

INVx1_ASAP7_75t_SL g5854 ( 
.A(n_5722),
.Y(n_5854)
);

NAND2x1p5_ASAP7_75t_L g5855 ( 
.A(n_5686),
.B(n_5441),
.Y(n_5855)
);

INVx2_ASAP7_75t_L g5856 ( 
.A(n_5741),
.Y(n_5856)
);

INVx1_ASAP7_75t_L g5857 ( 
.A(n_5816),
.Y(n_5857)
);

AND2x2_ASAP7_75t_L g5858 ( 
.A(n_5822),
.B(n_5718),
.Y(n_5858)
);

OAI21x1_ASAP7_75t_L g5859 ( 
.A1(n_5766),
.A2(n_5751),
.B(n_5806),
.Y(n_5859)
);

INVx2_ASAP7_75t_L g5860 ( 
.A(n_5764),
.Y(n_5860)
);

INVx1_ASAP7_75t_L g5861 ( 
.A(n_5817),
.Y(n_5861)
);

INVx2_ASAP7_75t_L g5862 ( 
.A(n_5764),
.Y(n_5862)
);

INVx2_ASAP7_75t_L g5863 ( 
.A(n_5799),
.Y(n_5863)
);

INVx1_ASAP7_75t_L g5864 ( 
.A(n_5788),
.Y(n_5864)
);

INVx1_ASAP7_75t_L g5865 ( 
.A(n_5793),
.Y(n_5865)
);

INVx1_ASAP7_75t_L g5866 ( 
.A(n_5736),
.Y(n_5866)
);

INVx2_ASAP7_75t_L g5867 ( 
.A(n_5727),
.Y(n_5867)
);

OAI22xp5_ASAP7_75t_L g5868 ( 
.A1(n_5828),
.A2(n_5593),
.B1(n_5672),
.B2(n_5620),
.Y(n_5868)
);

INVx1_ASAP7_75t_L g5869 ( 
.A(n_5838),
.Y(n_5869)
);

OA21x2_ASAP7_75t_L g5870 ( 
.A1(n_5842),
.A2(n_5629),
.B(n_5714),
.Y(n_5870)
);

INVx1_ASAP7_75t_L g5871 ( 
.A(n_5796),
.Y(n_5871)
);

INVx2_ASAP7_75t_L g5872 ( 
.A(n_5754),
.Y(n_5872)
);

OAI21x1_ASAP7_75t_L g5873 ( 
.A1(n_5747),
.A2(n_5721),
.B(n_5699),
.Y(n_5873)
);

AOI22xp33_ASAP7_75t_SL g5874 ( 
.A1(n_5828),
.A2(n_5720),
.B1(n_5472),
.B2(n_5031),
.Y(n_5874)
);

INVx1_ASAP7_75t_L g5875 ( 
.A(n_5738),
.Y(n_5875)
);

INVx1_ASAP7_75t_L g5876 ( 
.A(n_5745),
.Y(n_5876)
);

NAND2xp5_ASAP7_75t_L g5877 ( 
.A(n_5854),
.B(n_5635),
.Y(n_5877)
);

AND2x2_ASAP7_75t_L g5878 ( 
.A(n_5746),
.B(n_5472),
.Y(n_5878)
);

INVx1_ASAP7_75t_L g5879 ( 
.A(n_5748),
.Y(n_5879)
);

OAI22xp5_ASAP7_75t_L g5880 ( 
.A1(n_5725),
.A2(n_5677),
.B1(n_4897),
.B2(n_4868),
.Y(n_5880)
);

OR2x2_ASAP7_75t_L g5881 ( 
.A(n_5786),
.B(n_5226),
.Y(n_5881)
);

INVx1_ASAP7_75t_L g5882 ( 
.A(n_5757),
.Y(n_5882)
);

CKINVDCx5p33_ASAP7_75t_R g5883 ( 
.A(n_5734),
.Y(n_5883)
);

BUFx6f_ASAP7_75t_L g5884 ( 
.A(n_5743),
.Y(n_5884)
);

AND2x2_ASAP7_75t_L g5885 ( 
.A(n_5811),
.B(n_5202),
.Y(n_5885)
);

AO21x2_ASAP7_75t_L g5886 ( 
.A1(n_5852),
.A2(n_4786),
.B(n_4782),
.Y(n_5886)
);

INVx2_ASAP7_75t_L g5887 ( 
.A(n_5789),
.Y(n_5887)
);

AND2x2_ASAP7_75t_L g5888 ( 
.A(n_5818),
.B(n_5739),
.Y(n_5888)
);

INVx2_ASAP7_75t_L g5889 ( 
.A(n_5731),
.Y(n_5889)
);

INVx1_ASAP7_75t_L g5890 ( 
.A(n_5763),
.Y(n_5890)
);

INVx1_ASAP7_75t_L g5891 ( 
.A(n_5767),
.Y(n_5891)
);

INVx2_ASAP7_75t_SL g5892 ( 
.A(n_5744),
.Y(n_5892)
);

OAI21x1_ASAP7_75t_L g5893 ( 
.A1(n_5784),
.A2(n_4789),
.B(n_4787),
.Y(n_5893)
);

AOI22xp33_ASAP7_75t_L g5894 ( 
.A1(n_5829),
.A2(n_5716),
.B1(n_5049),
.B2(n_5044),
.Y(n_5894)
);

INVx1_ASAP7_75t_L g5895 ( 
.A(n_5771),
.Y(n_5895)
);

BUFx3_ASAP7_75t_L g5896 ( 
.A(n_5726),
.Y(n_5896)
);

INVx2_ASAP7_75t_L g5897 ( 
.A(n_5732),
.Y(n_5897)
);

AND2x4_ASAP7_75t_L g5898 ( 
.A(n_5839),
.B(n_5202),
.Y(n_5898)
);

BUFx2_ASAP7_75t_L g5899 ( 
.A(n_5725),
.Y(n_5899)
);

AND2x4_ASAP7_75t_L g5900 ( 
.A(n_5756),
.B(n_5226),
.Y(n_5900)
);

INVx3_ASAP7_75t_L g5901 ( 
.A(n_5823),
.Y(n_5901)
);

CKINVDCx5p33_ASAP7_75t_R g5902 ( 
.A(n_5752),
.Y(n_5902)
);

INVx1_ASAP7_75t_L g5903 ( 
.A(n_5773),
.Y(n_5903)
);

AOI22xp33_ASAP7_75t_SL g5904 ( 
.A1(n_5850),
.A2(n_4933),
.B1(n_5009),
.B2(n_5013),
.Y(n_5904)
);

AOI21x1_ASAP7_75t_L g5905 ( 
.A1(n_5805),
.A2(n_4797),
.B(n_4792),
.Y(n_5905)
);

AND2x2_ASAP7_75t_L g5906 ( 
.A(n_5783),
.B(n_4692),
.Y(n_5906)
);

INVx2_ASAP7_75t_L g5907 ( 
.A(n_5742),
.Y(n_5907)
);

INVx2_ASAP7_75t_L g5908 ( 
.A(n_5728),
.Y(n_5908)
);

INVx4_ASAP7_75t_L g5909 ( 
.A(n_5744),
.Y(n_5909)
);

AND2x2_ASAP7_75t_L g5910 ( 
.A(n_5753),
.B(n_4692),
.Y(n_5910)
);

AOI221xp5_ASAP7_75t_SL g5911 ( 
.A1(n_5730),
.A2(n_5010),
.B1(n_5255),
.B2(n_4908),
.C(n_5062),
.Y(n_5911)
);

INVx2_ASAP7_75t_L g5912 ( 
.A(n_5809),
.Y(n_5912)
);

OA21x2_ASAP7_75t_L g5913 ( 
.A1(n_5776),
.A2(n_4811),
.B(n_4818),
.Y(n_5913)
);

BUFx2_ASAP7_75t_L g5914 ( 
.A(n_5749),
.Y(n_5914)
);

INVx2_ASAP7_75t_L g5915 ( 
.A(n_5772),
.Y(n_5915)
);

INVx2_ASAP7_75t_L g5916 ( 
.A(n_5807),
.Y(n_5916)
);

OAI21x1_ASAP7_75t_L g5917 ( 
.A1(n_5832),
.A2(n_4825),
.B(n_4827),
.Y(n_5917)
);

INVx1_ASAP7_75t_L g5918 ( 
.A(n_5833),
.Y(n_5918)
);

INVx2_ASAP7_75t_L g5919 ( 
.A(n_5846),
.Y(n_5919)
);

INVx2_ASAP7_75t_L g5920 ( 
.A(n_5835),
.Y(n_5920)
);

BUFx3_ASAP7_75t_L g5921 ( 
.A(n_5779),
.Y(n_5921)
);

AND2x2_ASAP7_75t_L g5922 ( 
.A(n_5820),
.B(n_4692),
.Y(n_5922)
);

INVx2_ASAP7_75t_L g5923 ( 
.A(n_5840),
.Y(n_5923)
);

OA21x2_ASAP7_75t_L g5924 ( 
.A1(n_5825),
.A2(n_4943),
.B(n_4935),
.Y(n_5924)
);

HB1xp67_ASAP7_75t_L g5925 ( 
.A(n_5761),
.Y(n_5925)
);

AND2x2_ASAP7_75t_L g5926 ( 
.A(n_5791),
.B(n_5808),
.Y(n_5926)
);

OAI21x1_ASAP7_75t_L g5927 ( 
.A1(n_5765),
.A2(n_5310),
.B(n_5294),
.Y(n_5927)
);

INVx2_ASAP7_75t_L g5928 ( 
.A(n_5837),
.Y(n_5928)
);

INVx1_ASAP7_75t_L g5929 ( 
.A(n_5824),
.Y(n_5929)
);

AND2x2_ASAP7_75t_L g5930 ( 
.A(n_5791),
.B(n_5812),
.Y(n_5930)
);

INVx2_ASAP7_75t_L g5931 ( 
.A(n_5781),
.Y(n_5931)
);

OAI21xp5_ASAP7_75t_L g5932 ( 
.A1(n_5758),
.A2(n_5666),
.B(n_5693),
.Y(n_5932)
);

INVx1_ASAP7_75t_L g5933 ( 
.A(n_5802),
.Y(n_5933)
);

NOR2xp33_ASAP7_75t_L g5934 ( 
.A(n_5737),
.B(n_4901),
.Y(n_5934)
);

CKINVDCx5p33_ASAP7_75t_R g5935 ( 
.A(n_5782),
.Y(n_5935)
);

INVx2_ASAP7_75t_L g5936 ( 
.A(n_5781),
.Y(n_5936)
);

INVx2_ASAP7_75t_L g5937 ( 
.A(n_5853),
.Y(n_5937)
);

INVx2_ASAP7_75t_L g5938 ( 
.A(n_5815),
.Y(n_5938)
);

OA21x2_ASAP7_75t_L g5939 ( 
.A1(n_5815),
.A2(n_4955),
.B(n_4945),
.Y(n_5939)
);

INVx2_ASAP7_75t_L g5940 ( 
.A(n_5774),
.Y(n_5940)
);

INVx1_ASAP7_75t_L g5941 ( 
.A(n_5798),
.Y(n_5941)
);

OR2x2_ASAP7_75t_L g5942 ( 
.A(n_5803),
.B(n_5022),
.Y(n_5942)
);

INVx1_ASAP7_75t_L g5943 ( 
.A(n_5804),
.Y(n_5943)
);

INVx2_ASAP7_75t_L g5944 ( 
.A(n_5774),
.Y(n_5944)
);

HB1xp67_ASAP7_75t_L g5945 ( 
.A(n_5729),
.Y(n_5945)
);

BUFx2_ASAP7_75t_L g5946 ( 
.A(n_5755),
.Y(n_5946)
);

BUFx2_ASAP7_75t_L g5947 ( 
.A(n_5823),
.Y(n_5947)
);

AOI22xp5_ASAP7_75t_L g5948 ( 
.A1(n_5843),
.A2(n_4604),
.B1(n_4977),
.B2(n_4964),
.Y(n_5948)
);

AO21x1_ASAP7_75t_SL g5949 ( 
.A1(n_5813),
.A2(n_5036),
.B(n_4941),
.Y(n_5949)
);

HB1xp67_ASAP7_75t_L g5950 ( 
.A(n_5836),
.Y(n_5950)
);

INVx5_ASAP7_75t_SL g5951 ( 
.A(n_5735),
.Y(n_5951)
);

BUFx6f_ASAP7_75t_L g5952 ( 
.A(n_5760),
.Y(n_5952)
);

AOI22xp33_ASAP7_75t_L g5953 ( 
.A1(n_5850),
.A2(n_4810),
.B1(n_5065),
.B2(n_5058),
.Y(n_5953)
);

INVx1_ASAP7_75t_L g5954 ( 
.A(n_5800),
.Y(n_5954)
);

AOI22xp33_ASAP7_75t_SL g5955 ( 
.A1(n_5851),
.A2(n_4984),
.B1(n_4981),
.B2(n_4921),
.Y(n_5955)
);

OR2x2_ASAP7_75t_L g5956 ( 
.A(n_5762),
.B(n_4911),
.Y(n_5956)
);

INVx1_ASAP7_75t_L g5957 ( 
.A(n_5827),
.Y(n_5957)
);

INVx1_ASAP7_75t_SL g5958 ( 
.A(n_5760),
.Y(n_5958)
);

INVx1_ASAP7_75t_L g5959 ( 
.A(n_5849),
.Y(n_5959)
);

INVx1_ASAP7_75t_L g5960 ( 
.A(n_5848),
.Y(n_5960)
);

INVx2_ASAP7_75t_L g5961 ( 
.A(n_5855),
.Y(n_5961)
);

AND4x1_ASAP7_75t_L g5962 ( 
.A(n_5750),
.B(n_4791),
.C(n_4603),
.D(n_4842),
.Y(n_5962)
);

INVx1_ASAP7_75t_L g5963 ( 
.A(n_5801),
.Y(n_5963)
);

INVx4_ASAP7_75t_L g5964 ( 
.A(n_5780),
.Y(n_5964)
);

INVx1_ASAP7_75t_L g5965 ( 
.A(n_5847),
.Y(n_5965)
);

INVx1_ASAP7_75t_L g5966 ( 
.A(n_5847),
.Y(n_5966)
);

OR2x2_ASAP7_75t_L g5967 ( 
.A(n_5778),
.B(n_4814),
.Y(n_5967)
);

INVx3_ASAP7_75t_L g5968 ( 
.A(n_5834),
.Y(n_5968)
);

INVx1_ASAP7_75t_SL g5969 ( 
.A(n_5775),
.Y(n_5969)
);

INVx1_ASAP7_75t_SL g5970 ( 
.A(n_5770),
.Y(n_5970)
);

INVx1_ASAP7_75t_L g5971 ( 
.A(n_5740),
.Y(n_5971)
);

HB1xp67_ASAP7_75t_L g5972 ( 
.A(n_5830),
.Y(n_5972)
);

OR2x2_ASAP7_75t_L g5973 ( 
.A(n_5792),
.B(n_4815),
.Y(n_5973)
);

NAND2xp5_ASAP7_75t_L g5974 ( 
.A(n_5886),
.B(n_5841),
.Y(n_5974)
);

NAND2xp5_ASAP7_75t_L g5975 ( 
.A(n_5945),
.B(n_5831),
.Y(n_5975)
);

AO21x2_ASAP7_75t_L g5976 ( 
.A1(n_5965),
.A2(n_5845),
.B(n_5785),
.Y(n_5976)
);

INVx1_ASAP7_75t_L g5977 ( 
.A(n_5972),
.Y(n_5977)
);

INVx1_ASAP7_75t_L g5978 ( 
.A(n_5943),
.Y(n_5978)
);

AND2x2_ASAP7_75t_L g5979 ( 
.A(n_5899),
.B(n_5819),
.Y(n_5979)
);

INVx1_ASAP7_75t_L g5980 ( 
.A(n_5918),
.Y(n_5980)
);

AND2x2_ASAP7_75t_L g5981 ( 
.A(n_5925),
.B(n_5826),
.Y(n_5981)
);

INVx2_ASAP7_75t_SL g5982 ( 
.A(n_5921),
.Y(n_5982)
);

OR2x2_ASAP7_75t_L g5983 ( 
.A(n_5956),
.B(n_5787),
.Y(n_5983)
);

AO21x2_ASAP7_75t_L g5984 ( 
.A1(n_5965),
.A2(n_5795),
.B(n_5814),
.Y(n_5984)
);

AND2x2_ASAP7_75t_L g5985 ( 
.A(n_5964),
.B(n_5930),
.Y(n_5985)
);

OR2x2_ASAP7_75t_L g5986 ( 
.A(n_5881),
.B(n_5933),
.Y(n_5986)
);

NAND2xp5_ASAP7_75t_SL g5987 ( 
.A(n_5964),
.B(n_5733),
.Y(n_5987)
);

INVx1_ASAP7_75t_L g5988 ( 
.A(n_5941),
.Y(n_5988)
);

INVx2_ASAP7_75t_L g5989 ( 
.A(n_5914),
.Y(n_5989)
);

INVx1_ASAP7_75t_L g5990 ( 
.A(n_5857),
.Y(n_5990)
);

INVx1_ASAP7_75t_L g5991 ( 
.A(n_5861),
.Y(n_5991)
);

NAND2xp5_ASAP7_75t_L g5992 ( 
.A(n_5900),
.B(n_5844),
.Y(n_5992)
);

INVxp67_ASAP7_75t_L g5993 ( 
.A(n_5884),
.Y(n_5993)
);

HB1xp67_ASAP7_75t_L g5994 ( 
.A(n_5966),
.Y(n_5994)
);

AND2x2_ASAP7_75t_L g5995 ( 
.A(n_5947),
.B(n_5901),
.Y(n_5995)
);

OR2x2_ASAP7_75t_SL g5996 ( 
.A(n_5856),
.B(n_5821),
.Y(n_5996)
);

INVx1_ASAP7_75t_L g5997 ( 
.A(n_5954),
.Y(n_5997)
);

OA21x2_ASAP7_75t_L g5998 ( 
.A1(n_5859),
.A2(n_5777),
.B(n_5759),
.Y(n_5998)
);

INVx2_ASAP7_75t_L g5999 ( 
.A(n_5912),
.Y(n_5999)
);

INVx2_ASAP7_75t_L g6000 ( 
.A(n_5919),
.Y(n_6000)
);

INVx1_ASAP7_75t_L g6001 ( 
.A(n_5866),
.Y(n_6001)
);

INVx2_ASAP7_75t_L g6002 ( 
.A(n_5896),
.Y(n_6002)
);

NAND2x1p5_ASAP7_75t_L g6003 ( 
.A(n_5909),
.B(n_5768),
.Y(n_6003)
);

BUFx2_ASAP7_75t_L g6004 ( 
.A(n_5909),
.Y(n_6004)
);

INVx1_ASAP7_75t_L g6005 ( 
.A(n_5866),
.Y(n_6005)
);

INVx3_ASAP7_75t_L g6006 ( 
.A(n_5951),
.Y(n_6006)
);

INVx1_ASAP7_75t_L g6007 ( 
.A(n_5875),
.Y(n_6007)
);

HB1xp67_ASAP7_75t_L g6008 ( 
.A(n_5966),
.Y(n_6008)
);

AO21x2_ASAP7_75t_L g6009 ( 
.A1(n_5877),
.A2(n_5971),
.B(n_5932),
.Y(n_6009)
);

BUFx3_ASAP7_75t_L g6010 ( 
.A(n_5883),
.Y(n_6010)
);

INVx3_ASAP7_75t_L g6011 ( 
.A(n_5951),
.Y(n_6011)
);

OR2x6_ASAP7_75t_L g6012 ( 
.A(n_5884),
.B(n_5769),
.Y(n_6012)
);

BUFx3_ASAP7_75t_L g6013 ( 
.A(n_5884),
.Y(n_6013)
);

INVx1_ASAP7_75t_L g6014 ( 
.A(n_5876),
.Y(n_6014)
);

INVx2_ASAP7_75t_L g6015 ( 
.A(n_5938),
.Y(n_6015)
);

INVx2_ASAP7_75t_L g6016 ( 
.A(n_5907),
.Y(n_6016)
);

BUFx2_ASAP7_75t_L g6017 ( 
.A(n_5952),
.Y(n_6017)
);

OR2x2_ASAP7_75t_L g6018 ( 
.A(n_5871),
.B(n_5834),
.Y(n_6018)
);

AO21x2_ASAP7_75t_L g6019 ( 
.A1(n_5868),
.A2(n_5794),
.B(n_4971),
.Y(n_6019)
);

AO21x2_ASAP7_75t_L g6020 ( 
.A1(n_5929),
.A2(n_5794),
.B(n_4777),
.Y(n_6020)
);

BUFx3_ASAP7_75t_L g6021 ( 
.A(n_5952),
.Y(n_6021)
);

BUFx2_ASAP7_75t_L g6022 ( 
.A(n_5952),
.Y(n_6022)
);

INVx1_ASAP7_75t_L g6023 ( 
.A(n_5879),
.Y(n_6023)
);

INVx2_ASAP7_75t_L g6024 ( 
.A(n_5872),
.Y(n_6024)
);

NOR2xp33_ASAP7_75t_L g6025 ( 
.A(n_5902),
.B(n_5892),
.Y(n_6025)
);

BUFx2_ASAP7_75t_L g6026 ( 
.A(n_5901),
.Y(n_6026)
);

NOR2xp33_ASAP7_75t_L g6027 ( 
.A(n_5969),
.B(n_5790),
.Y(n_6027)
);

AND2x4_ASAP7_75t_L g6028 ( 
.A(n_5940),
.B(n_5810),
.Y(n_6028)
);

OA21x2_ASAP7_75t_L g6029 ( 
.A1(n_5873),
.A2(n_5797),
.B(n_5357),
.Y(n_6029)
);

INVxp67_ASAP7_75t_L g6030 ( 
.A(n_5934),
.Y(n_6030)
);

INVx1_ASAP7_75t_L g6031 ( 
.A(n_5882),
.Y(n_6031)
);

INVx2_ASAP7_75t_L g6032 ( 
.A(n_5887),
.Y(n_6032)
);

CKINVDCx6p67_ASAP7_75t_R g6033 ( 
.A(n_5970),
.Y(n_6033)
);

INVx2_ASAP7_75t_L g6034 ( 
.A(n_5867),
.Y(n_6034)
);

NAND2xp5_ASAP7_75t_L g6035 ( 
.A(n_5900),
.B(n_5910),
.Y(n_6035)
);

HB1xp67_ASAP7_75t_L g6036 ( 
.A(n_5950),
.Y(n_6036)
);

INVx2_ASAP7_75t_L g6037 ( 
.A(n_5860),
.Y(n_6037)
);

AND2x4_ASAP7_75t_L g6038 ( 
.A(n_5944),
.B(n_5371),
.Y(n_6038)
);

HB1xp67_ASAP7_75t_L g6039 ( 
.A(n_5928),
.Y(n_6039)
);

BUFx2_ASAP7_75t_SL g6040 ( 
.A(n_5958),
.Y(n_6040)
);

INVx2_ASAP7_75t_SL g6041 ( 
.A(n_5946),
.Y(n_6041)
);

INVx3_ASAP7_75t_L g6042 ( 
.A(n_5888),
.Y(n_6042)
);

AOI21xp5_ASAP7_75t_SL g6043 ( 
.A1(n_5924),
.A2(n_5002),
.B(n_4991),
.Y(n_6043)
);

INVx2_ASAP7_75t_L g6044 ( 
.A(n_5862),
.Y(n_6044)
);

INVx3_ASAP7_75t_L g6045 ( 
.A(n_5935),
.Y(n_6045)
);

INVx1_ASAP7_75t_L g6046 ( 
.A(n_5890),
.Y(n_6046)
);

INVx2_ASAP7_75t_SL g6047 ( 
.A(n_5878),
.Y(n_6047)
);

AND2x2_ASAP7_75t_L g6048 ( 
.A(n_5858),
.B(n_5020),
.Y(n_6048)
);

INVx1_ASAP7_75t_L g6049 ( 
.A(n_5891),
.Y(n_6049)
);

INVx1_ASAP7_75t_L g6050 ( 
.A(n_5895),
.Y(n_6050)
);

INVx2_ASAP7_75t_L g6051 ( 
.A(n_5863),
.Y(n_6051)
);

AND2x2_ASAP7_75t_L g6052 ( 
.A(n_5926),
.B(n_5020),
.Y(n_6052)
);

BUFx3_ASAP7_75t_L g6053 ( 
.A(n_5931),
.Y(n_6053)
);

INVx2_ASAP7_75t_L g6054 ( 
.A(n_5889),
.Y(n_6054)
);

INVx2_ASAP7_75t_L g6055 ( 
.A(n_5897),
.Y(n_6055)
);

INVx1_ASAP7_75t_L g6056 ( 
.A(n_5903),
.Y(n_6056)
);

NAND2xp5_ASAP7_75t_L g6057 ( 
.A(n_5939),
.B(n_5380),
.Y(n_6057)
);

INVx1_ASAP7_75t_L g6058 ( 
.A(n_5869),
.Y(n_6058)
);

INVx2_ASAP7_75t_L g6059 ( 
.A(n_5916),
.Y(n_6059)
);

INVx2_ASAP7_75t_L g6060 ( 
.A(n_5915),
.Y(n_6060)
);

AO21x2_ASAP7_75t_L g6061 ( 
.A1(n_5957),
.A2(n_5923),
.B(n_5959),
.Y(n_6061)
);

INVx3_ASAP7_75t_L g6062 ( 
.A(n_5936),
.Y(n_6062)
);

AO21x2_ASAP7_75t_L g6063 ( 
.A1(n_5905),
.A2(n_4794),
.B(n_4770),
.Y(n_6063)
);

INVx2_ASAP7_75t_L g6064 ( 
.A(n_5908),
.Y(n_6064)
);

BUFx6f_ASAP7_75t_L g6065 ( 
.A(n_5927),
.Y(n_6065)
);

INVx1_ASAP7_75t_L g6066 ( 
.A(n_5960),
.Y(n_6066)
);

BUFx2_ASAP7_75t_L g6067 ( 
.A(n_5870),
.Y(n_6067)
);

NAND2xp5_ASAP7_75t_L g6068 ( 
.A(n_5939),
.B(n_5380),
.Y(n_6068)
);

AND2x2_ASAP7_75t_L g6069 ( 
.A(n_5885),
.B(n_5020),
.Y(n_6069)
);

INVx2_ASAP7_75t_L g6070 ( 
.A(n_5864),
.Y(n_6070)
);

BUFx6f_ASAP7_75t_L g6071 ( 
.A(n_5949),
.Y(n_6071)
);

NAND2xp5_ASAP7_75t_L g6072 ( 
.A(n_5898),
.B(n_5924),
.Y(n_6072)
);

INVx3_ASAP7_75t_L g6073 ( 
.A(n_5961),
.Y(n_6073)
);

OR2x2_ASAP7_75t_L g6074 ( 
.A(n_5942),
.B(n_6),
.Y(n_6074)
);

INVx1_ASAP7_75t_L g6075 ( 
.A(n_5864),
.Y(n_6075)
);

INVx3_ASAP7_75t_L g6076 ( 
.A(n_5968),
.Y(n_6076)
);

INVx1_ASAP7_75t_L g6077 ( 
.A(n_5865),
.Y(n_6077)
);

INVx1_ASAP7_75t_L g6078 ( 
.A(n_5865),
.Y(n_6078)
);

INVx1_ASAP7_75t_L g6079 ( 
.A(n_5906),
.Y(n_6079)
);

AND2x2_ASAP7_75t_L g6080 ( 
.A(n_5922),
.B(n_5329),
.Y(n_6080)
);

INVx1_ASAP7_75t_L g6081 ( 
.A(n_5937),
.Y(n_6081)
);

AND2x2_ASAP7_75t_L g6082 ( 
.A(n_5963),
.B(n_5003),
.Y(n_6082)
);

INVx1_ASAP7_75t_L g6083 ( 
.A(n_5920),
.Y(n_6083)
);

INVx1_ASAP7_75t_L g6084 ( 
.A(n_5898),
.Y(n_6084)
);

AO21x2_ASAP7_75t_L g6085 ( 
.A1(n_5905),
.A2(n_4804),
.B(n_4798),
.Y(n_6085)
);

BUFx3_ASAP7_75t_L g6086 ( 
.A(n_5968),
.Y(n_6086)
);

AND2x4_ASAP7_75t_L g6087 ( 
.A(n_5893),
.B(n_4805),
.Y(n_6087)
);

AND2x2_ASAP7_75t_L g6088 ( 
.A(n_5870),
.B(n_5024),
.Y(n_6088)
);

INVx1_ASAP7_75t_L g6089 ( 
.A(n_5917),
.Y(n_6089)
);

AO21x2_ASAP7_75t_L g6090 ( 
.A1(n_5880),
.A2(n_4809),
.B(n_4808),
.Y(n_6090)
);

INVx2_ASAP7_75t_L g6091 ( 
.A(n_5973),
.Y(n_6091)
);

OR2x2_ASAP7_75t_L g6092 ( 
.A(n_5967),
.B(n_7),
.Y(n_6092)
);

AO21x2_ASAP7_75t_L g6093 ( 
.A1(n_5948),
.A2(n_4968),
.B(n_4892),
.Y(n_6093)
);

INVx1_ASAP7_75t_L g6094 ( 
.A(n_5913),
.Y(n_6094)
);

NOR2x1_ASAP7_75t_SL g6095 ( 
.A(n_5874),
.B(n_507),
.Y(n_6095)
);

HB1xp67_ASAP7_75t_L g6096 ( 
.A(n_5913),
.Y(n_6096)
);

AOI21xp5_ASAP7_75t_L g6097 ( 
.A1(n_5894),
.A2(n_4893),
.B(n_4890),
.Y(n_6097)
);

INVx3_ASAP7_75t_L g6098 ( 
.A(n_5962),
.Y(n_6098)
);

NOR2xp33_ASAP7_75t_L g6099 ( 
.A(n_5904),
.B(n_507),
.Y(n_6099)
);

BUFx3_ASAP7_75t_L g6100 ( 
.A(n_5955),
.Y(n_6100)
);

AO21x2_ASAP7_75t_L g6101 ( 
.A1(n_5953),
.A2(n_4927),
.B(n_4903),
.Y(n_6101)
);

INVx1_ASAP7_75t_L g6102 ( 
.A(n_5911),
.Y(n_6102)
);

INVx2_ASAP7_75t_L g6103 ( 
.A(n_5972),
.Y(n_6103)
);

INVx1_ASAP7_75t_L g6104 ( 
.A(n_5945),
.Y(n_6104)
);

AO21x2_ASAP7_75t_L g6105 ( 
.A1(n_5965),
.A2(n_4957),
.B(n_4928),
.Y(n_6105)
);

OA21x2_ASAP7_75t_L g6106 ( 
.A1(n_5859),
.A2(n_4826),
.B(n_4824),
.Y(n_6106)
);

OR2x6_ASAP7_75t_L g6107 ( 
.A(n_5909),
.B(n_508),
.Y(n_6107)
);

AND2x2_ASAP7_75t_L g6108 ( 
.A(n_5899),
.B(n_7),
.Y(n_6108)
);

AND2x2_ASAP7_75t_L g6109 ( 
.A(n_5899),
.B(n_7),
.Y(n_6109)
);

OR2x2_ASAP7_75t_L g6110 ( 
.A(n_5956),
.B(n_7),
.Y(n_6110)
);

INVx1_ASAP7_75t_L g6111 ( 
.A(n_5945),
.Y(n_6111)
);

AO21x2_ASAP7_75t_L g6112 ( 
.A1(n_5965),
.A2(n_8),
.B(n_9),
.Y(n_6112)
);

INVx1_ASAP7_75t_L g6113 ( 
.A(n_5945),
.Y(n_6113)
);

INVx1_ASAP7_75t_L g6114 ( 
.A(n_5945),
.Y(n_6114)
);

AND2x4_ASAP7_75t_L g6115 ( 
.A(n_5925),
.B(n_508),
.Y(n_6115)
);

INVx1_ASAP7_75t_L g6116 ( 
.A(n_5945),
.Y(n_6116)
);

HB1xp67_ASAP7_75t_L g6117 ( 
.A(n_5972),
.Y(n_6117)
);

INVx2_ASAP7_75t_SL g6118 ( 
.A(n_5921),
.Y(n_6118)
);

HB1xp67_ASAP7_75t_L g6119 ( 
.A(n_5972),
.Y(n_6119)
);

INVx2_ASAP7_75t_L g6120 ( 
.A(n_5972),
.Y(n_6120)
);

AO21x2_ASAP7_75t_L g6121 ( 
.A1(n_5965),
.A2(n_8),
.B(n_9),
.Y(n_6121)
);

AOI22xp33_ASAP7_75t_L g6122 ( 
.A1(n_5925),
.A2(n_510),
.B1(n_511),
.B2(n_509),
.Y(n_6122)
);

INVx1_ASAP7_75t_L g6123 ( 
.A(n_5945),
.Y(n_6123)
);

INVx2_ASAP7_75t_L g6124 ( 
.A(n_5972),
.Y(n_6124)
);

HB1xp67_ASAP7_75t_L g6125 ( 
.A(n_5972),
.Y(n_6125)
);

AOI21x1_ASAP7_75t_L g6126 ( 
.A1(n_5925),
.A2(n_8),
.B(n_9),
.Y(n_6126)
);

AOI22xp5_ASAP7_75t_L g6127 ( 
.A1(n_5868),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_6127)
);

INVx1_ASAP7_75t_L g6128 ( 
.A(n_5945),
.Y(n_6128)
);

OR2x6_ASAP7_75t_L g6129 ( 
.A(n_5909),
.B(n_509),
.Y(n_6129)
);

AOI22xp33_ASAP7_75t_L g6130 ( 
.A1(n_5925),
.A2(n_511),
.B1(n_512),
.B2(n_509),
.Y(n_6130)
);

OR2x2_ASAP7_75t_L g6131 ( 
.A(n_6079),
.B(n_10),
.Y(n_6131)
);

INVx2_ASAP7_75t_L g6132 ( 
.A(n_6103),
.Y(n_6132)
);

NAND2xp5_ASAP7_75t_L g6133 ( 
.A(n_6117),
.B(n_11),
.Y(n_6133)
);

AND2x4_ASAP7_75t_L g6134 ( 
.A(n_5985),
.B(n_512),
.Y(n_6134)
);

AND2x2_ASAP7_75t_L g6135 ( 
.A(n_6004),
.B(n_11),
.Y(n_6135)
);

AND2x4_ASAP7_75t_L g6136 ( 
.A(n_6004),
.B(n_512),
.Y(n_6136)
);

HB1xp67_ASAP7_75t_L g6137 ( 
.A(n_6119),
.Y(n_6137)
);

AND2x2_ASAP7_75t_L g6138 ( 
.A(n_6040),
.B(n_11),
.Y(n_6138)
);

AND2x2_ASAP7_75t_L g6139 ( 
.A(n_6040),
.B(n_11),
.Y(n_6139)
);

INVx1_ASAP7_75t_L g6140 ( 
.A(n_6125),
.Y(n_6140)
);

INVx2_ASAP7_75t_L g6141 ( 
.A(n_6120),
.Y(n_6141)
);

AND2x2_ASAP7_75t_L g6142 ( 
.A(n_5981),
.B(n_12),
.Y(n_6142)
);

AND2x4_ASAP7_75t_L g6143 ( 
.A(n_6013),
.B(n_513),
.Y(n_6143)
);

AND2x2_ASAP7_75t_L g6144 ( 
.A(n_5995),
.B(n_12),
.Y(n_6144)
);

INVx2_ASAP7_75t_SL g6145 ( 
.A(n_6003),
.Y(n_6145)
);

NAND2xp5_ASAP7_75t_L g6146 ( 
.A(n_5977),
.B(n_12),
.Y(n_6146)
);

AND2x2_ASAP7_75t_L g6147 ( 
.A(n_6021),
.B(n_13),
.Y(n_6147)
);

NAND3xp33_ASAP7_75t_L g6148 ( 
.A(n_6102),
.B(n_6127),
.C(n_6099),
.Y(n_6148)
);

INVx1_ASAP7_75t_L g6149 ( 
.A(n_5994),
.Y(n_6149)
);

AND2x2_ASAP7_75t_L g6150 ( 
.A(n_5979),
.B(n_6033),
.Y(n_6150)
);

INVx1_ASAP7_75t_L g6151 ( 
.A(n_6124),
.Y(n_6151)
);

INVx1_ASAP7_75t_L g6152 ( 
.A(n_6008),
.Y(n_6152)
);

HB1xp67_ASAP7_75t_L g6153 ( 
.A(n_6104),
.Y(n_6153)
);

INVx2_ASAP7_75t_L g6154 ( 
.A(n_6026),
.Y(n_6154)
);

INVx2_ASAP7_75t_L g6155 ( 
.A(n_6026),
.Y(n_6155)
);

AND2x2_ASAP7_75t_L g6156 ( 
.A(n_6012),
.B(n_6115),
.Y(n_6156)
);

INVx2_ASAP7_75t_L g6157 ( 
.A(n_6042),
.Y(n_6157)
);

INVx2_ASAP7_75t_L g6158 ( 
.A(n_6041),
.Y(n_6158)
);

INVx1_ASAP7_75t_L g6159 ( 
.A(n_6111),
.Y(n_6159)
);

BUFx3_ASAP7_75t_L g6160 ( 
.A(n_6010),
.Y(n_6160)
);

INVx3_ASAP7_75t_L g6161 ( 
.A(n_6006),
.Y(n_6161)
);

AND2x2_ASAP7_75t_L g6162 ( 
.A(n_6012),
.B(n_13),
.Y(n_6162)
);

OR2x2_ASAP7_75t_L g6163 ( 
.A(n_6113),
.B(n_13),
.Y(n_6163)
);

INVx2_ASAP7_75t_L g6164 ( 
.A(n_5989),
.Y(n_6164)
);

HB1xp67_ASAP7_75t_L g6165 ( 
.A(n_6114),
.Y(n_6165)
);

INVx1_ASAP7_75t_L g6166 ( 
.A(n_6116),
.Y(n_6166)
);

AOI21xp33_ASAP7_75t_L g6167 ( 
.A1(n_5993),
.A2(n_13),
.B(n_14),
.Y(n_6167)
);

INVx2_ASAP7_75t_L g6168 ( 
.A(n_6002),
.Y(n_6168)
);

AND2x2_ASAP7_75t_L g6169 ( 
.A(n_6115),
.B(n_14),
.Y(n_6169)
);

HB1xp67_ASAP7_75t_L g6170 ( 
.A(n_6123),
.Y(n_6170)
);

OAI222xp33_ASAP7_75t_L g6171 ( 
.A1(n_5974),
.A2(n_16),
.B1(n_18),
.B2(n_14),
.C1(n_15),
.C2(n_17),
.Y(n_6171)
);

HB1xp67_ASAP7_75t_L g6172 ( 
.A(n_6128),
.Y(n_6172)
);

INVxp67_ASAP7_75t_L g6173 ( 
.A(n_6027),
.Y(n_6173)
);

HB1xp67_ASAP7_75t_L g6174 ( 
.A(n_6036),
.Y(n_6174)
);

BUFx3_ASAP7_75t_L g6175 ( 
.A(n_6011),
.Y(n_6175)
);

AND2x2_ASAP7_75t_L g6176 ( 
.A(n_5982),
.B(n_14),
.Y(n_6176)
);

AND2x2_ASAP7_75t_L g6177 ( 
.A(n_6118),
.B(n_15),
.Y(n_6177)
);

AND2x2_ASAP7_75t_L g6178 ( 
.A(n_6028),
.B(n_15),
.Y(n_6178)
);

AOI211xp5_ASAP7_75t_L g6179 ( 
.A1(n_5987),
.A2(n_18),
.B(n_15),
.C(n_16),
.Y(n_6179)
);

AND2x2_ASAP7_75t_L g6180 ( 
.A(n_6028),
.B(n_16),
.Y(n_6180)
);

INVx3_ASAP7_75t_L g6181 ( 
.A(n_6045),
.Y(n_6181)
);

AND2x2_ASAP7_75t_L g6182 ( 
.A(n_6017),
.B(n_16),
.Y(n_6182)
);

INVx3_ASAP7_75t_L g6183 ( 
.A(n_6107),
.Y(n_6183)
);

AND2x2_ASAP7_75t_L g6184 ( 
.A(n_6017),
.B(n_6022),
.Y(n_6184)
);

BUFx6f_ASAP7_75t_L g6185 ( 
.A(n_6022),
.Y(n_6185)
);

INVx3_ASAP7_75t_L g6186 ( 
.A(n_6107),
.Y(n_6186)
);

AOI22xp33_ASAP7_75t_SL g6187 ( 
.A1(n_5998),
.A2(n_514),
.B1(n_515),
.B2(n_513),
.Y(n_6187)
);

OAI22xp5_ASAP7_75t_L g6188 ( 
.A1(n_5996),
.A2(n_5998),
.B1(n_5992),
.B2(n_6091),
.Y(n_6188)
);

INVx2_ASAP7_75t_L g6189 ( 
.A(n_6038),
.Y(n_6189)
);

NOR2xp67_ASAP7_75t_L g6190 ( 
.A(n_6098),
.B(n_18),
.Y(n_6190)
);

INVx2_ASAP7_75t_SL g6191 ( 
.A(n_6129),
.Y(n_6191)
);

INVxp67_ASAP7_75t_SL g6192 ( 
.A(n_6126),
.Y(n_6192)
);

AND2x2_ASAP7_75t_L g6193 ( 
.A(n_6025),
.B(n_18),
.Y(n_6193)
);

INVx2_ASAP7_75t_L g6194 ( 
.A(n_6038),
.Y(n_6194)
);

INVx2_ASAP7_75t_L g6195 ( 
.A(n_5999),
.Y(n_6195)
);

AND2x2_ASAP7_75t_L g6196 ( 
.A(n_6080),
.B(n_19),
.Y(n_6196)
);

INVx3_ASAP7_75t_L g6197 ( 
.A(n_6129),
.Y(n_6197)
);

INVx2_ASAP7_75t_L g6198 ( 
.A(n_6000),
.Y(n_6198)
);

NAND2xp5_ASAP7_75t_L g6199 ( 
.A(n_6030),
.B(n_19),
.Y(n_6199)
);

INVx1_ASAP7_75t_L g6200 ( 
.A(n_6108),
.Y(n_6200)
);

INVx1_ASAP7_75t_L g6201 ( 
.A(n_6109),
.Y(n_6201)
);

AND2x4_ASAP7_75t_L g6202 ( 
.A(n_6047),
.B(n_513),
.Y(n_6202)
);

INVx1_ASAP7_75t_L g6203 ( 
.A(n_5978),
.Y(n_6203)
);

INVx1_ASAP7_75t_L g6204 ( 
.A(n_5988),
.Y(n_6204)
);

AND2x2_ASAP7_75t_L g6205 ( 
.A(n_6053),
.B(n_19),
.Y(n_6205)
);

NAND2xp5_ASAP7_75t_L g6206 ( 
.A(n_6088),
.B(n_19),
.Y(n_6206)
);

AND2x2_ASAP7_75t_L g6207 ( 
.A(n_6073),
.B(n_20),
.Y(n_6207)
);

INVx1_ASAP7_75t_L g6208 ( 
.A(n_5997),
.Y(n_6208)
);

INVx1_ASAP7_75t_L g6209 ( 
.A(n_6007),
.Y(n_6209)
);

NOR2x1_ASAP7_75t_SL g6210 ( 
.A(n_6126),
.B(n_514),
.Y(n_6210)
);

BUFx3_ASAP7_75t_L g6211 ( 
.A(n_6071),
.Y(n_6211)
);

HB1xp67_ASAP7_75t_L g6212 ( 
.A(n_6112),
.Y(n_6212)
);

OR2x2_ASAP7_75t_L g6213 ( 
.A(n_5975),
.B(n_20),
.Y(n_6213)
);

INVx2_ASAP7_75t_L g6214 ( 
.A(n_6015),
.Y(n_6214)
);

AND2x2_ASAP7_75t_L g6215 ( 
.A(n_6052),
.B(n_6048),
.Y(n_6215)
);

INVx1_ASAP7_75t_SL g6216 ( 
.A(n_6071),
.Y(n_6216)
);

INVx2_ASAP7_75t_L g6217 ( 
.A(n_6037),
.Y(n_6217)
);

INVx2_ASAP7_75t_L g6218 ( 
.A(n_6044),
.Y(n_6218)
);

AND2x2_ASAP7_75t_L g6219 ( 
.A(n_6062),
.B(n_20),
.Y(n_6219)
);

AND2x4_ASAP7_75t_SL g6220 ( 
.A(n_6122),
.B(n_21),
.Y(n_6220)
);

OR2x6_ASAP7_75t_L g6221 ( 
.A(n_6100),
.B(n_515),
.Y(n_6221)
);

INVx1_ASAP7_75t_L g6222 ( 
.A(n_6075),
.Y(n_6222)
);

AND2x2_ASAP7_75t_L g6223 ( 
.A(n_6069),
.B(n_21),
.Y(n_6223)
);

NAND2xp5_ASAP7_75t_L g6224 ( 
.A(n_6101),
.B(n_22),
.Y(n_6224)
);

INVx2_ASAP7_75t_L g6225 ( 
.A(n_6016),
.Y(n_6225)
);

NAND2xp5_ASAP7_75t_L g6226 ( 
.A(n_6090),
.B(n_22),
.Y(n_6226)
);

OR2x2_ASAP7_75t_L g6227 ( 
.A(n_6035),
.B(n_22),
.Y(n_6227)
);

OR2x2_ASAP7_75t_L g6228 ( 
.A(n_5983),
.B(n_22),
.Y(n_6228)
);

AND2x2_ASAP7_75t_L g6229 ( 
.A(n_6084),
.B(n_23),
.Y(n_6229)
);

NAND2xp5_ASAP7_75t_L g6230 ( 
.A(n_6092),
.B(n_23),
.Y(n_6230)
);

HB1xp67_ASAP7_75t_L g6231 ( 
.A(n_6121),
.Y(n_6231)
);

INVx1_ASAP7_75t_L g6232 ( 
.A(n_6075),
.Y(n_6232)
);

NAND2x1_ASAP7_75t_L g6233 ( 
.A(n_6029),
.B(n_515),
.Y(n_6233)
);

NAND2xp5_ASAP7_75t_L g6234 ( 
.A(n_6094),
.B(n_23),
.Y(n_6234)
);

INVxp67_ASAP7_75t_L g6235 ( 
.A(n_6095),
.Y(n_6235)
);

INVx2_ASAP7_75t_L g6236 ( 
.A(n_6024),
.Y(n_6236)
);

INVxp67_ASAP7_75t_L g6237 ( 
.A(n_6095),
.Y(n_6237)
);

INVx2_ASAP7_75t_L g6238 ( 
.A(n_6032),
.Y(n_6238)
);

OAI21xp5_ASAP7_75t_L g6239 ( 
.A1(n_6043),
.A2(n_23),
.B(n_24),
.Y(n_6239)
);

BUFx3_ASAP7_75t_L g6240 ( 
.A(n_6086),
.Y(n_6240)
);

INVx2_ASAP7_75t_SL g6241 ( 
.A(n_6018),
.Y(n_6241)
);

AO221x2_ASAP7_75t_L g6242 ( 
.A1(n_6072),
.A2(n_519),
.B1(n_520),
.B2(n_517),
.C(n_516),
.Y(n_6242)
);

AND2x2_ASAP7_75t_SL g6243 ( 
.A(n_6029),
.B(n_516),
.Y(n_6243)
);

AOI22xp5_ASAP7_75t_L g6244 ( 
.A1(n_6087),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_6244)
);

INVx1_ASAP7_75t_L g6245 ( 
.A(n_6014),
.Y(n_6245)
);

NOR2xp33_ASAP7_75t_L g6246 ( 
.A(n_6110),
.B(n_24),
.Y(n_6246)
);

INVx1_ASAP7_75t_L g6247 ( 
.A(n_6023),
.Y(n_6247)
);

AND2x2_ASAP7_75t_L g6248 ( 
.A(n_6019),
.B(n_24),
.Y(n_6248)
);

INVx1_ASAP7_75t_L g6249 ( 
.A(n_6031),
.Y(n_6249)
);

AND2x2_ASAP7_75t_L g6250 ( 
.A(n_6106),
.B(n_25),
.Y(n_6250)
);

INVx2_ASAP7_75t_L g6251 ( 
.A(n_6054),
.Y(n_6251)
);

INVx1_ASAP7_75t_L g6252 ( 
.A(n_6046),
.Y(n_6252)
);

INVx2_ASAP7_75t_L g6253 ( 
.A(n_6055),
.Y(n_6253)
);

AND2x4_ASAP7_75t_L g6254 ( 
.A(n_6087),
.B(n_516),
.Y(n_6254)
);

INVx2_ASAP7_75t_L g6255 ( 
.A(n_6034),
.Y(n_6255)
);

HB1xp67_ASAP7_75t_L g6256 ( 
.A(n_5980),
.Y(n_6256)
);

INVx1_ASAP7_75t_L g6257 ( 
.A(n_6070),
.Y(n_6257)
);

AND2x2_ASAP7_75t_L g6258 ( 
.A(n_6106),
.B(n_25),
.Y(n_6258)
);

INVx2_ASAP7_75t_L g6259 ( 
.A(n_6051),
.Y(n_6259)
);

INVx1_ASAP7_75t_L g6260 ( 
.A(n_6049),
.Y(n_6260)
);

AND2x2_ASAP7_75t_L g6261 ( 
.A(n_6076),
.B(n_6082),
.Y(n_6261)
);

AND2x2_ASAP7_75t_L g6262 ( 
.A(n_6096),
.B(n_25),
.Y(n_6262)
);

INVx3_ASAP7_75t_L g6263 ( 
.A(n_6064),
.Y(n_6263)
);

INVx2_ASAP7_75t_L g6264 ( 
.A(n_6059),
.Y(n_6264)
);

AND2x2_ASAP7_75t_L g6265 ( 
.A(n_6089),
.B(n_26),
.Y(n_6265)
);

NAND4xp25_ASAP7_75t_L g6266 ( 
.A(n_6130),
.B(n_28),
.C(n_26),
.D(n_27),
.Y(n_6266)
);

AND2x4_ASAP7_75t_L g6267 ( 
.A(n_6050),
.B(n_517),
.Y(n_6267)
);

AND2x2_ASAP7_75t_L g6268 ( 
.A(n_5976),
.B(n_6060),
.Y(n_6268)
);

INVx2_ASAP7_75t_L g6269 ( 
.A(n_5980),
.Y(n_6269)
);

AND2x2_ASAP7_75t_L g6270 ( 
.A(n_6009),
.B(n_26),
.Y(n_6270)
);

NAND2xp5_ASAP7_75t_L g6271 ( 
.A(n_6056),
.B(n_27),
.Y(n_6271)
);

INVx1_ASAP7_75t_L g6272 ( 
.A(n_5990),
.Y(n_6272)
);

AND2x4_ASAP7_75t_L g6273 ( 
.A(n_6058),
.B(n_517),
.Y(n_6273)
);

HB1xp67_ASAP7_75t_L g6274 ( 
.A(n_5990),
.Y(n_6274)
);

AND2x2_ASAP7_75t_L g6275 ( 
.A(n_6074),
.B(n_27),
.Y(n_6275)
);

INVx2_ASAP7_75t_L g6276 ( 
.A(n_5991),
.Y(n_6276)
);

AND2x2_ASAP7_75t_L g6277 ( 
.A(n_6020),
.B(n_27),
.Y(n_6277)
);

INVx1_ASAP7_75t_L g6278 ( 
.A(n_5991),
.Y(n_6278)
);

INVx2_ASAP7_75t_L g6279 ( 
.A(n_6077),
.Y(n_6279)
);

AND2x2_ASAP7_75t_L g6280 ( 
.A(n_5984),
.B(n_5986),
.Y(n_6280)
);

NAND2xp5_ASAP7_75t_L g6281 ( 
.A(n_6063),
.B(n_28),
.Y(n_6281)
);

AND2x2_ASAP7_75t_L g6282 ( 
.A(n_6039),
.B(n_28),
.Y(n_6282)
);

INVx1_ASAP7_75t_L g6283 ( 
.A(n_6078),
.Y(n_6283)
);

NAND2xp5_ASAP7_75t_L g6284 ( 
.A(n_6085),
.B(n_29),
.Y(n_6284)
);

INVx2_ASAP7_75t_L g6285 ( 
.A(n_6081),
.Y(n_6285)
);

AND2x2_ASAP7_75t_L g6286 ( 
.A(n_6065),
.B(n_29),
.Y(n_6286)
);

NAND2xp5_ASAP7_75t_L g6287 ( 
.A(n_6093),
.B(n_29),
.Y(n_6287)
);

INVx3_ASAP7_75t_L g6288 ( 
.A(n_6065),
.Y(n_6288)
);

INVx1_ASAP7_75t_L g6289 ( 
.A(n_6001),
.Y(n_6289)
);

AND2x2_ASAP7_75t_L g6290 ( 
.A(n_6083),
.B(n_30),
.Y(n_6290)
);

AO21x2_ASAP7_75t_L g6291 ( 
.A1(n_6061),
.A2(n_31),
.B(n_32),
.Y(n_6291)
);

INVx3_ASAP7_75t_L g6292 ( 
.A(n_6067),
.Y(n_6292)
);

INVx2_ASAP7_75t_L g6293 ( 
.A(n_6005),
.Y(n_6293)
);

INVx1_ASAP7_75t_L g6294 ( 
.A(n_6066),
.Y(n_6294)
);

INVx2_ASAP7_75t_L g6295 ( 
.A(n_6067),
.Y(n_6295)
);

HB1xp67_ASAP7_75t_L g6296 ( 
.A(n_6057),
.Y(n_6296)
);

INVxp67_ASAP7_75t_R g6297 ( 
.A(n_6097),
.Y(n_6297)
);

AND2x2_ASAP7_75t_L g6298 ( 
.A(n_6068),
.B(n_31),
.Y(n_6298)
);

OR2x2_ASAP7_75t_L g6299 ( 
.A(n_6105),
.B(n_32),
.Y(n_6299)
);

INVx1_ASAP7_75t_L g6300 ( 
.A(n_6117),
.Y(n_6300)
);

NAND2xp5_ASAP7_75t_L g6301 ( 
.A(n_6117),
.B(n_32),
.Y(n_6301)
);

INVx1_ASAP7_75t_L g6302 ( 
.A(n_6117),
.Y(n_6302)
);

AND2x2_ASAP7_75t_L g6303 ( 
.A(n_5985),
.B(n_33),
.Y(n_6303)
);

INVx3_ASAP7_75t_L g6304 ( 
.A(n_6010),
.Y(n_6304)
);

NAND2xp5_ASAP7_75t_L g6305 ( 
.A(n_6117),
.B(n_33),
.Y(n_6305)
);

INVx1_ASAP7_75t_L g6306 ( 
.A(n_6117),
.Y(n_6306)
);

INVx1_ASAP7_75t_L g6307 ( 
.A(n_6117),
.Y(n_6307)
);

AND2x2_ASAP7_75t_L g6308 ( 
.A(n_5985),
.B(n_33),
.Y(n_6308)
);

BUFx3_ASAP7_75t_L g6309 ( 
.A(n_6160),
.Y(n_6309)
);

INVx2_ASAP7_75t_L g6310 ( 
.A(n_6168),
.Y(n_6310)
);

INVx4_ASAP7_75t_L g6311 ( 
.A(n_6304),
.Y(n_6311)
);

OR2x2_ASAP7_75t_L g6312 ( 
.A(n_6234),
.B(n_33),
.Y(n_6312)
);

BUFx3_ASAP7_75t_L g6313 ( 
.A(n_6211),
.Y(n_6313)
);

AND2x2_ASAP7_75t_L g6314 ( 
.A(n_6150),
.B(n_34),
.Y(n_6314)
);

INVx1_ASAP7_75t_L g6315 ( 
.A(n_6135),
.Y(n_6315)
);

NOR2xp33_ASAP7_75t_L g6316 ( 
.A(n_6173),
.B(n_34),
.Y(n_6316)
);

HB1xp67_ASAP7_75t_L g6317 ( 
.A(n_6137),
.Y(n_6317)
);

INVx1_ASAP7_75t_L g6318 ( 
.A(n_6182),
.Y(n_6318)
);

OR2x2_ASAP7_75t_L g6319 ( 
.A(n_6206),
.B(n_34),
.Y(n_6319)
);

AND2x4_ASAP7_75t_L g6320 ( 
.A(n_6175),
.B(n_35),
.Y(n_6320)
);

NAND2xp5_ASAP7_75t_L g6321 ( 
.A(n_6178),
.B(n_34),
.Y(n_6321)
);

INVx3_ASAP7_75t_L g6322 ( 
.A(n_6240),
.Y(n_6322)
);

BUFx6f_ASAP7_75t_L g6323 ( 
.A(n_6185),
.Y(n_6323)
);

OR2x2_ASAP7_75t_L g6324 ( 
.A(n_6300),
.B(n_35),
.Y(n_6324)
);

AND2x2_ASAP7_75t_L g6325 ( 
.A(n_6216),
.B(n_35),
.Y(n_6325)
);

AND2x2_ASAP7_75t_L g6326 ( 
.A(n_6161),
.B(n_36),
.Y(n_6326)
);

AND2x2_ASAP7_75t_L g6327 ( 
.A(n_6156),
.B(n_36),
.Y(n_6327)
);

OR2x2_ASAP7_75t_L g6328 ( 
.A(n_6307),
.B(n_36),
.Y(n_6328)
);

OR2x2_ASAP7_75t_L g6329 ( 
.A(n_6140),
.B(n_36),
.Y(n_6329)
);

NAND2xp5_ASAP7_75t_L g6330 ( 
.A(n_6180),
.B(n_37),
.Y(n_6330)
);

INVx3_ASAP7_75t_L g6331 ( 
.A(n_6185),
.Y(n_6331)
);

BUFx3_ASAP7_75t_L g6332 ( 
.A(n_6181),
.Y(n_6332)
);

INVx1_ASAP7_75t_L g6333 ( 
.A(n_6174),
.Y(n_6333)
);

HB1xp67_ASAP7_75t_L g6334 ( 
.A(n_6140),
.Y(n_6334)
);

AND2x2_ASAP7_75t_L g6335 ( 
.A(n_6145),
.B(n_37),
.Y(n_6335)
);

INVx5_ASAP7_75t_L g6336 ( 
.A(n_6185),
.Y(n_6336)
);

AND2x2_ASAP7_75t_L g6337 ( 
.A(n_6183),
.B(n_37),
.Y(n_6337)
);

AND2x2_ASAP7_75t_L g6338 ( 
.A(n_6186),
.B(n_38),
.Y(n_6338)
);

INVx2_ASAP7_75t_L g6339 ( 
.A(n_6136),
.Y(n_6339)
);

INVx2_ASAP7_75t_L g6340 ( 
.A(n_6136),
.Y(n_6340)
);

AND2x2_ASAP7_75t_L g6341 ( 
.A(n_6197),
.B(n_38),
.Y(n_6341)
);

INVx1_ASAP7_75t_L g6342 ( 
.A(n_6138),
.Y(n_6342)
);

INVx1_ASAP7_75t_L g6343 ( 
.A(n_6139),
.Y(n_6343)
);

BUFx12f_ASAP7_75t_L g6344 ( 
.A(n_6191),
.Y(n_6344)
);

INVx2_ASAP7_75t_L g6345 ( 
.A(n_6202),
.Y(n_6345)
);

NAND2xp5_ASAP7_75t_L g6346 ( 
.A(n_6270),
.B(n_38),
.Y(n_6346)
);

INVx1_ASAP7_75t_L g6347 ( 
.A(n_6302),
.Y(n_6347)
);

AOI22xp33_ASAP7_75t_L g6348 ( 
.A1(n_6241),
.A2(n_520),
.B1(n_521),
.B2(n_519),
.Y(n_6348)
);

AND2x2_ASAP7_75t_L g6349 ( 
.A(n_6158),
.B(n_38),
.Y(n_6349)
);

INVx3_ASAP7_75t_L g6350 ( 
.A(n_6202),
.Y(n_6350)
);

INVx2_ASAP7_75t_L g6351 ( 
.A(n_6154),
.Y(n_6351)
);

INVx1_ASAP7_75t_L g6352 ( 
.A(n_6302),
.Y(n_6352)
);

INVx1_ASAP7_75t_L g6353 ( 
.A(n_6306),
.Y(n_6353)
);

AND2x2_ASAP7_75t_L g6354 ( 
.A(n_6184),
.B(n_39),
.Y(n_6354)
);

INVx1_ASAP7_75t_SL g6355 ( 
.A(n_6176),
.Y(n_6355)
);

HB1xp67_ASAP7_75t_L g6356 ( 
.A(n_6306),
.Y(n_6356)
);

NOR2xp33_ASAP7_75t_L g6357 ( 
.A(n_6235),
.B(n_39),
.Y(n_6357)
);

NOR2x1_ASAP7_75t_L g6358 ( 
.A(n_6291),
.B(n_39),
.Y(n_6358)
);

AND2x2_ASAP7_75t_L g6359 ( 
.A(n_6261),
.B(n_6265),
.Y(n_6359)
);

AND2x4_ASAP7_75t_L g6360 ( 
.A(n_6162),
.B(n_521),
.Y(n_6360)
);

BUFx2_ASAP7_75t_L g6361 ( 
.A(n_6155),
.Y(n_6361)
);

INVx4_ASAP7_75t_L g6362 ( 
.A(n_6177),
.Y(n_6362)
);

INVx1_ASAP7_75t_L g6363 ( 
.A(n_6282),
.Y(n_6363)
);

HB1xp67_ASAP7_75t_L g6364 ( 
.A(n_6262),
.Y(n_6364)
);

AND2x2_ASAP7_75t_L g6365 ( 
.A(n_6196),
.B(n_40),
.Y(n_6365)
);

HB1xp67_ASAP7_75t_L g6366 ( 
.A(n_6153),
.Y(n_6366)
);

NOR2x1_ASAP7_75t_SL g6367 ( 
.A(n_6248),
.B(n_521),
.Y(n_6367)
);

INVxp67_ASAP7_75t_R g6368 ( 
.A(n_6286),
.Y(n_6368)
);

AND2x4_ASAP7_75t_L g6369 ( 
.A(n_6143),
.B(n_522),
.Y(n_6369)
);

AND2x2_ASAP7_75t_L g6370 ( 
.A(n_6142),
.B(n_40),
.Y(n_6370)
);

INVx1_ASAP7_75t_L g6371 ( 
.A(n_6165),
.Y(n_6371)
);

AND2x2_ASAP7_75t_L g6372 ( 
.A(n_6297),
.B(n_41),
.Y(n_6372)
);

NAND2xp5_ASAP7_75t_L g6373 ( 
.A(n_6223),
.B(n_41),
.Y(n_6373)
);

INVx1_ASAP7_75t_L g6374 ( 
.A(n_6170),
.Y(n_6374)
);

INVx2_ASAP7_75t_L g6375 ( 
.A(n_6210),
.Y(n_6375)
);

HB1xp67_ASAP7_75t_L g6376 ( 
.A(n_6172),
.Y(n_6376)
);

INVx1_ASAP7_75t_L g6377 ( 
.A(n_6295),
.Y(n_6377)
);

INVx1_ASAP7_75t_L g6378 ( 
.A(n_6133),
.Y(n_6378)
);

INVx2_ASAP7_75t_L g6379 ( 
.A(n_6210),
.Y(n_6379)
);

INVx1_ASAP7_75t_L g6380 ( 
.A(n_6301),
.Y(n_6380)
);

AND2x2_ASAP7_75t_L g6381 ( 
.A(n_6221),
.B(n_41),
.Y(n_6381)
);

INVx3_ASAP7_75t_SL g6382 ( 
.A(n_6143),
.Y(n_6382)
);

HB1xp67_ASAP7_75t_L g6383 ( 
.A(n_6151),
.Y(n_6383)
);

BUFx2_ASAP7_75t_L g6384 ( 
.A(n_6292),
.Y(n_6384)
);

BUFx2_ASAP7_75t_SL g6385 ( 
.A(n_6190),
.Y(n_6385)
);

INVx1_ASAP7_75t_L g6386 ( 
.A(n_6305),
.Y(n_6386)
);

AND2x4_ASAP7_75t_L g6387 ( 
.A(n_6157),
.B(n_522),
.Y(n_6387)
);

OR2x2_ASAP7_75t_L g6388 ( 
.A(n_6213),
.B(n_42),
.Y(n_6388)
);

INVx1_ASAP7_75t_L g6389 ( 
.A(n_6132),
.Y(n_6389)
);

BUFx3_ASAP7_75t_L g6390 ( 
.A(n_6147),
.Y(n_6390)
);

AND2x2_ASAP7_75t_L g6391 ( 
.A(n_6221),
.B(n_42),
.Y(n_6391)
);

INVx1_ASAP7_75t_L g6392 ( 
.A(n_6141),
.Y(n_6392)
);

HB1xp67_ASAP7_75t_L g6393 ( 
.A(n_6149),
.Y(n_6393)
);

BUFx2_ASAP7_75t_L g6394 ( 
.A(n_6164),
.Y(n_6394)
);

AND2x2_ASAP7_75t_L g6395 ( 
.A(n_6237),
.B(n_6193),
.Y(n_6395)
);

HB1xp67_ASAP7_75t_L g6396 ( 
.A(n_6149),
.Y(n_6396)
);

OR2x2_ASAP7_75t_L g6397 ( 
.A(n_6131),
.B(n_6228),
.Y(n_6397)
);

NAND2xp5_ASAP7_75t_L g6398 ( 
.A(n_6192),
.B(n_42),
.Y(n_6398)
);

INVx1_ASAP7_75t_L g6399 ( 
.A(n_6144),
.Y(n_6399)
);

AND2x2_ASAP7_75t_L g6400 ( 
.A(n_6303),
.B(n_42),
.Y(n_6400)
);

HB1xp67_ASAP7_75t_L g6401 ( 
.A(n_6152),
.Y(n_6401)
);

AND2x2_ASAP7_75t_L g6402 ( 
.A(n_6308),
.B(n_523),
.Y(n_6402)
);

INVx3_ASAP7_75t_L g6403 ( 
.A(n_6134),
.Y(n_6403)
);

AND2x2_ASAP7_75t_L g6404 ( 
.A(n_6200),
.B(n_523),
.Y(n_6404)
);

BUFx3_ASAP7_75t_L g6405 ( 
.A(n_6134),
.Y(n_6405)
);

INVx4_ASAP7_75t_L g6406 ( 
.A(n_6169),
.Y(n_6406)
);

INVx2_ASAP7_75t_L g6407 ( 
.A(n_6263),
.Y(n_6407)
);

AND2x2_ASAP7_75t_L g6408 ( 
.A(n_6201),
.B(n_523),
.Y(n_6408)
);

INVx1_ASAP7_75t_L g6409 ( 
.A(n_6290),
.Y(n_6409)
);

NAND2xp5_ASAP7_75t_L g6410 ( 
.A(n_6250),
.B(n_524),
.Y(n_6410)
);

AOI22xp5_ASAP7_75t_L g6411 ( 
.A1(n_6187),
.A2(n_6243),
.B1(n_6188),
.B2(n_6148),
.Y(n_6411)
);

NAND2xp5_ASAP7_75t_L g6412 ( 
.A(n_6258),
.B(n_524),
.Y(n_6412)
);

OR2x2_ASAP7_75t_L g6413 ( 
.A(n_6226),
.B(n_524),
.Y(n_6413)
);

AO21x2_ASAP7_75t_L g6414 ( 
.A1(n_6212),
.A2(n_6231),
.B(n_6277),
.Y(n_6414)
);

INVx2_ASAP7_75t_L g6415 ( 
.A(n_6214),
.Y(n_6415)
);

AND2x4_ASAP7_75t_L g6416 ( 
.A(n_6159),
.B(n_525),
.Y(n_6416)
);

INVx2_ASAP7_75t_L g6417 ( 
.A(n_6217),
.Y(n_6417)
);

OR2x6_ASAP7_75t_L g6418 ( 
.A(n_6199),
.B(n_525),
.Y(n_6418)
);

INVx2_ASAP7_75t_L g6419 ( 
.A(n_6218),
.Y(n_6419)
);

BUFx2_ASAP7_75t_L g6420 ( 
.A(n_6288),
.Y(n_6420)
);

INVx1_ASAP7_75t_L g6421 ( 
.A(n_6207),
.Y(n_6421)
);

INVx1_ASAP7_75t_L g6422 ( 
.A(n_6205),
.Y(n_6422)
);

INVx2_ASAP7_75t_L g6423 ( 
.A(n_6195),
.Y(n_6423)
);

INVxp67_ASAP7_75t_L g6424 ( 
.A(n_6246),
.Y(n_6424)
);

INVx2_ASAP7_75t_L g6425 ( 
.A(n_6198),
.Y(n_6425)
);

INVx1_ASAP7_75t_L g6426 ( 
.A(n_6219),
.Y(n_6426)
);

HB1xp67_ASAP7_75t_L g6427 ( 
.A(n_6256),
.Y(n_6427)
);

INVx1_ASAP7_75t_L g6428 ( 
.A(n_6229),
.Y(n_6428)
);

AND2x4_ASAP7_75t_L g6429 ( 
.A(n_6166),
.B(n_526),
.Y(n_6429)
);

OR2x2_ASAP7_75t_L g6430 ( 
.A(n_6227),
.B(n_526),
.Y(n_6430)
);

INVx3_ASAP7_75t_L g6431 ( 
.A(n_6189),
.Y(n_6431)
);

NOR2xp67_ASAP7_75t_L g6432 ( 
.A(n_6194),
.B(n_527),
.Y(n_6432)
);

BUFx3_ASAP7_75t_L g6433 ( 
.A(n_6267),
.Y(n_6433)
);

NAND2xp5_ASAP7_75t_L g6434 ( 
.A(n_6298),
.B(n_6244),
.Y(n_6434)
);

INVx2_ASAP7_75t_L g6435 ( 
.A(n_6225),
.Y(n_6435)
);

INVx2_ASAP7_75t_L g6436 ( 
.A(n_6236),
.Y(n_6436)
);

INVx1_ASAP7_75t_L g6437 ( 
.A(n_6274),
.Y(n_6437)
);

AND2x2_ASAP7_75t_L g6438 ( 
.A(n_6215),
.B(n_527),
.Y(n_6438)
);

AND2x2_ASAP7_75t_L g6439 ( 
.A(n_6254),
.B(n_527),
.Y(n_6439)
);

INVx1_ASAP7_75t_L g6440 ( 
.A(n_6267),
.Y(n_6440)
);

AOI22xp33_ASAP7_75t_L g6441 ( 
.A1(n_6254),
.A2(n_6296),
.B1(n_6239),
.B2(n_6233),
.Y(n_6441)
);

NAND2x1_ASAP7_75t_L g6442 ( 
.A(n_6238),
.B(n_528),
.Y(n_6442)
);

HB1xp67_ASAP7_75t_L g6443 ( 
.A(n_6299),
.Y(n_6443)
);

INVxp67_ASAP7_75t_SL g6444 ( 
.A(n_6146),
.Y(n_6444)
);

AND2x4_ASAP7_75t_L g6445 ( 
.A(n_6273),
.B(n_528),
.Y(n_6445)
);

OR2x2_ASAP7_75t_L g6446 ( 
.A(n_6163),
.B(n_6281),
.Y(n_6446)
);

NAND2xp5_ASAP7_75t_L g6447 ( 
.A(n_6242),
.B(n_528),
.Y(n_6447)
);

OR2x2_ASAP7_75t_L g6448 ( 
.A(n_6284),
.B(n_529),
.Y(n_6448)
);

BUFx3_ASAP7_75t_L g6449 ( 
.A(n_6273),
.Y(n_6449)
);

INVx1_ASAP7_75t_L g6450 ( 
.A(n_6242),
.Y(n_6450)
);

INVx3_ASAP7_75t_L g6451 ( 
.A(n_6251),
.Y(n_6451)
);

NOR2x1_ASAP7_75t_L g6452 ( 
.A(n_6233),
.B(n_529),
.Y(n_6452)
);

INVxp67_ASAP7_75t_L g6453 ( 
.A(n_6275),
.Y(n_6453)
);

AND2x2_ASAP7_75t_L g6454 ( 
.A(n_6253),
.B(n_529),
.Y(n_6454)
);

AND2x2_ASAP7_75t_L g6455 ( 
.A(n_6255),
.B(n_530),
.Y(n_6455)
);

INVx1_ASAP7_75t_L g6456 ( 
.A(n_6222),
.Y(n_6456)
);

CKINVDCx5p33_ASAP7_75t_R g6457 ( 
.A(n_6230),
.Y(n_6457)
);

AND2x2_ASAP7_75t_L g6458 ( 
.A(n_6259),
.B(n_6264),
.Y(n_6458)
);

AND2x2_ASAP7_75t_L g6459 ( 
.A(n_6285),
.B(n_530),
.Y(n_6459)
);

CKINVDCx5p33_ASAP7_75t_R g6460 ( 
.A(n_6271),
.Y(n_6460)
);

INVx2_ASAP7_75t_L g6461 ( 
.A(n_6257),
.Y(n_6461)
);

INVxp67_ASAP7_75t_SL g6462 ( 
.A(n_6179),
.Y(n_6462)
);

AND2x2_ASAP7_75t_L g6463 ( 
.A(n_6280),
.B(n_531),
.Y(n_6463)
);

AO22x1_ASAP7_75t_L g6464 ( 
.A1(n_6224),
.A2(n_1050),
.B1(n_1051),
.B2(n_1049),
.Y(n_6464)
);

AND2x2_ASAP7_75t_L g6465 ( 
.A(n_6268),
.B(n_531),
.Y(n_6465)
);

INVx2_ASAP7_75t_L g6466 ( 
.A(n_6257),
.Y(n_6466)
);

INVxp67_ASAP7_75t_SL g6467 ( 
.A(n_6287),
.Y(n_6467)
);

HB1xp67_ASAP7_75t_L g6468 ( 
.A(n_6269),
.Y(n_6468)
);

INVx2_ASAP7_75t_SL g6469 ( 
.A(n_6279),
.Y(n_6469)
);

INVx2_ASAP7_75t_SL g6470 ( 
.A(n_6293),
.Y(n_6470)
);

INVx2_ASAP7_75t_L g6471 ( 
.A(n_6276),
.Y(n_6471)
);

INVx2_ASAP7_75t_SL g6472 ( 
.A(n_6220),
.Y(n_6472)
);

INVx1_ASAP7_75t_L g6473 ( 
.A(n_6222),
.Y(n_6473)
);

AND2x2_ASAP7_75t_L g6474 ( 
.A(n_6203),
.B(n_532),
.Y(n_6474)
);

INVx1_ASAP7_75t_L g6475 ( 
.A(n_6232),
.Y(n_6475)
);

HB1xp67_ASAP7_75t_L g6476 ( 
.A(n_6204),
.Y(n_6476)
);

INVx1_ASAP7_75t_L g6477 ( 
.A(n_6232),
.Y(n_6477)
);

HB1xp67_ASAP7_75t_L g6478 ( 
.A(n_6208),
.Y(n_6478)
);

INVx1_ASAP7_75t_L g6479 ( 
.A(n_6283),
.Y(n_6479)
);

INVx4_ASAP7_75t_SL g6480 ( 
.A(n_6209),
.Y(n_6480)
);

AND2x2_ASAP7_75t_L g6481 ( 
.A(n_6245),
.B(n_532),
.Y(n_6481)
);

INVx1_ASAP7_75t_L g6482 ( 
.A(n_6283),
.Y(n_6482)
);

INVx1_ASAP7_75t_L g6483 ( 
.A(n_6335),
.Y(n_6483)
);

OR2x2_ASAP7_75t_L g6484 ( 
.A(n_6398),
.B(n_6294),
.Y(n_6484)
);

INVx1_ASAP7_75t_SL g6485 ( 
.A(n_6309),
.Y(n_6485)
);

INVx2_ASAP7_75t_L g6486 ( 
.A(n_6322),
.Y(n_6486)
);

INVx2_ASAP7_75t_L g6487 ( 
.A(n_6325),
.Y(n_6487)
);

OR2x2_ASAP7_75t_L g6488 ( 
.A(n_6329),
.B(n_6247),
.Y(n_6488)
);

INVx2_ASAP7_75t_L g6489 ( 
.A(n_6313),
.Y(n_6489)
);

NOR2x1_ASAP7_75t_L g6490 ( 
.A(n_6311),
.B(n_6452),
.Y(n_6490)
);

INVx1_ASAP7_75t_L g6491 ( 
.A(n_6337),
.Y(n_6491)
);

BUFx2_ASAP7_75t_L g6492 ( 
.A(n_6344),
.Y(n_6492)
);

AOI21xp5_ASAP7_75t_L g6493 ( 
.A1(n_6462),
.A2(n_6171),
.B(n_6249),
.Y(n_6493)
);

INVx6_ASAP7_75t_L g6494 ( 
.A(n_6336),
.Y(n_6494)
);

AOI21xp5_ASAP7_75t_L g6495 ( 
.A1(n_6434),
.A2(n_6260),
.B(n_6252),
.Y(n_6495)
);

INVx2_ASAP7_75t_L g6496 ( 
.A(n_6361),
.Y(n_6496)
);

AND2x2_ASAP7_75t_L g6497 ( 
.A(n_6368),
.B(n_6272),
.Y(n_6497)
);

AND2x2_ASAP7_75t_L g6498 ( 
.A(n_6368),
.B(n_6278),
.Y(n_6498)
);

BUFx2_ASAP7_75t_L g6499 ( 
.A(n_6332),
.Y(n_6499)
);

OR2x6_ASAP7_75t_L g6500 ( 
.A(n_6385),
.B(n_6289),
.Y(n_6500)
);

INVx1_ASAP7_75t_L g6501 ( 
.A(n_6338),
.Y(n_6501)
);

INVx2_ASAP7_75t_L g6502 ( 
.A(n_6361),
.Y(n_6502)
);

NAND4xp25_ASAP7_75t_L g6503 ( 
.A(n_6411),
.B(n_6441),
.C(n_6333),
.D(n_6463),
.Y(n_6503)
);

HB1xp67_ASAP7_75t_L g6504 ( 
.A(n_6317),
.Y(n_6504)
);

INVx1_ASAP7_75t_L g6505 ( 
.A(n_6341),
.Y(n_6505)
);

INVx2_ASAP7_75t_L g6506 ( 
.A(n_6394),
.Y(n_6506)
);

INVx2_ASAP7_75t_L g6507 ( 
.A(n_6394),
.Y(n_6507)
);

A2O1A1Ixp33_ASAP7_75t_L g6508 ( 
.A1(n_6450),
.A2(n_6167),
.B(n_6289),
.C(n_6266),
.Y(n_6508)
);

INVx1_ASAP7_75t_SL g6509 ( 
.A(n_6382),
.Y(n_6509)
);

AOI21xp5_ASAP7_75t_L g6510 ( 
.A1(n_6357),
.A2(n_532),
.B(n_533),
.Y(n_6510)
);

AND2x2_ASAP7_75t_L g6511 ( 
.A(n_6395),
.B(n_1051),
.Y(n_6511)
);

INVx1_ASAP7_75t_L g6512 ( 
.A(n_6354),
.Y(n_6512)
);

INVx2_ASAP7_75t_L g6513 ( 
.A(n_6320),
.Y(n_6513)
);

NAND2xp5_ASAP7_75t_L g6514 ( 
.A(n_6372),
.B(n_533),
.Y(n_6514)
);

INVx1_ASAP7_75t_L g6515 ( 
.A(n_6326),
.Y(n_6515)
);

INVx2_ASAP7_75t_L g6516 ( 
.A(n_6387),
.Y(n_6516)
);

A2O1A1Ixp33_ASAP7_75t_L g6517 ( 
.A1(n_6375),
.A2(n_535),
.B(n_533),
.C(n_534),
.Y(n_6517)
);

INVxp67_ASAP7_75t_L g6518 ( 
.A(n_6314),
.Y(n_6518)
);

INVx1_ASAP7_75t_L g6519 ( 
.A(n_6383),
.Y(n_6519)
);

OR2x2_ASAP7_75t_L g6520 ( 
.A(n_6364),
.B(n_534),
.Y(n_6520)
);

INVxp67_ASAP7_75t_SL g6521 ( 
.A(n_6331),
.Y(n_6521)
);

OAI21xp5_ASAP7_75t_SL g6522 ( 
.A1(n_6465),
.A2(n_534),
.B(n_535),
.Y(n_6522)
);

INVx1_ASAP7_75t_L g6523 ( 
.A(n_6366),
.Y(n_6523)
);

INVx1_ASAP7_75t_L g6524 ( 
.A(n_6376),
.Y(n_6524)
);

AOI21xp5_ASAP7_75t_L g6525 ( 
.A1(n_6472),
.A2(n_535),
.B(n_536),
.Y(n_6525)
);

INVx1_ASAP7_75t_L g6526 ( 
.A(n_6334),
.Y(n_6526)
);

INVx2_ASAP7_75t_L g6527 ( 
.A(n_6387),
.Y(n_6527)
);

INVx2_ASAP7_75t_L g6528 ( 
.A(n_6451),
.Y(n_6528)
);

AND2x2_ASAP7_75t_L g6529 ( 
.A(n_6359),
.B(n_1060),
.Y(n_6529)
);

INVx1_ASAP7_75t_L g6530 ( 
.A(n_6356),
.Y(n_6530)
);

BUFx2_ASAP7_75t_L g6531 ( 
.A(n_6390),
.Y(n_6531)
);

INVx2_ASAP7_75t_L g6532 ( 
.A(n_6310),
.Y(n_6532)
);

INVx2_ASAP7_75t_L g6533 ( 
.A(n_6350),
.Y(n_6533)
);

HB1xp67_ASAP7_75t_L g6534 ( 
.A(n_6393),
.Y(n_6534)
);

INVx1_ASAP7_75t_L g6535 ( 
.A(n_6327),
.Y(n_6535)
);

INVx3_ASAP7_75t_L g6536 ( 
.A(n_6323),
.Y(n_6536)
);

INVx2_ASAP7_75t_L g6537 ( 
.A(n_6458),
.Y(n_6537)
);

HB1xp67_ASAP7_75t_L g6538 ( 
.A(n_6396),
.Y(n_6538)
);

INVx1_ASAP7_75t_SL g6539 ( 
.A(n_6420),
.Y(n_6539)
);

HB1xp67_ASAP7_75t_L g6540 ( 
.A(n_6427),
.Y(n_6540)
);

INVx1_ASAP7_75t_L g6541 ( 
.A(n_6384),
.Y(n_6541)
);

AO21x2_ASAP7_75t_L g6542 ( 
.A1(n_6414),
.A2(n_537),
.B(n_538),
.Y(n_6542)
);

AND2x2_ASAP7_75t_L g6543 ( 
.A(n_6362),
.B(n_1060),
.Y(n_6543)
);

A2O1A1Ixp33_ASAP7_75t_L g6544 ( 
.A1(n_6379),
.A2(n_539),
.B(n_537),
.C(n_538),
.Y(n_6544)
);

INVx1_ASAP7_75t_L g6545 ( 
.A(n_6384),
.Y(n_6545)
);

INVx1_ASAP7_75t_SL g6546 ( 
.A(n_6420),
.Y(n_6546)
);

INVx2_ASAP7_75t_L g6547 ( 
.A(n_6351),
.Y(n_6547)
);

NAND4xp25_ASAP7_75t_L g6548 ( 
.A(n_6371),
.B(n_540),
.C(n_538),
.D(n_539),
.Y(n_6548)
);

INVxp67_ASAP7_75t_L g6549 ( 
.A(n_6316),
.Y(n_6549)
);

AOI21xp33_ASAP7_75t_L g6550 ( 
.A1(n_6323),
.A2(n_539),
.B(n_540),
.Y(n_6550)
);

INVx1_ASAP7_75t_L g6551 ( 
.A(n_6377),
.Y(n_6551)
);

OAI21xp5_ASAP7_75t_L g6552 ( 
.A1(n_6358),
.A2(n_540),
.B(n_541),
.Y(n_6552)
);

INVx2_ASAP7_75t_L g6553 ( 
.A(n_6339),
.Y(n_6553)
);

NAND2xp5_ASAP7_75t_L g6554 ( 
.A(n_6464),
.B(n_541),
.Y(n_6554)
);

INVx2_ASAP7_75t_L g6555 ( 
.A(n_6340),
.Y(n_6555)
);

INVx2_ASAP7_75t_L g6556 ( 
.A(n_6431),
.Y(n_6556)
);

AOI21xp5_ASAP7_75t_L g6557 ( 
.A1(n_6355),
.A2(n_6367),
.B(n_6442),
.Y(n_6557)
);

NOR3xp33_ASAP7_75t_SL g6558 ( 
.A(n_6457),
.B(n_542),
.C(n_543),
.Y(n_6558)
);

INVx2_ASAP7_75t_L g6559 ( 
.A(n_6345),
.Y(n_6559)
);

NOR2x1p5_ASAP7_75t_L g6560 ( 
.A(n_6467),
.B(n_542),
.Y(n_6560)
);

A2O1A1Ixp33_ASAP7_75t_L g6561 ( 
.A1(n_6405),
.A2(n_545),
.B(n_543),
.C(n_544),
.Y(n_6561)
);

BUFx2_ASAP7_75t_L g6562 ( 
.A(n_6433),
.Y(n_6562)
);

INVx1_ASAP7_75t_L g6563 ( 
.A(n_6349),
.Y(n_6563)
);

HB1xp67_ASAP7_75t_L g6564 ( 
.A(n_6389),
.Y(n_6564)
);

AO21x2_ASAP7_75t_L g6565 ( 
.A1(n_6347),
.A2(n_544),
.B(n_545),
.Y(n_6565)
);

NAND2xp5_ASAP7_75t_L g6566 ( 
.A(n_6438),
.B(n_544),
.Y(n_6566)
);

OR2x2_ASAP7_75t_L g6567 ( 
.A(n_6315),
.B(n_545),
.Y(n_6567)
);

AND2x4_ASAP7_75t_L g6568 ( 
.A(n_6449),
.B(n_546),
.Y(n_6568)
);

BUFx2_ASAP7_75t_L g6569 ( 
.A(n_6403),
.Y(n_6569)
);

AOI21xp5_ASAP7_75t_L g6570 ( 
.A1(n_6346),
.A2(n_546),
.B(n_547),
.Y(n_6570)
);

OA21x2_ASAP7_75t_L g6571 ( 
.A1(n_6424),
.A2(n_546),
.B(n_547),
.Y(n_6571)
);

INVx1_ASAP7_75t_L g6572 ( 
.A(n_6401),
.Y(n_6572)
);

AND2x2_ASAP7_75t_L g6573 ( 
.A(n_6406),
.B(n_1049),
.Y(n_6573)
);

A2O1A1Ixp33_ASAP7_75t_L g6574 ( 
.A1(n_6374),
.A2(n_550),
.B(n_547),
.C(n_549),
.Y(n_6574)
);

BUFx3_ASAP7_75t_L g6575 ( 
.A(n_6336),
.Y(n_6575)
);

INVx1_ASAP7_75t_L g6576 ( 
.A(n_6468),
.Y(n_6576)
);

A2O1A1Ixp33_ASAP7_75t_L g6577 ( 
.A1(n_6342),
.A2(n_551),
.B(n_549),
.C(n_550),
.Y(n_6577)
);

INVx4_ASAP7_75t_L g6578 ( 
.A(n_6336),
.Y(n_6578)
);

INVx1_ASAP7_75t_L g6579 ( 
.A(n_6392),
.Y(n_6579)
);

OA21x2_ASAP7_75t_L g6580 ( 
.A1(n_6352),
.A2(n_550),
.B(n_551),
.Y(n_6580)
);

INVx2_ASAP7_75t_SL g6581 ( 
.A(n_6407),
.Y(n_6581)
);

OA21x2_ASAP7_75t_L g6582 ( 
.A1(n_6353),
.A2(n_551),
.B(n_552),
.Y(n_6582)
);

CKINVDCx5p33_ASAP7_75t_R g6583 ( 
.A(n_6418),
.Y(n_6583)
);

OAI21xp5_ASAP7_75t_L g6584 ( 
.A1(n_6443),
.A2(n_6444),
.B(n_6343),
.Y(n_6584)
);

NAND2xp5_ASAP7_75t_L g6585 ( 
.A(n_6318),
.B(n_552),
.Y(n_6585)
);

INVxp67_ASAP7_75t_L g6586 ( 
.A(n_6381),
.Y(n_6586)
);

INVx2_ASAP7_75t_L g6587 ( 
.A(n_6415),
.Y(n_6587)
);

INVx1_ASAP7_75t_L g6588 ( 
.A(n_6391),
.Y(n_6588)
);

O2A1O1Ixp33_ASAP7_75t_L g6589 ( 
.A1(n_6447),
.A2(n_554),
.B(n_552),
.C(n_553),
.Y(n_6589)
);

INVx2_ASAP7_75t_L g6590 ( 
.A(n_6417),
.Y(n_6590)
);

INVx1_ASAP7_75t_L g6591 ( 
.A(n_6422),
.Y(n_6591)
);

INVx1_ASAP7_75t_SL g6592 ( 
.A(n_6369),
.Y(n_6592)
);

INVx1_ASAP7_75t_L g6593 ( 
.A(n_6416),
.Y(n_6593)
);

AND2x2_ASAP7_75t_L g6594 ( 
.A(n_6428),
.B(n_1061),
.Y(n_6594)
);

OAI21xp5_ASAP7_75t_L g6595 ( 
.A1(n_6453),
.A2(n_553),
.B(n_554),
.Y(n_6595)
);

AOI21xp5_ASAP7_75t_L g6596 ( 
.A1(n_6440),
.A2(n_553),
.B(n_554),
.Y(n_6596)
);

INVx2_ASAP7_75t_L g6597 ( 
.A(n_6419),
.Y(n_6597)
);

OAI21xp5_ASAP7_75t_L g6598 ( 
.A1(n_6432),
.A2(n_555),
.B(n_556),
.Y(n_6598)
);

INVx1_ASAP7_75t_L g6599 ( 
.A(n_6416),
.Y(n_6599)
);

OAI21x1_ASAP7_75t_L g6600 ( 
.A1(n_6437),
.A2(n_555),
.B(n_556),
.Y(n_6600)
);

NAND4xp25_ASAP7_75t_L g6601 ( 
.A(n_6348),
.B(n_557),
.C(n_555),
.D(n_556),
.Y(n_6601)
);

INVxp67_ASAP7_75t_SL g6602 ( 
.A(n_6410),
.Y(n_6602)
);

INVx2_ASAP7_75t_L g6603 ( 
.A(n_6423),
.Y(n_6603)
);

OA21x2_ASAP7_75t_L g6604 ( 
.A1(n_6460),
.A2(n_557),
.B(n_558),
.Y(n_6604)
);

AOI21xp5_ASAP7_75t_L g6605 ( 
.A1(n_6412),
.A2(n_558),
.B(n_559),
.Y(n_6605)
);

INVx1_ASAP7_75t_L g6606 ( 
.A(n_6429),
.Y(n_6606)
);

NAND3xp33_ASAP7_75t_L g6607 ( 
.A(n_6425),
.B(n_558),
.C(n_559),
.Y(n_6607)
);

AND2x6_ASAP7_75t_SL g6608 ( 
.A(n_6418),
.B(n_559),
.Y(n_6608)
);

INVx1_ASAP7_75t_L g6609 ( 
.A(n_6429),
.Y(n_6609)
);

AO21x2_ASAP7_75t_L g6610 ( 
.A1(n_6479),
.A2(n_560),
.B(n_561),
.Y(n_6610)
);

INVx2_ASAP7_75t_L g6611 ( 
.A(n_6435),
.Y(n_6611)
);

A2O1A1Ixp33_ASAP7_75t_L g6612 ( 
.A1(n_6363),
.A2(n_562),
.B(n_560),
.C(n_561),
.Y(n_6612)
);

NAND2x1_ASAP7_75t_L g6613 ( 
.A(n_6436),
.B(n_560),
.Y(n_6613)
);

INVx1_ASAP7_75t_L g6614 ( 
.A(n_6454),
.Y(n_6614)
);

INVx1_ASAP7_75t_L g6615 ( 
.A(n_6455),
.Y(n_6615)
);

AND2x2_ASAP7_75t_L g6616 ( 
.A(n_6399),
.B(n_1046),
.Y(n_6616)
);

INVx2_ASAP7_75t_L g6617 ( 
.A(n_6369),
.Y(n_6617)
);

INVx4_ASAP7_75t_L g6618 ( 
.A(n_6360),
.Y(n_6618)
);

AND2x4_ASAP7_75t_L g6619 ( 
.A(n_6360),
.B(n_561),
.Y(n_6619)
);

OAI21x1_ASAP7_75t_L g6620 ( 
.A1(n_6461),
.A2(n_562),
.B(n_563),
.Y(n_6620)
);

INVx1_ASAP7_75t_L g6621 ( 
.A(n_6388),
.Y(n_6621)
);

AO21x2_ASAP7_75t_L g6622 ( 
.A1(n_6482),
.A2(n_562),
.B(n_563),
.Y(n_6622)
);

NAND2xp5_ASAP7_75t_SL g6623 ( 
.A(n_6480),
.B(n_6446),
.Y(n_6623)
);

AOI21xp5_ASAP7_75t_L g6624 ( 
.A1(n_6373),
.A2(n_564),
.B(n_565),
.Y(n_6624)
);

INVx1_ASAP7_75t_L g6625 ( 
.A(n_6324),
.Y(n_6625)
);

NAND2xp5_ASAP7_75t_L g6626 ( 
.A(n_6409),
.B(n_564),
.Y(n_6626)
);

INVx2_ASAP7_75t_L g6627 ( 
.A(n_6445),
.Y(n_6627)
);

A2O1A1Ixp33_ASAP7_75t_L g6628 ( 
.A1(n_6378),
.A2(n_566),
.B(n_564),
.C(n_565),
.Y(n_6628)
);

BUFx6f_ASAP7_75t_L g6629 ( 
.A(n_6445),
.Y(n_6629)
);

INVx1_ASAP7_75t_L g6630 ( 
.A(n_6328),
.Y(n_6630)
);

INVx1_ASAP7_75t_L g6631 ( 
.A(n_6404),
.Y(n_6631)
);

AOI21xp5_ASAP7_75t_L g6632 ( 
.A1(n_6469),
.A2(n_566),
.B(n_567),
.Y(n_6632)
);

NAND2xp5_ASAP7_75t_L g6633 ( 
.A(n_6421),
.B(n_6426),
.Y(n_6633)
);

HB1xp67_ASAP7_75t_L g6634 ( 
.A(n_6476),
.Y(n_6634)
);

A2O1A1Ixp33_ASAP7_75t_L g6635 ( 
.A1(n_6380),
.A2(n_568),
.B(n_566),
.C(n_567),
.Y(n_6635)
);

INVx1_ASAP7_75t_L g6636 ( 
.A(n_6408),
.Y(n_6636)
);

INVx2_ASAP7_75t_L g6637 ( 
.A(n_6470),
.Y(n_6637)
);

HB1xp67_ASAP7_75t_L g6638 ( 
.A(n_6478),
.Y(n_6638)
);

OAI21x1_ASAP7_75t_L g6639 ( 
.A1(n_6466),
.A2(n_567),
.B(n_568),
.Y(n_6639)
);

INVx2_ASAP7_75t_SL g6640 ( 
.A(n_6459),
.Y(n_6640)
);

INVx1_ASAP7_75t_L g6641 ( 
.A(n_6413),
.Y(n_6641)
);

INVx1_ASAP7_75t_L g6642 ( 
.A(n_6312),
.Y(n_6642)
);

OAI21x1_ASAP7_75t_L g6643 ( 
.A1(n_6471),
.A2(n_6475),
.B(n_6473),
.Y(n_6643)
);

NAND2xp5_ASAP7_75t_L g6644 ( 
.A(n_6386),
.B(n_569),
.Y(n_6644)
);

A2O1A1Ixp33_ASAP7_75t_L g6645 ( 
.A1(n_6397),
.A2(n_571),
.B(n_569),
.C(n_570),
.Y(n_6645)
);

INVx1_ASAP7_75t_L g6646 ( 
.A(n_6448),
.Y(n_6646)
);

NAND2xp5_ASAP7_75t_L g6647 ( 
.A(n_6474),
.B(n_570),
.Y(n_6647)
);

INVx1_ASAP7_75t_L g6648 ( 
.A(n_6481),
.Y(n_6648)
);

AO21x1_ASAP7_75t_L g6649 ( 
.A1(n_6456),
.A2(n_572),
.B(n_571),
.Y(n_6649)
);

OAI21x1_ASAP7_75t_L g6650 ( 
.A1(n_6477),
.A2(n_570),
.B(n_572),
.Y(n_6650)
);

OR2x2_ASAP7_75t_L g6651 ( 
.A(n_6319),
.B(n_572),
.Y(n_6651)
);

AND2x2_ASAP7_75t_L g6652 ( 
.A(n_6400),
.B(n_6370),
.Y(n_6652)
);

INVxp67_ASAP7_75t_L g6653 ( 
.A(n_6365),
.Y(n_6653)
);

AOI21xp5_ASAP7_75t_L g6654 ( 
.A1(n_6321),
.A2(n_573),
.B(n_574),
.Y(n_6654)
);

BUFx3_ASAP7_75t_L g6655 ( 
.A(n_6402),
.Y(n_6655)
);

BUFx2_ASAP7_75t_L g6656 ( 
.A(n_6480),
.Y(n_6656)
);

INVx2_ASAP7_75t_SL g6657 ( 
.A(n_6439),
.Y(n_6657)
);

INVx3_ASAP7_75t_L g6658 ( 
.A(n_6430),
.Y(n_6658)
);

INVx1_ASAP7_75t_L g6659 ( 
.A(n_6330),
.Y(n_6659)
);

AO21x1_ASAP7_75t_L g6660 ( 
.A1(n_6311),
.A2(n_576),
.B(n_575),
.Y(n_6660)
);

INVxp67_ASAP7_75t_L g6661 ( 
.A(n_6309),
.Y(n_6661)
);

OAI21xp5_ASAP7_75t_L g6662 ( 
.A1(n_6411),
.A2(n_573),
.B(n_575),
.Y(n_6662)
);

INVx1_ASAP7_75t_L g6663 ( 
.A(n_6335),
.Y(n_6663)
);

INVx2_ASAP7_75t_L g6664 ( 
.A(n_6309),
.Y(n_6664)
);

HB1xp67_ASAP7_75t_L g6665 ( 
.A(n_6317),
.Y(n_6665)
);

HB1xp67_ASAP7_75t_L g6666 ( 
.A(n_6317),
.Y(n_6666)
);

INVx3_ASAP7_75t_SL g6667 ( 
.A(n_6311),
.Y(n_6667)
);

INVx1_ASAP7_75t_L g6668 ( 
.A(n_6335),
.Y(n_6668)
);

INVx2_ASAP7_75t_SL g6669 ( 
.A(n_6309),
.Y(n_6669)
);

OR2x2_ASAP7_75t_L g6670 ( 
.A(n_6398),
.B(n_573),
.Y(n_6670)
);

INVx1_ASAP7_75t_L g6671 ( 
.A(n_6335),
.Y(n_6671)
);

INVx1_ASAP7_75t_L g6672 ( 
.A(n_6335),
.Y(n_6672)
);

OA21x2_ASAP7_75t_L g6673 ( 
.A1(n_6398),
.A2(n_575),
.B(n_576),
.Y(n_6673)
);

INVx2_ASAP7_75t_L g6674 ( 
.A(n_6309),
.Y(n_6674)
);

OA21x2_ASAP7_75t_L g6675 ( 
.A1(n_6398),
.A2(n_576),
.B(n_577),
.Y(n_6675)
);

INVx1_ASAP7_75t_L g6676 ( 
.A(n_6335),
.Y(n_6676)
);

OA21x2_ASAP7_75t_L g6677 ( 
.A1(n_6398),
.A2(n_578),
.B(n_579),
.Y(n_6677)
);

OR2x2_ASAP7_75t_L g6678 ( 
.A(n_6398),
.B(n_578),
.Y(n_6678)
);

INVx4_ASAP7_75t_L g6679 ( 
.A(n_6309),
.Y(n_6679)
);

INVx1_ASAP7_75t_L g6680 ( 
.A(n_6335),
.Y(n_6680)
);

AND4x1_ASAP7_75t_L g6681 ( 
.A(n_6357),
.B(n_581),
.C(n_579),
.D(n_580),
.Y(n_6681)
);

INVx1_ASAP7_75t_L g6682 ( 
.A(n_6335),
.Y(n_6682)
);

AND2x4_ASAP7_75t_L g6683 ( 
.A(n_6309),
.B(n_580),
.Y(n_6683)
);

AO21x2_ASAP7_75t_L g6684 ( 
.A1(n_6411),
.A2(n_580),
.B(n_581),
.Y(n_6684)
);

AND2x2_ASAP7_75t_L g6685 ( 
.A(n_6492),
.B(n_581),
.Y(n_6685)
);

AND2x2_ASAP7_75t_L g6686 ( 
.A(n_6667),
.B(n_582),
.Y(n_6686)
);

AND2x2_ASAP7_75t_L g6687 ( 
.A(n_6679),
.B(n_582),
.Y(n_6687)
);

NOR3xp33_ASAP7_75t_L g6688 ( 
.A(n_6661),
.B(n_584),
.C(n_583),
.Y(n_6688)
);

INVx2_ASAP7_75t_SL g6689 ( 
.A(n_6664),
.Y(n_6689)
);

XNOR2x1_ASAP7_75t_L g6690 ( 
.A(n_6485),
.B(n_582),
.Y(n_6690)
);

AND2x2_ASAP7_75t_L g6691 ( 
.A(n_6669),
.B(n_583),
.Y(n_6691)
);

NOR2xp33_ASAP7_75t_L g6692 ( 
.A(n_6509),
.B(n_6674),
.Y(n_6692)
);

NAND3xp33_ASAP7_75t_L g6693 ( 
.A(n_6489),
.B(n_583),
.C(n_584),
.Y(n_6693)
);

NAND3xp33_ASAP7_75t_L g6694 ( 
.A(n_6578),
.B(n_585),
.C(n_586),
.Y(n_6694)
);

NAND3xp33_ASAP7_75t_L g6695 ( 
.A(n_6486),
.B(n_585),
.C(n_586),
.Y(n_6695)
);

XNOR2xp5_ASAP7_75t_L g6696 ( 
.A(n_6681),
.B(n_586),
.Y(n_6696)
);

NAND2xp5_ASAP7_75t_L g6697 ( 
.A(n_6539),
.B(n_6546),
.Y(n_6697)
);

AND2x2_ASAP7_75t_L g6698 ( 
.A(n_6499),
.B(n_587),
.Y(n_6698)
);

AOI22xp33_ASAP7_75t_L g6699 ( 
.A1(n_6562),
.A2(n_589),
.B1(n_587),
.B2(n_588),
.Y(n_6699)
);

AO21x2_ASAP7_75t_L g6700 ( 
.A1(n_6542),
.A2(n_587),
.B(n_588),
.Y(n_6700)
);

AND2x2_ASAP7_75t_L g6701 ( 
.A(n_6531),
.B(n_588),
.Y(n_6701)
);

INVx3_ASAP7_75t_L g6702 ( 
.A(n_6575),
.Y(n_6702)
);

OR2x2_ASAP7_75t_L g6703 ( 
.A(n_6520),
.B(n_589),
.Y(n_6703)
);

BUFx2_ASAP7_75t_L g6704 ( 
.A(n_6656),
.Y(n_6704)
);

INVx1_ASAP7_75t_L g6705 ( 
.A(n_6504),
.Y(n_6705)
);

NOR4xp25_ASAP7_75t_L g6706 ( 
.A(n_6503),
.B(n_1044),
.C(n_1045),
.D(n_1043),
.Y(n_6706)
);

OR2x2_ASAP7_75t_L g6707 ( 
.A(n_6541),
.B(n_590),
.Y(n_6707)
);

AOI22xp5_ASAP7_75t_L g6708 ( 
.A1(n_6583),
.A2(n_592),
.B1(n_590),
.B2(n_591),
.Y(n_6708)
);

INVx2_ASAP7_75t_L g6709 ( 
.A(n_6496),
.Y(n_6709)
);

NAND3xp33_ASAP7_75t_L g6710 ( 
.A(n_6662),
.B(n_590),
.C(n_591),
.Y(n_6710)
);

NOR2x1_ASAP7_75t_SL g6711 ( 
.A(n_6500),
.B(n_591),
.Y(n_6711)
);

NAND4xp25_ASAP7_75t_L g6712 ( 
.A(n_6490),
.B(n_594),
.C(n_592),
.D(n_593),
.Y(n_6712)
);

NAND2xp5_ASAP7_75t_L g6713 ( 
.A(n_6521),
.B(n_592),
.Y(n_6713)
);

AOI22xp33_ASAP7_75t_L g6714 ( 
.A1(n_6569),
.A2(n_6581),
.B1(n_6556),
.B2(n_6533),
.Y(n_6714)
);

AOI22xp33_ASAP7_75t_L g6715 ( 
.A1(n_6637),
.A2(n_596),
.B1(n_593),
.B2(n_595),
.Y(n_6715)
);

AOI22xp5_ASAP7_75t_L g6716 ( 
.A1(n_6537),
.A2(n_597),
.B1(n_595),
.B2(n_596),
.Y(n_6716)
);

AND2x2_ASAP7_75t_L g6717 ( 
.A(n_6652),
.B(n_596),
.Y(n_6717)
);

AND2x2_ASAP7_75t_SL g6718 ( 
.A(n_6618),
.B(n_597),
.Y(n_6718)
);

HB1xp67_ASAP7_75t_L g6719 ( 
.A(n_6665),
.Y(n_6719)
);

NOR2xp33_ASAP7_75t_L g6720 ( 
.A(n_6494),
.B(n_598),
.Y(n_6720)
);

INVx1_ASAP7_75t_L g6721 ( 
.A(n_6666),
.Y(n_6721)
);

AND2x2_ASAP7_75t_L g6722 ( 
.A(n_6511),
.B(n_598),
.Y(n_6722)
);

NAND3xp33_ASAP7_75t_L g6723 ( 
.A(n_6536),
.B(n_6545),
.C(n_6540),
.Y(n_6723)
);

AND2x2_ASAP7_75t_L g6724 ( 
.A(n_6529),
.B(n_598),
.Y(n_6724)
);

INVx2_ASAP7_75t_L g6725 ( 
.A(n_6502),
.Y(n_6725)
);

NOR2xp33_ASAP7_75t_L g6726 ( 
.A(n_6494),
.B(n_599),
.Y(n_6726)
);

OAI211xp5_ASAP7_75t_L g6727 ( 
.A1(n_6623),
.A2(n_601),
.B(n_599),
.C(n_600),
.Y(n_6727)
);

AOI22xp33_ASAP7_75t_SL g6728 ( 
.A1(n_6553),
.A2(n_601),
.B1(n_599),
.B2(n_600),
.Y(n_6728)
);

AND2x4_ASAP7_75t_SL g6729 ( 
.A(n_6513),
.B(n_600),
.Y(n_6729)
);

NAND3xp33_ASAP7_75t_L g6730 ( 
.A(n_6523),
.B(n_602),
.C(n_603),
.Y(n_6730)
);

AOI211x1_ASAP7_75t_L g6731 ( 
.A1(n_6493),
.A2(n_605),
.B(n_603),
.C(n_604),
.Y(n_6731)
);

NAND3xp33_ASAP7_75t_L g6732 ( 
.A(n_6524),
.B(n_6538),
.C(n_6534),
.Y(n_6732)
);

AND2x2_ASAP7_75t_L g6733 ( 
.A(n_6616),
.B(n_603),
.Y(n_6733)
);

NAND4xp75_ASAP7_75t_L g6734 ( 
.A(n_6584),
.B(n_612),
.C(n_620),
.D(n_604),
.Y(n_6734)
);

NOR3xp33_ASAP7_75t_L g6735 ( 
.A(n_6589),
.B(n_6607),
.C(n_6554),
.Y(n_6735)
);

INVx1_ASAP7_75t_L g6736 ( 
.A(n_6543),
.Y(n_6736)
);

NOR2x1_ASAP7_75t_L g6737 ( 
.A(n_6604),
.B(n_605),
.Y(n_6737)
);

OR2x2_ASAP7_75t_L g6738 ( 
.A(n_6547),
.B(n_605),
.Y(n_6738)
);

NOR3xp33_ASAP7_75t_L g6739 ( 
.A(n_6549),
.B(n_608),
.C(n_607),
.Y(n_6739)
);

INVx3_ASAP7_75t_L g6740 ( 
.A(n_6568),
.Y(n_6740)
);

AND2x4_ASAP7_75t_L g6741 ( 
.A(n_6555),
.B(n_606),
.Y(n_6741)
);

AOI21xp5_ASAP7_75t_SL g6742 ( 
.A1(n_6604),
.A2(n_1044),
.B(n_1043),
.Y(n_6742)
);

OA211x2_ASAP7_75t_L g6743 ( 
.A1(n_6613),
.A2(n_608),
.B(n_606),
.C(n_607),
.Y(n_6743)
);

HB1xp67_ASAP7_75t_L g6744 ( 
.A(n_6564),
.Y(n_6744)
);

NAND4xp75_ASAP7_75t_L g6745 ( 
.A(n_6572),
.B(n_616),
.C(n_624),
.D(n_608),
.Y(n_6745)
);

NAND3xp33_ASAP7_75t_L g6746 ( 
.A(n_6526),
.B(n_609),
.C(n_610),
.Y(n_6746)
);

AND2x2_ASAP7_75t_L g6747 ( 
.A(n_6594),
.B(n_609),
.Y(n_6747)
);

NAND3xp33_ASAP7_75t_L g6748 ( 
.A(n_6530),
.B(n_610),
.C(n_611),
.Y(n_6748)
);

AND2x4_ASAP7_75t_L g6749 ( 
.A(n_6559),
.B(n_610),
.Y(n_6749)
);

NAND3xp33_ASAP7_75t_L g6750 ( 
.A(n_6629),
.B(n_611),
.C(n_612),
.Y(n_6750)
);

NOR3xp33_ASAP7_75t_L g6751 ( 
.A(n_6508),
.B(n_614),
.C(n_613),
.Y(n_6751)
);

OR2x2_ASAP7_75t_SL g6752 ( 
.A(n_6506),
.B(n_612),
.Y(n_6752)
);

BUFx2_ASAP7_75t_L g6753 ( 
.A(n_6500),
.Y(n_6753)
);

NAND4xp25_ASAP7_75t_L g6754 ( 
.A(n_6557),
.B(n_615),
.C(n_613),
.D(n_614),
.Y(n_6754)
);

NAND2xp5_ASAP7_75t_L g6755 ( 
.A(n_6525),
.B(n_614),
.Y(n_6755)
);

INVx2_ASAP7_75t_L g6756 ( 
.A(n_6507),
.Y(n_6756)
);

NAND2xp5_ASAP7_75t_L g6757 ( 
.A(n_6573),
.B(n_615),
.Y(n_6757)
);

NOR3xp33_ASAP7_75t_L g6758 ( 
.A(n_6552),
.B(n_6548),
.C(n_6544),
.Y(n_6758)
);

AND2x2_ASAP7_75t_L g6759 ( 
.A(n_6655),
.B(n_615),
.Y(n_6759)
);

NAND2xp5_ASAP7_75t_SL g6760 ( 
.A(n_6660),
.B(n_616),
.Y(n_6760)
);

OAI221xp5_ASAP7_75t_L g6761 ( 
.A1(n_6518),
.A2(n_618),
.B1(n_616),
.B2(n_617),
.C(n_619),
.Y(n_6761)
);

OAI211xp5_ASAP7_75t_L g6762 ( 
.A1(n_6576),
.A2(n_619),
.B(n_617),
.C(n_618),
.Y(n_6762)
);

INVx1_ASAP7_75t_L g6763 ( 
.A(n_6634),
.Y(n_6763)
);

NOR2xp33_ASAP7_75t_L g6764 ( 
.A(n_6592),
.B(n_618),
.Y(n_6764)
);

INVx1_ASAP7_75t_L g6765 ( 
.A(n_6638),
.Y(n_6765)
);

AOI211xp5_ASAP7_75t_L g6766 ( 
.A1(n_6528),
.A2(n_621),
.B(n_619),
.C(n_620),
.Y(n_6766)
);

AOI211xp5_ASAP7_75t_L g6767 ( 
.A1(n_6519),
.A2(n_623),
.B(n_621),
.C(n_622),
.Y(n_6767)
);

NOR2xp33_ASAP7_75t_L g6768 ( 
.A(n_6608),
.B(n_621),
.Y(n_6768)
);

OR2x2_ASAP7_75t_L g6769 ( 
.A(n_6535),
.B(n_622),
.Y(n_6769)
);

NAND3xp33_ASAP7_75t_L g6770 ( 
.A(n_6629),
.B(n_622),
.C(n_623),
.Y(n_6770)
);

NOR2xp33_ASAP7_75t_L g6771 ( 
.A(n_6653),
.B(n_623),
.Y(n_6771)
);

INVx1_ASAP7_75t_L g6772 ( 
.A(n_6651),
.Y(n_6772)
);

NAND3xp33_ASAP7_75t_L g6773 ( 
.A(n_6571),
.B(n_624),
.C(n_625),
.Y(n_6773)
);

AND4x1_ASAP7_75t_L g6774 ( 
.A(n_6558),
.B(n_1048),
.C(n_1050),
.D(n_1047),
.Y(n_6774)
);

INVx1_ASAP7_75t_L g6775 ( 
.A(n_6532),
.Y(n_6775)
);

AND2x4_ASAP7_75t_L g6776 ( 
.A(n_6516),
.B(n_624),
.Y(n_6776)
);

NAND2xp5_ASAP7_75t_SL g6777 ( 
.A(n_6587),
.B(n_625),
.Y(n_6777)
);

OAI21xp5_ASAP7_75t_L g6778 ( 
.A1(n_6586),
.A2(n_626),
.B(n_627),
.Y(n_6778)
);

NAND4xp75_ASAP7_75t_L g6779 ( 
.A(n_6497),
.B(n_6498),
.C(n_6591),
.D(n_6551),
.Y(n_6779)
);

AOI22xp33_ASAP7_75t_L g6780 ( 
.A1(n_6641),
.A2(n_628),
.B1(n_626),
.B2(n_627),
.Y(n_6780)
);

AOI22xp33_ASAP7_75t_L g6781 ( 
.A1(n_6646),
.A2(n_629),
.B1(n_627),
.B2(n_628),
.Y(n_6781)
);

NAND3xp33_ASAP7_75t_L g6782 ( 
.A(n_6571),
.B(n_628),
.C(n_629),
.Y(n_6782)
);

NOR2xp33_ASAP7_75t_L g6783 ( 
.A(n_6483),
.B(n_629),
.Y(n_6783)
);

NOR2xp33_ASAP7_75t_L g6784 ( 
.A(n_6663),
.B(n_630),
.Y(n_6784)
);

OR2x2_ASAP7_75t_L g6785 ( 
.A(n_6567),
.B(n_630),
.Y(n_6785)
);

OR2x2_ASAP7_75t_L g6786 ( 
.A(n_6668),
.B(n_630),
.Y(n_6786)
);

AOI22xp33_ASAP7_75t_SL g6787 ( 
.A1(n_6684),
.A2(n_633),
.B1(n_631),
.B2(n_632),
.Y(n_6787)
);

BUFx3_ASAP7_75t_L g6788 ( 
.A(n_6683),
.Y(n_6788)
);

AND2x2_ASAP7_75t_L g6789 ( 
.A(n_6487),
.B(n_631),
.Y(n_6789)
);

NAND2xp5_ASAP7_75t_L g6790 ( 
.A(n_6632),
.B(n_631),
.Y(n_6790)
);

OA211x2_ASAP7_75t_L g6791 ( 
.A1(n_6595),
.A2(n_634),
.B(n_632),
.C(n_633),
.Y(n_6791)
);

NOR2xp33_ASAP7_75t_L g6792 ( 
.A(n_6671),
.B(n_633),
.Y(n_6792)
);

AOI22xp5_ASAP7_75t_L g6793 ( 
.A1(n_6672),
.A2(n_636),
.B1(n_634),
.B2(n_635),
.Y(n_6793)
);

NOR3xp33_ASAP7_75t_L g6794 ( 
.A(n_6517),
.B(n_636),
.C(n_635),
.Y(n_6794)
);

NAND4xp75_ASAP7_75t_L g6795 ( 
.A(n_6579),
.B(n_643),
.C(n_651),
.D(n_634),
.Y(n_6795)
);

OR2x2_ASAP7_75t_L g6796 ( 
.A(n_6676),
.B(n_636),
.Y(n_6796)
);

OAI211xp5_ASAP7_75t_SL g6797 ( 
.A1(n_6590),
.A2(n_639),
.B(n_637),
.C(n_638),
.Y(n_6797)
);

NAND4xp75_ASAP7_75t_L g6798 ( 
.A(n_6649),
.B(n_645),
.C(n_653),
.D(n_637),
.Y(n_6798)
);

AOI22xp5_ASAP7_75t_L g6799 ( 
.A1(n_6680),
.A2(n_639),
.B1(n_637),
.B2(n_638),
.Y(n_6799)
);

AOI211xp5_ASAP7_75t_L g6800 ( 
.A1(n_6621),
.A2(n_6599),
.B(n_6606),
.C(n_6593),
.Y(n_6800)
);

INVx2_ASAP7_75t_L g6801 ( 
.A(n_6597),
.Y(n_6801)
);

AND2x2_ASAP7_75t_L g6802 ( 
.A(n_6682),
.B(n_638),
.Y(n_6802)
);

NAND3xp33_ASAP7_75t_L g6803 ( 
.A(n_6574),
.B(n_640),
.C(n_641),
.Y(n_6803)
);

AND2x4_ASAP7_75t_L g6804 ( 
.A(n_6527),
.B(n_640),
.Y(n_6804)
);

OR2x6_ASAP7_75t_L g6805 ( 
.A(n_6617),
.B(n_640),
.Y(n_6805)
);

NAND3xp33_ASAP7_75t_L g6806 ( 
.A(n_6561),
.B(n_641),
.C(n_642),
.Y(n_6806)
);

AND2x2_ASAP7_75t_L g6807 ( 
.A(n_6627),
.B(n_642),
.Y(n_6807)
);

OA211x2_ASAP7_75t_L g6808 ( 
.A1(n_6626),
.A2(n_644),
.B(n_642),
.C(n_643),
.Y(n_6808)
);

INVx1_ASAP7_75t_L g6809 ( 
.A(n_6603),
.Y(n_6809)
);

AO21x2_ASAP7_75t_L g6810 ( 
.A1(n_6643),
.A2(n_644),
.B(n_645),
.Y(n_6810)
);

NAND2xp5_ASAP7_75t_L g6811 ( 
.A(n_6640),
.B(n_645),
.Y(n_6811)
);

AND2x2_ASAP7_75t_L g6812 ( 
.A(n_6491),
.B(n_646),
.Y(n_6812)
);

OAI211xp5_ASAP7_75t_L g6813 ( 
.A1(n_6602),
.A2(n_648),
.B(n_646),
.C(n_647),
.Y(n_6813)
);

INVx2_ASAP7_75t_SL g6814 ( 
.A(n_6611),
.Y(n_6814)
);

NOR3xp33_ASAP7_75t_L g6815 ( 
.A(n_6601),
.B(n_6550),
.C(n_6644),
.Y(n_6815)
);

NOR3xp33_ASAP7_75t_L g6816 ( 
.A(n_6628),
.B(n_649),
.C(n_648),
.Y(n_6816)
);

NOR3xp33_ASAP7_75t_L g6817 ( 
.A(n_6635),
.B(n_6645),
.C(n_6577),
.Y(n_6817)
);

AND2x2_ASAP7_75t_L g6818 ( 
.A(n_6501),
.B(n_647),
.Y(n_6818)
);

INVxp67_ASAP7_75t_SL g6819 ( 
.A(n_6514),
.Y(n_6819)
);

INVx1_ASAP7_75t_L g6820 ( 
.A(n_6582),
.Y(n_6820)
);

NAND2xp5_ASAP7_75t_L g6821 ( 
.A(n_6657),
.B(n_647),
.Y(n_6821)
);

OR2x2_ASAP7_75t_L g6822 ( 
.A(n_6512),
.B(n_648),
.Y(n_6822)
);

INVx4_ASAP7_75t_L g6823 ( 
.A(n_6619),
.Y(n_6823)
);

INVx1_ASAP7_75t_L g6824 ( 
.A(n_6582),
.Y(n_6824)
);

AOI22xp33_ASAP7_75t_L g6825 ( 
.A1(n_6658),
.A2(n_6642),
.B1(n_6659),
.B2(n_6609),
.Y(n_6825)
);

AO21x2_ASAP7_75t_L g6826 ( 
.A1(n_6495),
.A2(n_649),
.B(n_650),
.Y(n_6826)
);

AOI22xp33_ASAP7_75t_L g6827 ( 
.A1(n_6625),
.A2(n_651),
.B1(n_649),
.B2(n_650),
.Y(n_6827)
);

INVx1_ASAP7_75t_L g6828 ( 
.A(n_6600),
.Y(n_6828)
);

BUFx3_ASAP7_75t_L g6829 ( 
.A(n_6673),
.Y(n_6829)
);

INVx1_ASAP7_75t_L g6830 ( 
.A(n_6505),
.Y(n_6830)
);

AOI221xp5_ASAP7_75t_L g6831 ( 
.A1(n_6633),
.A2(n_653),
.B1(n_651),
.B2(n_652),
.C(n_654),
.Y(n_6831)
);

NAND4xp75_ASAP7_75t_L g6832 ( 
.A(n_6673),
.B(n_662),
.C(n_670),
.D(n_652),
.Y(n_6832)
);

NAND2xp5_ASAP7_75t_L g6833 ( 
.A(n_6563),
.B(n_654),
.Y(n_6833)
);

NAND2xp5_ASAP7_75t_L g6834 ( 
.A(n_6624),
.B(n_654),
.Y(n_6834)
);

AND2x2_ASAP7_75t_L g6835 ( 
.A(n_6515),
.B(n_655),
.Y(n_6835)
);

AOI22xp33_ASAP7_75t_L g6836 ( 
.A1(n_6630),
.A2(n_658),
.B1(n_656),
.B2(n_657),
.Y(n_6836)
);

NAND2xp33_ASAP7_75t_SL g6837 ( 
.A(n_6560),
.B(n_656),
.Y(n_6837)
);

AND2x2_ASAP7_75t_L g6838 ( 
.A(n_6631),
.B(n_657),
.Y(n_6838)
);

NAND3xp33_ASAP7_75t_L g6839 ( 
.A(n_6675),
.B(n_6677),
.C(n_6588),
.Y(n_6839)
);

OAI211xp5_ASAP7_75t_L g6840 ( 
.A1(n_6522),
.A2(n_661),
.B(n_657),
.C(n_660),
.Y(n_6840)
);

AND2x2_ASAP7_75t_SL g6841 ( 
.A(n_6580),
.B(n_660),
.Y(n_6841)
);

NOR2xp33_ASAP7_75t_L g6842 ( 
.A(n_6636),
.B(n_660),
.Y(n_6842)
);

NAND2xp5_ASAP7_75t_L g6843 ( 
.A(n_6596),
.B(n_661),
.Y(n_6843)
);

NAND3xp33_ASAP7_75t_L g6844 ( 
.A(n_6675),
.B(n_662),
.C(n_663),
.Y(n_6844)
);

OAI211xp5_ASAP7_75t_L g6845 ( 
.A1(n_6510),
.A2(n_665),
.B(n_662),
.C(n_664),
.Y(n_6845)
);

OR2x2_ASAP7_75t_L g6846 ( 
.A(n_6488),
.B(n_664),
.Y(n_6846)
);

CKINVDCx5p33_ASAP7_75t_R g6847 ( 
.A(n_6670),
.Y(n_6847)
);

INVx1_ASAP7_75t_L g6848 ( 
.A(n_6678),
.Y(n_6848)
);

AND2x2_ASAP7_75t_L g6849 ( 
.A(n_6614),
.B(n_664),
.Y(n_6849)
);

NOR2xp33_ASAP7_75t_L g6850 ( 
.A(n_6615),
.B(n_665),
.Y(n_6850)
);

NAND2xp5_ASAP7_75t_L g6851 ( 
.A(n_6654),
.B(n_665),
.Y(n_6851)
);

AND2x2_ASAP7_75t_L g6852 ( 
.A(n_6685),
.B(n_6648),
.Y(n_6852)
);

NAND2xp5_ASAP7_75t_L g6853 ( 
.A(n_6692),
.B(n_6570),
.Y(n_6853)
);

AND2x2_ASAP7_75t_L g6854 ( 
.A(n_6689),
.B(n_6677),
.Y(n_6854)
);

INVx1_ASAP7_75t_L g6855 ( 
.A(n_6686),
.Y(n_6855)
);

INVx1_ASAP7_75t_L g6856 ( 
.A(n_6687),
.Y(n_6856)
);

OAI21xp33_ASAP7_75t_L g6857 ( 
.A1(n_6714),
.A2(n_6484),
.B(n_6585),
.Y(n_6857)
);

OAI221xp5_ASAP7_75t_L g6858 ( 
.A1(n_6754),
.A2(n_6598),
.B1(n_6612),
.B2(n_6605),
.C(n_6647),
.Y(n_6858)
);

OAI31xp33_ASAP7_75t_L g6859 ( 
.A1(n_6837),
.A2(n_6566),
.A3(n_6565),
.B(n_6610),
.Y(n_6859)
);

NAND3xp33_ASAP7_75t_SL g6860 ( 
.A(n_6751),
.B(n_6622),
.C(n_6650),
.Y(n_6860)
);

NAND2xp5_ASAP7_75t_L g6861 ( 
.A(n_6704),
.B(n_6620),
.Y(n_6861)
);

NAND2xp5_ASAP7_75t_L g6862 ( 
.A(n_6698),
.B(n_6639),
.Y(n_6862)
);

OR2x2_ASAP7_75t_L g6863 ( 
.A(n_6697),
.B(n_666),
.Y(n_6863)
);

AND2x2_ASAP7_75t_L g6864 ( 
.A(n_6691),
.B(n_1070),
.Y(n_6864)
);

AOI22xp5_ASAP7_75t_L g6865 ( 
.A1(n_6758),
.A2(n_668),
.B1(n_666),
.B2(n_667),
.Y(n_6865)
);

AND2x2_ASAP7_75t_L g6866 ( 
.A(n_6717),
.B(n_1070),
.Y(n_6866)
);

AOI211xp5_ASAP7_75t_L g6867 ( 
.A1(n_6706),
.A2(n_668),
.B(n_666),
.C(n_667),
.Y(n_6867)
);

INVx2_ASAP7_75t_SL g6868 ( 
.A(n_6702),
.Y(n_6868)
);

AOI22xp33_ASAP7_75t_L g6869 ( 
.A1(n_6753),
.A2(n_671),
.B1(n_669),
.B2(n_670),
.Y(n_6869)
);

NAND2xp5_ASAP7_75t_L g6870 ( 
.A(n_6731),
.B(n_669),
.Y(n_6870)
);

AND2x2_ASAP7_75t_SL g6871 ( 
.A(n_6841),
.B(n_669),
.Y(n_6871)
);

INVx2_ASAP7_75t_L g6872 ( 
.A(n_6788),
.Y(n_6872)
);

INVx1_ASAP7_75t_L g6873 ( 
.A(n_6701),
.Y(n_6873)
);

INVx1_ASAP7_75t_L g6874 ( 
.A(n_6820),
.Y(n_6874)
);

AND2x2_ASAP7_75t_L g6875 ( 
.A(n_6759),
.B(n_671),
.Y(n_6875)
);

INVx1_ASAP7_75t_L g6876 ( 
.A(n_6824),
.Y(n_6876)
);

AND2x2_ASAP7_75t_L g6877 ( 
.A(n_6807),
.B(n_672),
.Y(n_6877)
);

INVx1_ASAP7_75t_L g6878 ( 
.A(n_6713),
.Y(n_6878)
);

NAND2xp5_ASAP7_75t_L g6879 ( 
.A(n_6768),
.B(n_672),
.Y(n_6879)
);

INVx2_ASAP7_75t_L g6880 ( 
.A(n_6709),
.Y(n_6880)
);

AND2x2_ASAP7_75t_L g6881 ( 
.A(n_6812),
.B(n_672),
.Y(n_6881)
);

AND2x2_ASAP7_75t_L g6882 ( 
.A(n_6818),
.B(n_673),
.Y(n_6882)
);

INVx1_ASAP7_75t_L g6883 ( 
.A(n_6829),
.Y(n_6883)
);

AND2x2_ASAP7_75t_L g6884 ( 
.A(n_6835),
.B(n_674),
.Y(n_6884)
);

INVx2_ASAP7_75t_SL g6885 ( 
.A(n_6725),
.Y(n_6885)
);

AOI221x1_ASAP7_75t_L g6886 ( 
.A1(n_6723),
.A2(n_677),
.B1(n_675),
.B2(n_676),
.C(n_678),
.Y(n_6886)
);

HB1xp67_ASAP7_75t_L g6887 ( 
.A(n_6719),
.Y(n_6887)
);

INVx1_ASAP7_75t_L g6888 ( 
.A(n_6744),
.Y(n_6888)
);

AOI22xp5_ASAP7_75t_L g6889 ( 
.A1(n_6735),
.A2(n_1062),
.B1(n_677),
.B2(n_675),
.Y(n_6889)
);

AOI22xp33_ASAP7_75t_SL g6890 ( 
.A1(n_6814),
.A2(n_678),
.B1(n_676),
.B2(n_677),
.Y(n_6890)
);

AND2x2_ASAP7_75t_L g6891 ( 
.A(n_6802),
.B(n_676),
.Y(n_6891)
);

AOI33xp33_ASAP7_75t_L g6892 ( 
.A1(n_6825),
.A2(n_680),
.A3(n_682),
.B1(n_678),
.B2(n_679),
.B3(n_681),
.Y(n_6892)
);

CKINVDCx5p33_ASAP7_75t_R g6893 ( 
.A(n_6696),
.Y(n_6893)
);

INVx1_ASAP7_75t_L g6894 ( 
.A(n_6741),
.Y(n_6894)
);

AND2x2_ASAP7_75t_L g6895 ( 
.A(n_6789),
.B(n_679),
.Y(n_6895)
);

INVx1_ASAP7_75t_L g6896 ( 
.A(n_6741),
.Y(n_6896)
);

HB1xp67_ASAP7_75t_L g6897 ( 
.A(n_6756),
.Y(n_6897)
);

INVx2_ASAP7_75t_L g6898 ( 
.A(n_6749),
.Y(n_6898)
);

AOI211xp5_ASAP7_75t_L g6899 ( 
.A1(n_6732),
.A2(n_681),
.B(n_679),
.C(n_680),
.Y(n_6899)
);

NAND5xp2_ASAP7_75t_SL g6900 ( 
.A(n_6847),
.B(n_683),
.C(n_680),
.D(n_682),
.E(n_684),
.Y(n_6900)
);

AOI211xp5_ASAP7_75t_L g6901 ( 
.A1(n_6712),
.A2(n_685),
.B(n_683),
.C(n_684),
.Y(n_6901)
);

OR2x2_ASAP7_75t_L g6902 ( 
.A(n_6805),
.B(n_684),
.Y(n_6902)
);

INVx1_ASAP7_75t_L g6903 ( 
.A(n_6749),
.Y(n_6903)
);

INVxp67_ASAP7_75t_SL g6904 ( 
.A(n_6711),
.Y(n_6904)
);

CKINVDCx16_ASAP7_75t_R g6905 ( 
.A(n_6823),
.Y(n_6905)
);

INVx2_ASAP7_75t_L g6906 ( 
.A(n_6740),
.Y(n_6906)
);

INVx3_ASAP7_75t_L g6907 ( 
.A(n_6823),
.Y(n_6907)
);

AND2x2_ASAP7_75t_L g6908 ( 
.A(n_6838),
.B(n_685),
.Y(n_6908)
);

INVx1_ASAP7_75t_SL g6909 ( 
.A(n_6729),
.Y(n_6909)
);

NAND2xp5_ASAP7_75t_SL g6910 ( 
.A(n_6737),
.B(n_686),
.Y(n_6910)
);

NAND3xp33_ASAP7_75t_L g6911 ( 
.A(n_6690),
.B(n_686),
.C(n_687),
.Y(n_6911)
);

NAND4xp25_ASAP7_75t_L g6912 ( 
.A(n_6800),
.B(n_688),
.C(n_686),
.D(n_687),
.Y(n_6912)
);

NAND2x1p5_ASAP7_75t_L g6913 ( 
.A(n_6720),
.B(n_687),
.Y(n_6913)
);

NOR2xp33_ASAP7_75t_L g6914 ( 
.A(n_6828),
.B(n_688),
.Y(n_6914)
);

AND2x2_ASAP7_75t_L g6915 ( 
.A(n_6849),
.B(n_689),
.Y(n_6915)
);

AND2x2_ASAP7_75t_L g6916 ( 
.A(n_6718),
.B(n_689),
.Y(n_6916)
);

OAI221xp5_ASAP7_75t_L g6917 ( 
.A1(n_6787),
.A2(n_691),
.B1(n_689),
.B2(n_690),
.C(n_692),
.Y(n_6917)
);

INVx1_ASAP7_75t_L g6918 ( 
.A(n_6776),
.Y(n_6918)
);

INVx1_ASAP7_75t_SL g6919 ( 
.A(n_6776),
.Y(n_6919)
);

AND2x2_ASAP7_75t_L g6920 ( 
.A(n_6764),
.B(n_690),
.Y(n_6920)
);

INVx2_ASAP7_75t_L g6921 ( 
.A(n_6804),
.Y(n_6921)
);

OR2x2_ASAP7_75t_L g6922 ( 
.A(n_6805),
.B(n_690),
.Y(n_6922)
);

AND2x4_ASAP7_75t_L g6923 ( 
.A(n_6804),
.B(n_691),
.Y(n_6923)
);

AND2x2_ASAP7_75t_L g6924 ( 
.A(n_6722),
.B(n_6724),
.Y(n_6924)
);

INVx2_ASAP7_75t_L g6925 ( 
.A(n_6801),
.Y(n_6925)
);

AND2x2_ASAP7_75t_L g6926 ( 
.A(n_6733),
.B(n_692),
.Y(n_6926)
);

INVx1_ASAP7_75t_L g6927 ( 
.A(n_6775),
.Y(n_6927)
);

AND2x2_ASAP7_75t_L g6928 ( 
.A(n_6747),
.B(n_6736),
.Y(n_6928)
);

INVx1_ASAP7_75t_L g6929 ( 
.A(n_6809),
.Y(n_6929)
);

AND2x2_ASAP7_75t_L g6930 ( 
.A(n_6815),
.B(n_692),
.Y(n_6930)
);

INVx1_ASAP7_75t_L g6931 ( 
.A(n_6707),
.Y(n_6931)
);

AND2x2_ASAP7_75t_L g6932 ( 
.A(n_6771),
.B(n_693),
.Y(n_6932)
);

AO31x2_ASAP7_75t_L g6933 ( 
.A1(n_6705),
.A2(n_695),
.A3(n_693),
.B(n_694),
.Y(n_6933)
);

AND2x2_ASAP7_75t_L g6934 ( 
.A(n_6772),
.B(n_693),
.Y(n_6934)
);

INVx1_ASAP7_75t_SL g6935 ( 
.A(n_6738),
.Y(n_6935)
);

HB1xp67_ASAP7_75t_L g6936 ( 
.A(n_6721),
.Y(n_6936)
);

INVx1_ASAP7_75t_L g6937 ( 
.A(n_6821),
.Y(n_6937)
);

INVx1_ASAP7_75t_L g6938 ( 
.A(n_6755),
.Y(n_6938)
);

AND2x2_ASAP7_75t_L g6939 ( 
.A(n_6783),
.B(n_694),
.Y(n_6939)
);

OAI33xp33_ASAP7_75t_L g6940 ( 
.A1(n_6763),
.A2(n_697),
.A3(n_699),
.B1(n_695),
.B2(n_696),
.B3(n_698),
.Y(n_6940)
);

AOI211xp5_ASAP7_75t_L g6941 ( 
.A1(n_6839),
.A2(n_698),
.B(n_696),
.C(n_697),
.Y(n_6941)
);

INVx1_ASAP7_75t_L g6942 ( 
.A(n_6811),
.Y(n_6942)
);

INVx1_ASAP7_75t_L g6943 ( 
.A(n_6694),
.Y(n_6943)
);

AOI221xp5_ASAP7_75t_L g6944 ( 
.A1(n_6765),
.A2(n_6830),
.B1(n_6817),
.B2(n_6819),
.C(n_6848),
.Y(n_6944)
);

AOI22xp33_ASAP7_75t_SL g6945 ( 
.A1(n_6810),
.A2(n_699),
.B1(n_696),
.B2(n_697),
.Y(n_6945)
);

INVx2_ASAP7_75t_L g6946 ( 
.A(n_6752),
.Y(n_6946)
);

INVx2_ASAP7_75t_SL g6947 ( 
.A(n_6703),
.Y(n_6947)
);

INVx2_ASAP7_75t_L g6948 ( 
.A(n_6745),
.Y(n_6948)
);

OAI31xp33_ASAP7_75t_L g6949 ( 
.A1(n_6727),
.A2(n_702),
.A3(n_700),
.B(n_701),
.Y(n_6949)
);

AO21x2_ASAP7_75t_L g6950 ( 
.A1(n_6742),
.A2(n_700),
.B(n_701),
.Y(n_6950)
);

AOI222xp33_ASAP7_75t_L g6951 ( 
.A1(n_6773),
.A2(n_703),
.B1(n_705),
.B2(n_700),
.C1(n_702),
.C2(n_704),
.Y(n_6951)
);

AND2x2_ASAP7_75t_L g6952 ( 
.A(n_6784),
.B(n_703),
.Y(n_6952)
);

OAI321xp33_ASAP7_75t_L g6953 ( 
.A1(n_6844),
.A2(n_706),
.A3(n_708),
.B1(n_704),
.B2(n_705),
.C(n_707),
.Y(n_6953)
);

INVxp67_ASAP7_75t_L g6954 ( 
.A(n_6726),
.Y(n_6954)
);

HB1xp67_ASAP7_75t_L g6955 ( 
.A(n_6795),
.Y(n_6955)
);

OAI31xp33_ASAP7_75t_L g6956 ( 
.A1(n_6840),
.A2(n_6782),
.A3(n_6813),
.B(n_6845),
.Y(n_6956)
);

NOR2xp33_ASAP7_75t_L g6957 ( 
.A(n_6779),
.B(n_704),
.Y(n_6957)
);

AND2x2_ASAP7_75t_L g6958 ( 
.A(n_6792),
.B(n_705),
.Y(n_6958)
);

HB1xp67_ASAP7_75t_L g6959 ( 
.A(n_6734),
.Y(n_6959)
);

AND2x2_ASAP7_75t_L g6960 ( 
.A(n_6850),
.B(n_706),
.Y(n_6960)
);

INVx2_ASAP7_75t_L g6961 ( 
.A(n_6785),
.Y(n_6961)
);

HB1xp67_ASAP7_75t_L g6962 ( 
.A(n_6832),
.Y(n_6962)
);

OAI31xp33_ASAP7_75t_L g6963 ( 
.A1(n_6762),
.A2(n_708),
.A3(n_706),
.B(n_707),
.Y(n_6963)
);

NAND2xp5_ASAP7_75t_L g6964 ( 
.A(n_6728),
.B(n_707),
.Y(n_6964)
);

INVx1_ASAP7_75t_SL g6965 ( 
.A(n_6786),
.Y(n_6965)
);

OAI33xp33_ASAP7_75t_L g6966 ( 
.A1(n_6760),
.A2(n_6846),
.A3(n_6777),
.B1(n_6796),
.B2(n_6833),
.B3(n_6769),
.Y(n_6966)
);

OAI211xp5_ASAP7_75t_L g6967 ( 
.A1(n_6715),
.A2(n_711),
.B(n_709),
.C(n_710),
.Y(n_6967)
);

AND2x2_ASAP7_75t_L g6968 ( 
.A(n_6842),
.B(n_709),
.Y(n_6968)
);

NAND2xp5_ASAP7_75t_L g6969 ( 
.A(n_6774),
.B(n_709),
.Y(n_6969)
);

INVx1_ASAP7_75t_SL g6970 ( 
.A(n_6822),
.Y(n_6970)
);

AND2x2_ASAP7_75t_L g6971 ( 
.A(n_6826),
.B(n_710),
.Y(n_6971)
);

INVx1_ASAP7_75t_L g6972 ( 
.A(n_6757),
.Y(n_6972)
);

HB1xp67_ASAP7_75t_L g6973 ( 
.A(n_6790),
.Y(n_6973)
);

AND2x2_ASAP7_75t_L g6974 ( 
.A(n_6778),
.B(n_711),
.Y(n_6974)
);

INVx2_ASAP7_75t_L g6975 ( 
.A(n_6743),
.Y(n_6975)
);

INVx1_ASAP7_75t_L g6976 ( 
.A(n_6693),
.Y(n_6976)
);

INVx2_ASAP7_75t_L g6977 ( 
.A(n_6798),
.Y(n_6977)
);

HB1xp67_ASAP7_75t_L g6978 ( 
.A(n_6700),
.Y(n_6978)
);

OAI22xp5_ASAP7_75t_L g6979 ( 
.A1(n_6710),
.A2(n_713),
.B1(n_711),
.B2(n_712),
.Y(n_6979)
);

OAI31xp33_ASAP7_75t_L g6980 ( 
.A1(n_6806),
.A2(n_6803),
.A3(n_6797),
.B(n_6695),
.Y(n_6980)
);

NAND2xp5_ASAP7_75t_L g6981 ( 
.A(n_6766),
.B(n_712),
.Y(n_6981)
);

NAND2xp5_ASAP7_75t_L g6982 ( 
.A(n_6699),
.B(n_712),
.Y(n_6982)
);

AND2x2_ASAP7_75t_L g6983 ( 
.A(n_6834),
.B(n_713),
.Y(n_6983)
);

HB1xp67_ASAP7_75t_L g6984 ( 
.A(n_6851),
.Y(n_6984)
);

AND2x2_ASAP7_75t_L g6985 ( 
.A(n_6793),
.B(n_713),
.Y(n_6985)
);

AOI33xp33_ASAP7_75t_L g6986 ( 
.A1(n_6780),
.A2(n_716),
.A3(n_718),
.B1(n_714),
.B2(n_715),
.B3(n_717),
.Y(n_6986)
);

INVx1_ASAP7_75t_L g6987 ( 
.A(n_6750),
.Y(n_6987)
);

INVx1_ASAP7_75t_L g6988 ( 
.A(n_6770),
.Y(n_6988)
);

INVx1_ASAP7_75t_L g6989 ( 
.A(n_6843),
.Y(n_6989)
);

AND2x4_ASAP7_75t_L g6990 ( 
.A(n_6730),
.B(n_714),
.Y(n_6990)
);

INVx5_ASAP7_75t_L g6991 ( 
.A(n_6808),
.Y(n_6991)
);

INVx1_ASAP7_75t_L g6992 ( 
.A(n_6716),
.Y(n_6992)
);

AND2x2_ASAP7_75t_L g6993 ( 
.A(n_6799),
.B(n_714),
.Y(n_6993)
);

INVx1_ASAP7_75t_L g6994 ( 
.A(n_6708),
.Y(n_6994)
);

INVx2_ASAP7_75t_L g6995 ( 
.A(n_6791),
.Y(n_6995)
);

INVx2_ASAP7_75t_L g6996 ( 
.A(n_6761),
.Y(n_6996)
);

AND2x4_ASAP7_75t_L g6997 ( 
.A(n_6746),
.B(n_715),
.Y(n_6997)
);

AND2x2_ASAP7_75t_L g6998 ( 
.A(n_6781),
.B(n_716),
.Y(n_6998)
);

AOI211xp5_ASAP7_75t_L g6999 ( 
.A1(n_6794),
.A2(n_719),
.B(n_717),
.C(n_718),
.Y(n_6999)
);

OAI22xp5_ASAP7_75t_L g7000 ( 
.A1(n_6748),
.A2(n_719),
.B1(n_717),
.B2(n_718),
.Y(n_7000)
);

AND2x2_ASAP7_75t_L g7001 ( 
.A(n_6827),
.B(n_719),
.Y(n_7001)
);

INVx2_ASAP7_75t_L g7002 ( 
.A(n_6767),
.Y(n_7002)
);

OR2x2_ASAP7_75t_L g7003 ( 
.A(n_6836),
.B(n_720),
.Y(n_7003)
);

INVx2_ASAP7_75t_L g7004 ( 
.A(n_6688),
.Y(n_7004)
);

INVx4_ASAP7_75t_L g7005 ( 
.A(n_6739),
.Y(n_7005)
);

OAI211xp5_ASAP7_75t_L g7006 ( 
.A1(n_6831),
.A2(n_1061),
.B(n_722),
.C(n_720),
.Y(n_7006)
);

AND2x2_ASAP7_75t_L g7007 ( 
.A(n_6816),
.B(n_720),
.Y(n_7007)
);

BUFx3_ASAP7_75t_L g7008 ( 
.A(n_6702),
.Y(n_7008)
);

AOI21x1_ASAP7_75t_L g7009 ( 
.A1(n_6820),
.A2(n_721),
.B(n_722),
.Y(n_7009)
);

OAI31xp33_ASAP7_75t_L g7010 ( 
.A1(n_6754),
.A2(n_724),
.A3(n_721),
.B(n_723),
.Y(n_7010)
);

OR2x2_ASAP7_75t_L g7011 ( 
.A(n_6697),
.B(n_721),
.Y(n_7011)
);

INVx1_ASAP7_75t_L g7012 ( 
.A(n_6685),
.Y(n_7012)
);

AND2x2_ASAP7_75t_L g7013 ( 
.A(n_6685),
.B(n_723),
.Y(n_7013)
);

AND2x4_ASAP7_75t_L g7014 ( 
.A(n_6689),
.B(n_724),
.Y(n_7014)
);

INVx2_ASAP7_75t_L g7015 ( 
.A(n_6689),
.Y(n_7015)
);

INVx2_ASAP7_75t_SL g7016 ( 
.A(n_6702),
.Y(n_7016)
);

INVx1_ASAP7_75t_L g7017 ( 
.A(n_6685),
.Y(n_7017)
);

AND2x2_ASAP7_75t_L g7018 ( 
.A(n_6685),
.B(n_724),
.Y(n_7018)
);

AND2x2_ASAP7_75t_L g7019 ( 
.A(n_6685),
.B(n_725),
.Y(n_7019)
);

INVx1_ASAP7_75t_L g7020 ( 
.A(n_6685),
.Y(n_7020)
);

OAI221xp5_ASAP7_75t_L g7021 ( 
.A1(n_6754),
.A2(n_728),
.B1(n_726),
.B2(n_727),
.C(n_729),
.Y(n_7021)
);

INVx1_ASAP7_75t_L g7022 ( 
.A(n_6685),
.Y(n_7022)
);

AND2x2_ASAP7_75t_L g7023 ( 
.A(n_6685),
.B(n_726),
.Y(n_7023)
);

INVx2_ASAP7_75t_L g7024 ( 
.A(n_7008),
.Y(n_7024)
);

INVx1_ASAP7_75t_L g7025 ( 
.A(n_6874),
.Y(n_7025)
);

INVx1_ASAP7_75t_L g7026 ( 
.A(n_6876),
.Y(n_7026)
);

INVx1_ASAP7_75t_L g7027 ( 
.A(n_7009),
.Y(n_7027)
);

INVx1_ASAP7_75t_L g7028 ( 
.A(n_6883),
.Y(n_7028)
);

INVx1_ASAP7_75t_L g7029 ( 
.A(n_6897),
.Y(n_7029)
);

AND2x2_ASAP7_75t_L g7030 ( 
.A(n_6905),
.B(n_726),
.Y(n_7030)
);

NAND2xp33_ASAP7_75t_R g7031 ( 
.A(n_6907),
.B(n_727),
.Y(n_7031)
);

OR2x2_ASAP7_75t_L g7032 ( 
.A(n_7015),
.B(n_728),
.Y(n_7032)
);

NAND2xp5_ASAP7_75t_L g7033 ( 
.A(n_6868),
.B(n_728),
.Y(n_7033)
);

CKINVDCx5p33_ASAP7_75t_R g7034 ( 
.A(n_6893),
.Y(n_7034)
);

INVx2_ASAP7_75t_L g7035 ( 
.A(n_7016),
.Y(n_7035)
);

INVx1_ASAP7_75t_L g7036 ( 
.A(n_7014),
.Y(n_7036)
);

INVx1_ASAP7_75t_L g7037 ( 
.A(n_7014),
.Y(n_7037)
);

INVx1_ASAP7_75t_L g7038 ( 
.A(n_6854),
.Y(n_7038)
);

AND2x2_ASAP7_75t_L g7039 ( 
.A(n_6872),
.B(n_729),
.Y(n_7039)
);

INVx1_ASAP7_75t_L g7040 ( 
.A(n_6864),
.Y(n_7040)
);

INVx2_ASAP7_75t_L g7041 ( 
.A(n_6885),
.Y(n_7041)
);

HB1xp67_ASAP7_75t_L g7042 ( 
.A(n_6880),
.Y(n_7042)
);

O2A1O1Ixp5_ASAP7_75t_L g7043 ( 
.A1(n_6904),
.A2(n_731),
.B(n_729),
.C(n_730),
.Y(n_7043)
);

INVx2_ASAP7_75t_L g7044 ( 
.A(n_6906),
.Y(n_7044)
);

OR2x2_ASAP7_75t_L g7045 ( 
.A(n_6969),
.B(n_730),
.Y(n_7045)
);

INVx1_ASAP7_75t_L g7046 ( 
.A(n_6877),
.Y(n_7046)
);

INVx1_ASAP7_75t_L g7047 ( 
.A(n_6875),
.Y(n_7047)
);

INVx1_ASAP7_75t_L g7048 ( 
.A(n_6902),
.Y(n_7048)
);

AND2x2_ASAP7_75t_L g7049 ( 
.A(n_6909),
.B(n_7013),
.Y(n_7049)
);

OR2x2_ASAP7_75t_L g7050 ( 
.A(n_6919),
.B(n_730),
.Y(n_7050)
);

AOI32xp33_ASAP7_75t_L g7051 ( 
.A1(n_6977),
.A2(n_733),
.A3(n_731),
.B1(n_732),
.B2(n_734),
.Y(n_7051)
);

INVx1_ASAP7_75t_L g7052 ( 
.A(n_6922),
.Y(n_7052)
);

INVx1_ASAP7_75t_L g7053 ( 
.A(n_6933),
.Y(n_7053)
);

OR2x2_ASAP7_75t_L g7054 ( 
.A(n_6853),
.B(n_731),
.Y(n_7054)
);

NAND2xp5_ASAP7_75t_L g7055 ( 
.A(n_6991),
.B(n_732),
.Y(n_7055)
);

AND2x2_ASAP7_75t_L g7056 ( 
.A(n_7018),
.B(n_733),
.Y(n_7056)
);

HB1xp67_ASAP7_75t_L g7057 ( 
.A(n_6933),
.Y(n_7057)
);

INVx2_ASAP7_75t_L g7058 ( 
.A(n_6925),
.Y(n_7058)
);

AND2x2_ASAP7_75t_L g7059 ( 
.A(n_7019),
.B(n_733),
.Y(n_7059)
);

INVx1_ASAP7_75t_L g7060 ( 
.A(n_6933),
.Y(n_7060)
);

AND2x4_ASAP7_75t_L g7061 ( 
.A(n_6921),
.B(n_734),
.Y(n_7061)
);

AND2x4_ASAP7_75t_L g7062 ( 
.A(n_6898),
.B(n_734),
.Y(n_7062)
);

INVx1_ASAP7_75t_L g7063 ( 
.A(n_6887),
.Y(n_7063)
);

AOI22xp5_ASAP7_75t_L g7064 ( 
.A1(n_6995),
.A2(n_737),
.B1(n_735),
.B2(n_736),
.Y(n_7064)
);

INVx1_ASAP7_75t_L g7065 ( 
.A(n_6895),
.Y(n_7065)
);

AND2x2_ASAP7_75t_L g7066 ( 
.A(n_7023),
.B(n_736),
.Y(n_7066)
);

NAND2xp5_ASAP7_75t_L g7067 ( 
.A(n_6991),
.B(n_737),
.Y(n_7067)
);

INVx1_ASAP7_75t_L g7068 ( 
.A(n_6923),
.Y(n_7068)
);

NAND4xp25_ASAP7_75t_L g7069 ( 
.A(n_6956),
.B(n_740),
.C(n_738),
.D(n_739),
.Y(n_7069)
);

AND2x2_ASAP7_75t_L g7070 ( 
.A(n_6924),
.B(n_738),
.Y(n_7070)
);

INVx1_ASAP7_75t_L g7071 ( 
.A(n_6923),
.Y(n_7071)
);

AND2x4_ASAP7_75t_L g7072 ( 
.A(n_6918),
.B(n_738),
.Y(n_7072)
);

INVx1_ASAP7_75t_L g7073 ( 
.A(n_6916),
.Y(n_7073)
);

INVx2_ASAP7_75t_L g7074 ( 
.A(n_6894),
.Y(n_7074)
);

AND2x2_ASAP7_75t_L g7075 ( 
.A(n_6866),
.B(n_739),
.Y(n_7075)
);

AND2x2_ASAP7_75t_L g7076 ( 
.A(n_6920),
.B(n_6881),
.Y(n_7076)
);

INVx1_ASAP7_75t_SL g7077 ( 
.A(n_6896),
.Y(n_7077)
);

AND2x2_ASAP7_75t_L g7078 ( 
.A(n_6882),
.B(n_740),
.Y(n_7078)
);

INVx2_ASAP7_75t_L g7079 ( 
.A(n_6903),
.Y(n_7079)
);

AND2x2_ASAP7_75t_L g7080 ( 
.A(n_6884),
.B(n_741),
.Y(n_7080)
);

OAI211xp5_ASAP7_75t_L g7081 ( 
.A1(n_6941),
.A2(n_743),
.B(n_741),
.C(n_742),
.Y(n_7081)
);

NAND2xp5_ASAP7_75t_L g7082 ( 
.A(n_6991),
.B(n_742),
.Y(n_7082)
);

NAND2xp5_ASAP7_75t_L g7083 ( 
.A(n_6971),
.B(n_743),
.Y(n_7083)
);

INVx1_ASAP7_75t_L g7084 ( 
.A(n_6863),
.Y(n_7084)
);

INVx2_ASAP7_75t_SL g7085 ( 
.A(n_6927),
.Y(n_7085)
);

AO21x1_ASAP7_75t_L g7086 ( 
.A1(n_6957),
.A2(n_743),
.B(n_744),
.Y(n_7086)
);

NAND2xp5_ASAP7_75t_L g7087 ( 
.A(n_6890),
.B(n_744),
.Y(n_7087)
);

AND2x2_ASAP7_75t_L g7088 ( 
.A(n_6891),
.B(n_744),
.Y(n_7088)
);

INVx1_ASAP7_75t_L g7089 ( 
.A(n_7011),
.Y(n_7089)
);

AND2x2_ASAP7_75t_L g7090 ( 
.A(n_6908),
.B(n_745),
.Y(n_7090)
);

OR2x2_ASAP7_75t_L g7091 ( 
.A(n_7003),
.B(n_745),
.Y(n_7091)
);

INVx1_ASAP7_75t_L g7092 ( 
.A(n_6936),
.Y(n_7092)
);

AND2x2_ASAP7_75t_L g7093 ( 
.A(n_6915),
.B(n_745),
.Y(n_7093)
);

OR2x2_ASAP7_75t_L g7094 ( 
.A(n_6879),
.B(n_746),
.Y(n_7094)
);

INVx2_ASAP7_75t_L g7095 ( 
.A(n_6929),
.Y(n_7095)
);

OR2x2_ASAP7_75t_L g7096 ( 
.A(n_6861),
.B(n_746),
.Y(n_7096)
);

AND2x4_ASAP7_75t_L g7097 ( 
.A(n_6975),
.B(n_746),
.Y(n_7097)
);

AND2x4_ASAP7_75t_L g7098 ( 
.A(n_6987),
.B(n_747),
.Y(n_7098)
);

OR2x2_ASAP7_75t_L g7099 ( 
.A(n_6964),
.B(n_747),
.Y(n_7099)
);

INVx2_ASAP7_75t_L g7100 ( 
.A(n_6888),
.Y(n_7100)
);

A2O1A1Ixp33_ASAP7_75t_L g7101 ( 
.A1(n_6963),
.A2(n_749),
.B(n_747),
.C(n_748),
.Y(n_7101)
);

INVx2_ASAP7_75t_L g7102 ( 
.A(n_6913),
.Y(n_7102)
);

HB1xp67_ASAP7_75t_L g7103 ( 
.A(n_6926),
.Y(n_7103)
);

AND2x2_ASAP7_75t_L g7104 ( 
.A(n_6934),
.B(n_748),
.Y(n_7104)
);

OR2x2_ASAP7_75t_L g7105 ( 
.A(n_6912),
.B(n_748),
.Y(n_7105)
);

INVx2_ASAP7_75t_L g7106 ( 
.A(n_6988),
.Y(n_7106)
);

INVx1_ASAP7_75t_L g7107 ( 
.A(n_6983),
.Y(n_7107)
);

INVx1_ASAP7_75t_L g7108 ( 
.A(n_6974),
.Y(n_7108)
);

OR2x2_ASAP7_75t_L g7109 ( 
.A(n_6982),
.B(n_750),
.Y(n_7109)
);

INVxp67_ASAP7_75t_SL g7110 ( 
.A(n_6962),
.Y(n_7110)
);

INVx3_ASAP7_75t_L g7111 ( 
.A(n_6990),
.Y(n_7111)
);

INVx1_ASAP7_75t_L g7112 ( 
.A(n_6892),
.Y(n_7112)
);

OR2x2_ASAP7_75t_L g7113 ( 
.A(n_6910),
.B(n_750),
.Y(n_7113)
);

OR2x2_ASAP7_75t_L g7114 ( 
.A(n_6948),
.B(n_750),
.Y(n_7114)
);

INVx2_ASAP7_75t_SL g7115 ( 
.A(n_6961),
.Y(n_7115)
);

NOR2xp33_ASAP7_75t_L g7116 ( 
.A(n_6966),
.B(n_751),
.Y(n_7116)
);

NAND2xp5_ASAP7_75t_L g7117 ( 
.A(n_6945),
.B(n_751),
.Y(n_7117)
);

OR2x2_ASAP7_75t_L g7118 ( 
.A(n_6870),
.B(n_751),
.Y(n_7118)
);

NAND2xp5_ASAP7_75t_L g7119 ( 
.A(n_6867),
.B(n_752),
.Y(n_7119)
);

OR2x2_ASAP7_75t_L g7120 ( 
.A(n_7022),
.B(n_752),
.Y(n_7120)
);

NAND2x1p5_ASAP7_75t_L g7121 ( 
.A(n_6930),
.B(n_7005),
.Y(n_7121)
);

AND2x2_ASAP7_75t_L g7122 ( 
.A(n_6852),
.B(n_6932),
.Y(n_7122)
);

INVx2_ASAP7_75t_L g7123 ( 
.A(n_6947),
.Y(n_7123)
);

INVx1_ASAP7_75t_L g7124 ( 
.A(n_6856),
.Y(n_7124)
);

INVx2_ASAP7_75t_L g7125 ( 
.A(n_6935),
.Y(n_7125)
);

INVx1_ASAP7_75t_L g7126 ( 
.A(n_6914),
.Y(n_7126)
);

AND2x2_ASAP7_75t_L g7127 ( 
.A(n_6928),
.B(n_6939),
.Y(n_7127)
);

AOI22xp5_ASAP7_75t_L g7128 ( 
.A1(n_6996),
.A2(n_754),
.B1(n_752),
.B2(n_753),
.Y(n_7128)
);

INVxp67_ASAP7_75t_L g7129 ( 
.A(n_6959),
.Y(n_7129)
);

INVxp33_ASAP7_75t_L g7130 ( 
.A(n_6955),
.Y(n_7130)
);

INVx2_ASAP7_75t_L g7131 ( 
.A(n_6950),
.Y(n_7131)
);

NAND2xp5_ASAP7_75t_L g7132 ( 
.A(n_7010),
.B(n_753),
.Y(n_7132)
);

INVx1_ASAP7_75t_L g7133 ( 
.A(n_6855),
.Y(n_7133)
);

NAND2x1_ASAP7_75t_L g7134 ( 
.A(n_6946),
.B(n_753),
.Y(n_7134)
);

INVx1_ASAP7_75t_L g7135 ( 
.A(n_6998),
.Y(n_7135)
);

AND2x4_ASAP7_75t_L g7136 ( 
.A(n_6990),
.B(n_754),
.Y(n_7136)
);

INVx2_ASAP7_75t_L g7137 ( 
.A(n_6997),
.Y(n_7137)
);

NAND2xp5_ASAP7_75t_L g7138 ( 
.A(n_6871),
.B(n_754),
.Y(n_7138)
);

AND2x2_ASAP7_75t_L g7139 ( 
.A(n_6952),
.B(n_755),
.Y(n_7139)
);

AOI21xp33_ASAP7_75t_SL g7140 ( 
.A1(n_6949),
.A2(n_1058),
.B(n_755),
.Y(n_7140)
);

INVx1_ASAP7_75t_SL g7141 ( 
.A(n_6965),
.Y(n_7141)
);

INVx1_ASAP7_75t_L g7142 ( 
.A(n_7001),
.Y(n_7142)
);

OR2x2_ASAP7_75t_L g7143 ( 
.A(n_7012),
.B(n_755),
.Y(n_7143)
);

INVx1_ASAP7_75t_L g7144 ( 
.A(n_6985),
.Y(n_7144)
);

NAND2xp5_ASAP7_75t_L g7145 ( 
.A(n_6901),
.B(n_756),
.Y(n_7145)
);

INVx1_ASAP7_75t_L g7146 ( 
.A(n_6993),
.Y(n_7146)
);

NAND2xp5_ASAP7_75t_L g7147 ( 
.A(n_6951),
.B(n_756),
.Y(n_7147)
);

INVx1_ASAP7_75t_L g7148 ( 
.A(n_6986),
.Y(n_7148)
);

INVx2_ASAP7_75t_L g7149 ( 
.A(n_6997),
.Y(n_7149)
);

NOR2xp33_ASAP7_75t_R g7150 ( 
.A(n_6900),
.B(n_756),
.Y(n_7150)
);

NOR2xp33_ASAP7_75t_L g7151 ( 
.A(n_6940),
.B(n_757),
.Y(n_7151)
);

NAND2xp5_ASAP7_75t_L g7152 ( 
.A(n_6899),
.B(n_757),
.Y(n_7152)
);

INVx1_ASAP7_75t_SL g7153 ( 
.A(n_6970),
.Y(n_7153)
);

NOR2xp33_ASAP7_75t_L g7154 ( 
.A(n_6860),
.B(n_757),
.Y(n_7154)
);

OR2x2_ASAP7_75t_L g7155 ( 
.A(n_7017),
.B(n_758),
.Y(n_7155)
);

INVx1_ASAP7_75t_L g7156 ( 
.A(n_6976),
.Y(n_7156)
);

INVx1_ASAP7_75t_L g7157 ( 
.A(n_6943),
.Y(n_7157)
);

AOI22xp5_ASAP7_75t_L g7158 ( 
.A1(n_7034),
.A2(n_7002),
.B1(n_6857),
.B2(n_6911),
.Y(n_7158)
);

NAND2xp5_ASAP7_75t_L g7159 ( 
.A(n_7097),
.B(n_6869),
.Y(n_7159)
);

AND2x2_ASAP7_75t_L g7160 ( 
.A(n_7030),
.B(n_7049),
.Y(n_7160)
);

HB1xp67_ASAP7_75t_L g7161 ( 
.A(n_7097),
.Y(n_7161)
);

INVx1_ASAP7_75t_L g7162 ( 
.A(n_7055),
.Y(n_7162)
);

OAI22xp5_ASAP7_75t_L g7163 ( 
.A1(n_7128),
.A2(n_6994),
.B1(n_6992),
.B2(n_6954),
.Y(n_7163)
);

AND2x2_ASAP7_75t_L g7164 ( 
.A(n_7024),
.B(n_6958),
.Y(n_7164)
);

INVx1_ASAP7_75t_L g7165 ( 
.A(n_7067),
.Y(n_7165)
);

AND2x2_ASAP7_75t_L g7166 ( 
.A(n_7035),
.B(n_6960),
.Y(n_7166)
);

AND2x2_ASAP7_75t_L g7167 ( 
.A(n_7070),
.B(n_6968),
.Y(n_7167)
);

INVx1_ASAP7_75t_L g7168 ( 
.A(n_7082),
.Y(n_7168)
);

NOR2xp33_ASAP7_75t_L g7169 ( 
.A(n_7069),
.B(n_6858),
.Y(n_7169)
);

INVx1_ASAP7_75t_L g7170 ( 
.A(n_7039),
.Y(n_7170)
);

AND2x2_ASAP7_75t_L g7171 ( 
.A(n_7127),
.B(n_7020),
.Y(n_7171)
);

NOR2xp33_ASAP7_75t_L g7172 ( 
.A(n_7038),
.B(n_6873),
.Y(n_7172)
);

AOI21xp5_ASAP7_75t_L g7173 ( 
.A1(n_7132),
.A2(n_6981),
.B(n_6953),
.Y(n_7173)
);

INVx1_ASAP7_75t_L g7174 ( 
.A(n_7042),
.Y(n_7174)
);

INVx2_ASAP7_75t_SL g7175 ( 
.A(n_7044),
.Y(n_7175)
);

INVx1_ASAP7_75t_L g7176 ( 
.A(n_7136),
.Y(n_7176)
);

NAND2xp5_ASAP7_75t_L g7177 ( 
.A(n_7027),
.B(n_7007),
.Y(n_7177)
);

INVx1_ASAP7_75t_L g7178 ( 
.A(n_7136),
.Y(n_7178)
);

OAI211xp5_ASAP7_75t_L g7179 ( 
.A1(n_7140),
.A2(n_6944),
.B(n_6980),
.C(n_6889),
.Y(n_7179)
);

OAI221xp5_ASAP7_75t_L g7180 ( 
.A1(n_7101),
.A2(n_6859),
.B1(n_6999),
.B2(n_7021),
.C(n_6865),
.Y(n_7180)
);

INVx1_ASAP7_75t_L g7181 ( 
.A(n_7050),
.Y(n_7181)
);

NAND2xp5_ASAP7_75t_L g7182 ( 
.A(n_7151),
.B(n_6886),
.Y(n_7182)
);

INVx2_ASAP7_75t_L g7183 ( 
.A(n_7041),
.Y(n_7183)
);

INVxp67_ASAP7_75t_L g7184 ( 
.A(n_7031),
.Y(n_7184)
);

NOR2xp33_ASAP7_75t_L g7185 ( 
.A(n_7130),
.B(n_6862),
.Y(n_7185)
);

OR2x2_ASAP7_75t_L g7186 ( 
.A(n_7058),
.B(n_6931),
.Y(n_7186)
);

OAI22xp33_ASAP7_75t_SL g7187 ( 
.A1(n_7134),
.A2(n_6938),
.B1(n_6989),
.B2(n_6972),
.Y(n_7187)
);

INVx2_ASAP7_75t_L g7188 ( 
.A(n_7029),
.Y(n_7188)
);

INVx1_ASAP7_75t_L g7189 ( 
.A(n_7061),
.Y(n_7189)
);

NAND2xp5_ASAP7_75t_L g7190 ( 
.A(n_7062),
.B(n_7000),
.Y(n_7190)
);

AND2x2_ASAP7_75t_SL g7191 ( 
.A(n_7154),
.B(n_7004),
.Y(n_7191)
);

XNOR2x1_ASAP7_75t_L g7192 ( 
.A(n_7105),
.B(n_6979),
.Y(n_7192)
);

NAND2xp5_ASAP7_75t_L g7193 ( 
.A(n_7110),
.B(n_6967),
.Y(n_7193)
);

NOR2xp33_ASAP7_75t_L g7194 ( 
.A(n_7036),
.B(n_6973),
.Y(n_7194)
);

NAND4xp25_ASAP7_75t_L g7195 ( 
.A(n_7116),
.B(n_6878),
.C(n_6942),
.D(n_6937),
.Y(n_7195)
);

OAI32xp33_ASAP7_75t_L g7196 ( 
.A1(n_7112),
.A2(n_6984),
.A3(n_6978),
.B1(n_6917),
.B2(n_7006),
.Y(n_7196)
);

INVx1_ASAP7_75t_SL g7197 ( 
.A(n_7077),
.Y(n_7197)
);

INVx1_ASAP7_75t_L g7198 ( 
.A(n_7033),
.Y(n_7198)
);

OR2x2_ASAP7_75t_L g7199 ( 
.A(n_7037),
.B(n_758),
.Y(n_7199)
);

NAND2xp5_ASAP7_75t_L g7200 ( 
.A(n_7104),
.B(n_758),
.Y(n_7200)
);

AOI22xp5_ASAP7_75t_L g7201 ( 
.A1(n_7148),
.A2(n_761),
.B1(n_759),
.B2(n_760),
.Y(n_7201)
);

OAI21xp33_ASAP7_75t_L g7202 ( 
.A1(n_7115),
.A2(n_759),
.B(n_760),
.Y(n_7202)
);

AOI22xp5_ASAP7_75t_L g7203 ( 
.A1(n_7129),
.A2(n_7141),
.B1(n_7153),
.B2(n_7125),
.Y(n_7203)
);

INVx1_ASAP7_75t_L g7204 ( 
.A(n_7032),
.Y(n_7204)
);

HB1xp67_ASAP7_75t_L g7205 ( 
.A(n_7072),
.Y(n_7205)
);

INVx2_ASAP7_75t_SL g7206 ( 
.A(n_7123),
.Y(n_7206)
);

INVx1_ASAP7_75t_L g7207 ( 
.A(n_7043),
.Y(n_7207)
);

INVx1_ASAP7_75t_L g7208 ( 
.A(n_7054),
.Y(n_7208)
);

OAI22xp5_ASAP7_75t_L g7209 ( 
.A1(n_7147),
.A2(n_761),
.B1(n_759),
.B2(n_760),
.Y(n_7209)
);

INVx2_ASAP7_75t_L g7210 ( 
.A(n_7098),
.Y(n_7210)
);

NAND2xp5_ASAP7_75t_L g7211 ( 
.A(n_7078),
.B(n_762),
.Y(n_7211)
);

AND2x4_ASAP7_75t_L g7212 ( 
.A(n_7028),
.B(n_762),
.Y(n_7212)
);

OAI22xp33_ASAP7_75t_R g7213 ( 
.A1(n_7118),
.A2(n_764),
.B1(n_762),
.B2(n_763),
.Y(n_7213)
);

OAI32xp33_ASAP7_75t_L g7214 ( 
.A1(n_7096),
.A2(n_765),
.A3(n_763),
.B1(n_764),
.B2(n_766),
.Y(n_7214)
);

INVx1_ASAP7_75t_L g7215 ( 
.A(n_7114),
.Y(n_7215)
);

AOI22xp5_ASAP7_75t_L g7216 ( 
.A1(n_7135),
.A2(n_765),
.B1(n_763),
.B2(n_764),
.Y(n_7216)
);

OR2x2_ASAP7_75t_L g7217 ( 
.A(n_7083),
.B(n_765),
.Y(n_7217)
);

BUFx2_ASAP7_75t_L g7218 ( 
.A(n_7150),
.Y(n_7218)
);

AOI211xp5_ASAP7_75t_L g7219 ( 
.A1(n_7081),
.A2(n_768),
.B(n_766),
.C(n_767),
.Y(n_7219)
);

NAND2xp5_ASAP7_75t_L g7220 ( 
.A(n_7080),
.B(n_766),
.Y(n_7220)
);

AND2x2_ASAP7_75t_L g7221 ( 
.A(n_7122),
.B(n_7088),
.Y(n_7221)
);

INVx1_ASAP7_75t_L g7222 ( 
.A(n_7064),
.Y(n_7222)
);

NOR2xp33_ASAP7_75t_L g7223 ( 
.A(n_7111),
.B(n_768),
.Y(n_7223)
);

INVx1_ASAP7_75t_L g7224 ( 
.A(n_7120),
.Y(n_7224)
);

AOI22xp33_ASAP7_75t_L g7225 ( 
.A1(n_7063),
.A2(n_770),
.B1(n_768),
.B2(n_769),
.Y(n_7225)
);

NOR2xp33_ASAP7_75t_L g7226 ( 
.A(n_7142),
.B(n_769),
.Y(n_7226)
);

INVx1_ASAP7_75t_L g7227 ( 
.A(n_7143),
.Y(n_7227)
);

OAI22xp5_ASAP7_75t_L g7228 ( 
.A1(n_7092),
.A2(n_771),
.B1(n_769),
.B2(n_770),
.Y(n_7228)
);

INVx2_ASAP7_75t_L g7229 ( 
.A(n_7098),
.Y(n_7229)
);

OAI322xp33_ASAP7_75t_L g7230 ( 
.A1(n_7156),
.A2(n_775),
.A3(n_774),
.B1(n_772),
.B2(n_770),
.C1(n_771),
.C2(n_773),
.Y(n_7230)
);

OAI31xp33_ASAP7_75t_L g7231 ( 
.A1(n_7121),
.A2(n_775),
.A3(n_773),
.B(n_774),
.Y(n_7231)
);

INVx1_ASAP7_75t_L g7232 ( 
.A(n_7155),
.Y(n_7232)
);

XOR2x2_ASAP7_75t_L g7233 ( 
.A(n_7145),
.B(n_773),
.Y(n_7233)
);

OAI21xp5_ASAP7_75t_L g7234 ( 
.A1(n_7119),
.A2(n_775),
.B(n_776),
.Y(n_7234)
);

NAND2xp5_ASAP7_75t_L g7235 ( 
.A(n_7090),
.B(n_776),
.Y(n_7235)
);

NAND2x1p5_ASAP7_75t_L g7236 ( 
.A(n_7074),
.B(n_776),
.Y(n_7236)
);

INVx1_ASAP7_75t_L g7237 ( 
.A(n_7075),
.Y(n_7237)
);

AOI321xp33_ASAP7_75t_L g7238 ( 
.A1(n_7157),
.A2(n_7079),
.A3(n_7100),
.B1(n_7106),
.B2(n_7133),
.C(n_7124),
.Y(n_7238)
);

AOI321xp33_ASAP7_75t_L g7239 ( 
.A1(n_7137),
.A2(n_779),
.A3(n_781),
.B1(n_777),
.B2(n_778),
.C(n_780),
.Y(n_7239)
);

INVx1_ASAP7_75t_L g7240 ( 
.A(n_7045),
.Y(n_7240)
);

AND2x2_ASAP7_75t_L g7241 ( 
.A(n_7093),
.B(n_778),
.Y(n_7241)
);

INVx1_ASAP7_75t_L g7242 ( 
.A(n_7139),
.Y(n_7242)
);

OAI22xp5_ASAP7_75t_L g7243 ( 
.A1(n_7138),
.A2(n_781),
.B1(n_779),
.B2(n_780),
.Y(n_7243)
);

NAND2xp5_ASAP7_75t_L g7244 ( 
.A(n_7056),
.B(n_781),
.Y(n_7244)
);

OAI22xp5_ASAP7_75t_L g7245 ( 
.A1(n_7117),
.A2(n_7149),
.B1(n_7113),
.B2(n_7091),
.Y(n_7245)
);

INVx1_ASAP7_75t_L g7246 ( 
.A(n_7059),
.Y(n_7246)
);

INVx1_ASAP7_75t_L g7247 ( 
.A(n_7066),
.Y(n_7247)
);

NAND2xp5_ASAP7_75t_L g7248 ( 
.A(n_7051),
.B(n_782),
.Y(n_7248)
);

INVx2_ASAP7_75t_L g7249 ( 
.A(n_7102),
.Y(n_7249)
);

OAI32xp33_ASAP7_75t_L g7250 ( 
.A1(n_7073),
.A2(n_7071),
.A3(n_7068),
.B1(n_7146),
.B2(n_7144),
.Y(n_7250)
);

INVx1_ASAP7_75t_L g7251 ( 
.A(n_7087),
.Y(n_7251)
);

INVx1_ASAP7_75t_L g7252 ( 
.A(n_7094),
.Y(n_7252)
);

INVxp67_ASAP7_75t_L g7253 ( 
.A(n_7103),
.Y(n_7253)
);

O2A1O1Ixp33_ASAP7_75t_L g7254 ( 
.A1(n_7152),
.A2(n_784),
.B(n_782),
.C(n_783),
.Y(n_7254)
);

INVx1_ASAP7_75t_L g7255 ( 
.A(n_7076),
.Y(n_7255)
);

AOI22xp33_ASAP7_75t_SL g7256 ( 
.A1(n_7085),
.A2(n_784),
.B1(n_782),
.B2(n_783),
.Y(n_7256)
);

AOI22xp33_ASAP7_75t_SL g7257 ( 
.A1(n_7108),
.A2(n_785),
.B1(n_783),
.B2(n_784),
.Y(n_7257)
);

AOI21xp5_ASAP7_75t_L g7258 ( 
.A1(n_7086),
.A2(n_786),
.B(n_787),
.Y(n_7258)
);

NAND2xp5_ASAP7_75t_L g7259 ( 
.A(n_7107),
.B(n_786),
.Y(n_7259)
);

XOR2x2_ASAP7_75t_L g7260 ( 
.A(n_7099),
.B(n_786),
.Y(n_7260)
);

INVx1_ASAP7_75t_L g7261 ( 
.A(n_7109),
.Y(n_7261)
);

AND2x4_ASAP7_75t_L g7262 ( 
.A(n_7095),
.B(n_787),
.Y(n_7262)
);

INVx1_ASAP7_75t_L g7263 ( 
.A(n_7047),
.Y(n_7263)
);

INVx2_ASAP7_75t_L g7264 ( 
.A(n_7048),
.Y(n_7264)
);

INVx1_ASAP7_75t_L g7265 ( 
.A(n_7040),
.Y(n_7265)
);

AO21x1_ASAP7_75t_L g7266 ( 
.A1(n_7053),
.A2(n_787),
.B(n_788),
.Y(n_7266)
);

INVx2_ASAP7_75t_L g7267 ( 
.A(n_7052),
.Y(n_7267)
);

OR2x2_ASAP7_75t_L g7268 ( 
.A(n_7046),
.B(n_788),
.Y(n_7268)
);

INVx1_ASAP7_75t_L g7269 ( 
.A(n_7065),
.Y(n_7269)
);

INVx1_ASAP7_75t_L g7270 ( 
.A(n_7057),
.Y(n_7270)
);

AO21x1_ASAP7_75t_L g7271 ( 
.A1(n_7060),
.A2(n_788),
.B(n_789),
.Y(n_7271)
);

NAND2xp5_ASAP7_75t_L g7272 ( 
.A(n_7084),
.B(n_789),
.Y(n_7272)
);

INVxp67_ASAP7_75t_L g7273 ( 
.A(n_7089),
.Y(n_7273)
);

OR2x2_ASAP7_75t_L g7274 ( 
.A(n_7025),
.B(n_7026),
.Y(n_7274)
);

INVx2_ASAP7_75t_L g7275 ( 
.A(n_7131),
.Y(n_7275)
);

INVx1_ASAP7_75t_L g7276 ( 
.A(n_7126),
.Y(n_7276)
);

AOI222xp33_ASAP7_75t_L g7277 ( 
.A1(n_7038),
.A2(n_792),
.B1(n_794),
.B2(n_790),
.C1(n_791),
.C2(n_793),
.Y(n_7277)
);

INVx1_ASAP7_75t_L g7278 ( 
.A(n_7030),
.Y(n_7278)
);

NAND2xp5_ASAP7_75t_L g7279 ( 
.A(n_7097),
.B(n_790),
.Y(n_7279)
);

INVx1_ASAP7_75t_L g7280 ( 
.A(n_7030),
.Y(n_7280)
);

OR2x2_ASAP7_75t_L g7281 ( 
.A(n_7024),
.B(n_790),
.Y(n_7281)
);

OR2x2_ASAP7_75t_L g7282 ( 
.A(n_7024),
.B(n_791),
.Y(n_7282)
);

INVx1_ASAP7_75t_L g7283 ( 
.A(n_7030),
.Y(n_7283)
);

INVx1_ASAP7_75t_L g7284 ( 
.A(n_7030),
.Y(n_7284)
);

NOR3xp33_ASAP7_75t_L g7285 ( 
.A(n_7055),
.B(n_791),
.C(n_792),
.Y(n_7285)
);

AOI21xp33_ASAP7_75t_L g7286 ( 
.A1(n_7130),
.A2(n_793),
.B(n_794),
.Y(n_7286)
);

AND2x4_ASAP7_75t_L g7287 ( 
.A(n_7024),
.B(n_794),
.Y(n_7287)
);

INVx1_ASAP7_75t_L g7288 ( 
.A(n_7030),
.Y(n_7288)
);

INVx1_ASAP7_75t_L g7289 ( 
.A(n_7030),
.Y(n_7289)
);

NAND2xp5_ASAP7_75t_L g7290 ( 
.A(n_7097),
.B(n_795),
.Y(n_7290)
);

AND2x4_ASAP7_75t_L g7291 ( 
.A(n_7024),
.B(n_795),
.Y(n_7291)
);

AND2x2_ASAP7_75t_L g7292 ( 
.A(n_7030),
.B(n_795),
.Y(n_7292)
);

INVx2_ASAP7_75t_L g7293 ( 
.A(n_7024),
.Y(n_7293)
);

INVx2_ASAP7_75t_L g7294 ( 
.A(n_7024),
.Y(n_7294)
);

INVx1_ASAP7_75t_L g7295 ( 
.A(n_7030),
.Y(n_7295)
);

AND2x2_ASAP7_75t_L g7296 ( 
.A(n_7030),
.B(n_796),
.Y(n_7296)
);

INVx2_ASAP7_75t_L g7297 ( 
.A(n_7024),
.Y(n_7297)
);

OAI22xp5_ASAP7_75t_L g7298 ( 
.A1(n_7203),
.A2(n_798),
.B1(n_796),
.B2(n_797),
.Y(n_7298)
);

HB1xp67_ASAP7_75t_L g7299 ( 
.A(n_7297),
.Y(n_7299)
);

INVx2_ASAP7_75t_L g7300 ( 
.A(n_7293),
.Y(n_7300)
);

AND2x2_ASAP7_75t_L g7301 ( 
.A(n_7160),
.B(n_1058),
.Y(n_7301)
);

INVx1_ASAP7_75t_SL g7302 ( 
.A(n_7197),
.Y(n_7302)
);

INVx1_ASAP7_75t_L g7303 ( 
.A(n_7161),
.Y(n_7303)
);

INVxp67_ASAP7_75t_SL g7304 ( 
.A(n_7279),
.Y(n_7304)
);

AOI22xp33_ASAP7_75t_L g7305 ( 
.A1(n_7294),
.A2(n_799),
.B1(n_797),
.B2(n_798),
.Y(n_7305)
);

INVx2_ASAP7_75t_L g7306 ( 
.A(n_7183),
.Y(n_7306)
);

INVx1_ASAP7_75t_L g7307 ( 
.A(n_7290),
.Y(n_7307)
);

NAND2xp5_ASAP7_75t_L g7308 ( 
.A(n_7291),
.B(n_797),
.Y(n_7308)
);

INVx1_ASAP7_75t_L g7309 ( 
.A(n_7291),
.Y(n_7309)
);

AND2x2_ASAP7_75t_L g7310 ( 
.A(n_7221),
.B(n_799),
.Y(n_7310)
);

INVx2_ASAP7_75t_L g7311 ( 
.A(n_7175),
.Y(n_7311)
);

INVx2_ASAP7_75t_L g7312 ( 
.A(n_7206),
.Y(n_7312)
);

OAI22xp5_ASAP7_75t_L g7313 ( 
.A1(n_7207),
.A2(n_801),
.B1(n_799),
.B2(n_800),
.Y(n_7313)
);

NAND2xp5_ASAP7_75t_L g7314 ( 
.A(n_7287),
.B(n_800),
.Y(n_7314)
);

NAND2x1_ASAP7_75t_SL g7315 ( 
.A(n_7292),
.B(n_800),
.Y(n_7315)
);

AND2x2_ASAP7_75t_L g7316 ( 
.A(n_7296),
.B(n_801),
.Y(n_7316)
);

NAND2xp5_ASAP7_75t_L g7317 ( 
.A(n_7262),
.B(n_801),
.Y(n_7317)
);

NAND2xp5_ASAP7_75t_L g7318 ( 
.A(n_7262),
.B(n_802),
.Y(n_7318)
);

AOI22xp33_ASAP7_75t_L g7319 ( 
.A1(n_7218),
.A2(n_804),
.B1(n_802),
.B2(n_803),
.Y(n_7319)
);

INVx1_ASAP7_75t_L g7320 ( 
.A(n_7164),
.Y(n_7320)
);

NAND2x1p5_ASAP7_75t_L g7321 ( 
.A(n_7249),
.B(n_802),
.Y(n_7321)
);

NAND2x1p5_ASAP7_75t_L g7322 ( 
.A(n_7210),
.B(n_803),
.Y(n_7322)
);

INVx1_ASAP7_75t_L g7323 ( 
.A(n_7166),
.Y(n_7323)
);

OR2x2_ASAP7_75t_L g7324 ( 
.A(n_7199),
.B(n_803),
.Y(n_7324)
);

INVx2_ASAP7_75t_L g7325 ( 
.A(n_7174),
.Y(n_7325)
);

INVx1_ASAP7_75t_L g7326 ( 
.A(n_7212),
.Y(n_7326)
);

NAND2xp5_ASAP7_75t_L g7327 ( 
.A(n_7258),
.B(n_804),
.Y(n_7327)
);

AOI21xp5_ASAP7_75t_L g7328 ( 
.A1(n_7196),
.A2(n_805),
.B(n_806),
.Y(n_7328)
);

AOI22xp33_ASAP7_75t_L g7329 ( 
.A1(n_7169),
.A2(n_807),
.B1(n_805),
.B2(n_806),
.Y(n_7329)
);

BUFx3_ASAP7_75t_L g7330 ( 
.A(n_7229),
.Y(n_7330)
);

HB1xp67_ASAP7_75t_L g7331 ( 
.A(n_7212),
.Y(n_7331)
);

INVx1_ASAP7_75t_SL g7332 ( 
.A(n_7186),
.Y(n_7332)
);

AND2x2_ASAP7_75t_L g7333 ( 
.A(n_7241),
.B(n_1053),
.Y(n_7333)
);

NAND2xp5_ASAP7_75t_SL g7334 ( 
.A(n_7238),
.B(n_1053),
.Y(n_7334)
);

INVx1_ASAP7_75t_L g7335 ( 
.A(n_7205),
.Y(n_7335)
);

AOI22xp33_ASAP7_75t_L g7336 ( 
.A1(n_7188),
.A2(n_808),
.B1(n_806),
.B2(n_807),
.Y(n_7336)
);

HB1xp67_ASAP7_75t_L g7337 ( 
.A(n_7236),
.Y(n_7337)
);

NOR2x1_ASAP7_75t_R g7338 ( 
.A(n_7176),
.B(n_7178),
.Y(n_7338)
);

INVx1_ASAP7_75t_SL g7339 ( 
.A(n_7281),
.Y(n_7339)
);

INVx3_ASAP7_75t_L g7340 ( 
.A(n_7282),
.Y(n_7340)
);

NAND2xp5_ASAP7_75t_L g7341 ( 
.A(n_7256),
.B(n_7277),
.Y(n_7341)
);

INVx1_ASAP7_75t_SL g7342 ( 
.A(n_7189),
.Y(n_7342)
);

OR2x2_ASAP7_75t_L g7343 ( 
.A(n_7159),
.B(n_808),
.Y(n_7343)
);

NAND3xp33_ASAP7_75t_L g7344 ( 
.A(n_7225),
.B(n_809),
.C(n_810),
.Y(n_7344)
);

INVx2_ASAP7_75t_SL g7345 ( 
.A(n_7264),
.Y(n_7345)
);

AND2x2_ASAP7_75t_L g7346 ( 
.A(n_7171),
.B(n_1053),
.Y(n_7346)
);

INVx1_ASAP7_75t_L g7347 ( 
.A(n_7266),
.Y(n_7347)
);

INVx1_ASAP7_75t_L g7348 ( 
.A(n_7271),
.Y(n_7348)
);

INVx1_ASAP7_75t_L g7349 ( 
.A(n_7211),
.Y(n_7349)
);

INVx1_ASAP7_75t_L g7350 ( 
.A(n_7220),
.Y(n_7350)
);

AND2x4_ASAP7_75t_L g7351 ( 
.A(n_7267),
.B(n_810),
.Y(n_7351)
);

AND2x2_ASAP7_75t_L g7352 ( 
.A(n_7167),
.B(n_1052),
.Y(n_7352)
);

HB1xp67_ASAP7_75t_L g7353 ( 
.A(n_7255),
.Y(n_7353)
);

AND2x2_ASAP7_75t_L g7354 ( 
.A(n_7253),
.B(n_7184),
.Y(n_7354)
);

INVx2_ASAP7_75t_L g7355 ( 
.A(n_7275),
.Y(n_7355)
);

INVx1_ASAP7_75t_L g7356 ( 
.A(n_7235),
.Y(n_7356)
);

INVxp67_ASAP7_75t_SL g7357 ( 
.A(n_7223),
.Y(n_7357)
);

INVx1_ASAP7_75t_L g7358 ( 
.A(n_7244),
.Y(n_7358)
);

INVx1_ASAP7_75t_SL g7359 ( 
.A(n_7190),
.Y(n_7359)
);

AND2x4_ASAP7_75t_L g7360 ( 
.A(n_7215),
.B(n_811),
.Y(n_7360)
);

AND2x4_ASAP7_75t_SL g7361 ( 
.A(n_7170),
.B(n_811),
.Y(n_7361)
);

INVx2_ASAP7_75t_SL g7362 ( 
.A(n_7192),
.Y(n_7362)
);

AOI22xp33_ASAP7_75t_L g7363 ( 
.A1(n_7285),
.A2(n_813),
.B1(n_811),
.B2(n_812),
.Y(n_7363)
);

NAND2xp5_ASAP7_75t_L g7364 ( 
.A(n_7257),
.B(n_812),
.Y(n_7364)
);

INVx1_ASAP7_75t_L g7365 ( 
.A(n_7200),
.Y(n_7365)
);

INVx1_ASAP7_75t_L g7366 ( 
.A(n_7268),
.Y(n_7366)
);

NAND2xp5_ASAP7_75t_L g7367 ( 
.A(n_7219),
.B(n_812),
.Y(n_7367)
);

INVx1_ASAP7_75t_L g7368 ( 
.A(n_7248),
.Y(n_7368)
);

AND2x4_ASAP7_75t_L g7369 ( 
.A(n_7204),
.B(n_813),
.Y(n_7369)
);

INVx1_ASAP7_75t_L g7370 ( 
.A(n_7228),
.Y(n_7370)
);

AOI22x1_ASAP7_75t_L g7371 ( 
.A1(n_7173),
.A2(n_815),
.B1(n_813),
.B2(n_814),
.Y(n_7371)
);

NAND2xp5_ASAP7_75t_L g7372 ( 
.A(n_7201),
.B(n_814),
.Y(n_7372)
);

AOI22xp33_ASAP7_75t_SL g7373 ( 
.A1(n_7179),
.A2(n_817),
.B1(n_815),
.B2(n_816),
.Y(n_7373)
);

INVx1_ASAP7_75t_L g7374 ( 
.A(n_7202),
.Y(n_7374)
);

INVx1_ASAP7_75t_L g7375 ( 
.A(n_7272),
.Y(n_7375)
);

AOI22xp33_ASAP7_75t_L g7376 ( 
.A1(n_7185),
.A2(n_818),
.B1(n_816),
.B2(n_817),
.Y(n_7376)
);

INVx1_ASAP7_75t_L g7377 ( 
.A(n_7217),
.Y(n_7377)
);

INVx1_ASAP7_75t_L g7378 ( 
.A(n_7278),
.Y(n_7378)
);

INVx2_ASAP7_75t_L g7379 ( 
.A(n_7181),
.Y(n_7379)
);

NAND2xp5_ASAP7_75t_L g7380 ( 
.A(n_7226),
.B(n_816),
.Y(n_7380)
);

INVx1_ASAP7_75t_L g7381 ( 
.A(n_7280),
.Y(n_7381)
);

OR2x2_ASAP7_75t_L g7382 ( 
.A(n_7302),
.B(n_7283),
.Y(n_7382)
);

AOI221xp5_ASAP7_75t_L g7383 ( 
.A1(n_7313),
.A2(n_7286),
.B1(n_7250),
.B2(n_7214),
.C(n_7163),
.Y(n_7383)
);

OAI32xp33_ASAP7_75t_L g7384 ( 
.A1(n_7332),
.A2(n_7193),
.A3(n_7182),
.B1(n_7177),
.B2(n_7222),
.Y(n_7384)
);

INVx1_ASAP7_75t_L g7385 ( 
.A(n_7299),
.Y(n_7385)
);

INVx2_ASAP7_75t_L g7386 ( 
.A(n_7300),
.Y(n_7386)
);

AOI21xp5_ASAP7_75t_L g7387 ( 
.A1(n_7334),
.A2(n_7254),
.B(n_7213),
.Y(n_7387)
);

AOI22xp5_ASAP7_75t_L g7388 ( 
.A1(n_7312),
.A2(n_7172),
.B1(n_7194),
.B2(n_7180),
.Y(n_7388)
);

BUFx2_ASAP7_75t_L g7389 ( 
.A(n_7351),
.Y(n_7389)
);

AND2x2_ASAP7_75t_L g7390 ( 
.A(n_7346),
.B(n_7284),
.Y(n_7390)
);

INVxp67_ASAP7_75t_L g7391 ( 
.A(n_7338),
.Y(n_7391)
);

INVx1_ASAP7_75t_SL g7392 ( 
.A(n_7306),
.Y(n_7392)
);

OAI211xp5_ASAP7_75t_SL g7393 ( 
.A1(n_7373),
.A2(n_7158),
.B(n_7273),
.C(n_7231),
.Y(n_7393)
);

INVx1_ASAP7_75t_L g7394 ( 
.A(n_7308),
.Y(n_7394)
);

OAI22xp5_ASAP7_75t_L g7395 ( 
.A1(n_7311),
.A2(n_7288),
.B1(n_7295),
.B2(n_7289),
.Y(n_7395)
);

INVx1_ASAP7_75t_L g7396 ( 
.A(n_7317),
.Y(n_7396)
);

NAND3xp33_ASAP7_75t_SL g7397 ( 
.A(n_7328),
.B(n_7216),
.C(n_7239),
.Y(n_7397)
);

CKINVDCx20_ASAP7_75t_R g7398 ( 
.A(n_7330),
.Y(n_7398)
);

AND2x2_ASAP7_75t_L g7399 ( 
.A(n_7310),
.B(n_7237),
.Y(n_7399)
);

NAND2xp5_ASAP7_75t_L g7400 ( 
.A(n_7351),
.B(n_7246),
.Y(n_7400)
);

AND2x2_ASAP7_75t_L g7401 ( 
.A(n_7301),
.B(n_7247),
.Y(n_7401)
);

NAND3xp33_ASAP7_75t_L g7402 ( 
.A(n_7371),
.B(n_7209),
.C(n_7243),
.Y(n_7402)
);

NAND2xp5_ASAP7_75t_SL g7403 ( 
.A(n_7355),
.B(n_7187),
.Y(n_7403)
);

NAND2xp5_ASAP7_75t_L g7404 ( 
.A(n_7352),
.B(n_7242),
.Y(n_7404)
);

INVx2_ASAP7_75t_L g7405 ( 
.A(n_7325),
.Y(n_7405)
);

OR2x6_ASAP7_75t_L g7406 ( 
.A(n_7345),
.B(n_7234),
.Y(n_7406)
);

INVx1_ASAP7_75t_L g7407 ( 
.A(n_7318),
.Y(n_7407)
);

INVx1_ASAP7_75t_L g7408 ( 
.A(n_7353),
.Y(n_7408)
);

INVx1_ASAP7_75t_L g7409 ( 
.A(n_7314),
.Y(n_7409)
);

INVx2_ASAP7_75t_L g7410 ( 
.A(n_7335),
.Y(n_7410)
);

AOI222xp33_ASAP7_75t_L g7411 ( 
.A1(n_7359),
.A2(n_7270),
.B1(n_7269),
.B2(n_7265),
.C1(n_7263),
.C2(n_7251),
.Y(n_7411)
);

INVx1_ASAP7_75t_L g7412 ( 
.A(n_7322),
.Y(n_7412)
);

OAI321xp33_ASAP7_75t_L g7413 ( 
.A1(n_7341),
.A2(n_7195),
.A3(n_7245),
.B1(n_7208),
.B2(n_7165),
.C(n_7168),
.Y(n_7413)
);

A2O1A1Ixp33_ASAP7_75t_L g7414 ( 
.A1(n_7320),
.A2(n_7162),
.B(n_7227),
.C(n_7224),
.Y(n_7414)
);

OR2x2_ASAP7_75t_L g7415 ( 
.A(n_7323),
.B(n_7274),
.Y(n_7415)
);

AOI21xp33_ASAP7_75t_SL g7416 ( 
.A1(n_7327),
.A2(n_7259),
.B(n_7232),
.Y(n_7416)
);

INVx1_ASAP7_75t_L g7417 ( 
.A(n_7331),
.Y(n_7417)
);

OAI322xp33_ASAP7_75t_L g7418 ( 
.A1(n_7342),
.A2(n_7240),
.A3(n_7261),
.B1(n_7252),
.B2(n_7276),
.C1(n_7198),
.C2(n_7191),
.Y(n_7418)
);

OAI22xp33_ASAP7_75t_SL g7419 ( 
.A1(n_7364),
.A2(n_7260),
.B1(n_7233),
.B2(n_7230),
.Y(n_7419)
);

INVxp67_ASAP7_75t_SL g7420 ( 
.A(n_7321),
.Y(n_7420)
);

INVx1_ASAP7_75t_L g7421 ( 
.A(n_7360),
.Y(n_7421)
);

INVx2_ASAP7_75t_L g7422 ( 
.A(n_7309),
.Y(n_7422)
);

NAND2xp5_ASAP7_75t_L g7423 ( 
.A(n_7316),
.B(n_817),
.Y(n_7423)
);

NAND4xp25_ASAP7_75t_L g7424 ( 
.A(n_7354),
.B(n_7363),
.C(n_7376),
.D(n_7329),
.Y(n_7424)
);

NAND2xp5_ASAP7_75t_L g7425 ( 
.A(n_7360),
.B(n_818),
.Y(n_7425)
);

AOI22xp5_ASAP7_75t_L g7426 ( 
.A1(n_7303),
.A2(n_821),
.B1(n_819),
.B2(n_820),
.Y(n_7426)
);

OAI322xp33_ASAP7_75t_L g7427 ( 
.A1(n_7343),
.A2(n_819),
.A3(n_820),
.B1(n_821),
.B2(n_822),
.C1(n_823),
.C2(n_824),
.Y(n_7427)
);

AND2x2_ASAP7_75t_L g7428 ( 
.A(n_7333),
.B(n_819),
.Y(n_7428)
);

INVx2_ASAP7_75t_L g7429 ( 
.A(n_7379),
.Y(n_7429)
);

AOI222xp33_ASAP7_75t_L g7430 ( 
.A1(n_7347),
.A2(n_823),
.B1(n_825),
.B2(n_821),
.C1(n_822),
.C2(n_824),
.Y(n_7430)
);

NAND2xp5_ASAP7_75t_L g7431 ( 
.A(n_7369),
.B(n_822),
.Y(n_7431)
);

AOI21xp5_ASAP7_75t_L g7432 ( 
.A1(n_7367),
.A2(n_823),
.B(n_824),
.Y(n_7432)
);

INVx2_ASAP7_75t_L g7433 ( 
.A(n_7369),
.Y(n_7433)
);

OAI21xp5_ASAP7_75t_SL g7434 ( 
.A1(n_7319),
.A2(n_825),
.B(n_826),
.Y(n_7434)
);

INVx1_ASAP7_75t_SL g7435 ( 
.A(n_7339),
.Y(n_7435)
);

OAI221xp5_ASAP7_75t_L g7436 ( 
.A1(n_7305),
.A2(n_827),
.B1(n_825),
.B2(n_826),
.C(n_828),
.Y(n_7436)
);

NAND2xp5_ASAP7_75t_L g7437 ( 
.A(n_7348),
.B(n_826),
.Y(n_7437)
);

AOI21xp33_ASAP7_75t_SL g7438 ( 
.A1(n_7298),
.A2(n_827),
.B(n_828),
.Y(n_7438)
);

NAND3xp33_ASAP7_75t_L g7439 ( 
.A(n_7336),
.B(n_829),
.C(n_830),
.Y(n_7439)
);

AOI22xp5_ASAP7_75t_L g7440 ( 
.A1(n_7362),
.A2(n_831),
.B1(n_829),
.B2(n_830),
.Y(n_7440)
);

NAND2xp5_ASAP7_75t_L g7441 ( 
.A(n_7326),
.B(n_831),
.Y(n_7441)
);

AOI222xp33_ASAP7_75t_L g7442 ( 
.A1(n_7361),
.A2(n_834),
.B1(n_836),
.B2(n_832),
.C1(n_833),
.C2(n_835),
.Y(n_7442)
);

INVx1_ASAP7_75t_L g7443 ( 
.A(n_7324),
.Y(n_7443)
);

AOI22xp5_ASAP7_75t_L g7444 ( 
.A1(n_7374),
.A2(n_834),
.B1(n_832),
.B2(n_833),
.Y(n_7444)
);

HB1xp67_ASAP7_75t_L g7445 ( 
.A(n_7337),
.Y(n_7445)
);

INVx1_ASAP7_75t_L g7446 ( 
.A(n_7315),
.Y(n_7446)
);

OR2x2_ASAP7_75t_L g7447 ( 
.A(n_7372),
.B(n_832),
.Y(n_7447)
);

O2A1O1Ixp33_ASAP7_75t_L g7448 ( 
.A1(n_7380),
.A2(n_836),
.B(n_834),
.C(n_835),
.Y(n_7448)
);

NAND2xp5_ASAP7_75t_L g7449 ( 
.A(n_7340),
.B(n_7357),
.Y(n_7449)
);

OR2x2_ASAP7_75t_L g7450 ( 
.A(n_7340),
.B(n_836),
.Y(n_7450)
);

OAI32xp33_ASAP7_75t_L g7451 ( 
.A1(n_7370),
.A2(n_7381),
.A3(n_7378),
.B1(n_7366),
.B2(n_7368),
.Y(n_7451)
);

INVxp67_ASAP7_75t_L g7452 ( 
.A(n_7344),
.Y(n_7452)
);

OAI22xp33_ASAP7_75t_SL g7453 ( 
.A1(n_7377),
.A2(n_839),
.B1(n_837),
.B2(n_838),
.Y(n_7453)
);

AOI22xp33_ASAP7_75t_L g7454 ( 
.A1(n_7307),
.A2(n_839),
.B1(n_837),
.B2(n_838),
.Y(n_7454)
);

INVx1_ASAP7_75t_SL g7455 ( 
.A(n_7349),
.Y(n_7455)
);

INVxp67_ASAP7_75t_SL g7456 ( 
.A(n_7304),
.Y(n_7456)
);

INVx1_ASAP7_75t_SL g7457 ( 
.A(n_7350),
.Y(n_7457)
);

O2A1O1Ixp33_ASAP7_75t_L g7458 ( 
.A1(n_7356),
.A2(n_841),
.B(n_839),
.C(n_840),
.Y(n_7458)
);

INVx1_ASAP7_75t_L g7459 ( 
.A(n_7358),
.Y(n_7459)
);

NAND2xp5_ASAP7_75t_L g7460 ( 
.A(n_7365),
.B(n_840),
.Y(n_7460)
);

AND2x2_ASAP7_75t_L g7461 ( 
.A(n_7375),
.B(n_840),
.Y(n_7461)
);

AND2x2_ASAP7_75t_L g7462 ( 
.A(n_7346),
.B(n_841),
.Y(n_7462)
);

AOI21xp5_ASAP7_75t_L g7463 ( 
.A1(n_7334),
.A2(n_842),
.B(n_843),
.Y(n_7463)
);

INVx1_ASAP7_75t_L g7464 ( 
.A(n_7299),
.Y(n_7464)
);

INVx2_ASAP7_75t_L g7465 ( 
.A(n_7300),
.Y(n_7465)
);

INVx1_ASAP7_75t_L g7466 ( 
.A(n_7299),
.Y(n_7466)
);

O2A1O1Ixp33_ASAP7_75t_L g7467 ( 
.A1(n_7313),
.A2(n_844),
.B(n_842),
.C(n_843),
.Y(n_7467)
);

NAND2xp5_ASAP7_75t_L g7468 ( 
.A(n_7300),
.B(n_844),
.Y(n_7468)
);

INVx2_ASAP7_75t_L g7469 ( 
.A(n_7300),
.Y(n_7469)
);

INVxp67_ASAP7_75t_SL g7470 ( 
.A(n_7299),
.Y(n_7470)
);

OA21x2_ASAP7_75t_L g7471 ( 
.A1(n_7328),
.A2(n_845),
.B(n_846),
.Y(n_7471)
);

INVx1_ASAP7_75t_L g7472 ( 
.A(n_7299),
.Y(n_7472)
);

INVx1_ASAP7_75t_L g7473 ( 
.A(n_7299),
.Y(n_7473)
);

INVx2_ASAP7_75t_SL g7474 ( 
.A(n_7300),
.Y(n_7474)
);

OAI21xp33_ASAP7_75t_L g7475 ( 
.A1(n_7302),
.A2(n_845),
.B(n_846),
.Y(n_7475)
);

AND2x2_ASAP7_75t_L g7476 ( 
.A(n_7346),
.B(n_847),
.Y(n_7476)
);

INVx1_ASAP7_75t_L g7477 ( 
.A(n_7470),
.Y(n_7477)
);

INVx1_ASAP7_75t_L g7478 ( 
.A(n_7398),
.Y(n_7478)
);

NAND2xp5_ASAP7_75t_L g7479 ( 
.A(n_7392),
.B(n_847),
.Y(n_7479)
);

INVx1_ASAP7_75t_L g7480 ( 
.A(n_7386),
.Y(n_7480)
);

OR2x2_ASAP7_75t_L g7481 ( 
.A(n_7465),
.B(n_1052),
.Y(n_7481)
);

NAND2xp5_ASAP7_75t_L g7482 ( 
.A(n_7474),
.B(n_847),
.Y(n_7482)
);

NAND2xp5_ASAP7_75t_L g7483 ( 
.A(n_7469),
.B(n_848),
.Y(n_7483)
);

AOI21xp33_ASAP7_75t_L g7484 ( 
.A1(n_7430),
.A2(n_849),
.B(n_850),
.Y(n_7484)
);

HB1xp67_ASAP7_75t_L g7485 ( 
.A(n_7445),
.Y(n_7485)
);

OAI22xp5_ASAP7_75t_L g7486 ( 
.A1(n_7388),
.A2(n_851),
.B1(n_849),
.B2(n_850),
.Y(n_7486)
);

INVx1_ASAP7_75t_L g7487 ( 
.A(n_7425),
.Y(n_7487)
);

INVx1_ASAP7_75t_SL g7488 ( 
.A(n_7382),
.Y(n_7488)
);

INVx1_ASAP7_75t_L g7489 ( 
.A(n_7431),
.Y(n_7489)
);

AND2x4_ASAP7_75t_L g7490 ( 
.A(n_7385),
.B(n_849),
.Y(n_7490)
);

INVx2_ASAP7_75t_L g7491 ( 
.A(n_7429),
.Y(n_7491)
);

AOI22xp5_ASAP7_75t_L g7492 ( 
.A1(n_7391),
.A2(n_1052),
.B1(n_853),
.B2(n_851),
.Y(n_7492)
);

A2O1A1Ixp33_ASAP7_75t_L g7493 ( 
.A1(n_7458),
.A2(n_853),
.B(n_851),
.C(n_852),
.Y(n_7493)
);

NAND2xp5_ASAP7_75t_SL g7494 ( 
.A(n_7453),
.B(n_852),
.Y(n_7494)
);

INVx1_ASAP7_75t_L g7495 ( 
.A(n_7415),
.Y(n_7495)
);

OAI22xp33_ASAP7_75t_L g7496 ( 
.A1(n_7440),
.A2(n_854),
.B1(n_852),
.B2(n_853),
.Y(n_7496)
);

INVx1_ASAP7_75t_L g7497 ( 
.A(n_7464),
.Y(n_7497)
);

OR2x2_ASAP7_75t_L g7498 ( 
.A(n_7466),
.B(n_1051),
.Y(n_7498)
);

AOI22xp5_ASAP7_75t_L g7499 ( 
.A1(n_7472),
.A2(n_7473),
.B1(n_7417),
.B2(n_7397),
.Y(n_7499)
);

OR2x2_ASAP7_75t_L g7500 ( 
.A(n_7405),
.B(n_854),
.Y(n_7500)
);

INVx1_ASAP7_75t_L g7501 ( 
.A(n_7441),
.Y(n_7501)
);

NAND2xp5_ASAP7_75t_L g7502 ( 
.A(n_7462),
.B(n_7476),
.Y(n_7502)
);

AOI22xp5_ASAP7_75t_L g7503 ( 
.A1(n_7435),
.A2(n_1050),
.B1(n_857),
.B2(n_855),
.Y(n_7503)
);

AOI22xp33_ASAP7_75t_L g7504 ( 
.A1(n_7410),
.A2(n_857),
.B1(n_855),
.B2(n_856),
.Y(n_7504)
);

HB1xp67_ASAP7_75t_L g7505 ( 
.A(n_7450),
.Y(n_7505)
);

NAND2xp33_ASAP7_75t_R g7506 ( 
.A(n_7471),
.B(n_7389),
.Y(n_7506)
);

INVx2_ASAP7_75t_L g7507 ( 
.A(n_7433),
.Y(n_7507)
);

AOI22xp33_ASAP7_75t_SL g7508 ( 
.A1(n_7456),
.A2(n_858),
.B1(n_856),
.B2(n_857),
.Y(n_7508)
);

INVx1_ASAP7_75t_L g7509 ( 
.A(n_7468),
.Y(n_7509)
);

NAND2xp5_ASAP7_75t_L g7510 ( 
.A(n_7428),
.B(n_856),
.Y(n_7510)
);

OR2x2_ASAP7_75t_L g7511 ( 
.A(n_7408),
.B(n_1048),
.Y(n_7511)
);

AOI21xp5_ASAP7_75t_L g7512 ( 
.A1(n_7403),
.A2(n_7423),
.B(n_7437),
.Y(n_7512)
);

OAI321xp33_ASAP7_75t_L g7513 ( 
.A1(n_7393),
.A2(n_858),
.A3(n_859),
.B1(n_860),
.B2(n_861),
.C(n_862),
.Y(n_7513)
);

INVx1_ASAP7_75t_L g7514 ( 
.A(n_7461),
.Y(n_7514)
);

AND2x2_ASAP7_75t_L g7515 ( 
.A(n_7399),
.B(n_7401),
.Y(n_7515)
);

AOI221xp5_ASAP7_75t_L g7516 ( 
.A1(n_7384),
.A2(n_860),
.B1(n_858),
.B2(n_859),
.C(n_862),
.Y(n_7516)
);

INVx2_ASAP7_75t_SL g7517 ( 
.A(n_7422),
.Y(n_7517)
);

AND2x2_ASAP7_75t_L g7518 ( 
.A(n_7390),
.B(n_859),
.Y(n_7518)
);

AND2x2_ASAP7_75t_L g7519 ( 
.A(n_7421),
.B(n_862),
.Y(n_7519)
);

INVx1_ASAP7_75t_L g7520 ( 
.A(n_7400),
.Y(n_7520)
);

AOI221x1_ASAP7_75t_L g7521 ( 
.A1(n_7395),
.A2(n_865),
.B1(n_863),
.B2(n_864),
.C(n_866),
.Y(n_7521)
);

INVx2_ASAP7_75t_SL g7522 ( 
.A(n_7412),
.Y(n_7522)
);

NAND2xp5_ASAP7_75t_L g7523 ( 
.A(n_7471),
.B(n_7442),
.Y(n_7523)
);

AOI22xp33_ASAP7_75t_SL g7524 ( 
.A1(n_7485),
.A2(n_7480),
.B1(n_7477),
.B2(n_7522),
.Y(n_7524)
);

INVxp67_ASAP7_75t_L g7525 ( 
.A(n_7478),
.Y(n_7525)
);

AND2x2_ASAP7_75t_L g7526 ( 
.A(n_7515),
.B(n_7420),
.Y(n_7526)
);

AND2x2_ASAP7_75t_L g7527 ( 
.A(n_7491),
.B(n_7406),
.Y(n_7527)
);

HB1xp67_ASAP7_75t_L g7528 ( 
.A(n_7490),
.Y(n_7528)
);

NAND2xp5_ASAP7_75t_L g7529 ( 
.A(n_7490),
.B(n_7454),
.Y(n_7529)
);

INVx2_ASAP7_75t_L g7530 ( 
.A(n_7507),
.Y(n_7530)
);

INVx1_ASAP7_75t_L g7531 ( 
.A(n_7519),
.Y(n_7531)
);

INVx1_ASAP7_75t_L g7532 ( 
.A(n_7518),
.Y(n_7532)
);

INVx2_ASAP7_75t_L g7533 ( 
.A(n_7517),
.Y(n_7533)
);

OR2x2_ASAP7_75t_L g7534 ( 
.A(n_7488),
.B(n_7449),
.Y(n_7534)
);

AOI22xp5_ASAP7_75t_L g7535 ( 
.A1(n_7495),
.A2(n_7452),
.B1(n_7457),
.B2(n_7455),
.Y(n_7535)
);

INVx1_ASAP7_75t_L g7536 ( 
.A(n_7483),
.Y(n_7536)
);

AND2x2_ASAP7_75t_L g7537 ( 
.A(n_7497),
.B(n_7406),
.Y(n_7537)
);

INVx1_ASAP7_75t_L g7538 ( 
.A(n_7479),
.Y(n_7538)
);

INVx2_ASAP7_75t_SL g7539 ( 
.A(n_7481),
.Y(n_7539)
);

INVx1_ASAP7_75t_L g7540 ( 
.A(n_7498),
.Y(n_7540)
);

NAND2xp5_ASAP7_75t_L g7541 ( 
.A(n_7516),
.B(n_7444),
.Y(n_7541)
);

INVx1_ASAP7_75t_L g7542 ( 
.A(n_7511),
.Y(n_7542)
);

INVx2_ASAP7_75t_L g7543 ( 
.A(n_7520),
.Y(n_7543)
);

INVx1_ASAP7_75t_L g7544 ( 
.A(n_7482),
.Y(n_7544)
);

AND2x2_ASAP7_75t_L g7545 ( 
.A(n_7505),
.B(n_7443),
.Y(n_7545)
);

OR2x2_ASAP7_75t_L g7546 ( 
.A(n_7502),
.B(n_7404),
.Y(n_7546)
);

INVx2_ASAP7_75t_SL g7547 ( 
.A(n_7500),
.Y(n_7547)
);

NAND2x1p5_ASAP7_75t_L g7548 ( 
.A(n_7499),
.B(n_7459),
.Y(n_7548)
);

INVx1_ASAP7_75t_L g7549 ( 
.A(n_7523),
.Y(n_7549)
);

AND2x2_ASAP7_75t_L g7550 ( 
.A(n_7514),
.B(n_7411),
.Y(n_7550)
);

INVx1_ASAP7_75t_L g7551 ( 
.A(n_7510),
.Y(n_7551)
);

INVx1_ASAP7_75t_L g7552 ( 
.A(n_7503),
.Y(n_7552)
);

NOR2xp33_ASAP7_75t_L g7553 ( 
.A(n_7513),
.B(n_7413),
.Y(n_7553)
);

NAND2xp5_ASAP7_75t_L g7554 ( 
.A(n_7508),
.B(n_7504),
.Y(n_7554)
);

AND2x2_ASAP7_75t_L g7555 ( 
.A(n_7501),
.B(n_7446),
.Y(n_7555)
);

INVx1_ASAP7_75t_L g7556 ( 
.A(n_7494),
.Y(n_7556)
);

INVx1_ASAP7_75t_SL g7557 ( 
.A(n_7509),
.Y(n_7557)
);

INVx1_ASAP7_75t_SL g7558 ( 
.A(n_7487),
.Y(n_7558)
);

NAND2xp5_ASAP7_75t_L g7559 ( 
.A(n_7492),
.B(n_7426),
.Y(n_7559)
);

OR2x2_ASAP7_75t_L g7560 ( 
.A(n_7486),
.B(n_7460),
.Y(n_7560)
);

AND2x4_ASAP7_75t_L g7561 ( 
.A(n_7489),
.B(n_7414),
.Y(n_7561)
);

INVx2_ASAP7_75t_L g7562 ( 
.A(n_7506),
.Y(n_7562)
);

OR2x2_ASAP7_75t_L g7563 ( 
.A(n_7493),
.B(n_7447),
.Y(n_7563)
);

NOR2xp33_ASAP7_75t_L g7564 ( 
.A(n_7484),
.B(n_7418),
.Y(n_7564)
);

NOR2xp33_ASAP7_75t_L g7565 ( 
.A(n_7496),
.B(n_7451),
.Y(n_7565)
);

AND2x2_ASAP7_75t_L g7566 ( 
.A(n_7512),
.B(n_7394),
.Y(n_7566)
);

BUFx2_ASAP7_75t_L g7567 ( 
.A(n_7521),
.Y(n_7567)
);

INVx1_ASAP7_75t_L g7568 ( 
.A(n_7485),
.Y(n_7568)
);

INVx2_ASAP7_75t_L g7569 ( 
.A(n_7491),
.Y(n_7569)
);

INVx1_ASAP7_75t_SL g7570 ( 
.A(n_7488),
.Y(n_7570)
);

AND2x2_ASAP7_75t_L g7571 ( 
.A(n_7485),
.B(n_7396),
.Y(n_7571)
);

AND2x2_ASAP7_75t_L g7572 ( 
.A(n_7485),
.B(n_7407),
.Y(n_7572)
);

NAND2xp5_ASAP7_75t_L g7573 ( 
.A(n_7485),
.B(n_7475),
.Y(n_7573)
);

INVx1_ASAP7_75t_L g7574 ( 
.A(n_7485),
.Y(n_7574)
);

INVx1_ASAP7_75t_L g7575 ( 
.A(n_7485),
.Y(n_7575)
);

HB1xp67_ASAP7_75t_L g7576 ( 
.A(n_7485),
.Y(n_7576)
);

NAND3xp33_ASAP7_75t_L g7577 ( 
.A(n_7524),
.B(n_7383),
.C(n_7463),
.Y(n_7577)
);

NAND2xp5_ASAP7_75t_L g7578 ( 
.A(n_7526),
.B(n_7530),
.Y(n_7578)
);

NOR3xp33_ASAP7_75t_L g7579 ( 
.A(n_7549),
.B(n_7427),
.C(n_7436),
.Y(n_7579)
);

NAND2x1_ASAP7_75t_L g7580 ( 
.A(n_7569),
.B(n_7409),
.Y(n_7580)
);

NAND2xp5_ASAP7_75t_SL g7581 ( 
.A(n_7535),
.B(n_7419),
.Y(n_7581)
);

AOI221xp5_ASAP7_75t_L g7582 ( 
.A1(n_7553),
.A2(n_7438),
.B1(n_7467),
.B2(n_7448),
.C(n_7416),
.Y(n_7582)
);

OAI21xp5_ASAP7_75t_L g7583 ( 
.A1(n_7525),
.A2(n_7387),
.B(n_7432),
.Y(n_7583)
);

NAND3xp33_ASAP7_75t_L g7584 ( 
.A(n_7564),
.B(n_7439),
.C(n_7424),
.Y(n_7584)
);

NOR3xp33_ASAP7_75t_L g7585 ( 
.A(n_7570),
.B(n_7434),
.C(n_7402),
.Y(n_7585)
);

INVx1_ASAP7_75t_L g7586 ( 
.A(n_7534),
.Y(n_7586)
);

INVx1_ASAP7_75t_L g7587 ( 
.A(n_7576),
.Y(n_7587)
);

NOR2xp33_ASAP7_75t_L g7588 ( 
.A(n_7568),
.B(n_863),
.Y(n_7588)
);

INVx1_ASAP7_75t_L g7589 ( 
.A(n_7527),
.Y(n_7589)
);

NOR2x1_ASAP7_75t_L g7590 ( 
.A(n_7574),
.B(n_863),
.Y(n_7590)
);

AOI31xp33_ASAP7_75t_L g7591 ( 
.A1(n_7528),
.A2(n_866),
.A3(n_864),
.B(n_865),
.Y(n_7591)
);

NAND2xp5_ASAP7_75t_L g7592 ( 
.A(n_7575),
.B(n_7533),
.Y(n_7592)
);

NAND2xp5_ASAP7_75t_L g7593 ( 
.A(n_7543),
.B(n_864),
.Y(n_7593)
);

NAND2xp5_ASAP7_75t_SL g7594 ( 
.A(n_7562),
.B(n_7561),
.Y(n_7594)
);

NAND4xp25_ASAP7_75t_L g7595 ( 
.A(n_7546),
.B(n_867),
.C(n_865),
.D(n_866),
.Y(n_7595)
);

NAND2xp5_ASAP7_75t_SL g7596 ( 
.A(n_7561),
.B(n_7537),
.Y(n_7596)
);

INVx1_ASAP7_75t_L g7597 ( 
.A(n_7545),
.Y(n_7597)
);

OR2x2_ASAP7_75t_L g7598 ( 
.A(n_7548),
.B(n_867),
.Y(n_7598)
);

OAI21xp33_ASAP7_75t_L g7599 ( 
.A1(n_7573),
.A2(n_867),
.B(n_868),
.Y(n_7599)
);

OAI211xp5_ASAP7_75t_L g7600 ( 
.A1(n_7565),
.A2(n_870),
.B(n_868),
.C(n_869),
.Y(n_7600)
);

NOR3xp33_ASAP7_75t_SL g7601 ( 
.A(n_7556),
.B(n_7552),
.C(n_7554),
.Y(n_7601)
);

NAND4xp25_ASAP7_75t_L g7602 ( 
.A(n_7532),
.B(n_871),
.C(n_869),
.D(n_870),
.Y(n_7602)
);

INVx1_ASAP7_75t_L g7603 ( 
.A(n_7571),
.Y(n_7603)
);

NOR3xp33_ASAP7_75t_L g7604 ( 
.A(n_7572),
.B(n_1048),
.C(n_869),
.Y(n_7604)
);

NOR3xp33_ASAP7_75t_L g7605 ( 
.A(n_7550),
.B(n_1047),
.C(n_870),
.Y(n_7605)
);

AOI21xp5_ASAP7_75t_L g7606 ( 
.A1(n_7541),
.A2(n_872),
.B(n_873),
.Y(n_7606)
);

NAND2xp5_ASAP7_75t_SL g7607 ( 
.A(n_7558),
.B(n_872),
.Y(n_7607)
);

OAI21xp33_ASAP7_75t_SL g7608 ( 
.A1(n_7529),
.A2(n_873),
.B(n_874),
.Y(n_7608)
);

AND2x2_ASAP7_75t_L g7609 ( 
.A(n_7531),
.B(n_873),
.Y(n_7609)
);

NOR3xp33_ASAP7_75t_L g7610 ( 
.A(n_7566),
.B(n_1046),
.C(n_874),
.Y(n_7610)
);

NOR2xp33_ASAP7_75t_L g7611 ( 
.A(n_7557),
.B(n_874),
.Y(n_7611)
);

NAND3xp33_ASAP7_75t_L g7612 ( 
.A(n_7578),
.B(n_7542),
.C(n_7540),
.Y(n_7612)
);

OAI21xp33_ASAP7_75t_L g7613 ( 
.A1(n_7586),
.A2(n_7555),
.B(n_7547),
.Y(n_7613)
);

NAND3xp33_ASAP7_75t_L g7614 ( 
.A(n_7579),
.B(n_7605),
.C(n_7585),
.Y(n_7614)
);

NOR3xp33_ASAP7_75t_L g7615 ( 
.A(n_7577),
.B(n_7538),
.C(n_7536),
.Y(n_7615)
);

INVx2_ASAP7_75t_SL g7616 ( 
.A(n_7589),
.Y(n_7616)
);

NAND2xp5_ASAP7_75t_SL g7617 ( 
.A(n_7582),
.B(n_7567),
.Y(n_7617)
);

AND2x2_ASAP7_75t_L g7618 ( 
.A(n_7603),
.B(n_7539),
.Y(n_7618)
);

INVx1_ASAP7_75t_L g7619 ( 
.A(n_7592),
.Y(n_7619)
);

O2A1O1Ixp33_ASAP7_75t_L g7620 ( 
.A1(n_7591),
.A2(n_7559),
.B(n_7536),
.C(n_7563),
.Y(n_7620)
);

NAND3xp33_ASAP7_75t_SL g7621 ( 
.A(n_7604),
.B(n_7560),
.C(n_7544),
.Y(n_7621)
);

AOI221xp5_ASAP7_75t_L g7622 ( 
.A1(n_7599),
.A2(n_7551),
.B1(n_877),
.B2(n_875),
.C(n_876),
.Y(n_7622)
);

AND2x2_ASAP7_75t_L g7623 ( 
.A(n_7597),
.B(n_875),
.Y(n_7623)
);

OAI21xp33_ASAP7_75t_SL g7624 ( 
.A1(n_7581),
.A2(n_875),
.B(n_876),
.Y(n_7624)
);

INVx1_ASAP7_75t_L g7625 ( 
.A(n_7609),
.Y(n_7625)
);

AND2x4_ASAP7_75t_L g7626 ( 
.A(n_7587),
.B(n_876),
.Y(n_7626)
);

NAND3xp33_ASAP7_75t_L g7627 ( 
.A(n_7610),
.B(n_877),
.C(n_878),
.Y(n_7627)
);

NAND2xp5_ASAP7_75t_SL g7628 ( 
.A(n_7606),
.B(n_877),
.Y(n_7628)
);

CKINVDCx14_ASAP7_75t_R g7629 ( 
.A(n_7598),
.Y(n_7629)
);

INVx1_ASAP7_75t_L g7630 ( 
.A(n_7593),
.Y(n_7630)
);

NOR2xp33_ASAP7_75t_L g7631 ( 
.A(n_7594),
.B(n_878),
.Y(n_7631)
);

NAND3xp33_ASAP7_75t_L g7632 ( 
.A(n_7601),
.B(n_7588),
.C(n_7584),
.Y(n_7632)
);

INVx1_ASAP7_75t_L g7633 ( 
.A(n_7590),
.Y(n_7633)
);

INVx1_ASAP7_75t_L g7634 ( 
.A(n_7580),
.Y(n_7634)
);

NOR2x1_ASAP7_75t_L g7635 ( 
.A(n_7596),
.B(n_878),
.Y(n_7635)
);

AND3x2_ASAP7_75t_L g7636 ( 
.A(n_7611),
.B(n_7583),
.C(n_7608),
.Y(n_7636)
);

NAND2xp5_ASAP7_75t_L g7637 ( 
.A(n_7600),
.B(n_879),
.Y(n_7637)
);

AOI22xp5_ASAP7_75t_L g7638 ( 
.A1(n_7602),
.A2(n_881),
.B1(n_879),
.B2(n_880),
.Y(n_7638)
);

NOR3xp33_ASAP7_75t_SL g7639 ( 
.A(n_7595),
.B(n_879),
.C(n_880),
.Y(n_7639)
);

NAND4xp25_ASAP7_75t_L g7640 ( 
.A(n_7607),
.B(n_882),
.C(n_880),
.D(n_881),
.Y(n_7640)
);

INVx2_ASAP7_75t_SL g7641 ( 
.A(n_7578),
.Y(n_7641)
);

NOR3xp33_ASAP7_75t_L g7642 ( 
.A(n_7578),
.B(n_881),
.C(n_882),
.Y(n_7642)
);

INVx2_ASAP7_75t_L g7643 ( 
.A(n_7578),
.Y(n_7643)
);

NAND2xp5_ASAP7_75t_L g7644 ( 
.A(n_7578),
.B(n_1046),
.Y(n_7644)
);

NAND4xp25_ASAP7_75t_L g7645 ( 
.A(n_7578),
.B(n_884),
.C(n_882),
.D(n_883),
.Y(n_7645)
);

NOR3x1_ASAP7_75t_L g7646 ( 
.A(n_7578),
.B(n_883),
.C(n_884),
.Y(n_7646)
);

AOI21xp5_ASAP7_75t_L g7647 ( 
.A1(n_7578),
.A2(n_883),
.B(n_884),
.Y(n_7647)
);

INVxp67_ASAP7_75t_L g7648 ( 
.A(n_7578),
.Y(n_7648)
);

INVx1_ASAP7_75t_L g7649 ( 
.A(n_7578),
.Y(n_7649)
);

NOR3xp33_ASAP7_75t_L g7650 ( 
.A(n_7578),
.B(n_885),
.C(n_886),
.Y(n_7650)
);

AOI221xp5_ASAP7_75t_L g7651 ( 
.A1(n_7591),
.A2(n_887),
.B1(n_885),
.B2(n_886),
.C(n_888),
.Y(n_7651)
);

AOI21xp5_ASAP7_75t_L g7652 ( 
.A1(n_7578),
.A2(n_886),
.B(n_887),
.Y(n_7652)
);

NAND4xp25_ASAP7_75t_L g7653 ( 
.A(n_7578),
.B(n_889),
.C(n_887),
.D(n_888),
.Y(n_7653)
);

NAND2xp5_ASAP7_75t_L g7654 ( 
.A(n_7578),
.B(n_888),
.Y(n_7654)
);

INVx1_ASAP7_75t_L g7655 ( 
.A(n_7578),
.Y(n_7655)
);

NAND2xp5_ASAP7_75t_SL g7656 ( 
.A(n_7578),
.B(n_889),
.Y(n_7656)
);

XOR2x2_ASAP7_75t_L g7657 ( 
.A(n_7612),
.B(n_889),
.Y(n_7657)
);

INVx1_ASAP7_75t_L g7658 ( 
.A(n_7643),
.Y(n_7658)
);

AND2x2_ASAP7_75t_L g7659 ( 
.A(n_7649),
.B(n_7655),
.Y(n_7659)
);

AOI22xp33_ASAP7_75t_L g7660 ( 
.A1(n_7641),
.A2(n_892),
.B1(n_890),
.B2(n_891),
.Y(n_7660)
);

NOR2x1_ASAP7_75t_L g7661 ( 
.A(n_7614),
.B(n_890),
.Y(n_7661)
);

OAI22xp33_ASAP7_75t_L g7662 ( 
.A1(n_7648),
.A2(n_893),
.B1(n_890),
.B2(n_891),
.Y(n_7662)
);

BUFx6f_ASAP7_75t_L g7663 ( 
.A(n_7616),
.Y(n_7663)
);

NAND2xp5_ASAP7_75t_L g7664 ( 
.A(n_7626),
.B(n_891),
.Y(n_7664)
);

AND2x2_ASAP7_75t_L g7665 ( 
.A(n_7623),
.B(n_893),
.Y(n_7665)
);

INVx1_ASAP7_75t_L g7666 ( 
.A(n_7626),
.Y(n_7666)
);

NAND3xp33_ASAP7_75t_L g7667 ( 
.A(n_7651),
.B(n_7650),
.C(n_7642),
.Y(n_7667)
);

AOI22xp5_ASAP7_75t_L g7668 ( 
.A1(n_7619),
.A2(n_896),
.B1(n_894),
.B2(n_895),
.Y(n_7668)
);

NOR2x1p5_ASAP7_75t_L g7669 ( 
.A(n_7644),
.B(n_894),
.Y(n_7669)
);

OAI21xp5_ASAP7_75t_L g7670 ( 
.A1(n_7631),
.A2(n_895),
.B(n_896),
.Y(n_7670)
);

OAI22xp33_ASAP7_75t_SL g7671 ( 
.A1(n_7654),
.A2(n_1045),
.B1(n_897),
.B2(n_895),
.Y(n_7671)
);

OAI22xp5_ASAP7_75t_L g7672 ( 
.A1(n_7632),
.A2(n_898),
.B1(n_896),
.B2(n_897),
.Y(n_7672)
);

NOR3xp33_ASAP7_75t_L g7673 ( 
.A(n_7613),
.B(n_897),
.C(n_898),
.Y(n_7673)
);

OAI221xp5_ASAP7_75t_L g7674 ( 
.A1(n_7645),
.A2(n_7653),
.B1(n_7638),
.B2(n_7622),
.C(n_7624),
.Y(n_7674)
);

OAI221xp5_ASAP7_75t_L g7675 ( 
.A1(n_7634),
.A2(n_900),
.B1(n_898),
.B2(n_899),
.C(n_901),
.Y(n_7675)
);

O2A1O1Ixp33_ASAP7_75t_L g7676 ( 
.A1(n_7617),
.A2(n_901),
.B(n_899),
.C(n_900),
.Y(n_7676)
);

NOR3xp33_ASAP7_75t_L g7677 ( 
.A(n_7621),
.B(n_899),
.C(n_900),
.Y(n_7677)
);

INVx1_ASAP7_75t_L g7678 ( 
.A(n_7637),
.Y(n_7678)
);

NAND3xp33_ASAP7_75t_L g7679 ( 
.A(n_7615),
.B(n_901),
.C(n_902),
.Y(n_7679)
);

OAI221xp5_ASAP7_75t_L g7680 ( 
.A1(n_7640),
.A2(n_904),
.B1(n_902),
.B2(n_903),
.C(n_905),
.Y(n_7680)
);

INVx1_ASAP7_75t_L g7681 ( 
.A(n_7618),
.Y(n_7681)
);

INVx1_ASAP7_75t_SL g7682 ( 
.A(n_7625),
.Y(n_7682)
);

AND2x2_ASAP7_75t_SL g7683 ( 
.A(n_7646),
.B(n_1045),
.Y(n_7683)
);

NAND2xp5_ASAP7_75t_L g7684 ( 
.A(n_7647),
.B(n_903),
.Y(n_7684)
);

XNOR2x1_ASAP7_75t_L g7685 ( 
.A(n_7636),
.B(n_903),
.Y(n_7685)
);

AOI21xp5_ASAP7_75t_L g7686 ( 
.A1(n_7652),
.A2(n_904),
.B(n_905),
.Y(n_7686)
);

AOI22xp5_ASAP7_75t_L g7687 ( 
.A1(n_7629),
.A2(n_908),
.B1(n_906),
.B2(n_907),
.Y(n_7687)
);

INVx1_ASAP7_75t_L g7688 ( 
.A(n_7635),
.Y(n_7688)
);

INVx1_ASAP7_75t_L g7689 ( 
.A(n_7627),
.Y(n_7689)
);

NAND2xp5_ASAP7_75t_SL g7690 ( 
.A(n_7620),
.B(n_907),
.Y(n_7690)
);

XNOR2xp5_ASAP7_75t_L g7691 ( 
.A(n_7639),
.B(n_907),
.Y(n_7691)
);

INVx1_ASAP7_75t_L g7692 ( 
.A(n_7656),
.Y(n_7692)
);

INVx1_ASAP7_75t_L g7693 ( 
.A(n_7628),
.Y(n_7693)
);

XNOR2xp5_ASAP7_75t_L g7694 ( 
.A(n_7630),
.B(n_908),
.Y(n_7694)
);

OAI21xp5_ASAP7_75t_L g7695 ( 
.A1(n_7633),
.A2(n_908),
.B(n_909),
.Y(n_7695)
);

OAI22xp5_ASAP7_75t_L g7696 ( 
.A1(n_7648),
.A2(n_911),
.B1(n_909),
.B2(n_910),
.Y(n_7696)
);

INVx1_ASAP7_75t_L g7697 ( 
.A(n_7643),
.Y(n_7697)
);

NAND4xp25_ASAP7_75t_L g7698 ( 
.A(n_7681),
.B(n_912),
.C(n_910),
.D(n_911),
.Y(n_7698)
);

NOR4xp25_ASAP7_75t_L g7699 ( 
.A(n_7658),
.B(n_913),
.C(n_910),
.D(n_911),
.Y(n_7699)
);

NOR2x1_ASAP7_75t_L g7700 ( 
.A(n_7697),
.B(n_913),
.Y(n_7700)
);

INVx1_ASAP7_75t_L g7701 ( 
.A(n_7659),
.Y(n_7701)
);

INVx2_ASAP7_75t_L g7702 ( 
.A(n_7685),
.Y(n_7702)
);

AOI22xp5_ASAP7_75t_L g7703 ( 
.A1(n_7682),
.A2(n_916),
.B1(n_914),
.B2(n_915),
.Y(n_7703)
);

NOR2x1_ASAP7_75t_L g7704 ( 
.A(n_7661),
.B(n_914),
.Y(n_7704)
);

NAND4xp25_ASAP7_75t_SL g7705 ( 
.A(n_7677),
.B(n_917),
.C(n_915),
.D(n_916),
.Y(n_7705)
);

INVx1_ASAP7_75t_L g7706 ( 
.A(n_7694),
.Y(n_7706)
);

INVx1_ASAP7_75t_L g7707 ( 
.A(n_7691),
.Y(n_7707)
);

NOR4xp25_ASAP7_75t_L g7708 ( 
.A(n_7690),
.B(n_7676),
.C(n_7680),
.D(n_7675),
.Y(n_7708)
);

AO22x2_ASAP7_75t_L g7709 ( 
.A1(n_7666),
.A2(n_1042),
.B1(n_918),
.B2(n_915),
.Y(n_7709)
);

INVx1_ASAP7_75t_L g7710 ( 
.A(n_7672),
.Y(n_7710)
);

AOI22xp33_ASAP7_75t_SL g7711 ( 
.A1(n_7665),
.A2(n_919),
.B1(n_917),
.B2(n_918),
.Y(n_7711)
);

NAND2xp5_ASAP7_75t_L g7712 ( 
.A(n_7660),
.B(n_917),
.Y(n_7712)
);

OAI22xp5_ASAP7_75t_SL g7713 ( 
.A1(n_7674),
.A2(n_920),
.B1(n_918),
.B2(n_919),
.Y(n_7713)
);

OAI22xp5_ASAP7_75t_SL g7714 ( 
.A1(n_7683),
.A2(n_921),
.B1(n_919),
.B2(n_920),
.Y(n_7714)
);

INVx1_ASAP7_75t_L g7715 ( 
.A(n_7668),
.Y(n_7715)
);

AOI22xp5_ASAP7_75t_L g7716 ( 
.A1(n_7657),
.A2(n_922),
.B1(n_920),
.B2(n_921),
.Y(n_7716)
);

INVx1_ASAP7_75t_L g7717 ( 
.A(n_7687),
.Y(n_7717)
);

NOR2xp33_ASAP7_75t_SL g7718 ( 
.A(n_7667),
.B(n_922),
.Y(n_7718)
);

AOI22xp5_ASAP7_75t_L g7719 ( 
.A1(n_7663),
.A2(n_925),
.B1(n_923),
.B2(n_924),
.Y(n_7719)
);

AOI22xp5_ASAP7_75t_L g7720 ( 
.A1(n_7663),
.A2(n_925),
.B1(n_923),
.B2(n_924),
.Y(n_7720)
);

INVxp67_ASAP7_75t_L g7721 ( 
.A(n_7664),
.Y(n_7721)
);

INVx1_ASAP7_75t_L g7722 ( 
.A(n_7679),
.Y(n_7722)
);

NOR4xp25_ASAP7_75t_L g7723 ( 
.A(n_7689),
.B(n_927),
.C(n_924),
.D(n_926),
.Y(n_7723)
);

OAI22xp5_ASAP7_75t_L g7724 ( 
.A1(n_7684),
.A2(n_928),
.B1(n_926),
.B2(n_927),
.Y(n_7724)
);

NAND2xp5_ASAP7_75t_SL g7725 ( 
.A(n_7671),
.B(n_926),
.Y(n_7725)
);

AOI22xp5_ASAP7_75t_L g7726 ( 
.A1(n_7663),
.A2(n_930),
.B1(n_928),
.B2(n_929),
.Y(n_7726)
);

INVx1_ASAP7_75t_L g7727 ( 
.A(n_7709),
.Y(n_7727)
);

OR2x2_ASAP7_75t_L g7728 ( 
.A(n_7701),
.B(n_7698),
.Y(n_7728)
);

HB1xp67_ASAP7_75t_L g7729 ( 
.A(n_7700),
.Y(n_7729)
);

OAI21xp33_ASAP7_75t_L g7730 ( 
.A1(n_7718),
.A2(n_7678),
.B(n_7693),
.Y(n_7730)
);

AND2x2_ASAP7_75t_L g7731 ( 
.A(n_7716),
.B(n_7669),
.Y(n_7731)
);

INVxp67_ASAP7_75t_SL g7732 ( 
.A(n_7713),
.Y(n_7732)
);

INVx1_ASAP7_75t_L g7733 ( 
.A(n_7709),
.Y(n_7733)
);

CKINVDCx16_ASAP7_75t_R g7734 ( 
.A(n_7714),
.Y(n_7734)
);

INVx1_ASAP7_75t_SL g7735 ( 
.A(n_7712),
.Y(n_7735)
);

INVx1_ASAP7_75t_SL g7736 ( 
.A(n_7704),
.Y(n_7736)
);

AND2x2_ASAP7_75t_L g7737 ( 
.A(n_7707),
.B(n_7688),
.Y(n_7737)
);

INVx1_ASAP7_75t_L g7738 ( 
.A(n_7703),
.Y(n_7738)
);

AND2x2_ASAP7_75t_L g7739 ( 
.A(n_7710),
.B(n_7692),
.Y(n_7739)
);

INVx1_ASAP7_75t_L g7740 ( 
.A(n_7719),
.Y(n_7740)
);

AOI22xp33_ASAP7_75t_L g7741 ( 
.A1(n_7717),
.A2(n_7673),
.B1(n_7670),
.B2(n_7686),
.Y(n_7741)
);

INVx1_ASAP7_75t_SL g7742 ( 
.A(n_7725),
.Y(n_7742)
);

NAND2xp5_ASAP7_75t_L g7743 ( 
.A(n_7711),
.B(n_7662),
.Y(n_7743)
);

INVx1_ASAP7_75t_L g7744 ( 
.A(n_7720),
.Y(n_7744)
);

AND3x1_ASAP7_75t_L g7745 ( 
.A(n_7708),
.B(n_7695),
.C(n_7696),
.Y(n_7745)
);

NAND2xp5_ASAP7_75t_L g7746 ( 
.A(n_7723),
.B(n_7699),
.Y(n_7746)
);

INVx1_ASAP7_75t_L g7747 ( 
.A(n_7726),
.Y(n_7747)
);

NAND3xp33_ASAP7_75t_SL g7748 ( 
.A(n_7739),
.B(n_7706),
.C(n_7702),
.Y(n_7748)
);

AND4x1_ASAP7_75t_L g7749 ( 
.A(n_7741),
.B(n_7715),
.C(n_7722),
.D(n_7721),
.Y(n_7749)
);

NOR3xp33_ASAP7_75t_L g7750 ( 
.A(n_7728),
.B(n_7705),
.C(n_7724),
.Y(n_7750)
);

AND2x4_ASAP7_75t_L g7751 ( 
.A(n_7737),
.B(n_929),
.Y(n_7751)
);

INVx1_ASAP7_75t_L g7752 ( 
.A(n_7727),
.Y(n_7752)
);

OAI211xp5_ASAP7_75t_SL g7753 ( 
.A1(n_7746),
.A2(n_7730),
.B(n_7732),
.C(n_7733),
.Y(n_7753)
);

NOR3xp33_ASAP7_75t_L g7754 ( 
.A(n_7734),
.B(n_929),
.C(n_930),
.Y(n_7754)
);

NOR3xp33_ASAP7_75t_L g7755 ( 
.A(n_7735),
.B(n_930),
.C(n_931),
.Y(n_7755)
);

NAND3xp33_ASAP7_75t_SL g7756 ( 
.A(n_7742),
.B(n_931),
.C(n_932),
.Y(n_7756)
);

NOR3xp33_ASAP7_75t_L g7757 ( 
.A(n_7738),
.B(n_931),
.C(n_933),
.Y(n_7757)
);

NOR3xp33_ASAP7_75t_SL g7758 ( 
.A(n_7743),
.B(n_933),
.C(n_934),
.Y(n_7758)
);

INVx1_ASAP7_75t_L g7759 ( 
.A(n_7745),
.Y(n_7759)
);

NAND4xp25_ASAP7_75t_L g7760 ( 
.A(n_7731),
.B(n_935),
.C(n_933),
.D(n_934),
.Y(n_7760)
);

NOR3xp33_ASAP7_75t_L g7761 ( 
.A(n_7729),
.B(n_934),
.C(n_936),
.Y(n_7761)
);

NOR2x1_ASAP7_75t_L g7762 ( 
.A(n_7753),
.B(n_7736),
.Y(n_7762)
);

NAND2xp5_ASAP7_75t_L g7763 ( 
.A(n_7749),
.B(n_7740),
.Y(n_7763)
);

INVx1_ASAP7_75t_L g7764 ( 
.A(n_7759),
.Y(n_7764)
);

NAND4xp25_ASAP7_75t_L g7765 ( 
.A(n_7750),
.B(n_7744),
.C(n_7747),
.D(n_938),
.Y(n_7765)
);

XNOR2x1_ASAP7_75t_L g7766 ( 
.A(n_7762),
.B(n_7752),
.Y(n_7766)
);

OAI22xp5_ASAP7_75t_L g7767 ( 
.A1(n_7766),
.A2(n_7763),
.B1(n_7764),
.B2(n_7748),
.Y(n_7767)
);

OA22x2_ASAP7_75t_L g7768 ( 
.A1(n_7766),
.A2(n_7765),
.B1(n_7751),
.B2(n_7758),
.Y(n_7768)
);

XNOR2x1_ASAP7_75t_L g7769 ( 
.A(n_7767),
.B(n_7768),
.Y(n_7769)
);

NAND2xp5_ASAP7_75t_L g7770 ( 
.A(n_7767),
.B(n_7754),
.Y(n_7770)
);

HB1xp67_ASAP7_75t_L g7771 ( 
.A(n_7770),
.Y(n_7771)
);

INVx1_ASAP7_75t_L g7772 ( 
.A(n_7769),
.Y(n_7772)
);

INVx1_ASAP7_75t_L g7773 ( 
.A(n_7771),
.Y(n_7773)
);

INVx1_ASAP7_75t_L g7774 ( 
.A(n_7773),
.Y(n_7774)
);

XOR2xp5_ASAP7_75t_L g7775 ( 
.A(n_7774),
.B(n_7772),
.Y(n_7775)
);

AOI21xp5_ASAP7_75t_L g7776 ( 
.A1(n_7775),
.A2(n_7751),
.B(n_7757),
.Y(n_7776)
);

OAI22xp5_ASAP7_75t_L g7777 ( 
.A1(n_7776),
.A2(n_7761),
.B1(n_7755),
.B2(n_7756),
.Y(n_7777)
);

OAI222xp33_ASAP7_75t_L g7778 ( 
.A1(n_7777),
.A2(n_7760),
.B1(n_937),
.B2(n_938),
.C1(n_939),
.C2(n_940),
.Y(n_7778)
);

NAND2xp5_ASAP7_75t_L g7779 ( 
.A(n_7778),
.B(n_936),
.Y(n_7779)
);

AOI22xp33_ASAP7_75t_L g7780 ( 
.A1(n_7779),
.A2(n_938),
.B1(n_936),
.B2(n_937),
.Y(n_7780)
);

OAI221xp5_ASAP7_75t_R g7781 ( 
.A1(n_7780),
.A2(n_937),
.B1(n_939),
.B2(n_940),
.C(n_941),
.Y(n_7781)
);

AOI22xp33_ASAP7_75t_L g7782 ( 
.A1(n_7781),
.A2(n_941),
.B1(n_939),
.B2(n_940),
.Y(n_7782)
);

AOI211xp5_ASAP7_75t_L g7783 ( 
.A1(n_7782),
.A2(n_944),
.B(n_942),
.C(n_943),
.Y(n_7783)
);


endmodule