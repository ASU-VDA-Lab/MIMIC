module fake_jpeg_31330_n_177 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_177);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_14),
.B(n_6),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_48),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx8_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_20),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_11),
.A2(n_9),
.B(n_8),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_62),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_77),
.A2(n_76),
.B1(n_71),
.B2(n_62),
.Y(n_94)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_81),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_1),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_85),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_58),
.B(n_3),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_3),
.Y(n_98)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_73),
.C(n_54),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_4),
.Y(n_119)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_99),
.B1(n_65),
.B2(n_59),
.Y(n_104)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_4),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_82),
.A2(n_64),
.B1(n_71),
.B2(n_74),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_69),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_100),
.B(n_51),
.Y(n_111)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_90),
.A2(n_65),
.B1(n_59),
.B2(n_61),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_109),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_116),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_85),
.B1(n_61),
.B2(n_74),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_105),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_106),
.B(n_108),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_70),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_100),
.A2(n_51),
.B1(n_75),
.B2(n_53),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_76),
.B(n_60),
.C(n_67),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_5),
.B(n_6),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_115),
.Y(n_140)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_118),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_66),
.B1(n_56),
.B2(n_55),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_68),
.B1(n_21),
.B2(n_23),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_68),
.B1(n_18),
.B2(n_24),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_120),
.Y(n_128)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_14),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_89),
.A2(n_16),
.B1(n_47),
.B2(n_41),
.Y(n_120)
);

AND2x6_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_50),
.Y(n_121)
);

AOI32xp33_ASAP7_75t_L g125 ( 
.A1(n_121),
.A2(n_40),
.A3(n_38),
.B1(n_37),
.B2(n_33),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_7),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_130),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_129),
.A2(n_134),
.B1(n_142),
.B2(n_131),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_30),
.C(n_28),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_142),
.C(n_144),
.Y(n_158)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_135),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_9),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_138),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_11),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_12),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_139),
.B(n_143),
.Y(n_151)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_12),
.C(n_13),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_13),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_145),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_15),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_136),
.A2(n_15),
.B1(n_118),
.B2(n_140),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_148),
.Y(n_166)
);

NOR4xp25_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_149),
.C(n_158),
.D(n_155),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_SL g155 ( 
.A1(n_129),
.A2(n_134),
.B(n_126),
.C(n_128),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_156),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_145),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_146),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_124),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_159),
.B(n_124),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_126),
.C(n_128),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_147),
.C(n_151),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_161),
.B(n_164),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_163),
.Y(n_169)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_165),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_168),
.A2(n_165),
.B(n_166),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_170),
.B(n_171),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_169),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_167),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_155),
.B(n_154),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_175),
.A2(n_155),
.B(n_150),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_153),
.Y(n_177)
);


endmodule