module fake_jpeg_16433_n_30 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_30);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_30;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_29;
wire n_12;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_4),
.Y(n_8)
);

AOI22xp33_ASAP7_75t_L g9 ( 
.A1(n_4),
.A2(n_5),
.B1(n_1),
.B2(n_0),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_2),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_10),
.A2(n_2),
.B1(n_6),
.B2(n_11),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_19),
.C(n_20),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_14),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_8),
.A2(n_9),
.B(n_13),
.Y(n_21)
);

MAJx2_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_22),
.C(n_23),
.Y(n_26)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_13),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_26),
.B(n_19),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_28),
.Y(n_29)
);

NAND2x1_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_18),
.Y(n_28)
);

AOI322xp5_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_28),
.A3(n_25),
.B1(n_18),
.B2(n_23),
.C1(n_12),
.C2(n_15),
.Y(n_30)
);


endmodule