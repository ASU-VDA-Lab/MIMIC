module fake_netlist_5_2234_n_80 (n_16, n_0, n_12, n_9, n_18, n_22, n_1, n_8, n_10, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_20, n_5, n_14, n_2, n_23, n_13, n_3, n_6, n_80);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_22;
input n_1;
input n_8;
input n_10;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_20;
input n_5;
input n_14;
input n_2;
input n_23;
input n_13;
input n_3;
input n_6;

output n_80;

wire n_24;
wire n_61;
wire n_75;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_37;
wire n_31;
wire n_66;
wire n_60;
wire n_43;
wire n_58;
wire n_69;
wire n_42;
wire n_45;
wire n_46;
wire n_38;
wire n_35;
wire n_73;
wire n_30;
wire n_33;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_71;
wire n_59;
wire n_26;
wire n_55;
wire n_49;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_27;
wire n_64;
wire n_77;
wire n_28;
wire n_70;
wire n_68;
wire n_72;
wire n_32;
wire n_41;
wire n_56;
wire n_51;
wire n_63;
wire n_48;
wire n_50;
wire n_52;

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_11),
.B(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_19),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_12),
.B(n_10),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_4),
.B(n_9),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

OA21x2_ASAP7_75t_L g35 ( 
.A1(n_1),
.A2(n_16),
.B(n_21),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVxp67_ASAP7_75t_SL g39 ( 
.A(n_27),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_0),
.Y(n_42)
);

O2A1O1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_6),
.B(n_8),
.C(n_13),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_38),
.B(n_14),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_18),
.Y(n_45)
);

NOR2xp67_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_22),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_35),
.B1(n_37),
.B2(n_26),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_36),
.B(n_25),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_25),
.B(n_37),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_30),
.B1(n_33),
.B2(n_29),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_35),
.B1(n_28),
.B2(n_24),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_41),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

OAI21x1_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_32),
.B(n_30),
.Y(n_58)
);

NAND2x1_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_30),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

AND2x4_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_39),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_50),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_53),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_52),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_69),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_60),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_66),
.B(n_69),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_SL g73 ( 
.A1(n_71),
.A2(n_45),
.B(n_44),
.C(n_42),
.Y(n_73)
);

NOR3x1_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_40),
.C(n_60),
.Y(n_74)
);

NAND3x1_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_67),
.C(n_61),
.Y(n_75)
);

NOR3xp33_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_73),
.C(n_43),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_75),
.A2(n_30),
.B1(n_76),
.B2(n_57),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_46),
.B1(n_47),
.B2(n_57),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_77),
.B1(n_49),
.B2(n_63),
.Y(n_80)
);


endmodule