module real_aes_9113_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_119;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_212;
wire n_210;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g565 ( .A1(n_0), .A2(n_203), .B(n_566), .C(n_569), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_1), .B(n_554), .Y(n_570) );
INVx1_ASAP7_75t_L g114 ( .A(n_2), .Y(n_114) );
AOI22xp5_ASAP7_75t_L g131 ( .A1(n_3), .A2(n_132), .B1(n_133), .B2(n_136), .Y(n_131) );
INVx1_ASAP7_75t_L g136 ( .A(n_3), .Y(n_136) );
INVx1_ASAP7_75t_L g221 ( .A(n_4), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_5), .B(n_192), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_6), .A2(n_469), .B(n_548), .Y(n_547) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_7), .A2(n_168), .B(n_516), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_8), .A2(n_38), .B1(n_148), .B2(n_157), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_9), .B(n_168), .Y(n_232) );
AND2x6_ASAP7_75t_L g166 ( .A(n_10), .B(n_167), .Y(n_166) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_11), .A2(n_166), .B(n_472), .C(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g111 ( .A(n_12), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_12), .B(n_39), .Y(n_129) );
INVx1_ASAP7_75t_L g164 ( .A(n_13), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_14), .B(n_155), .Y(n_175) );
INVx1_ASAP7_75t_L g213 ( .A(n_15), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_16), .B(n_192), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_17), .B(n_169), .Y(n_237) );
AO32x2_ASAP7_75t_L g200 ( .A1(n_18), .A2(n_165), .A3(n_168), .B1(n_201), .B2(n_205), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_19), .B(n_157), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_20), .B(n_169), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_21), .A2(n_55), .B1(n_148), .B2(n_157), .Y(n_204) );
AOI22xp33_ASAP7_75t_SL g154 ( .A1(n_22), .A2(n_83), .B1(n_155), .B2(n_157), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_23), .B(n_157), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_L g471 ( .A1(n_24), .A2(n_165), .B(n_472), .C(n_474), .Y(n_471) );
AOI222xp33_ASAP7_75t_L g450 ( .A1(n_25), .A2(n_451), .B1(n_755), .B2(n_756), .C1(n_765), .C2(n_769), .Y(n_450) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_26), .A2(n_165), .B(n_472), .C(n_519), .Y(n_518) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_27), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_28), .B(n_160), .Y(n_257) );
OAI22xp5_ASAP7_75t_SL g759 ( .A1(n_29), .A2(n_760), .B1(n_763), .B2(n_764), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_29), .Y(n_764) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_30), .A2(n_469), .B(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_31), .B(n_160), .Y(n_198) );
INVx2_ASAP7_75t_L g150 ( .A(n_32), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_33), .A2(n_493), .B(n_502), .C(n_504), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_34), .B(n_157), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_35), .B(n_160), .Y(n_182) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_36), .A2(n_76), .B1(n_761), .B2(n_762), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_36), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_37), .B(n_177), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_39), .B(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_40), .B(n_468), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_41), .A2(n_757), .B1(n_758), .B2(n_759), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_41), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_42), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_43), .B(n_192), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_44), .B(n_469), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_45), .A2(n_493), .B(n_502), .C(n_539), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_46), .A2(n_81), .B1(n_443), .B2(n_444), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_46), .Y(n_443) );
OAI22xp5_ASAP7_75t_SL g453 ( .A1(n_46), .A2(n_443), .B1(n_454), .B2(n_455), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_47), .B(n_157), .Y(n_227) );
INVx1_ASAP7_75t_L g567 ( .A(n_48), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g147 ( .A1(n_49), .A2(n_91), .B1(n_148), .B2(n_151), .Y(n_147) );
INVx1_ASAP7_75t_L g540 ( .A(n_50), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_51), .B(n_157), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_52), .B(n_157), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_53), .B(n_469), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_54), .B(n_219), .Y(n_231) );
AOI22xp33_ASAP7_75t_SL g241 ( .A1(n_56), .A2(n_60), .B1(n_155), .B2(n_157), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_57), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_58), .B(n_157), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_59), .B(n_157), .Y(n_256) );
INVx1_ASAP7_75t_L g167 ( .A(n_61), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_62), .B(n_469), .Y(n_495) );
OAI22xp5_ASAP7_75t_SL g133 ( .A1(n_63), .A2(n_100), .B1(n_134), .B2(n_135), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_63), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_63), .B(n_554), .Y(n_553) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_64), .A2(n_216), .B(n_219), .C(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_65), .B(n_157), .Y(n_222) );
INVx1_ASAP7_75t_L g163 ( .A(n_66), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_67), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_68), .B(n_192), .Y(n_506) );
AO32x2_ASAP7_75t_L g145 ( .A1(n_69), .A2(n_146), .A3(n_159), .B1(n_165), .B2(n_168), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_70), .B(n_158), .Y(n_530) );
INVx1_ASAP7_75t_L g255 ( .A(n_71), .Y(n_255) );
INVx1_ASAP7_75t_L g190 ( .A(n_72), .Y(n_190) );
CKINVDCx16_ASAP7_75t_R g564 ( .A(n_73), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_74), .B(n_476), .Y(n_475) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_75), .A2(n_472), .B(n_489), .C(n_493), .Y(n_488) );
INVx1_ASAP7_75t_L g762 ( .A(n_76), .Y(n_762) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_77), .B(n_155), .Y(n_191) );
CKINVDCx16_ASAP7_75t_R g549 ( .A(n_78), .Y(n_549) );
INVx1_ASAP7_75t_L g118 ( .A(n_79), .Y(n_118) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_80), .A2(n_106), .B1(n_119), .B2(n_774), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_81), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_82), .B(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_84), .B(n_148), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_85), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_86), .B(n_155), .Y(n_195) );
INVx2_ASAP7_75t_L g161 ( .A(n_87), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_88), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_89), .B(n_152), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_90), .B(n_155), .Y(n_228) );
INVx2_ASAP7_75t_L g115 ( .A(n_92), .Y(n_115) );
OR2x2_ASAP7_75t_L g126 ( .A(n_92), .B(n_127), .Y(n_126) );
OR2x2_ASAP7_75t_L g458 ( .A(n_92), .B(n_128), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_93), .A2(n_104), .B1(n_155), .B2(n_156), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_94), .B(n_469), .Y(n_500) );
INVx1_ASAP7_75t_L g505 ( .A(n_95), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_96), .B(n_447), .Y(n_446) );
INVxp67_ASAP7_75t_L g552 ( .A(n_97), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_98), .B(n_155), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_99), .B(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g134 ( .A(n_100), .Y(n_134) );
INVx1_ASAP7_75t_L g490 ( .A(n_101), .Y(n_490) );
INVx1_ASAP7_75t_L g526 ( .A(n_102), .Y(n_526) );
AND2x2_ASAP7_75t_L g542 ( .A(n_103), .B(n_160), .Y(n_542) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g776 ( .A(n_108), .Y(n_776) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_112), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
CKINVDCx14_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
NAND3xp33_ASAP7_75t_SL g113 ( .A(n_114), .B(n_115), .C(n_116), .Y(n_113) );
AND2x2_ASAP7_75t_L g128 ( .A(n_114), .B(n_129), .Y(n_128) );
OR2x2_ASAP7_75t_L g754 ( .A(n_115), .B(n_128), .Y(n_754) );
NOR2x2_ASAP7_75t_L g771 ( .A(n_115), .B(n_127), .Y(n_771) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
OA21x2_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_124), .B(n_449), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g773 ( .A(n_122), .Y(n_773) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI21xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_130), .B(n_446), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_126), .Y(n_448) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AOI22xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_137), .B1(n_138), .B2(n_445), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_131), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
XOR2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_442), .Y(n_138) );
INVx2_ASAP7_75t_L g454 ( .A(n_139), .Y(n_454) );
AND3x1_ASAP7_75t_L g139 ( .A(n_140), .B(n_362), .C(n_410), .Y(n_139) );
NOR4xp25_ASAP7_75t_L g140 ( .A(n_141), .B(n_290), .C(n_335), .D(n_349), .Y(n_140) );
OAI311xp33_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_206), .A3(n_233), .B1(n_243), .C1(n_258), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_170), .Y(n_142) );
OAI21xp33_ASAP7_75t_L g243 ( .A1(n_143), .A2(n_244), .B(n_246), .Y(n_243) );
AND2x2_ASAP7_75t_L g351 ( .A(n_143), .B(n_278), .Y(n_351) );
AND2x2_ASAP7_75t_L g408 ( .A(n_143), .B(n_294), .Y(n_408) );
BUFx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g301 ( .A(n_144), .B(n_199), .Y(n_301) );
AND2x2_ASAP7_75t_L g358 ( .A(n_144), .B(n_306), .Y(n_358) );
INVx1_ASAP7_75t_L g399 ( .A(n_144), .Y(n_399) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
BUFx6f_ASAP7_75t_L g267 ( .A(n_145), .Y(n_267) );
AND2x2_ASAP7_75t_L g308 ( .A(n_145), .B(n_199), .Y(n_308) );
AND2x2_ASAP7_75t_L g312 ( .A(n_145), .B(n_200), .Y(n_312) );
INVx1_ASAP7_75t_L g324 ( .A(n_145), .Y(n_324) );
OAI22xp5_ASAP7_75t_SL g146 ( .A1(n_147), .A2(n_152), .B1(n_154), .B2(n_158), .Y(n_146) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx3_ASAP7_75t_L g151 ( .A(n_149), .Y(n_151) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_149), .Y(n_157) );
AND2x6_ASAP7_75t_L g472 ( .A(n_149), .B(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g156 ( .A(n_150), .Y(n_156) );
INVx1_ASAP7_75t_L g220 ( .A(n_150), .Y(n_220) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_151), .Y(n_507) );
INVx2_ASAP7_75t_L g569 ( .A(n_151), .Y(n_569) );
INVx2_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
OAI22xp5_ASAP7_75t_L g201 ( .A1(n_152), .A2(n_202), .B1(n_203), .B2(n_204), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g239 ( .A1(n_152), .A2(n_203), .B1(n_240), .B2(n_241), .Y(n_239) );
INVx4_ASAP7_75t_L g568 ( .A(n_152), .Y(n_568) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx3_ASAP7_75t_L g158 ( .A(n_153), .Y(n_158) );
INVx1_ASAP7_75t_L g177 ( .A(n_153), .Y(n_177) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_153), .Y(n_197) );
AND2x2_ASAP7_75t_L g470 ( .A(n_153), .B(n_220), .Y(n_470) );
INVx1_ASAP7_75t_L g473 ( .A(n_153), .Y(n_473) );
INVx2_ASAP7_75t_L g214 ( .A(n_155), .Y(n_214) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx3_ASAP7_75t_L g189 ( .A(n_157), .Y(n_189) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_157), .Y(n_492) );
INVx5_ASAP7_75t_L g192 ( .A(n_158), .Y(n_192) );
INVx1_ASAP7_75t_L g479 ( .A(n_159), .Y(n_479) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
OA21x2_ASAP7_75t_L g171 ( .A1(n_160), .A2(n_172), .B(n_182), .Y(n_171) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_160), .A2(n_187), .B(n_198), .Y(n_186) );
INVx1_ASAP7_75t_L g482 ( .A(n_160), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_160), .A2(n_500), .B(n_501), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_160), .A2(n_537), .B(n_538), .Y(n_536) );
AND2x2_ASAP7_75t_SL g160 ( .A(n_161), .B(n_162), .Y(n_160) );
AND2x2_ASAP7_75t_L g169 ( .A(n_161), .B(n_162), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
NAND3xp33_ASAP7_75t_L g238 ( .A(n_165), .B(n_239), .C(n_242), .Y(n_238) );
OAI21xp5_ASAP7_75t_L g250 ( .A1(n_165), .A2(n_251), .B(n_254), .Y(n_250) );
BUFx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
OAI21xp5_ASAP7_75t_L g172 ( .A1(n_166), .A2(n_173), .B(n_178), .Y(n_172) );
OAI21xp5_ASAP7_75t_L g187 ( .A1(n_166), .A2(n_188), .B(n_193), .Y(n_187) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_166), .A2(n_212), .B(n_217), .Y(n_211) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_166), .A2(n_226), .B(n_229), .Y(n_225) );
AND2x4_ASAP7_75t_L g469 ( .A(n_166), .B(n_470), .Y(n_469) );
INVx4_ASAP7_75t_SL g494 ( .A(n_166), .Y(n_494) );
NAND2x1p5_ASAP7_75t_L g527 ( .A(n_166), .B(n_470), .Y(n_527) );
OA21x2_ASAP7_75t_L g224 ( .A1(n_168), .A2(n_225), .B(n_232), .Y(n_224) );
INVx4_ASAP7_75t_L g242 ( .A(n_168), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_168), .A2(n_517), .B(n_518), .Y(n_516) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_168), .Y(n_546) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g205 ( .A(n_169), .Y(n_205) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_183), .Y(n_170) );
AND2x2_ASAP7_75t_L g245 ( .A(n_171), .B(n_199), .Y(n_245) );
INVx2_ASAP7_75t_L g279 ( .A(n_171), .Y(n_279) );
AND2x2_ASAP7_75t_L g294 ( .A(n_171), .B(n_200), .Y(n_294) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_171), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_171), .B(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g314 ( .A(n_171), .B(n_277), .Y(n_314) );
INVx1_ASAP7_75t_L g326 ( .A(n_171), .Y(n_326) );
INVx1_ASAP7_75t_L g367 ( .A(n_171), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_171), .B(n_267), .Y(n_420) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_176), .Y(n_173) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_181), .Y(n_178) );
O2A1O1Ixp5_ASAP7_75t_L g254 ( .A1(n_181), .A2(n_218), .B(n_255), .C(n_256), .Y(n_254) );
NOR2xp67_ASAP7_75t_L g183 ( .A(n_184), .B(n_199), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g244 ( .A(n_185), .B(n_245), .Y(n_244) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_185), .Y(n_272) );
AND2x2_ASAP7_75t_SL g325 ( .A(n_185), .B(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g329 ( .A(n_185), .B(n_199), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_185), .B(n_324), .Y(n_387) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g277 ( .A(n_186), .Y(n_277) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_186), .Y(n_293) );
OR2x2_ASAP7_75t_L g366 ( .A(n_186), .B(n_367), .Y(n_366) );
O2A1O1Ixp5_ASAP7_75t_SL g188 ( .A1(n_189), .A2(n_190), .B(n_191), .C(n_192), .Y(n_188) );
INVx2_ASAP7_75t_L g203 ( .A(n_192), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_192), .A2(n_227), .B(n_228), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_192), .A2(n_252), .B(n_253), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_192), .B(n_552), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_196), .Y(n_193) );
INVx1_ASAP7_75t_L g216 ( .A(n_196), .Y(n_216) );
INVx4_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx2_ASAP7_75t_L g476 ( .A(n_197), .Y(n_476) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
BUFx2_ASAP7_75t_L g273 ( .A(n_200), .Y(n_273) );
AND2x2_ASAP7_75t_L g278 ( .A(n_200), .B(n_279), .Y(n_278) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_203), .A2(n_218), .B(n_221), .C(n_222), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_203), .A2(n_230), .B(n_231), .Y(n_229) );
INVx2_ASAP7_75t_L g210 ( .A(n_205), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_205), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_206), .B(n_261), .Y(n_424) );
INVx1_ASAP7_75t_SL g206 ( .A(n_207), .Y(n_206) );
OR2x2_ASAP7_75t_L g394 ( .A(n_207), .B(n_235), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_208), .B(n_224), .Y(n_207) );
AND2x2_ASAP7_75t_L g270 ( .A(n_208), .B(n_261), .Y(n_270) );
INVx2_ASAP7_75t_L g282 ( .A(n_208), .Y(n_282) );
AND2x2_ASAP7_75t_L g316 ( .A(n_208), .B(n_264), .Y(n_316) );
AND2x2_ASAP7_75t_L g383 ( .A(n_208), .B(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_209), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g263 ( .A(n_209), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g303 ( .A(n_209), .B(n_224), .Y(n_303) );
AND2x2_ASAP7_75t_L g320 ( .A(n_209), .B(n_321), .Y(n_320) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_223), .Y(n_209) );
OA21x2_ASAP7_75t_L g249 ( .A1(n_210), .A2(n_250), .B(n_257), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_215), .C(n_216), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_214), .A2(n_520), .B(n_521), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_214), .A2(n_530), .B(n_531), .Y(n_529) );
O2A1O1Ixp33_ASAP7_75t_L g489 ( .A1(n_216), .A2(n_490), .B(n_491), .C(n_492), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_218), .A2(n_475), .B(n_477), .Y(n_474) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g246 ( .A(n_224), .B(n_247), .Y(n_246) );
INVx3_ASAP7_75t_L g264 ( .A(n_224), .Y(n_264) );
AND2x2_ASAP7_75t_L g269 ( .A(n_224), .B(n_249), .Y(n_269) );
AND2x2_ASAP7_75t_L g342 ( .A(n_224), .B(n_321), .Y(n_342) );
AND2x2_ASAP7_75t_L g407 ( .A(n_224), .B(n_397), .Y(n_407) );
OAI311xp33_ASAP7_75t_L g290 ( .A1(n_233), .A2(n_291), .A3(n_295), .B1(n_297), .C1(n_317), .Y(n_290) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g302 ( .A(n_234), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g361 ( .A(n_234), .B(n_269), .Y(n_361) );
AND2x2_ASAP7_75t_L g435 ( .A(n_234), .B(n_316), .Y(n_435) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_235), .B(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g370 ( .A(n_235), .Y(n_370) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx3_ASAP7_75t_L g261 ( .A(n_236), .Y(n_261) );
NOR2x1_ASAP7_75t_L g333 ( .A(n_236), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g390 ( .A(n_236), .B(n_264), .Y(n_390) );
AND2x4_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
INVx1_ASAP7_75t_L g287 ( .A(n_237), .Y(n_287) );
AO21x1_ASAP7_75t_L g286 ( .A1(n_239), .A2(n_242), .B(n_287), .Y(n_286) );
AO21x2_ASAP7_75t_L g486 ( .A1(n_242), .A2(n_487), .B(n_496), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_242), .B(n_497), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_242), .B(n_509), .Y(n_508) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_242), .A2(n_525), .B(n_532), .Y(n_524) );
INVx3_ASAP7_75t_L g554 ( .A(n_242), .Y(n_554) );
AND2x2_ASAP7_75t_L g265 ( .A(n_245), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g318 ( .A(n_245), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g398 ( .A(n_245), .B(n_399), .Y(n_398) );
AOI221xp5_ASAP7_75t_L g297 ( .A1(n_246), .A2(n_278), .B1(n_298), .B2(n_302), .C(n_304), .Y(n_297) );
INVx1_ASAP7_75t_L g422 ( .A(n_247), .Y(n_422) );
OR2x2_ASAP7_75t_L g388 ( .A(n_248), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g283 ( .A(n_249), .B(n_264), .Y(n_283) );
OR2x2_ASAP7_75t_L g285 ( .A(n_249), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g310 ( .A(n_249), .Y(n_310) );
INVx2_ASAP7_75t_L g321 ( .A(n_249), .Y(n_321) );
AND2x2_ASAP7_75t_L g348 ( .A(n_249), .B(n_286), .Y(n_348) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_249), .Y(n_377) );
AOI221xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_265), .B1(n_268), .B2(n_271), .C(n_274), .Y(n_258) );
INVx1_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
AND2x2_ASAP7_75t_L g359 ( .A(n_261), .B(n_269), .Y(n_359) );
AND2x2_ASAP7_75t_L g409 ( .A(n_261), .B(n_263), .Y(n_409) );
INVx2_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g296 ( .A(n_263), .B(n_267), .Y(n_296) );
AND2x2_ASAP7_75t_L g375 ( .A(n_263), .B(n_348), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_264), .B(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g334 ( .A(n_264), .Y(n_334) );
OAI21xp33_ASAP7_75t_L g344 ( .A1(n_265), .A2(n_345), .B(n_347), .Y(n_344) );
OR2x2_ASAP7_75t_L g288 ( .A(n_266), .B(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g354 ( .A(n_266), .B(n_314), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_266), .B(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g331 ( .A(n_267), .B(n_300), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_267), .B(n_414), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_268), .B(n_294), .Y(n_404) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
AND2x2_ASAP7_75t_L g327 ( .A(n_269), .B(n_282), .Y(n_327) );
INVx1_ASAP7_75t_L g343 ( .A(n_270), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_280), .B1(n_284), .B2(n_288), .Y(n_274) );
INVx2_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx2_ASAP7_75t_L g306 ( .A(n_277), .Y(n_306) );
INVx1_ASAP7_75t_L g319 ( .A(n_277), .Y(n_319) );
INVx1_ASAP7_75t_L g289 ( .A(n_278), .Y(n_289) );
AND2x2_ASAP7_75t_L g360 ( .A(n_278), .B(n_306), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_278), .B(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
OR2x2_ASAP7_75t_L g284 ( .A(n_281), .B(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_281), .B(n_397), .Y(n_396) );
NOR2xp67_ASAP7_75t_L g428 ( .A(n_281), .B(n_429), .Y(n_428) );
INVx3_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g431 ( .A(n_283), .B(n_383), .Y(n_431) );
INVx1_ASAP7_75t_SL g397 ( .A(n_285), .Y(n_397) );
AND2x2_ASAP7_75t_L g337 ( .A(n_286), .B(n_321), .Y(n_337) );
INVx1_ASAP7_75t_L g384 ( .A(n_286), .Y(n_384) );
OAI222xp33_ASAP7_75t_L g425 ( .A1(n_291), .A2(n_381), .B1(n_426), .B2(n_427), .C1(n_430), .C2(n_432), .Y(n_425) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx1_ASAP7_75t_L g346 ( .A(n_293), .Y(n_346) );
AND2x2_ASAP7_75t_L g357 ( .A(n_294), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_SL g426 ( .A(n_294), .B(n_399), .Y(n_426) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_296), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g401 ( .A(n_298), .Y(n_401) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_SL g339 ( .A(n_301), .Y(n_339) );
AND2x2_ASAP7_75t_L g418 ( .A(n_301), .B(n_379), .Y(n_418) );
AND2x2_ASAP7_75t_L g441 ( .A(n_301), .B(n_325), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_303), .B(n_337), .Y(n_336) );
OAI32xp33_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_307), .A3(n_309), .B1(n_311), .B2(n_315), .Y(n_304) );
BUFx2_ASAP7_75t_L g379 ( .A(n_306), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_307), .B(n_325), .Y(n_406) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g345 ( .A(n_308), .B(n_346), .Y(n_345) );
AND2x4_ASAP7_75t_L g413 ( .A(n_308), .B(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g402 ( .A(n_309), .B(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
AND2x2_ASAP7_75t_L g373 ( .A(n_312), .B(n_346), .Y(n_373) );
INVx2_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
OAI221xp5_ASAP7_75t_SL g335 ( .A1(n_314), .A2(n_336), .B1(n_338), .B2(n_340), .C(n_344), .Y(n_335) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g347 ( .A(n_316), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g353 ( .A(n_316), .B(n_337), .Y(n_353) );
AOI221xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_320), .B1(n_322), .B2(n_327), .C(n_328), .Y(n_317) );
INVx1_ASAP7_75t_L g436 ( .A(n_318), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_319), .B(n_413), .Y(n_412) );
NAND2x1p5_ASAP7_75t_L g332 ( .A(n_320), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_325), .B(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g391 ( .A(n_325), .Y(n_391) );
BUFx3_ASAP7_75t_L g414 ( .A(n_326), .Y(n_414) );
INVx1_ASAP7_75t_SL g355 ( .A(n_327), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_327), .B(n_369), .Y(n_368) );
AOI21xp33_ASAP7_75t_SL g328 ( .A1(n_329), .A2(n_330), .B(n_332), .Y(n_328) );
OAI221xp5_ASAP7_75t_L g433 ( .A1(n_329), .A2(n_430), .B1(n_434), .B2(n_436), .C(n_437), .Y(n_433) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g376 ( .A(n_334), .B(n_337), .Y(n_376) );
INVx1_ASAP7_75t_L g440 ( .A(n_334), .Y(n_440) );
INVx2_ASAP7_75t_L g429 ( .A(n_337), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_337), .B(n_440), .Y(n_439) );
OR2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g382 ( .A(n_342), .B(n_383), .Y(n_382) );
OAI221xp5_ASAP7_75t_SL g349 ( .A1(n_350), .A2(n_352), .B1(n_354), .B2(n_355), .C(n_356), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_359), .B1(n_360), .B2(n_361), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_358), .A2(n_420), .B1(n_421), .B2(n_423), .Y(n_419) );
OAI21xp5_ASAP7_75t_L g437 ( .A1(n_361), .A2(n_438), .B(n_441), .Y(n_437) );
NOR4xp25_ASAP7_75t_SL g362 ( .A(n_363), .B(n_371), .C(n_380), .D(n_400), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_364), .B(n_368), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_374), .B1(n_377), .B2(n_378), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
INVx1_ASAP7_75t_L g416 ( .A(n_376), .Y(n_416) );
OAI221xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_385), .B1(n_388), .B2(n_391), .C(n_392), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g403 ( .A(n_383), .Y(n_403) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OAI21xp5_ASAP7_75t_SL g392 ( .A1(n_393), .A2(n_395), .B(n_398), .Y(n_392) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OAI211xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B(n_404), .C(n_405), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_407), .B1(n_408), .B2(n_409), .Y(n_405) );
CKINVDCx14_ASAP7_75t_R g415 ( .A(n_409), .Y(n_415) );
NOR3xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_425), .C(n_433), .Y(n_410) );
OAI221xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_415), .B1(n_416), .B2(n_417), .C(n_419), .Y(n_411) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
CKINVDCx16_ASAP7_75t_R g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NAND3xp33_ASAP7_75t_L g449 ( .A(n_446), .B(n_450), .C(n_772), .Y(n_449) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OAI22xp5_ASAP7_75t_SL g451 ( .A1(n_452), .A2(n_456), .B1(n_459), .B2(n_752), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OAI22xp5_ASAP7_75t_SL g765 ( .A1(n_453), .A2(n_766), .B1(n_767), .B2(n_768), .Y(n_765) );
INVx2_ASAP7_75t_L g455 ( .A(n_454), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g766 ( .A(n_457), .Y(n_766) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g767 ( .A(n_460), .Y(n_767) );
AND3x1_ASAP7_75t_L g460 ( .A(n_461), .B(n_656), .C(n_713), .Y(n_460) );
NOR3xp33_ASAP7_75t_L g461 ( .A(n_462), .B(n_601), .C(n_637), .Y(n_461) );
OAI211xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_510), .B(n_556), .C(n_588), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_483), .Y(n_463) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x4_ASAP7_75t_L g559 ( .A(n_465), .B(n_560), .Y(n_559) );
INVx5_ASAP7_75t_L g587 ( .A(n_465), .Y(n_587) );
AND2x2_ASAP7_75t_L g660 ( .A(n_465), .B(n_576), .Y(n_660) );
AND2x2_ASAP7_75t_L g698 ( .A(n_465), .B(n_604), .Y(n_698) );
AND2x2_ASAP7_75t_L g718 ( .A(n_465), .B(n_561), .Y(n_718) );
OR2x6_ASAP7_75t_L g465 ( .A(n_466), .B(n_480), .Y(n_465) );
AOI21xp5_ASAP7_75t_SL g466 ( .A1(n_467), .A2(n_471), .B(n_479), .Y(n_466) );
BUFx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx5_ASAP7_75t_L g503 ( .A(n_472), .Y(n_503) );
INVx2_ASAP7_75t_L g478 ( .A(n_476), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g504 ( .A1(n_478), .A2(n_505), .B(n_506), .C(n_507), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_L g539 ( .A1(n_478), .A2(n_507), .B(n_540), .C(n_541), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_483), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_498), .Y(n_483) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_484), .Y(n_599) );
AND2x2_ASAP7_75t_L g613 ( .A(n_484), .B(n_560), .Y(n_613) );
INVx1_ASAP7_75t_L g636 ( .A(n_484), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_484), .B(n_587), .Y(n_675) );
OR2x2_ASAP7_75t_L g712 ( .A(n_484), .B(n_558), .Y(n_712) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_485), .Y(n_648) );
AND2x2_ASAP7_75t_L g655 ( .A(n_485), .B(n_561), .Y(n_655) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g576 ( .A(n_486), .B(n_561), .Y(n_576) );
BUFx2_ASAP7_75t_L g604 ( .A(n_486), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_488), .B(n_495), .Y(n_487) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_L g548 ( .A1(n_494), .A2(n_503), .B(n_549), .C(n_550), .Y(n_548) );
O2A1O1Ixp33_ASAP7_75t_SL g563 ( .A1(n_494), .A2(n_503), .B(n_564), .C(n_565), .Y(n_563) );
INVx5_ASAP7_75t_L g558 ( .A(n_498), .Y(n_558) );
BUFx2_ASAP7_75t_L g580 ( .A(n_498), .Y(n_580) );
AND2x2_ASAP7_75t_L g737 ( .A(n_498), .B(n_591), .Y(n_737) );
OR2x6_ASAP7_75t_L g498 ( .A(n_499), .B(n_508), .Y(n_498) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NAND2xp33_ASAP7_75t_L g511 ( .A(n_512), .B(n_543), .Y(n_511) );
OAI221xp5_ASAP7_75t_L g637 ( .A1(n_512), .A2(n_638), .B1(n_645), .B2(n_646), .C(n_649), .Y(n_637) );
OR2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_522), .Y(n_512) );
AND2x2_ASAP7_75t_L g544 ( .A(n_513), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_513), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g572 ( .A(n_514), .B(n_523), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_514), .B(n_524), .Y(n_582) );
OR2x2_ASAP7_75t_L g593 ( .A(n_514), .B(n_545), .Y(n_593) );
AND2x2_ASAP7_75t_L g596 ( .A(n_514), .B(n_584), .Y(n_596) );
AND2x2_ASAP7_75t_L g612 ( .A(n_514), .B(n_534), .Y(n_612) );
OR2x2_ASAP7_75t_L g628 ( .A(n_514), .B(n_524), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_514), .B(n_545), .Y(n_690) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_515), .B(n_534), .Y(n_682) );
AND2x2_ASAP7_75t_L g685 ( .A(n_515), .B(n_524), .Y(n_685) );
OR2x2_ASAP7_75t_L g606 ( .A(n_522), .B(n_593), .Y(n_606) );
INVx2_ASAP7_75t_L g632 ( .A(n_522), .Y(n_632) );
OR2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_534), .Y(n_522) );
AND2x2_ASAP7_75t_L g555 ( .A(n_523), .B(n_535), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_523), .B(n_545), .Y(n_611) );
OR2x2_ASAP7_75t_L g622 ( .A(n_523), .B(n_535), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_523), .B(n_584), .Y(n_681) );
OAI221xp5_ASAP7_75t_L g714 ( .A1(n_523), .A2(n_715), .B1(n_717), .B2(n_719), .C(n_722), .Y(n_714) );
INVx5_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_524), .B(n_545), .Y(n_653) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_527), .B(n_528), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_534), .B(n_584), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_534), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g600 ( .A(n_534), .B(n_572), .Y(n_600) );
OR2x2_ASAP7_75t_L g644 ( .A(n_534), .B(n_545), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_534), .B(n_596), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_534), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g709 ( .A(n_534), .B(n_710), .Y(n_709) );
INVx5_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_SL g573 ( .A(n_535), .B(n_544), .Y(n_573) );
O2A1O1Ixp33_ASAP7_75t_SL g577 ( .A1(n_535), .A2(n_578), .B(n_581), .C(n_585), .Y(n_577) );
OR2x2_ASAP7_75t_L g615 ( .A(n_535), .B(n_611), .Y(n_615) );
OR2x2_ASAP7_75t_L g651 ( .A(n_535), .B(n_593), .Y(n_651) );
OAI311xp33_ASAP7_75t_L g657 ( .A1(n_535), .A2(n_596), .A3(n_658), .B1(n_661), .C1(n_668), .Y(n_657) );
AND2x2_ASAP7_75t_L g708 ( .A(n_535), .B(n_545), .Y(n_708) );
AND2x2_ASAP7_75t_L g716 ( .A(n_535), .B(n_571), .Y(n_716) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_535), .Y(n_734) );
AND2x2_ASAP7_75t_L g751 ( .A(n_535), .B(n_572), .Y(n_751) );
OR2x6_ASAP7_75t_L g535 ( .A(n_536), .B(n_542), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_555), .Y(n_543) );
AND2x2_ASAP7_75t_L g579 ( .A(n_544), .B(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g735 ( .A(n_544), .Y(n_735) );
AND2x2_ASAP7_75t_L g571 ( .A(n_545), .B(n_572), .Y(n_571) );
INVx3_ASAP7_75t_L g584 ( .A(n_545), .Y(n_584) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_545), .Y(n_627) );
INVxp67_ASAP7_75t_L g666 ( .A(n_545), .Y(n_666) );
OA21x2_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .B(n_553), .Y(n_545) );
OA21x2_ASAP7_75t_L g561 ( .A1(n_554), .A2(n_562), .B(n_570), .Y(n_561) );
AND2x2_ASAP7_75t_L g744 ( .A(n_555), .B(n_592), .Y(n_744) );
AOI221xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_571), .B1(n_573), .B2(n_574), .C(n_577), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_558), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g597 ( .A(n_558), .B(n_587), .Y(n_597) );
AND2x2_ASAP7_75t_L g605 ( .A(n_558), .B(n_560), .Y(n_605) );
OR2x2_ASAP7_75t_L g617 ( .A(n_558), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g635 ( .A(n_558), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g659 ( .A(n_558), .B(n_660), .Y(n_659) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_558), .Y(n_679) );
AND2x2_ASAP7_75t_L g731 ( .A(n_558), .B(n_655), .Y(n_731) );
OAI31xp33_ASAP7_75t_L g739 ( .A1(n_558), .A2(n_608), .A3(n_707), .B(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_559), .B(n_635), .Y(n_634) );
INVx1_ASAP7_75t_SL g703 ( .A(n_559), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_559), .B(n_712), .Y(n_711) );
AND2x4_ASAP7_75t_L g591 ( .A(n_560), .B(n_587), .Y(n_591) );
INVx1_ASAP7_75t_L g678 ( .A(n_560), .Y(n_678) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g728 ( .A(n_561), .B(n_587), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx1_ASAP7_75t_SL g738 ( .A(n_571), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_572), .B(n_643), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_573), .A2(n_685), .B1(n_723), .B2(n_726), .Y(n_722) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g586 ( .A(n_576), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g645 ( .A(n_576), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_576), .B(n_597), .Y(n_750) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g720 ( .A(n_579), .B(n_721), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_580), .A2(n_639), .B(n_641), .Y(n_638) );
OR2x2_ASAP7_75t_L g646 ( .A(n_580), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g667 ( .A(n_580), .B(n_655), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_580), .B(n_678), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_580), .B(n_718), .Y(n_717) );
OAI221xp5_ASAP7_75t_SL g694 ( .A1(n_581), .A2(n_695), .B1(n_700), .B2(n_703), .C(n_704), .Y(n_694) );
OR2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
OR2x2_ASAP7_75t_L g671 ( .A(n_582), .B(n_644), .Y(n_671) );
INVx1_ASAP7_75t_L g710 ( .A(n_582), .Y(n_710) );
INVx2_ASAP7_75t_L g686 ( .A(n_583), .Y(n_686) );
INVx1_ASAP7_75t_L g620 ( .A(n_584), .Y(n_620) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g625 ( .A(n_587), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_587), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g654 ( .A(n_587), .B(n_655), .Y(n_654) );
OR2x2_ASAP7_75t_L g742 ( .A(n_587), .B(n_712), .Y(n_742) );
AOI222xp33_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_592), .B1(n_594), .B2(n_597), .C1(n_598), .C2(n_600), .Y(n_588) );
INVxp67_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g598 ( .A(n_591), .B(n_599), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_591), .A2(n_641), .B1(n_669), .B2(n_670), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_591), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
OAI21xp33_ASAP7_75t_SL g629 ( .A1(n_600), .A2(n_630), .B(n_633), .Y(n_629) );
OAI211xp5_ASAP7_75t_SL g601 ( .A1(n_602), .A2(n_606), .B(n_607), .C(n_629), .Y(n_601) );
INVxp67_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
AOI221xp5_ASAP7_75t_L g607 ( .A1(n_605), .A2(n_608), .B1(n_613), .B2(n_614), .C(n_616), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_605), .B(n_693), .Y(n_692) );
INVxp67_ASAP7_75t_L g699 ( .A(n_605), .Y(n_699) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_612), .Y(n_609) );
AND2x2_ASAP7_75t_L g701 ( .A(n_610), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g618 ( .A(n_613), .Y(n_618) );
AND2x2_ASAP7_75t_L g624 ( .A(n_613), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_619), .B1(n_623), .B2(n_626), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_620), .B(n_632), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_621), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g721 ( .A(n_625), .Y(n_721) );
AND2x2_ASAP7_75t_L g740 ( .A(n_625), .B(n_655), .Y(n_740) );
OR2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_632), .B(n_689), .Y(n_748) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_635), .B(n_703), .Y(n_746) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g669 ( .A(n_647), .Y(n_669) );
BUFx2_ASAP7_75t_L g693 ( .A(n_648), .Y(n_693) );
OAI21xp5_ASAP7_75t_SL g649 ( .A1(n_650), .A2(n_652), .B(n_654), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NOR3xp33_ASAP7_75t_L g656 ( .A(n_657), .B(n_672), .C(n_694), .Y(n_656) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OAI21xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_664), .B(n_667), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
A2O1A1Ixp33_ASAP7_75t_SL g672 ( .A1(n_673), .A2(n_676), .B(n_680), .C(n_683), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_673), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NOR2xp67_ASAP7_75t_SL g677 ( .A(n_678), .B(n_679), .Y(n_677) );
OR2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
INVx1_ASAP7_75t_SL g702 ( .A(n_682), .Y(n_702) );
OAI21xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_687), .B(n_691), .Y(n_683) );
AND2x4_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
AND2x2_ASAP7_75t_L g707 ( .A(n_685), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_697), .B(n_699), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_707), .B1(n_709), .B2(n_711), .Y(n_704) );
INVx2_ASAP7_75t_SL g725 ( .A(n_712), .Y(n_725) );
NOR3xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_729), .C(n_741), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVxp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVxp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_725), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OAI221xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_732), .B1(n_736), .B2(n_738), .C(n_739), .Y(n_729) );
A2O1A1Ixp33_ASAP7_75t_L g741 ( .A1(n_730), .A2(n_742), .B(n_743), .C(n_745), .Y(n_741) );
INVx1_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
INVxp67_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_747), .B1(n_749), .B2(n_751), .Y(n_745) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g768 ( .A(n_753), .Y(n_768) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g763 ( .A(n_760), .Y(n_763) );
INVx1_ASAP7_75t_SL g769 ( .A(n_770), .Y(n_769) );
INVx3_ASAP7_75t_SL g770 ( .A(n_771), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
endmodule