module real_jpeg_16044_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_0),
.B(n_22),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_1),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_1),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_1),
.B(n_110),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_1),
.B(n_125),
.Y(n_214)
);

AND2x2_ASAP7_75t_SL g263 ( 
.A(n_1),
.B(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_2),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_2),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_3),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_3),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_3),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_3),
.B(n_165),
.Y(n_164)
);

NAND2xp67_ASAP7_75t_L g204 ( 
.A(n_3),
.B(n_202),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_3),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_3),
.B(n_256),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_3),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_4),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_4),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_4),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_5),
.B(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_5),
.B(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g288 ( 
.A(n_5),
.B(n_289),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_5),
.B(n_87),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_6),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_6),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_6),
.B(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_7),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_7),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_7),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_8),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_8),
.Y(n_238)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_8),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_9),
.A2(n_19),
.B(n_21),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_10),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_10),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_10),
.B(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_10),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_10),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_10),
.B(n_161),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_10),
.B(n_190),
.Y(n_189)
);

AND2x2_ASAP7_75t_SL g201 ( 
.A(n_10),
.B(n_202),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_11),
.B(n_27),
.Y(n_26)
);

NAND2x1_ASAP7_75t_L g32 ( 
.A(n_11),
.B(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_11),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_11),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_11),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_11),
.B(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_11),
.B(n_222),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_11),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_12),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_12),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_12),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_12),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_12),
.B(n_179),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_12),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_12),
.B(n_356),
.Y(n_355)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_13),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_13),
.Y(n_94)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_13),
.Y(n_298)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_14),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_14),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_14),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_14),
.B(n_27),
.Y(n_262)
);

AND2x2_ASAP7_75t_SL g327 ( 
.A(n_14),
.B(n_328),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_15),
.Y(n_83)
);

BUFx4f_ASAP7_75t_L g130 ( 
.A(n_16),
.Y(n_130)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_16),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_16),
.Y(n_192)
);

BUFx8_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_17),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g349 ( 
.A(n_17),
.Y(n_349)
);

BUFx12f_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

O2A1O1Ixp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_115),
.B(n_346),
.C(n_415),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_39),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_24),
.A2(n_25),
.B1(n_60),
.B2(n_72),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.C(n_36),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_26),
.A2(n_30),
.B1(n_31),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_26),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_26),
.B(n_53),
.C(n_55),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_26),
.A2(n_46),
.B1(n_55),
.B2(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_26),
.B(n_197),
.C(n_201),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_26),
.A2(n_46),
.B1(n_197),
.B2(n_198),
.Y(n_272)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_29),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_30),
.A2(n_68),
.B(n_71),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_30),
.B(n_68),
.Y(n_71)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_31),
.A2(n_32),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_32),
.Y(n_211)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_34),
.Y(n_326)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_35),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_36),
.B(n_354),
.Y(n_353)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_37),
.Y(n_200)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_38),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_73),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_40),
.B(n_73),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_59),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_47),
.C(n_52),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_SL g74 ( 
.A(n_42),
.B(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_43),
.B(n_201),
.C(n_358),
.Y(n_378)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_48),
.B1(n_52),
.B2(n_76),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx12_ASAP7_75t_R g76 ( 
.A(n_52),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_53),
.B(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_104),
.C(n_107),
.Y(n_103)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_55),
.B(n_157),
.C(n_160),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_55),
.A2(n_104),
.B1(n_114),
.B2(n_320),
.Y(n_376)
);

OR2x2_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_58),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_66),
.B2(n_67),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_61),
.A2(n_62),
.B1(n_386),
.B2(n_387),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_79),
.C(n_85),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_62),
.B(n_71),
.Y(n_415)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_64),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_65),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_68),
.B(n_220),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_68),
.B(n_193),
.C(n_224),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.C(n_100),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_74),
.B(n_77),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_89),
.C(n_95),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_78),
.B(n_102),
.Y(n_101)
);

INVxp33_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_80),
.B(n_85),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_82),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_83),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_83),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_84),
.B(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_85),
.A2(n_86),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_85),
.B(n_204),
.C(n_206),
.Y(n_216)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_88),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_90),
.B1(n_95),
.B2(n_96),
.Y(n_102)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_96),
.A2(n_97),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

MAJx2_ASAP7_75t_L g342 ( 
.A(n_96),
.B(n_215),
.C(n_216),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_96),
.B(n_346),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_96),
.B(n_346),
.C(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_100),
.B(n_391),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.C(n_112),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_101),
.B(n_373),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_103),
.B(n_112),
.Y(n_373)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_104),
.B(n_262),
.C(n_263),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_104),
.A2(n_262),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_104),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_104),
.A2(n_221),
.B1(n_224),
.B2(n_320),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_SL g377 ( 
.A(n_104),
.B(n_224),
.C(n_361),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_106),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_107),
.B(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_114),
.B(n_284),
.Y(n_283)
);

O2A1O1Ixp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_369),
.B(n_409),
.C(n_414),
.Y(n_115)
);

A2O1A1O1Ixp25_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_276),
.B(n_331),
.C(n_332),
.D(n_368),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_243),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_119),
.B(n_243),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_180),
.Y(n_119)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_120),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_154),
.C(n_173),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_122),
.B(n_246),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_134),
.C(n_143),
.Y(n_122)
);

XNOR2x1_ASAP7_75t_SL g299 ( 
.A(n_123),
.B(n_300),
.Y(n_299)
);

XNOR2x2_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_124),
.B(n_127),
.C(n_131),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_133),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_134),
.A2(n_135),
.B1(n_143),
.B2(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_135),
.A2(n_136),
.B(n_140),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_140),
.Y(n_135)
);

INVx4_ASAP7_75t_SL g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_143),
.Y(n_301)
);

MAJx3_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.C(n_152),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_144),
.B(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_148),
.B(n_152),
.Y(n_251)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_151),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_155),
.A2(n_173),
.B1(n_174),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_155),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_164),
.C(n_167),
.Y(n_155)
);

XNOR2x2_ASAP7_75t_SL g268 ( 
.A(n_156),
.B(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_157),
.B(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_160),
.B(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_160),
.Y(n_284)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_164),
.B(n_167),
.Y(n_269)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

MAJx2_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_178),
.C(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_218),
.B1(n_241),
.B2(n_242),
.Y(n_180)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_181),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_208),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_182),
.B(n_209),
.C(n_217),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_196),
.C(n_203),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_183),
.B(n_196),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g227 ( 
.A1(n_184),
.A2(n_189),
.B(n_193),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_193),
.B2(n_195),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_188),
.A2(n_189),
.B1(n_254),
.B2(n_255),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_193),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_189),
.B(n_254),
.Y(n_253)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_193),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_193),
.A2(n_195),
.B1(n_221),
.B2(n_224),
.Y(n_220)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_201),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_201),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_201),
.A2(n_273),
.B1(n_355),
.B2(n_358),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_202),
.Y(n_328)
);

XOR2x2_ASAP7_75t_L g274 ( 
.A(n_203),
.B(n_275),
.Y(n_274)
);

XNOR2x1_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_206),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_212),
.B2(n_217),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_212),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_216),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_214),
.Y(n_215)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_218),
.B(n_241),
.C(n_335),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_225),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_219),
.B(n_226),
.C(n_229),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_221),
.Y(n_224)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_229),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_228),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_235),
.B1(n_239),
.B2(n_240),
.Y(n_230)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_231),
.Y(n_240)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_235),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_235),
.B(n_240),
.C(n_284),
.Y(n_352)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_248),
.C(n_274),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_244),
.A2(n_245),
.B1(n_274),
.B2(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_248),
.B(n_303),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_268),
.C(n_270),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_280),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.C(n_261),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_250),
.B(n_314),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_252),
.A2(n_253),
.B1(n_261),
.B2(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_257),
.Y(n_256)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_261),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_262),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_263),
.B(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_270),
.Y(n_280)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_274),
.Y(n_304)
);

AOI21x1_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_305),
.B(n_330),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_302),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_278),
.B(n_302),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_281),
.C(n_299),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_279),
.B(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_281),
.B(n_299),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_285),
.C(n_286),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_282),
.B(n_285),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.C(n_292),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_308),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_312),
.C(n_316),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_321),
.C(n_322),
.Y(n_316)
);

MAJx2_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_327),
.C(n_329),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_336),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_334),
.B(n_336),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_337),
.B(n_339),
.C(n_350),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_350),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_340),
.B(n_342),
.C(n_343),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

XNOR2x1_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_344),
.Y(n_389)
);

INVx3_ASAP7_75t_SL g347 ( 
.A(n_348),
.Y(n_347)
);

INVx8_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_359),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_352),
.B(n_359),
.C(n_383),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_353),
.Y(n_383)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_355),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

NAND3xp33_ASAP7_75t_SL g369 ( 
.A(n_370),
.B(n_392),
.C(n_404),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_370),
.A2(n_410),
.B(n_413),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_390),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_371),
.B(n_390),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_374),
.C(n_379),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_372),
.B(n_374),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_377),
.C(n_378),
.Y(n_374)
);

XNOR2x2_ASAP7_75t_L g397 ( 
.A(n_375),
.B(n_398),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_377),
.B(n_378),
.Y(n_398)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_380),
.B(n_407),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_384),
.C(n_388),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_401),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_384),
.A2(n_385),
.B1(n_388),
.B2(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_388),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_394),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_393),
.B(n_394),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_403),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_397),
.B1(n_399),
.B2(n_400),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_397),
.B(n_399),
.C(n_403),
.Y(n_408)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_405),
.A2(n_411),
.B(n_412),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_SL g405 ( 
.A(n_406),
.B(n_408),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_406),
.B(n_408),
.Y(n_412)
);


endmodule