module fake_ibex_1145_n_4398 (n_151, n_85, n_599, n_778, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_781, n_421, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_739, n_755, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_598, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_168, n_526, n_785, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_789, n_654, n_656, n_724, n_437, n_731, n_602, n_355, n_767, n_474, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_793, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_772, n_810, n_768, n_338, n_173, n_696, n_796, n_797, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_257, n_77, n_718, n_801, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_803, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_776, n_409, n_582, n_653, n_214, n_238, n_579, n_332, n_799, n_517, n_211, n_744, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_217, n_324, n_391, n_537, n_728, n_78, n_805, n_670, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_668, n_779, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_232, n_380, n_749, n_281, n_559, n_425, n_4398);

input n_151;
input n_85;
input n_599;
input n_778;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_781;
input n_421;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_739;
input n_755;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_168;
input n_526;
input n_785;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_789;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_355;
input n_767;
input n_474;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_772;
input n_810;
input n_768;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_718;
input n_801;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_217;
input n_324;
input n_391;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_668;
input n_779;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_232;
input n_380;
input n_749;
input n_281;
input n_559;
input n_425;

output n_4398;

wire n_1084;
wire n_4368;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_4234;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_4146;
wire n_2835;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_4158;
wire n_845;
wire n_4095;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_4204;
wire n_4364;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_3812;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_3750;
wire n_3838;
wire n_957;
wire n_3255;
wire n_3674;
wire n_3272;
wire n_4249;
wire n_1652;
wire n_969;
wire n_1859;
wire n_2183;
wire n_1954;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_4159;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_2640;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_930;
wire n_4372;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_4343;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_4353;
wire n_1722;
wire n_4371;
wire n_3931;
wire n_911;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_4179;
wire n_3340;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_4360;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_3904;
wire n_4378;
wire n_850;
wire n_4169;
wire n_3175;
wire n_3729;
wire n_4239;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_3984;
wire n_4233;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_3721;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_4172;
wire n_1730;
wire n_4277;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_3479;
wire n_1840;
wire n_2837;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_3982;
wire n_2605;
wire n_2343;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_4201;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_4285;
wire n_1681;
wire n_2921;
wire n_4031;
wire n_3724;
wire n_939;
wire n_1636;
wire n_1687;
wire n_4120;
wire n_3192;
wire n_3533;
wire n_3896;
wire n_3753;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_4155;
wire n_1922;
wire n_3890;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_2311;
wire n_1937;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_3839;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3472;
wire n_3509;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_3976;
wire n_824;
wire n_4304;
wire n_4348;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_4160;
wire n_4382;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_4002;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_3969;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_4311;
wire n_2432;
wire n_3043;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_4144;
wire n_2273;
wire n_3298;
wire n_852;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_4211;
wire n_3264;
wire n_3204;
wire n_4119;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_3747;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3881;
wire n_3884;
wire n_3507;
wire n_3949;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2436;
wire n_2333;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_857;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_4389;
wire n_2846;
wire n_2685;
wire n_3197;
wire n_3699;
wire n_1955;
wire n_3668;
wire n_4312;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_3766;
wire n_4014;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_4217;
wire n_3973;
wire n_1313;
wire n_4214;
wire n_4223;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3977;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_4221;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_3943;
wire n_3809;
wire n_979;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_4295;
wire n_1716;
wire n_4238;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_3667;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_3822;
wire n_4171;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_3858;
wire n_4182;
wire n_1401;
wire n_4173;
wire n_3764;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_4166;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_4259;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_4188;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_4060;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_1653;
wire n_4067;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_4124;
wire n_971;
wire n_1326;
wire n_1350;
wire n_3627;
wire n_906;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_4393;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_1506;
wire n_881;
wire n_2987;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_4078;
wire n_4283;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_4174;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_4392;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_4054;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4129;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_4352;
wire n_3530;
wire n_1613;
wire n_820;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_4258;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_4290;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2660;
wire n_4252;
wire n_2661;
wire n_4079;
wire n_4219;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_4248;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2625;
wire n_2350;
wire n_1742;
wire n_2444;
wire n_4240;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_4055;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2646;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_3241;
wire n_2746;
wire n_2256;
wire n_3317;
wire n_3800;
wire n_3887;
wire n_3963;
wire n_3461;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_4103;
wire n_3583;
wire n_2019;
wire n_4126;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_889;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_4359;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_4331;
wire n_2602;
wire n_4090;
wire n_1441;
wire n_4105;
wire n_4206;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_4136;
wire n_1924;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_819;
wire n_3950;
wire n_4177;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_4156;
wire n_3754;
wire n_1964;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_4074;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_4355;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_4308;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_4271;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3788;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3634;
wire n_1377;
wire n_2473;
wire n_4096;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_3054;
wire n_2924;
wire n_2264;
wire n_2076;
wire n_2599;
wire n_974;
wire n_1036;
wire n_1831;
wire n_3626;
wire n_3733;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_4293;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_4039;
wire n_4253;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_4122;
wire n_2622;
wire n_3232;
wire n_4250;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_4374;
wire n_1140;
wire n_1985;
wire n_4375;
wire n_4205;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1421;
wire n_1203;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2880;
wire n_2390;
wire n_2573;
wire n_2423;
wire n_4230;
wire n_859;
wire n_3849;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_4333;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_4070;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_4134;
wire n_1051;
wire n_4180;
wire n_4131;
wire n_1008;
wire n_3065;
wire n_2964;
wire n_2375;
wire n_4062;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_4330;
wire n_1656;
wire n_1207;
wire n_4040;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_4232;
wire n_1589;
wire n_2717;
wire n_4199;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_3855;
wire n_4033;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_1236;
wire n_3364;
wire n_4384;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_4231;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1477;
wire n_1184;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_4323;
wire n_4184;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1890;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_4073;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_4325;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_4113;
wire n_1229;
wire n_4337;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_4292;
wire n_4187;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_4261;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_4063;
wire n_1464;
wire n_1566;
wire n_4362;
wire n_3568;
wire n_944;
wire n_3312;
wire n_4128;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_3331;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_4114;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_4347;
wire n_1852;
wire n_4191;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_827;
wire n_4209;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_4011;
wire n_4190;
wire n_2954;
wire n_4307;
wire n_3526;
wire n_2102;
wire n_4356;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_4151;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_4170;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_4097;
wire n_1436;
wire n_3239;
wire n_4137;
wire n_2600;
wire n_1485;
wire n_1069;
wire n_2239;
wire n_4152;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_4365;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_1345;
wire n_4215;
wire n_4315;
wire n_2434;
wire n_837;
wire n_1590;
wire n_2971;
wire n_2332;
wire n_954;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3797;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3584;
wire n_1395;
wire n_1729;
wire n_998;
wire n_1115;
wire n_2551;
wire n_3281;
wire n_2823;
wire n_3274;
wire n_4064;
wire n_4110;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_4379;
wire n_3397;
wire n_2934;
wire n_4145;
wire n_2807;
wire n_4047;
wire n_882;
wire n_4157;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_4042;
wire n_2525;
wire n_814;
wire n_3829;
wire n_1864;
wire n_943;
wire n_4317;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1523;
wire n_1086;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_4041;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_4297;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_2570;
wire n_4051;
wire n_4321;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_3948;
wire n_1599;
wire n_1400;
wire n_1539;
wire n_1806;
wire n_2842;
wire n_3070;
wire n_2711;
wire n_3477;
wire n_2635;
wire n_3646;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_4077;
wire n_3897;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_2193;
wire n_817;
wire n_2612;
wire n_3034;
wire n_4010;
wire n_4255;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_4059;
wire n_4130;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_4361;
wire n_3974;
wire n_1574;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_4237;
wire n_1746;
wire n_2716;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_3495;
wire n_863;
wire n_2185;
wire n_4141;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_4035;
wire n_2781;
wire n_4291;
wire n_3419;
wire n_3629;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_3999;
wire n_4117;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_4087;
wire n_3167;
wire n_3687;
wire n_997;
wire n_4154;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_4318;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_4385;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_4052;
wire n_2463;
wire n_2654;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_4072;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_4245;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_4100;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_4195;
wire n_836;
wire n_1475;
wire n_3316;
wire n_2465;
wire n_1263;
wire n_3337;
wire n_3925;
wire n_4089;
wire n_4176;
wire n_1185;
wire n_1683;
wire n_4256;
wire n_3575;
wire n_4175;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_4278;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_2948;
wire n_916;
wire n_4322;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_2936;
wire n_895;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_4227;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_4030;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_4276;
wire n_831;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1845;
wire n_1104;
wire n_2205;
wire n_1011;
wire n_2875;
wire n_2684;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_3902;
wire n_3927;
wire n_2422;
wire n_4185;
wire n_4203;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_4381;
wire n_1917;
wire n_4314;
wire n_1444;
wire n_4133;
wire n_920;
wire n_4316;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_4083;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_4306;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_3064;
wire n_2896;
wire n_4228;
wire n_2997;
wire n_3314;
wire n_1349;
wire n_1331;
wire n_961;
wire n_991;
wire n_1223;
wire n_2127;
wire n_3735;
wire n_1323;
wire n_3891;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_4254;
wire n_3420;
wire n_1432;
wire n_4192;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_4388;
wire n_996;
wire n_3914;
wire n_3632;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_4138;
wire n_3552;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_4116;
wire n_4164;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1601;
wire n_1294;
wire n_900;
wire n_4142;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_4118;
wire n_4183;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_4284;
wire n_1458;
wire n_1694;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_4066;
wire n_3990;
wire n_3673;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_4044;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3269;
wire n_3029;
wire n_3609;
wire n_4135;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_2223;
wire n_1850;
wire n_1660;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4000;
wire n_3154;
wire n_4123;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_4305;
wire n_2902;
wire n_4048;
wire n_4084;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3960;
wire n_4007;
wire n_3608;
wire n_4339;
wire n_4269;
wire n_4085;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_3878;
wire n_4016;
wire n_2849;
wire n_2947;
wire n_4080;
wire n_1754;
wire n_4286;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_4028;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_4289;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_4163;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3778;
wire n_3912;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_3047;
wire n_1625;
wire n_2959;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_4001;
wire n_1348;
wire n_1289;
wire n_838;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_3356;
wire n_1191;
wire n_2004;
wire n_4099;
wire n_4377;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_4264;
wire n_1942;
wire n_4326;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_3899;
wire n_3930;
wire n_1587;
wire n_2330;
wire n_2639;
wire n_2555;
wire n_4149;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_4101;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_4057;
wire n_2410;
wire n_3760;
wire n_4319;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_4021;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_4383;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3462;
wire n_3745;
wire n_3424;
wire n_4373;
wire n_2437;
wire n_2351;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_4132;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_851;
wire n_4202;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_4287;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_4300;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_4022;
wire n_4212;
wire n_1241;
wire n_3645;
wire n_4262;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_4019;
wire n_2736;
wire n_4320;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_826;
wire n_2154;
wire n_1976;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_3162;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_1647;
wire n_1901;
wire n_4357;
wire n_3096;
wire n_3333;
wire n_839;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_3276;
wire n_4366;
wire n_1006;
wire n_2956;
wire n_1415;
wire n_1238;
wire n_3959;
wire n_3743;
wire n_976;
wire n_1710;
wire n_4139;
wire n_3021;
wire n_1063;
wire n_4068;
wire n_4288;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_4340;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_3860;
wire n_2137;
wire n_1455;
wire n_1871;
wire n_1642;
wire n_2182;
wire n_3044;
wire n_2868;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_3784;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_4034;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_4082;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_3273;
wire n_4367;
wire n_950;
wire n_2700;
wire n_3139;
wire n_1222;
wire n_4282;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_4222;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3538;
wire n_1261;
wire n_2299;
wire n_3393;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_818;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_4029;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_3454;
wire n_4334;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_4143;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_2608;
wire n_4270;
wire n_3384;
wire n_2983;
wire n_4273;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_4338;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3604;
wire n_833;
wire n_3649;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_4198;
wire n_1513;
wire n_3740;
wire n_4397;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_4186;
wire n_2093;
wire n_2348;
wire n_2675;
wire n_2417;
wire n_2576;
wire n_2043;
wire n_3601;
wire n_4344;
wire n_2366;
wire n_4229;
wire n_4294;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_4351;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_4111;
wire n_4162;
wire n_4200;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_4341;
wire n_4328;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_4127;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_4076;
wire n_4189;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_4390;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_4058;
wire n_1275;
wire n_985;
wire n_1165;
wire n_4148;
wire n_1622;
wire n_897;
wire n_2757;
wire n_3066;
wire n_2714;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_4032;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_4268;
wire n_1507;
wire n_1809;
wire n_1206;
wire n_855;
wire n_2367;
wire n_3236;
wire n_3576;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3271;
wire n_3013;
wire n_2667;
wire n_1050;
wire n_2218;
wire n_2553;
wire n_4265;
wire n_3062;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_4260;
wire n_3391;
wire n_4017;
wire n_1547;
wire n_946;
wire n_1586;
wire n_1362;
wire n_1542;
wire n_3497;
wire n_4178;
wire n_4324;
wire n_1097;
wire n_3354;
wire n_4069;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_4236;
wire n_3012;
wire n_4313;
wire n_4140;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3586;
wire n_956;
wire n_3561;
wire n_4125;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_2574;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_4242;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_4243;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_4053;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_4279;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1584;
wire n_1481;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_4235;
wire n_1438;
wire n_3774;
wire n_3972;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_4036;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1518;
wire n_1366;
wire n_4350;
wire n_4380;
wire n_1361;
wire n_1187;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_3173;
wire n_2872;
wire n_3102;
wire n_4281;
wire n_4345;
wire n_2411;
wire n_4332;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_3844;
wire n_883;
wire n_2207;
wire n_4210;
wire n_4049;
wire n_2044;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_1572;
wire n_1635;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_3163;
wire n_2929;
wire n_3343;
wire n_3752;
wire n_4310;
wire n_3786;
wire n_4061;
wire n_1329;
wire n_2637;
wire n_2409;
wire n_2337;
wire n_4045;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3543;
wire n_3791;
wire n_3742;
wire n_3655;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_2323;
wire n_3532;
wire n_4257;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_4263;
wire n_3725;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_4363;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_4196;
wire n_4335;
wire n_2371;
wire n_914;
wire n_3992;
wire n_4147;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_4218;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_4301;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_4161;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_4267;
wire n_4386;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_2942;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_4193;
wire n_2296;
wire n_4342;
wire n_3782;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_4302;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_2310;
wire n_3318;
wire n_3223;
wire n_4013;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1488;
wire n_1193;
wire n_849;
wire n_980;
wire n_3067;
wire n_2928;
wire n_2227;
wire n_2652;
wire n_3225;
wire n_1074;
wire n_3557;
wire n_3380;
wire n_3207;
wire n_3596;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_4086;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_4112;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_4207;
wire n_960;
wire n_1022;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_4266;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3286;
wire n_3124;
wire n_1092;
wire n_4038;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_4102;
wire n_3612;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1385;
wire n_1142;
wire n_2927;
wire n_4274;
wire n_1062;
wire n_4395;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_3893;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_4272;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2303;
wire n_2357;
wire n_2618;
wire n_2653;
wire n_2855;
wire n_3938;
wire n_4354;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_4296;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_4088;
wire n_2136;
wire n_4309;
wire n_3617;
wire n_4027;
wire n_3602;
wire n_4298;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2560;
wire n_2453;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_4208;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2802;
wire n_2443;
wire n_3052;
wire n_3189;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_2066;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_4046;
wire n_4275;
wire n_2770;
wire n_2961;
wire n_2704;
wire n_2996;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_2168;
wire n_1948;
wire n_3247;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_4094;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_3613;
wire n_1383;
wire n_990;
wire n_4108;
wire n_1968;
wire n_3675;
wire n_2057;
wire n_2609;
wire n_4018;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_3715;
wire n_4194;
wire n_1059;
wire n_2969;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_3933;
wire n_955;
wire n_1916;
wire n_1333;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_3873;
wire n_3738;
wire n_2073;
wire n_4093;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_4226;
wire n_1551;
wire n_3793;
wire n_4153;
wire n_1533;
wire n_1145;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_4329;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_3988;
wire n_4327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_4168;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_4396;
wire n_2039;
wire n_1696;
wire n_1277;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_3691;
wire n_2544;
wire n_856;
wire n_3193;
wire n_3501;
wire n_3635;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_3258;
wire n_2932;
wire n_1335;
wire n_3266;
wire n_4280;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_4394;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1678;
wire n_1780;
wire n_1091;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_4220;
wire n_4075;
wire n_860;
wire n_1525;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_4224;
wire n_970;
wire n_3654;
wire n_3980;
wire n_2673;
wire n_2676;
wire n_921;
wire n_2430;
wire n_3515;
wire n_3489;
wire n_4213;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_4387;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_1655;
wire n_984;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_866;
wire n_2658;

INVx1_ASAP7_75t_L g814 ( 
.A(n_629),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_759),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_716),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_283),
.Y(n_817)
);

INVx1_ASAP7_75t_SL g818 ( 
.A(n_199),
.Y(n_818)
);

CKINVDCx14_ASAP7_75t_R g819 ( 
.A(n_219),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_194),
.Y(n_820)
);

BUFx2_ASAP7_75t_SL g821 ( 
.A(n_788),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_387),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_483),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_218),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_198),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_375),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_511),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_251),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_564),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_252),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_418),
.Y(n_831)
);

INVxp67_ASAP7_75t_L g832 ( 
.A(n_504),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_616),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_670),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_727),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_265),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_213),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_494),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_40),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_296),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_538),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_234),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_49),
.Y(n_843)
);

CKINVDCx20_ASAP7_75t_R g844 ( 
.A(n_602),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_579),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_412),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_248),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_432),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_260),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_333),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_778),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_49),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_85),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_624),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_265),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_665),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_238),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_282),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_617),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_791),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_346),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_563),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_676),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_92),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_222),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_792),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_804),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_607),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_222),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_700),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_361),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_593),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_537),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_367),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_537),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_768),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_242),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_248),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_277),
.Y(n_879)
);

CKINVDCx14_ASAP7_75t_R g880 ( 
.A(n_676),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_768),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_538),
.Y(n_882)
);

INVxp67_ASAP7_75t_SL g883 ( 
.A(n_258),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_305),
.Y(n_884)
);

BUFx2_ASAP7_75t_L g885 ( 
.A(n_19),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_48),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_170),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_562),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_13),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_777),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_512),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_241),
.Y(n_892)
);

INVx1_ASAP7_75t_SL g893 ( 
.A(n_667),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_91),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_477),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_530),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_636),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_794),
.Y(n_898)
);

CKINVDCx16_ASAP7_75t_R g899 ( 
.A(n_2),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_302),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_269),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_437),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_291),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_645),
.Y(n_904)
);

CKINVDCx20_ASAP7_75t_R g905 ( 
.A(n_40),
.Y(n_905)
);

INVxp67_ASAP7_75t_L g906 ( 
.A(n_454),
.Y(n_906)
);

INVxp67_ASAP7_75t_L g907 ( 
.A(n_235),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_772),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_33),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_124),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_566),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_30),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_458),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_747),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_785),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_16),
.Y(n_916)
);

CKINVDCx20_ASAP7_75t_R g917 ( 
.A(n_30),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_804),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_632),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_799),
.Y(n_920)
);

BUFx3_ASAP7_75t_L g921 ( 
.A(n_402),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_762),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_221),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_172),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_729),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_770),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_151),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_774),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_435),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_794),
.Y(n_930)
);

CKINVDCx20_ASAP7_75t_R g931 ( 
.A(n_101),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_188),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_425),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_784),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_240),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_713),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_495),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_162),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_327),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_765),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_578),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_731),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_781),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_61),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_576),
.Y(n_945)
);

CKINVDCx20_ASAP7_75t_R g946 ( 
.A(n_365),
.Y(n_946)
);

INVx1_ASAP7_75t_SL g947 ( 
.A(n_70),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_626),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_391),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_545),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_45),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_478),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_284),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_180),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_578),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_254),
.Y(n_956)
);

INVx2_ASAP7_75t_SL g957 ( 
.A(n_363),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_563),
.Y(n_958)
);

INVxp67_ASAP7_75t_SL g959 ( 
.A(n_263),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_105),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_221),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_746),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_294),
.Y(n_963)
);

BUFx5_ASAP7_75t_L g964 ( 
.A(n_712),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_750),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_230),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_800),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_157),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_807),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_57),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_725),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_322),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_704),
.Y(n_973)
);

BUFx2_ASAP7_75t_SL g974 ( 
.A(n_769),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_417),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_448),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_80),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_76),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_566),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_677),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_169),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_796),
.Y(n_982)
);

CKINVDCx16_ASAP7_75t_R g983 ( 
.A(n_362),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_780),
.Y(n_984)
);

CKINVDCx16_ASAP7_75t_R g985 ( 
.A(n_346),
.Y(n_985)
);

CKINVDCx20_ASAP7_75t_R g986 ( 
.A(n_251),
.Y(n_986)
);

CKINVDCx16_ASAP7_75t_R g987 ( 
.A(n_700),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_659),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_416),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_8),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_603),
.Y(n_991)
);

INVx2_ASAP7_75t_SL g992 ( 
.A(n_740),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_677),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_667),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_648),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_665),
.Y(n_996)
);

CKINVDCx20_ASAP7_75t_R g997 ( 
.A(n_13),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_678),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_793),
.Y(n_999)
);

BUFx10_ASAP7_75t_L g1000 ( 
.A(n_521),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_362),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_421),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_779),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_547),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_795),
.Y(n_1005)
);

BUFx2_ASAP7_75t_L g1006 ( 
.A(n_232),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_339),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_195),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_523),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_114),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_675),
.Y(n_1011)
);

BUFx5_ASAP7_75t_L g1012 ( 
.A(n_728),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_767),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_242),
.Y(n_1014)
);

BUFx3_ASAP7_75t_L g1015 ( 
.A(n_619),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_96),
.Y(n_1016)
);

INVx1_ASAP7_75t_SL g1017 ( 
.A(n_607),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_510),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_697),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_775),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_251),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_104),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_37),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_151),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_661),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_772),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_334),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_777),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_53),
.Y(n_1029)
);

CKINVDCx16_ASAP7_75t_R g1030 ( 
.A(n_249),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_778),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_356),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_72),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_43),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_15),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_773),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_7),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_471),
.Y(n_1038)
);

INVx2_ASAP7_75t_SL g1039 ( 
.A(n_543),
.Y(n_1039)
);

BUFx10_ASAP7_75t_L g1040 ( 
.A(n_322),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_618),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_273),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_385),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_31),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_29),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_710),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_519),
.Y(n_1047)
);

INVx1_ASAP7_75t_SL g1048 ( 
.A(n_551),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_76),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_342),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_151),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_41),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_686),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_686),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_76),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_357),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_44),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_724),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_357),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_735),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_419),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_526),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_801),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_144),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_438),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_770),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_507),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_526),
.Y(n_1068)
);

BUFx8_ASAP7_75t_SL g1069 ( 
.A(n_758),
.Y(n_1069)
);

BUFx10_ASAP7_75t_L g1070 ( 
.A(n_639),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_633),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_78),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_270),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_28),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_654),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_642),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_283),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_735),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_629),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_299),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_93),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_152),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_444),
.Y(n_1083)
);

CKINVDCx20_ASAP7_75t_R g1084 ( 
.A(n_253),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_542),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_388),
.Y(n_1086)
);

INVx1_ASAP7_75t_SL g1087 ( 
.A(n_28),
.Y(n_1087)
);

BUFx10_ASAP7_75t_L g1088 ( 
.A(n_143),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_691),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_766),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_714),
.Y(n_1091)
);

CKINVDCx16_ASAP7_75t_R g1092 ( 
.A(n_440),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_397),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_267),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_195),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_224),
.Y(n_1096)
);

INVx2_ASAP7_75t_SL g1097 ( 
.A(n_634),
.Y(n_1097)
);

BUFx10_ASAP7_75t_L g1098 ( 
.A(n_812),
.Y(n_1098)
);

CKINVDCx20_ASAP7_75t_R g1099 ( 
.A(n_503),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_675),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_57),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_776),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_424),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_28),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_267),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_482),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_672),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_340),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_456),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_117),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_790),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_334),
.Y(n_1112)
);

BUFx10_ASAP7_75t_L g1113 ( 
.A(n_207),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_608),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_783),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_159),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_703),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_298),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_73),
.Y(n_1119)
);

BUFx10_ASAP7_75t_L g1120 ( 
.A(n_354),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_52),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_785),
.Y(n_1122)
);

CKINVDCx6p67_ASAP7_75t_R g1123 ( 
.A(n_781),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_129),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_25),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_763),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_307),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_392),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_596),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_197),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_417),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_448),
.Y(n_1132)
);

BUFx10_ASAP7_75t_L g1133 ( 
.A(n_314),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_782),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_549),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_680),
.Y(n_1136)
);

CKINVDCx20_ASAP7_75t_R g1137 ( 
.A(n_95),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_332),
.Y(n_1138)
);

CKINVDCx20_ASAP7_75t_R g1139 ( 
.A(n_241),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_587),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_732),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_771),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_173),
.Y(n_1143)
);

CKINVDCx20_ASAP7_75t_R g1144 ( 
.A(n_271),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_789),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_467),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_313),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_568),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_662),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_237),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_600),
.Y(n_1151)
);

INVxp67_ASAP7_75t_L g1152 ( 
.A(n_46),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_524),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_418),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_750),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_732),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_476),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_305),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_98),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_806),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_644),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_185),
.Y(n_1162)
);

INVx1_ASAP7_75t_SL g1163 ( 
.A(n_788),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_644),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_443),
.Y(n_1165)
);

BUFx3_ASAP7_75t_L g1166 ( 
.A(n_83),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_84),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_562),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_543),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_161),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_116),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_119),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_453),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_521),
.Y(n_1174)
);

INVx2_ASAP7_75t_SL g1175 ( 
.A(n_674),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_747),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_632),
.Y(n_1177)
);

CKINVDCx20_ASAP7_75t_R g1178 ( 
.A(n_385),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_322),
.Y(n_1179)
);

INVxp67_ASAP7_75t_SL g1180 ( 
.A(n_613),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_370),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_725),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_402),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_500),
.Y(n_1184)
);

CKINVDCx20_ASAP7_75t_R g1185 ( 
.A(n_313),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_601),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_111),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_734),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_550),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_805),
.Y(n_1190)
);

BUFx5_ASAP7_75t_L g1191 ( 
.A(n_27),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_716),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_110),
.Y(n_1193)
);

CKINVDCx20_ASAP7_75t_R g1194 ( 
.A(n_787),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_808),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_365),
.Y(n_1196)
);

HB1xp67_ASAP7_75t_L g1197 ( 
.A(n_446),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_592),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_589),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_217),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_390),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_5),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_773),
.Y(n_1203)
);

CKINVDCx16_ASAP7_75t_R g1204 ( 
.A(n_389),
.Y(n_1204)
);

CKINVDCx16_ASAP7_75t_R g1205 ( 
.A(n_9),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_398),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_406),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_797),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_630),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_141),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_282),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_302),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_399),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_319),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_167),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_599),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_809),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_338),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_802),
.Y(n_1219)
);

CKINVDCx16_ASAP7_75t_R g1220 ( 
.A(n_786),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_317),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_214),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_454),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_314),
.Y(n_1224)
);

CKINVDCx20_ASAP7_75t_R g1225 ( 
.A(n_397),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_456),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_208),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_285),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_246),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_328),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_114),
.Y(n_1231)
);

CKINVDCx20_ASAP7_75t_R g1232 ( 
.A(n_672),
.Y(n_1232)
);

CKINVDCx20_ASAP7_75t_R g1233 ( 
.A(n_803),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_789),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_473),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_472),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_568),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_108),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_147),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_443),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_764),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_547),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_458),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_121),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_745),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_100),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_574),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_697),
.Y(n_1248)
);

INVx2_ASAP7_75t_SL g1249 ( 
.A(n_186),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_649),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_807),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_197),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_492),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_357),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_414),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_246),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_179),
.Y(n_1257)
);

CKINVDCx16_ASAP7_75t_R g1258 ( 
.A(n_55),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_757),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_484),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_22),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_595),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_515),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_757),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_533),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_341),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_699),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_541),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_315),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_393),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_523),
.Y(n_1271)
);

BUFx10_ASAP7_75t_L g1272 ( 
.A(n_6),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_34),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_611),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_690),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_188),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_798),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_352),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_355),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_121),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_129),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_679),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_23),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_613),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_268),
.Y(n_1285)
);

INVx1_ASAP7_75t_SL g1286 ( 
.A(n_430),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_14),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_714),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_296),
.Y(n_1289)
);

INVxp67_ASAP7_75t_L g1290 ( 
.A(n_703),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_306),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_437),
.Y(n_1292)
);

BUFx5_ASAP7_75t_L g1293 ( 
.A(n_84),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_655),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_343),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1190),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_819),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_820),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1190),
.Y(n_1299)
);

INVxp67_ASAP7_75t_SL g1300 ( 
.A(n_858),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_820),
.Y(n_1301)
);

CKINVDCx20_ASAP7_75t_R g1302 ( 
.A(n_899),
.Y(n_1302)
);

NOR2xp67_ASAP7_75t_L g1303 ( 
.A(n_1190),
.B(n_0),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_858),
.Y(n_1304)
);

CKINVDCx20_ASAP7_75t_R g1305 ( 
.A(n_983),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_858),
.Y(n_1306)
);

INVxp67_ASAP7_75t_L g1307 ( 
.A(n_885),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_822),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1006),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_985),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_817),
.Y(n_1311)
);

CKINVDCx20_ASAP7_75t_R g1312 ( 
.A(n_905),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1124),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1077),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_924),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_924),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1030),
.B(n_0),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_822),
.Y(n_1318)
);

CKINVDCx20_ASAP7_75t_R g1319 ( 
.A(n_1204),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_826),
.Y(n_1320)
);

INVxp33_ASAP7_75t_SL g1321 ( 
.A(n_955),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_L g1322 ( 
.A(n_1153),
.B(n_0),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_826),
.Y(n_1323)
);

CKINVDCx20_ASAP7_75t_R g1324 ( 
.A(n_917),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_964),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_957),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1205),
.B(n_1),
.Y(n_1327)
);

INVxp67_ASAP7_75t_SL g1328 ( 
.A(n_921),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_828),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_957),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1214),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1214),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1249),
.Y(n_1333)
);

INVxp67_ASAP7_75t_SL g1334 ( 
.A(n_921),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1249),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_875),
.Y(n_1336)
);

INVxp67_ASAP7_75t_SL g1337 ( 
.A(n_1112),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1245),
.B(n_1),
.Y(n_1338)
);

CKINVDCx16_ASAP7_75t_R g1339 ( 
.A(n_1258),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_931),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_875),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_946),
.Y(n_1342)
);

BUFx6f_ASAP7_75t_SL g1343 ( 
.A(n_1040),
.Y(n_1343)
);

INVxp67_ASAP7_75t_L g1344 ( 
.A(n_1062),
.Y(n_1344)
);

CKINVDCx20_ASAP7_75t_R g1345 ( 
.A(n_986),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_828),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_836),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_964),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_992),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_992),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1039),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_997),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1197),
.B(n_1),
.Y(n_1353)
);

INVxp33_ASAP7_75t_SL g1354 ( 
.A(n_1282),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_839),
.B(n_2),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1039),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_839),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1097),
.Y(n_1358)
);

INVx1_ASAP7_75t_SL g1359 ( 
.A(n_840),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1097),
.Y(n_1360)
);

INVxp67_ASAP7_75t_SL g1361 ( 
.A(n_1112),
.Y(n_1361)
);

CKINVDCx14_ASAP7_75t_R g1362 ( 
.A(n_880),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_840),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_843),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_1084),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_843),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_846),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1175),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_846),
.Y(n_1369)
);

CKINVDCx20_ASAP7_75t_R g1370 ( 
.A(n_1137),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_1139),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_865),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1166),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_847),
.B(n_2),
.Y(n_1374)
);

BUFx3_ASAP7_75t_L g1375 ( 
.A(n_1166),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_831),
.B(n_3),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1175),
.Y(n_1377)
);

CKINVDCx20_ASAP7_75t_R g1378 ( 
.A(n_1144),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_824),
.Y(n_1379)
);

CKINVDCx20_ASAP7_75t_R g1380 ( 
.A(n_1178),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_825),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_849),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_849),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_830),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_850),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_832),
.B(n_3),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_850),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_964),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_852),
.Y(n_1389)
);

CKINVDCx20_ASAP7_75t_R g1390 ( 
.A(n_1185),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_852),
.Y(n_1391)
);

CKINVDCx20_ASAP7_75t_R g1392 ( 
.A(n_1225),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_842),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_853),
.Y(n_1394)
);

INVxp67_ASAP7_75t_L g1395 ( 
.A(n_1040),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_857),
.Y(n_1396)
);

CKINVDCx20_ASAP7_75t_R g1397 ( 
.A(n_1291),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_857),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_855),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_869),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_879),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_884),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_900),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_923),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_906),
.B(n_3),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_935),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_1290),
.B(n_4),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_939),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_1295),
.Y(n_1409)
);

CKINVDCx20_ASAP7_75t_R g1410 ( 
.A(n_987),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_861),
.B(n_4),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_864),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_864),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_951),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_956),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_960),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_871),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_871),
.Y(n_1418)
);

INVxp67_ASAP7_75t_SL g1419 ( 
.A(n_1183),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_972),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_874),
.Y(n_1421)
);

CKINVDCx20_ASAP7_75t_R g1422 ( 
.A(n_1092),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_981),
.Y(n_1423)
);

CKINVDCx20_ASAP7_75t_R g1424 ( 
.A(n_1220),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_874),
.B(n_4),
.Y(n_1425)
);

NOR2xp67_ASAP7_75t_L g1426 ( 
.A(n_1001),
.B(n_5),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_877),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_877),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1027),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1037),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1300),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1328),
.B(n_1191),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1307),
.B(n_1040),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1298),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_SL g1435 ( 
.A(n_1395),
.B(n_1191),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1315),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1336),
.B(n_1123),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1316),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1372),
.Y(n_1439)
);

INVx3_ASAP7_75t_L g1440 ( 
.A(n_1373),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1334),
.B(n_1191),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1326),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1330),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1337),
.B(n_1191),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1375),
.Y(n_1445)
);

OR2x6_ASAP7_75t_L g1446 ( 
.A(n_1327),
.B(n_821),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1344),
.B(n_878),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1309),
.B(n_925),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_1301),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1331),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1318),
.B(n_1088),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1361),
.B(n_1191),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_SL g1453 ( 
.A(n_1314),
.B(n_1191),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1332),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1419),
.B(n_1191),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1296),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1333),
.Y(n_1457)
);

BUFx6f_ASAP7_75t_L g1458 ( 
.A(n_1372),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1335),
.Y(n_1459)
);

INVx3_ASAP7_75t_L g1460 ( 
.A(n_1341),
.Y(n_1460)
);

INVxp67_ASAP7_75t_L g1461 ( 
.A(n_1367),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_1343),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1372),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1349),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1350),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1351),
.Y(n_1466)
);

BUFx6f_ASAP7_75t_L g1467 ( 
.A(n_1372),
.Y(n_1467)
);

NAND2xp33_ASAP7_75t_SL g1468 ( 
.A(n_1343),
.B(n_878),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1304),
.B(n_1191),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1356),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1299),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_SL g1472 ( 
.A(n_1359),
.B(n_1293),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1358),
.B(n_1123),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1360),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1306),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1368),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1325),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1383),
.B(n_1088),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1325),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1377),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1297),
.B(n_1293),
.Y(n_1481)
);

BUFx6f_ASAP7_75t_L g1482 ( 
.A(n_1348),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1379),
.Y(n_1483)
);

AND2x6_ASAP7_75t_L g1484 ( 
.A(n_1313),
.B(n_1183),
.Y(n_1484)
);

BUFx6f_ASAP7_75t_L g1485 ( 
.A(n_1348),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1381),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1303),
.B(n_925),
.Y(n_1487)
);

INVx6_ASAP7_75t_L g1488 ( 
.A(n_1339),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1308),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1384),
.B(n_1293),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1393),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1388),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1320),
.B(n_973),
.Y(n_1493)
);

BUFx6f_ASAP7_75t_L g1494 ( 
.A(n_1388),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1323),
.B(n_1293),
.Y(n_1495)
);

INVx3_ASAP7_75t_L g1496 ( 
.A(n_1394),
.Y(n_1496)
);

AND2x6_ASAP7_75t_L g1497 ( 
.A(n_1322),
.B(n_865),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1399),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1400),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_L g1500 ( 
.A(n_1430),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1329),
.B(n_973),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1401),
.Y(n_1502)
);

INVxp67_ASAP7_75t_L g1503 ( 
.A(n_1346),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1402),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1403),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1404),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1406),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1408),
.B(n_1293),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1414),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1429),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1347),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1415),
.Y(n_1512)
);

CKINVDCx20_ASAP7_75t_R g1513 ( 
.A(n_1340),
.Y(n_1513)
);

BUFx2_ASAP7_75t_L g1514 ( 
.A(n_1357),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1416),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1420),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1423),
.Y(n_1517)
);

AND2x2_ASAP7_75t_SL g1518 ( 
.A(n_1317),
.B(n_895),
.Y(n_1518)
);

CKINVDCx16_ASAP7_75t_R g1519 ( 
.A(n_1362),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1428),
.B(n_1293),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1426),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1363),
.B(n_982),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_1364),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1362),
.B(n_907),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1353),
.Y(n_1525)
);

INVx3_ASAP7_75t_L g1526 ( 
.A(n_1427),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1355),
.Y(n_1527)
);

BUFx6f_ASAP7_75t_L g1528 ( 
.A(n_1374),
.Y(n_1528)
);

CKINVDCx20_ASAP7_75t_R g1529 ( 
.A(n_1340),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1411),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1425),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_L g1532 ( 
.A(n_1376),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1366),
.B(n_1293),
.Y(n_1533)
);

BUFx6f_ASAP7_75t_L g1534 ( 
.A(n_1386),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1405),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1407),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1338),
.Y(n_1537)
);

NAND2xp33_ASAP7_75t_R g1538 ( 
.A(n_1369),
.B(n_887),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1382),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1385),
.B(n_1293),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1387),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_SL g1542 ( 
.A1(n_1342),
.A2(n_1352),
.B1(n_1365),
.B2(n_1345),
.Y(n_1542)
);

BUFx6f_ASAP7_75t_L g1543 ( 
.A(n_1389),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1391),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1396),
.Y(n_1545)
);

BUFx6f_ASAP7_75t_L g1546 ( 
.A(n_1398),
.Y(n_1546)
);

BUFx6f_ASAP7_75t_L g1547 ( 
.A(n_1412),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1413),
.B(n_1417),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1418),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1421),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_SL g1551 ( 
.A(n_1321),
.B(n_1113),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1302),
.B(n_1113),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1305),
.Y(n_1553)
);

OA21x2_ASAP7_75t_L g1554 ( 
.A1(n_1354),
.A2(n_886),
.B(n_837),
.Y(n_1554)
);

BUFx6f_ASAP7_75t_L g1555 ( 
.A(n_1305),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1310),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1310),
.Y(n_1557)
);

INVx4_ASAP7_75t_L g1558 ( 
.A(n_1319),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1319),
.B(n_1113),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1410),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_L g1561 ( 
.A(n_1422),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1422),
.B(n_964),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1424),
.B(n_1015),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1424),
.B(n_964),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1311),
.B(n_964),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_SL g1566 ( 
.A(n_1312),
.B(n_1120),
.Y(n_1566)
);

BUFx6f_ASAP7_75t_L g1567 ( 
.A(n_1409),
.Y(n_1567)
);

INVxp67_ASAP7_75t_L g1568 ( 
.A(n_1324),
.Y(n_1568)
);

INVxp67_ASAP7_75t_L g1569 ( 
.A(n_1397),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_1378),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1380),
.Y(n_1571)
);

INVx4_ASAP7_75t_L g1572 ( 
.A(n_1390),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1342),
.B(n_964),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1345),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1352),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1365),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1392),
.B(n_1120),
.Y(n_1577)
);

AOI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1370),
.A2(n_1283),
.B1(n_1285),
.B2(n_1281),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1392),
.B(n_1120),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1370),
.Y(n_1580)
);

BUFx6f_ASAP7_75t_L g1581 ( 
.A(n_1371),
.Y(n_1581)
);

INVx4_ASAP7_75t_L g1582 ( 
.A(n_1371),
.Y(n_1582)
);

INVxp67_ASAP7_75t_L g1583 ( 
.A(n_1318),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1373),
.Y(n_1584)
);

INVx3_ASAP7_75t_L g1585 ( 
.A(n_1373),
.Y(n_1585)
);

CKINVDCx20_ASAP7_75t_R g1586 ( 
.A(n_1340),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1300),
.B(n_964),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1300),
.Y(n_1588)
);

BUFx6f_ASAP7_75t_L g1589 ( 
.A(n_1372),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1307),
.B(n_887),
.Y(n_1590)
);

BUFx2_ASAP7_75t_L g1591 ( 
.A(n_1298),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1300),
.B(n_1012),
.Y(n_1592)
);

BUFx2_ASAP7_75t_L g1593 ( 
.A(n_1298),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1300),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1300),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1300),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1373),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1300),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1300),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1300),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1373),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1300),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1300),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_SL g1604 ( 
.A(n_1343),
.B(n_1133),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1300),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1300),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_SL g1607 ( 
.A(n_1343),
.B(n_1133),
.Y(n_1607)
);

INVx4_ASAP7_75t_L g1608 ( 
.A(n_1343),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1343),
.Y(n_1609)
);

BUFx6f_ASAP7_75t_L g1610 ( 
.A(n_1372),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1309),
.B(n_1015),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_SL g1612 ( 
.A(n_1395),
.B(n_1133),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1300),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1300),
.B(n_1012),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1300),
.B(n_1012),
.Y(n_1615)
);

BUFx6f_ASAP7_75t_L g1616 ( 
.A(n_1372),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1300),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1309),
.B(n_1041),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1372),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1373),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1318),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1307),
.B(n_1272),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1300),
.Y(n_1623)
);

INVxp67_ASAP7_75t_L g1624 ( 
.A(n_1318),
.Y(n_1624)
);

INVx3_ASAP7_75t_L g1625 ( 
.A(n_1373),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1300),
.Y(n_1626)
);

BUFx8_ASAP7_75t_L g1627 ( 
.A(n_1343),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1307),
.B(n_1272),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1373),
.Y(n_1629)
);

BUFx6f_ASAP7_75t_L g1630 ( 
.A(n_1372),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1300),
.Y(n_1631)
);

AND2x6_ASAP7_75t_L g1632 ( 
.A(n_1314),
.B(n_865),
.Y(n_1632)
);

BUFx6f_ASAP7_75t_L g1633 ( 
.A(n_1372),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1300),
.Y(n_1634)
);

BUFx6f_ASAP7_75t_L g1635 ( 
.A(n_1372),
.Y(n_1635)
);

AOI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1327),
.A2(n_1287),
.B1(n_889),
.B2(n_1050),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1300),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1300),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1373),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1307),
.B(n_1272),
.Y(n_1640)
);

BUFx4f_ASAP7_75t_L g1641 ( 
.A(n_1488),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1440),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1440),
.Y(n_1643)
);

BUFx2_ASAP7_75t_L g1644 ( 
.A(n_1449),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1531),
.A2(n_1527),
.B1(n_1530),
.B2(n_1626),
.Y(n_1645)
);

OAI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1636),
.A2(n_892),
.B1(n_1050),
.B2(n_889),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1460),
.Y(n_1647)
);

INVx4_ASAP7_75t_L g1648 ( 
.A(n_1608),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_L g1649 ( 
.A(n_1535),
.B(n_1152),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1447),
.B(n_892),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1536),
.B(n_1055),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1585),
.Y(n_1652)
);

NAND2xp33_ASAP7_75t_L g1653 ( 
.A(n_1484),
.B(n_1012),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1460),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1466),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1585),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1625),
.Y(n_1657)
);

BUFx3_ASAP7_75t_L g1658 ( 
.A(n_1627),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1525),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1625),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1496),
.B(n_1509),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1604),
.B(n_1055),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1461),
.B(n_1238),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1466),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1496),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1445),
.Y(n_1666)
);

BUFx6f_ASAP7_75t_SL g1667 ( 
.A(n_1558),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1604),
.B(n_1238),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1509),
.Y(n_1669)
);

NOR2x1p5_ASAP7_75t_L g1670 ( 
.A(n_1608),
.B(n_1558),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1512),
.Y(n_1671)
);

INVx5_ASAP7_75t_L g1672 ( 
.A(n_1632),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1512),
.Y(n_1673)
);

INVx1_ASAP7_75t_SL g1674 ( 
.A(n_1590),
.Y(n_1674)
);

INVx3_ASAP7_75t_L g1675 ( 
.A(n_1528),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1436),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1461),
.B(n_1256),
.Y(n_1677)
);

BUFx2_ASAP7_75t_L g1678 ( 
.A(n_1514),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1438),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1442),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1578),
.B(n_1276),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_SL g1682 ( 
.A(n_1607),
.B(n_1256),
.Y(n_1682)
);

INVx6_ASAP7_75t_L g1683 ( 
.A(n_1627),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1483),
.B(n_1257),
.Y(n_1684)
);

AND2x6_ASAP7_75t_L g1685 ( 
.A(n_1451),
.B(n_837),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1443),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1450),
.Y(n_1687)
);

INVxp33_ASAP7_75t_L g1688 ( 
.A(n_1577),
.Y(n_1688)
);

INVx1_ASAP7_75t_SL g1689 ( 
.A(n_1591),
.Y(n_1689)
);

INVx3_ASAP7_75t_L g1690 ( 
.A(n_1528),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1584),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1454),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1457),
.Y(n_1693)
);

INVxp67_ASAP7_75t_SL g1694 ( 
.A(n_1432),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1597),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1537),
.B(n_1257),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1554),
.A2(n_1049),
.B1(n_1051),
.B2(n_1042),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1459),
.Y(n_1698)
);

INVx6_ASAP7_75t_L g1699 ( 
.A(n_1528),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_SL g1700 ( 
.A(n_1607),
.B(n_1261),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1554),
.A2(n_1059),
.B1(n_1082),
.B2(n_1052),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_SL g1702 ( 
.A(n_1525),
.B(n_1261),
.Y(n_1702)
);

INVx3_ASAP7_75t_L g1703 ( 
.A(n_1500),
.Y(n_1703)
);

BUFx6f_ASAP7_75t_SL g1704 ( 
.A(n_1556),
.Y(n_1704)
);

NOR2x1p5_ASAP7_75t_L g1705 ( 
.A(n_1462),
.B(n_1278),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_SL g1706 ( 
.A(n_1525),
.B(n_1270),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1601),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1464),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1465),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1620),
.Y(n_1710)
);

NAND2xp33_ASAP7_75t_L g1711 ( 
.A(n_1484),
.B(n_1012),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1470),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1474),
.Y(n_1713)
);

INVx2_ASAP7_75t_SL g1714 ( 
.A(n_1478),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1612),
.B(n_1270),
.Y(n_1715)
);

INVx3_ASAP7_75t_L g1716 ( 
.A(n_1500),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1486),
.B(n_1281),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1476),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1491),
.B(n_1283),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1431),
.A2(n_1094),
.B1(n_1101),
.B2(n_1093),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1583),
.B(n_1279),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1480),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1532),
.B(n_1279),
.Y(n_1723)
);

INVx3_ASAP7_75t_L g1724 ( 
.A(n_1500),
.Y(n_1724)
);

BUFx4f_ASAP7_75t_L g1725 ( 
.A(n_1488),
.Y(n_1725)
);

INVxp33_ASAP7_75t_SL g1726 ( 
.A(n_1578),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1456),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1532),
.B(n_1285),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1629),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1471),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1499),
.B(n_1287),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1433),
.A2(n_909),
.B1(n_910),
.B2(n_903),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_L g1733 ( 
.A(n_1588),
.B(n_916),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_SL g1734 ( 
.A(n_1532),
.B(n_886),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1639),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1475),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1441),
.Y(n_1737)
);

INVxp33_ASAP7_75t_L g1738 ( 
.A(n_1579),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1441),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1583),
.B(n_1000),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1505),
.B(n_1012),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1506),
.B(n_1012),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1510),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1444),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1510),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1594),
.B(n_927),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1444),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1510),
.Y(n_1748)
);

OR2x6_ASAP7_75t_L g1749 ( 
.A(n_1446),
.B(n_974),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1452),
.Y(n_1750)
);

NOR3xp33_ASAP7_75t_L g1751 ( 
.A(n_1573),
.B(n_901),
.C(n_818),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_L g1752 ( 
.A1(n_1595),
.A2(n_1118),
.B1(n_1119),
.B2(n_1105),
.Y(n_1752)
);

INVx4_ASAP7_75t_L g1753 ( 
.A(n_1484),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1452),
.Y(n_1754)
);

OR2x6_ASAP7_75t_L g1755 ( 
.A(n_1446),
.B(n_895),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1477),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1455),
.Y(n_1757)
);

NOR3xp33_ASAP7_75t_L g1758 ( 
.A(n_1573),
.B(n_1087),
.C(n_947),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1580),
.B(n_829),
.Y(n_1759)
);

INVx2_ASAP7_75t_SL g1760 ( 
.A(n_1622),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_SL g1761 ( 
.A(n_1534),
.B(n_894),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_SL g1762 ( 
.A(n_1534),
.B(n_894),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1628),
.A2(n_938),
.B1(n_944),
.B2(n_932),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1455),
.Y(n_1764)
);

INVx4_ASAP7_75t_L g1765 ( 
.A(n_1484),
.Y(n_1765)
);

INVx2_ASAP7_75t_SL g1766 ( 
.A(n_1640),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1517),
.B(n_1012),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1596),
.B(n_949),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1621),
.B(n_1000),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1621),
.B(n_1000),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1598),
.A2(n_1147),
.B1(n_1158),
.B2(n_1143),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1599),
.B(n_953),
.Y(n_1772)
);

INVx3_ASAP7_75t_L g1773 ( 
.A(n_1487),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_SL g1774 ( 
.A(n_1534),
.B(n_912),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1600),
.B(n_954),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1602),
.B(n_961),
.Y(n_1776)
);

INVx5_ASAP7_75t_L g1777 ( 
.A(n_1632),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1603),
.B(n_963),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_SL g1779 ( 
.A1(n_1518),
.A2(n_883),
.B1(n_959),
.B2(n_844),
.Y(n_1779)
);

NOR2xp33_ASAP7_75t_L g1780 ( 
.A(n_1605),
.B(n_968),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1606),
.B(n_970),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1613),
.B(n_977),
.Y(n_1782)
);

BUFx10_ASAP7_75t_L g1783 ( 
.A(n_1609),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1617),
.B(n_978),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1623),
.B(n_1631),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1634),
.B(n_990),
.Y(n_1786)
);

BUFx6f_ASAP7_75t_SL g1787 ( 
.A(n_1572),
.Y(n_1787)
);

BUFx6f_ASAP7_75t_L g1788 ( 
.A(n_1632),
.Y(n_1788)
);

AND2x6_ASAP7_75t_L g1789 ( 
.A(n_1523),
.B(n_912),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1477),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1477),
.Y(n_1791)
);

XOR2x2_ASAP7_75t_SL g1792 ( 
.A(n_1636),
.B(n_1075),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_SL g1793 ( 
.A(n_1548),
.B(n_1010),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1482),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1637),
.Y(n_1795)
);

INVx2_ASAP7_75t_SL g1796 ( 
.A(n_1493),
.Y(n_1796)
);

INVx2_ASAP7_75t_SL g1797 ( 
.A(n_1493),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1638),
.Y(n_1798)
);

INVx3_ASAP7_75t_L g1799 ( 
.A(n_1487),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_SL g1800 ( 
.A(n_1548),
.B(n_1010),
.Y(n_1800)
);

AOI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1624),
.A2(n_1008),
.B1(n_1014),
.B2(n_1007),
.Y(n_1801)
);

NAND2xp33_ASAP7_75t_L g1802 ( 
.A(n_1497),
.B(n_865),
.Y(n_1802)
);

INVx1_ASAP7_75t_SL g1803 ( 
.A(n_1593),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1587),
.Y(n_1804)
);

INVx5_ASAP7_75t_L g1805 ( 
.A(n_1632),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1592),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1520),
.B(n_1016),
.Y(n_1807)
);

AOI22xp33_ASAP7_75t_L g1808 ( 
.A1(n_1498),
.A2(n_1167),
.B1(n_1171),
.B2(n_1159),
.Y(n_1808)
);

INVx4_ASAP7_75t_L g1809 ( 
.A(n_1523),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1502),
.A2(n_1196),
.B1(n_1200),
.B2(n_1193),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1482),
.Y(n_1811)
);

INVx4_ASAP7_75t_L g1812 ( 
.A(n_1526),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1482),
.Y(n_1813)
);

OR2x6_ASAP7_75t_L g1814 ( 
.A(n_1446),
.B(n_897),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1592),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1624),
.B(n_1070),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1614),
.Y(n_1817)
);

BUFx2_ASAP7_75t_L g1818 ( 
.A(n_1503),
.Y(n_1818)
);

BUFx2_ASAP7_75t_L g1819 ( 
.A(n_1503),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1614),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_SL g1821 ( 
.A(n_1497),
.B(n_1021),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1520),
.B(n_1023),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1615),
.Y(n_1823)
);

INVx2_ASAP7_75t_SL g1824 ( 
.A(n_1501),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1533),
.B(n_1540),
.Y(n_1825)
);

AND2x6_ASAP7_75t_L g1826 ( 
.A(n_1526),
.B(n_1045),
.Y(n_1826)
);

INVx2_ASAP7_75t_SL g1827 ( 
.A(n_1501),
.Y(n_1827)
);

NOR2xp33_ASAP7_75t_L g1828 ( 
.A(n_1524),
.B(n_1539),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1615),
.Y(n_1829)
);

NAND2xp33_ASAP7_75t_L g1830 ( 
.A(n_1497),
.B(n_865),
.Y(n_1830)
);

CKINVDCx20_ASAP7_75t_R g1831 ( 
.A(n_1513),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_SL g1832 ( 
.A(n_1541),
.B(n_1045),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1485),
.Y(n_1833)
);

BUFx3_ASAP7_75t_L g1834 ( 
.A(n_1543),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1580),
.B(n_1552),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1533),
.B(n_1022),
.Y(n_1836)
);

NOR3xp33_ASAP7_75t_L g1837 ( 
.A(n_1565),
.B(n_1029),
.C(n_1024),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1469),
.Y(n_1838)
);

BUFx6f_ASAP7_75t_L g1839 ( 
.A(n_1485),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1469),
.Y(n_1840)
);

INVxp67_ASAP7_75t_SL g1841 ( 
.A(n_1490),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1485),
.Y(n_1842)
);

CKINVDCx20_ASAP7_75t_R g1843 ( 
.A(n_1529),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1504),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_1586),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1507),
.Y(n_1846)
);

INVx3_ASAP7_75t_L g1847 ( 
.A(n_1515),
.Y(n_1847)
);

INVxp33_ASAP7_75t_L g1848 ( 
.A(n_1555),
.Y(n_1848)
);

INVxp67_ASAP7_75t_SL g1849 ( 
.A(n_1490),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1516),
.Y(n_1850)
);

BUFx2_ASAP7_75t_L g1851 ( 
.A(n_1434),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1508),
.Y(n_1852)
);

AOI22xp5_ASAP7_75t_SL g1853 ( 
.A1(n_1582),
.A2(n_1134),
.B1(n_1194),
.B2(n_1099),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1494),
.Y(n_1854)
);

BUFx2_ASAP7_75t_L g1855 ( 
.A(n_1489),
.Y(n_1855)
);

OAI21xp33_ASAP7_75t_SL g1856 ( 
.A1(n_1540),
.A2(n_1521),
.B(n_1453),
.Y(n_1856)
);

BUFx6f_ASAP7_75t_L g1857 ( 
.A(n_1494),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1511),
.B(n_1070),
.Y(n_1858)
);

INVx2_ASAP7_75t_SL g1859 ( 
.A(n_1522),
.Y(n_1859)
);

BUFx3_ASAP7_75t_L g1860 ( 
.A(n_1543),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1550),
.B(n_1070),
.Y(n_1861)
);

INVx4_ASAP7_75t_SL g1862 ( 
.A(n_1497),
.Y(n_1862)
);

AO22x2_ASAP7_75t_L g1863 ( 
.A1(n_1563),
.A2(n_1180),
.B1(n_823),
.B2(n_827),
.Y(n_1863)
);

INVx4_ASAP7_75t_L g1864 ( 
.A(n_1550),
.Y(n_1864)
);

BUFx4f_ASAP7_75t_L g1865 ( 
.A(n_1543),
.Y(n_1865)
);

CKINVDCx5p33_ASAP7_75t_R g1866 ( 
.A(n_1538),
.Y(n_1866)
);

AOI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1551),
.A2(n_1034),
.B1(n_1035),
.B2(n_1032),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1522),
.Y(n_1868)
);

INVx1_ASAP7_75t_SL g1869 ( 
.A(n_1563),
.Y(n_1869)
);

INVx3_ASAP7_75t_L g1870 ( 
.A(n_1448),
.Y(n_1870)
);

INVx3_ASAP7_75t_L g1871 ( 
.A(n_1448),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1508),
.B(n_1043),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1437),
.B(n_1044),
.Y(n_1873)
);

AND2x6_ASAP7_75t_L g1874 ( 
.A(n_1546),
.B(n_1116),
.Y(n_1874)
);

INVx3_ASAP7_75t_L g1875 ( 
.A(n_1611),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1611),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1544),
.B(n_1056),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1618),
.Y(n_1878)
);

INVx3_ASAP7_75t_L g1879 ( 
.A(n_1618),
.Y(n_1879)
);

AND2x6_ASAP7_75t_L g1880 ( 
.A(n_1546),
.B(n_1547),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1562),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1479),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1545),
.B(n_1057),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1492),
.Y(n_1884)
);

BUFx10_ASAP7_75t_L g1885 ( 
.A(n_1473),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1435),
.B(n_1072),
.Y(n_1886)
);

NAND2xp33_ASAP7_75t_R g1887 ( 
.A(n_1570),
.B(n_829),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_SL g1888 ( 
.A(n_1549),
.B(n_1116),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_1542),
.Y(n_1889)
);

NOR2xp33_ASAP7_75t_SL g1890 ( 
.A(n_1519),
.B(n_1073),
.Y(n_1890)
);

INVx4_ASAP7_75t_L g1891 ( 
.A(n_1547),
.Y(n_1891)
);

INVx4_ASAP7_75t_L g1892 ( 
.A(n_1547),
.Y(n_1892)
);

NOR2xp33_ASAP7_75t_L g1893 ( 
.A(n_1481),
.B(n_1074),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_SL g1894 ( 
.A(n_1468),
.B(n_1172),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1565),
.B(n_1098),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1562),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1472),
.Y(n_1897)
);

AOI22xp33_ASAP7_75t_L g1898 ( 
.A1(n_1564),
.A2(n_1212),
.B1(n_1222),
.B2(n_1218),
.Y(n_1898)
);

INVx3_ASAP7_75t_L g1899 ( 
.A(n_1439),
.Y(n_1899)
);

INVx2_ASAP7_75t_SL g1900 ( 
.A(n_1555),
.Y(n_1900)
);

AOI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1559),
.A2(n_1081),
.B1(n_1086),
.B2(n_1080),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1495),
.B(n_1095),
.Y(n_1902)
);

OR2x6_ASAP7_75t_L g1903 ( 
.A(n_1555),
.B(n_897),
.Y(n_1903)
);

INVx4_ASAP7_75t_L g1904 ( 
.A(n_1561),
.Y(n_1904)
);

INVx2_ASAP7_75t_SL g1905 ( 
.A(n_1561),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1566),
.B(n_1098),
.Y(n_1906)
);

BUFx10_ASAP7_75t_L g1907 ( 
.A(n_1560),
.Y(n_1907)
);

INVx3_ASAP7_75t_L g1908 ( 
.A(n_1458),
.Y(n_1908)
);

AND2x4_ASAP7_75t_L g1909 ( 
.A(n_1553),
.B(n_1041),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1458),
.Y(n_1910)
);

AOI22xp33_ASAP7_75t_L g1911 ( 
.A1(n_1557),
.A2(n_1224),
.B1(n_1244),
.B2(n_1239),
.Y(n_1911)
);

AOI21x1_ASAP7_75t_L g1912 ( 
.A1(n_1463),
.A2(n_1252),
.B(n_1246),
.Y(n_1912)
);

OR2x6_ASAP7_75t_L g1913 ( 
.A(n_1572),
.B(n_967),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_1542),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_L g1915 ( 
.A(n_1561),
.B(n_1096),
.Y(n_1915)
);

BUFx3_ASAP7_75t_L g1916 ( 
.A(n_1567),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_SL g1917 ( 
.A(n_1582),
.B(n_1221),
.Y(n_1917)
);

NAND3xp33_ASAP7_75t_L g1918 ( 
.A(n_1463),
.B(n_1108),
.C(n_1104),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1463),
.Y(n_1919)
);

NOR2xp33_ASAP7_75t_L g1920 ( 
.A(n_1674),
.B(n_1575),
.Y(n_1920)
);

AOI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1674),
.A2(n_1121),
.B1(n_1125),
.B2(n_1110),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1694),
.B(n_1127),
.Y(n_1922)
);

AND2x2_ASAP7_75t_SL g1923 ( 
.A(n_1890),
.B(n_1567),
.Y(n_1923)
);

BUFx6f_ASAP7_75t_L g1924 ( 
.A(n_1788),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1675),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1694),
.B(n_1841),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_SL g1927 ( 
.A(n_1753),
.B(n_1170),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1661),
.Y(n_1928)
);

NOR2xp33_ASAP7_75t_L g1929 ( 
.A(n_1760),
.B(n_1568),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1841),
.B(n_1201),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_SL g1931 ( 
.A(n_1753),
.B(n_1202),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1849),
.B(n_1215),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1690),
.Y(n_1933)
);

AOI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1751),
.A2(n_1107),
.B1(n_1265),
.B2(n_1046),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_SL g1935 ( 
.A(n_1765),
.B(n_1230),
.Y(n_1935)
);

NOR2xp67_ASAP7_75t_L g1936 ( 
.A(n_1658),
.B(n_1568),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_SL g1937 ( 
.A(n_1765),
.B(n_1231),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1849),
.B(n_1130),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1804),
.B(n_1138),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_L g1940 ( 
.A(n_1766),
.B(n_1569),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1689),
.B(n_1581),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1661),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1714),
.B(n_1571),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1659),
.Y(n_1944)
);

NOR2xp33_ASAP7_75t_L g1945 ( 
.A(n_1688),
.B(n_1574),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1738),
.B(n_1576),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_SL g1947 ( 
.A(n_1809),
.B(n_1150),
.Y(n_1947)
);

BUFx8_ASAP7_75t_L g1948 ( 
.A(n_1667),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_L g1949 ( 
.A(n_1650),
.B(n_1581),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1659),
.Y(n_1950)
);

AOI22xp33_ASAP7_75t_L g1951 ( 
.A1(n_1758),
.A2(n_1275),
.B1(n_1181),
.B2(n_1187),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1795),
.Y(n_1952)
);

O2A1O1Ixp33_ASAP7_75t_L g1953 ( 
.A1(n_1646),
.A2(n_1269),
.B(n_1280),
.C(n_1254),
.Y(n_1953)
);

BUFx10_ASAP7_75t_L g1954 ( 
.A(n_1683),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1806),
.B(n_1179),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_SL g1956 ( 
.A(n_1809),
.B(n_1206),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1645),
.B(n_1207),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1647),
.Y(n_1958)
);

HB1xp67_ASAP7_75t_L g1959 ( 
.A(n_1689),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1645),
.B(n_1210),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1684),
.B(n_1211),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1684),
.B(n_1213),
.Y(n_1962)
);

INVx2_ASAP7_75t_SL g1963 ( 
.A(n_1803),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1654),
.Y(n_1964)
);

AOI22xp5_ASAP7_75t_L g1965 ( 
.A1(n_1663),
.A2(n_1228),
.B1(n_1229),
.B2(n_1227),
.Y(n_1965)
);

INVx3_ASAP7_75t_L g1966 ( 
.A(n_1699),
.Y(n_1966)
);

O2A1O1Ixp5_ASAP7_75t_L g1967 ( 
.A1(n_1793),
.A2(n_1289),
.B(n_993),
.C(n_1011),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1717),
.B(n_835),
.Y(n_1968)
);

NAND2xp33_ASAP7_75t_L g1969 ( 
.A(n_1789),
.B(n_835),
.Y(n_1969)
);

INVx2_ASAP7_75t_SL g1970 ( 
.A(n_1803),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1717),
.B(n_1719),
.Y(n_1971)
);

INVxp67_ASAP7_75t_L g1972 ( 
.A(n_1644),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1719),
.B(n_838),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1677),
.B(n_1581),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1731),
.B(n_838),
.Y(n_1975)
);

BUFx6f_ASAP7_75t_L g1976 ( 
.A(n_1788),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_L g1977 ( 
.A(n_1721),
.B(n_1567),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_SL g1978 ( 
.A(n_1812),
.B(n_841),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1798),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_SL g1980 ( 
.A(n_1812),
.B(n_841),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_SL g1981 ( 
.A(n_1864),
.B(n_1818),
.Y(n_1981)
);

NAND3xp33_ASAP7_75t_L g1982 ( 
.A(n_1758),
.B(n_1292),
.C(n_1284),
.Y(n_1982)
);

BUFx3_ASAP7_75t_L g1983 ( 
.A(n_1683),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1676),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1679),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1788),
.Y(n_1986)
);

OAI22xp5_ASAP7_75t_L g1987 ( 
.A1(n_1697),
.A2(n_1701),
.B1(n_1771),
.B2(n_1898),
.Y(n_1987)
);

HB1xp67_ASAP7_75t_L g1988 ( 
.A(n_1678),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1680),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_SL g1990 ( 
.A(n_1864),
.B(n_845),
.Y(n_1990)
);

BUFx6f_ASAP7_75t_L g1991 ( 
.A(n_1672),
.Y(n_1991)
);

AOI22xp33_ASAP7_75t_L g1992 ( 
.A1(n_1837),
.A2(n_1275),
.B1(n_1033),
.B2(n_1064),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_SL g1993 ( 
.A(n_1819),
.B(n_845),
.Y(n_1993)
);

INVx3_ASAP7_75t_L g1994 ( 
.A(n_1699),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1686),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1655),
.Y(n_1996)
);

BUFx8_ASAP7_75t_L g1997 ( 
.A(n_1667),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1687),
.Y(n_1998)
);

NOR2xp33_ASAP7_75t_L g1999 ( 
.A(n_1740),
.B(n_1069),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1731),
.B(n_848),
.Y(n_2000)
);

INVx2_ASAP7_75t_SL g2001 ( 
.A(n_1851),
.Y(n_2001)
);

CKINVDCx5p33_ASAP7_75t_R g2002 ( 
.A(n_1831),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1815),
.B(n_848),
.Y(n_2003)
);

BUFx5_ASAP7_75t_L g2004 ( 
.A(n_1880),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_L g2005 ( 
.A(n_1769),
.B(n_851),
.Y(n_2005)
);

INVxp67_ASAP7_75t_L g2006 ( 
.A(n_1855),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1817),
.B(n_851),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_L g2008 ( 
.A(n_1770),
.B(n_856),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_SL g2009 ( 
.A(n_1821),
.B(n_856),
.Y(n_2009)
);

NOR2xp33_ASAP7_75t_L g2010 ( 
.A(n_1816),
.B(n_859),
.Y(n_2010)
);

INVxp67_ASAP7_75t_L g2011 ( 
.A(n_1890),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1664),
.Y(n_2012)
);

AND2x2_ASAP7_75t_SL g2013 ( 
.A(n_1641),
.B(n_1232),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1692),
.Y(n_2014)
);

NAND2xp33_ASAP7_75t_L g2015 ( 
.A(n_1789),
.B(n_859),
.Y(n_2015)
);

A2O1A1Ixp33_ASAP7_75t_L g2016 ( 
.A1(n_1651),
.A2(n_833),
.B(n_834),
.C(n_814),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1820),
.B(n_860),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1665),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1693),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_SL g2020 ( 
.A(n_1821),
.B(n_860),
.Y(n_2020)
);

NOR2xp67_ASAP7_75t_L g2021 ( 
.A(n_1646),
.B(n_5),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1823),
.B(n_866),
.Y(n_2022)
);

NOR2xp33_ASAP7_75t_L g2023 ( 
.A(n_1858),
.B(n_866),
.Y(n_2023)
);

INVx2_ASAP7_75t_SL g2024 ( 
.A(n_1641),
.Y(n_2024)
);

BUFx8_ASAP7_75t_L g2025 ( 
.A(n_1787),
.Y(n_2025)
);

BUFx2_ASAP7_75t_L g2026 ( 
.A(n_1755),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1698),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1708),
.Y(n_2028)
);

OAI221xp5_ASAP7_75t_L g2029 ( 
.A1(n_1779),
.A2(n_867),
.B1(n_881),
.B2(n_876),
.C(n_872),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1669),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1829),
.B(n_867),
.Y(n_2031)
);

OAI22xp5_ASAP7_75t_L g2032 ( 
.A1(n_1771),
.A2(n_862),
.B1(n_863),
.B2(n_854),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1681),
.B(n_1779),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1709),
.Y(n_2034)
);

AOI22xp33_ASAP7_75t_L g2035 ( 
.A1(n_1837),
.A2(n_1033),
.B1(n_1064),
.B2(n_966),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1737),
.B(n_1292),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_SL g2037 ( 
.A(n_1872),
.B(n_1852),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_SL g2038 ( 
.A(n_1872),
.B(n_872),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_SL g2039 ( 
.A(n_1739),
.B(n_876),
.Y(n_2039)
);

AOI22xp5_ASAP7_75t_L g2040 ( 
.A1(n_1685),
.A2(n_882),
.B1(n_888),
.B2(n_881),
.Y(n_2040)
);

BUFx3_ASAP7_75t_L g2041 ( 
.A(n_1683),
.Y(n_2041)
);

NOR2xp33_ASAP7_75t_SL g2042 ( 
.A(n_1672),
.B(n_1233),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1671),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1712),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1673),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1744),
.B(n_882),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1747),
.B(n_888),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_1750),
.B(n_1754),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1847),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1757),
.B(n_891),
.Y(n_2050)
);

INVx2_ASAP7_75t_SL g2051 ( 
.A(n_1725),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1764),
.B(n_891),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1713),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_SL g2054 ( 
.A(n_1838),
.B(n_1053),
.Y(n_2054)
);

OAI22xp33_ASAP7_75t_L g2055 ( 
.A1(n_1726),
.A2(n_1255),
.B1(n_1234),
.B2(n_1235),
.Y(n_2055)
);

NOR2xp67_ASAP7_75t_L g2056 ( 
.A(n_1648),
.B(n_6),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1847),
.Y(n_2057)
);

AND2x4_ASAP7_75t_SL g2058 ( 
.A(n_1648),
.B(n_1098),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_SL g2059 ( 
.A(n_1840),
.B(n_1053),
.Y(n_2059)
);

NOR2xp33_ASAP7_75t_L g2060 ( 
.A(n_1732),
.B(n_1234),
.Y(n_2060)
);

NOR3xp33_ASAP7_75t_L g2061 ( 
.A(n_1835),
.B(n_1017),
.C(n_893),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1696),
.B(n_1768),
.Y(n_2062)
);

NOR2xp33_ASAP7_75t_L g2063 ( 
.A(n_1763),
.B(n_1235),
.Y(n_2063)
);

OAI22xp5_ASAP7_75t_L g2064 ( 
.A1(n_1881),
.A2(n_870),
.B1(n_873),
.B2(n_868),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1768),
.B(n_1236),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_SL g2066 ( 
.A(n_1896),
.B(n_1236),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1772),
.B(n_1240),
.Y(n_2067)
);

OR2x2_ASAP7_75t_L g2068 ( 
.A(n_1759),
.B(n_1294),
.Y(n_2068)
);

AOI22xp33_ASAP7_75t_L g2069 ( 
.A1(n_1685),
.A2(n_1033),
.B1(n_1064),
.B2(n_966),
.Y(n_2069)
);

BUFx3_ASAP7_75t_L g2070 ( 
.A(n_1916),
.Y(n_2070)
);

INVx1_ASAP7_75t_SL g2071 ( 
.A(n_1699),
.Y(n_2071)
);

NOR2x1p5_ASAP7_75t_L g2072 ( 
.A(n_1866),
.B(n_1241),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1718),
.Y(n_2073)
);

OR2x6_ASAP7_75t_L g2074 ( 
.A(n_1749),
.B(n_1755),
.Y(n_2074)
);

INVx2_ASAP7_75t_SL g2075 ( 
.A(n_1725),
.Y(n_2075)
);

OR2x6_ASAP7_75t_L g2076 ( 
.A(n_1749),
.B(n_967),
.Y(n_2076)
);

AOI21xp5_ASAP7_75t_L g2077 ( 
.A1(n_1825),
.A2(n_1589),
.B(n_1467),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_1825),
.B(n_1241),
.Y(n_2078)
);

INVx2_ASAP7_75t_SL g2079 ( 
.A(n_1907),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1722),
.Y(n_2080)
);

NOR3xp33_ASAP7_75t_L g2081 ( 
.A(n_1889),
.B(n_1102),
.C(n_1048),
.Y(n_2081)
);

OAI22xp5_ASAP7_75t_L g2082 ( 
.A1(n_1911),
.A2(n_902),
.B1(n_911),
.B2(n_890),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_1775),
.B(n_1274),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_1863),
.B(n_1242),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1785),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1666),
.Y(n_2086)
);

INVx2_ASAP7_75t_SL g2087 ( 
.A(n_1907),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1775),
.B(n_1274),
.Y(n_2088)
);

INVx2_ASAP7_75t_SL g2089 ( 
.A(n_1913),
.Y(n_2089)
);

NOR2xp33_ASAP7_75t_L g2090 ( 
.A(n_1828),
.B(n_1873),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1785),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1691),
.Y(n_2092)
);

NAND2xp33_ASAP7_75t_L g2093 ( 
.A(n_1789),
.B(n_1826),
.Y(n_2093)
);

INVx2_ASAP7_75t_SL g2094 ( 
.A(n_1913),
.Y(n_2094)
);

NOR2xp67_ASAP7_75t_L g2095 ( 
.A(n_1901),
.B(n_1801),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_1863),
.B(n_1242),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_SL g2097 ( 
.A(n_1776),
.B(n_1248),
.Y(n_2097)
);

AOI22xp5_ASAP7_75t_L g2098 ( 
.A1(n_1685),
.A2(n_1250),
.B1(n_1251),
.B2(n_1248),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_SL g2099 ( 
.A(n_1776),
.B(n_1250),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1876),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1778),
.B(n_1294),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1878),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1870),
.Y(n_2103)
);

INVx2_ASAP7_75t_SL g2104 ( 
.A(n_1913),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1784),
.B(n_1253),
.Y(n_2105)
);

INVx5_ASAP7_75t_L g2106 ( 
.A(n_1789),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1870),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_1784),
.B(n_1253),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1786),
.B(n_1259),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_SL g2110 ( 
.A(n_1786),
.B(n_1259),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1871),
.Y(n_2111)
);

OR2x6_ASAP7_75t_L g2112 ( 
.A(n_1749),
.B(n_993),
.Y(n_2112)
);

NOR2xp67_ASAP7_75t_L g2113 ( 
.A(n_1867),
.B(n_6),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1871),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1695),
.Y(n_2115)
);

INVx2_ASAP7_75t_SL g2116 ( 
.A(n_1865),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_SL g2117 ( 
.A(n_1807),
.B(n_1260),
.Y(n_2117)
);

NOR2xp33_ASAP7_75t_SL g2118 ( 
.A(n_1672),
.B(n_1260),
.Y(n_2118)
);

AND2x4_ASAP7_75t_L g2119 ( 
.A(n_1670),
.B(n_918),
.Y(n_2119)
);

AOI22xp5_ASAP7_75t_L g2120 ( 
.A1(n_1685),
.A2(n_1264),
.B1(n_1267),
.B2(n_1262),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1875),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_1863),
.B(n_1262),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1807),
.B(n_1264),
.Y(n_2123)
);

NOR2xp33_ASAP7_75t_L g2124 ( 
.A(n_1873),
.B(n_1869),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1822),
.B(n_1267),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1822),
.B(n_1268),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_1707),
.Y(n_2127)
);

NOR2xp33_ASAP7_75t_L g2128 ( 
.A(n_1869),
.B(n_1268),
.Y(n_2128)
);

OAI22xp5_ASAP7_75t_L g2129 ( 
.A1(n_1911),
.A2(n_919),
.B1(n_930),
.B2(n_928),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1875),
.Y(n_2130)
);

NAND3xp33_ASAP7_75t_L g2131 ( 
.A(n_1915),
.B(n_1284),
.C(n_1271),
.Y(n_2131)
);

A2O1A1Ixp33_ASAP7_75t_L g2132 ( 
.A1(n_1649),
.A2(n_936),
.B(n_942),
.C(n_934),
.Y(n_2132)
);

AOI21xp5_ASAP7_75t_L g2133 ( 
.A1(n_1836),
.A2(n_1589),
.B(n_1467),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1710),
.Y(n_2134)
);

NOR2xp33_ASAP7_75t_L g2135 ( 
.A(n_1868),
.B(n_815),
.Y(n_2135)
);

NOR2xp33_ASAP7_75t_L g2136 ( 
.A(n_1868),
.B(n_816),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_SL g2137 ( 
.A(n_1865),
.B(n_896),
.Y(n_2137)
);

O2A1O1Ixp33_ASAP7_75t_L g2138 ( 
.A1(n_1702),
.A2(n_952),
.B(n_976),
.C(n_948),
.Y(n_2138)
);

INVx2_ASAP7_75t_SL g2139 ( 
.A(n_1903),
.Y(n_2139)
);

INVx2_ASAP7_75t_SL g2140 ( 
.A(n_1903),
.Y(n_2140)
);

NAND2xp33_ASAP7_75t_L g2141 ( 
.A(n_1826),
.B(n_898),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1879),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1729),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_1755),
.B(n_1163),
.Y(n_2144)
);

NOR2xp33_ASAP7_75t_L g2145 ( 
.A(n_1796),
.B(n_904),
.Y(n_2145)
);

AOI22xp33_ASAP7_75t_L g2146 ( 
.A1(n_1733),
.A2(n_1128),
.B1(n_1162),
.B2(n_966),
.Y(n_2146)
);

INVx2_ASAP7_75t_SL g2147 ( 
.A(n_1903),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1879),
.Y(n_2148)
);

CKINVDCx5p33_ASAP7_75t_R g2149 ( 
.A(n_1843),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1720),
.B(n_908),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_1814),
.B(n_1286),
.Y(n_2151)
);

NOR2x1p5_ASAP7_75t_L g2152 ( 
.A(n_1845),
.B(n_1914),
.Y(n_2152)
);

INVxp67_ASAP7_75t_SL g2153 ( 
.A(n_1792),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1735),
.Y(n_2154)
);

INVx1_ASAP7_75t_SL g2155 ( 
.A(n_1826),
.Y(n_2155)
);

AND2x4_ASAP7_75t_L g2156 ( 
.A(n_1814),
.B(n_979),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_1642),
.Y(n_2157)
);

OAI22xp33_ASAP7_75t_L g2158 ( 
.A1(n_1814),
.A2(n_914),
.B1(n_920),
.B2(n_915),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_1895),
.B(n_922),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_1746),
.B(n_926),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1780),
.B(n_929),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1844),
.Y(n_2162)
);

AOI22xp33_ASAP7_75t_L g2163 ( 
.A1(n_1781),
.A2(n_1162),
.B1(n_1266),
.B2(n_1128),
.Y(n_2163)
);

OR2x6_ASAP7_75t_L g2164 ( 
.A(n_1797),
.B(n_1011),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_1861),
.B(n_937),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1643),
.Y(n_2166)
);

NOR2xp33_ASAP7_75t_L g2167 ( 
.A(n_1824),
.B(n_1827),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_1853),
.B(n_940),
.Y(n_2168)
);

BUFx6f_ASAP7_75t_L g2169 ( 
.A(n_1672),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_1652),
.Y(n_2170)
);

INVxp67_ASAP7_75t_L g2171 ( 
.A(n_1887),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1846),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1850),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_SL g2174 ( 
.A(n_1893),
.B(n_950),
.Y(n_2174)
);

AOI22xp5_ASAP7_75t_L g2175 ( 
.A1(n_1715),
.A2(n_962),
.B1(n_965),
.B2(n_958),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_1656),
.Y(n_2176)
);

BUFx6f_ASAP7_75t_L g2177 ( 
.A(n_1777),
.Y(n_2177)
);

INVxp67_ASAP7_75t_SL g2178 ( 
.A(n_1653),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_1782),
.B(n_969),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_1752),
.B(n_971),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1773),
.Y(n_2181)
);

INVx8_ASAP7_75t_L g2182 ( 
.A(n_1826),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_1727),
.B(n_1730),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1773),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_1736),
.B(n_975),
.Y(n_2185)
);

NAND3xp33_ASAP7_75t_SL g2186 ( 
.A(n_1662),
.B(n_984),
.C(n_980),
.Y(n_2186)
);

AND2x4_ASAP7_75t_SL g2187 ( 
.A(n_1783),
.B(n_1028),
.Y(n_2187)
);

NOR2xp33_ASAP7_75t_L g2188 ( 
.A(n_1859),
.B(n_1917),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_1808),
.B(n_1810),
.Y(n_2189)
);

INVxp67_ASAP7_75t_L g2190 ( 
.A(n_1706),
.Y(n_2190)
);

BUFx5_ASAP7_75t_L g2191 ( 
.A(n_1880),
.Y(n_2191)
);

AOI22xp33_ASAP7_75t_L g2192 ( 
.A1(n_1799),
.A2(n_1162),
.B1(n_1266),
.B2(n_1128),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_1657),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_SL g2194 ( 
.A(n_1877),
.B(n_988),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_1741),
.B(n_991),
.Y(n_2195)
);

BUFx6f_ASAP7_75t_L g2196 ( 
.A(n_1777),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_1741),
.B(n_995),
.Y(n_2197)
);

INVx8_ASAP7_75t_L g2198 ( 
.A(n_1787),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1799),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_1800),
.B(n_999),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1742),
.Y(n_2201)
);

NOR2xp33_ASAP7_75t_L g2202 ( 
.A(n_1885),
.B(n_1002),
.Y(n_2202)
);

INVx2_ASAP7_75t_SL g2203 ( 
.A(n_1834),
.Y(n_2203)
);

NOR2xp33_ASAP7_75t_L g2204 ( 
.A(n_1885),
.B(n_1003),
.Y(n_2204)
);

OAI22xp33_ASAP7_75t_L g2205 ( 
.A1(n_1848),
.A2(n_1020),
.B1(n_1026),
.B2(n_1009),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1767),
.Y(n_2206)
);

AO221x1_ASAP7_75t_L g2207 ( 
.A1(n_1703),
.A2(n_1266),
.B1(n_1273),
.B2(n_1162),
.C(n_1128),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1767),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_1883),
.B(n_1038),
.Y(n_2209)
);

NOR2xp33_ASAP7_75t_L g2210 ( 
.A(n_1904),
.B(n_1054),
.Y(n_2210)
);

AOI22xp33_ASAP7_75t_SL g2211 ( 
.A1(n_1704),
.A2(n_1061),
.B1(n_1063),
.B2(n_1060),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_1723),
.B(n_1066),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_SL g2213 ( 
.A(n_1777),
.B(n_1068),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_SL g2214 ( 
.A(n_1805),
.B(n_1902),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_1728),
.B(n_1078),
.Y(n_2215)
);

BUFx6f_ASAP7_75t_SL g2216 ( 
.A(n_1783),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_1660),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_SL g2218 ( 
.A(n_1805),
.B(n_1085),
.Y(n_2218)
);

NOR2xp33_ASAP7_75t_L g2219 ( 
.A(n_1904),
.B(n_1100),
.Y(n_2219)
);

AOI22xp5_ASAP7_75t_L g2220 ( 
.A1(n_1906),
.A2(n_1103),
.B1(n_1111),
.B2(n_1091),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_SL g2221 ( 
.A(n_1805),
.B(n_1114),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_1902),
.B(n_1117),
.Y(n_2222)
);

INVx2_ASAP7_75t_SL g2223 ( 
.A(n_1860),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_1909),
.B(n_1122),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_1909),
.B(n_1131),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_1886),
.B(n_1135),
.Y(n_2226)
);

OR2x2_ASAP7_75t_L g2227 ( 
.A(n_1900),
.B(n_1136),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_1886),
.B(n_1140),
.Y(n_2228)
);

NOR2xp33_ASAP7_75t_L g2229 ( 
.A(n_1891),
.B(n_1141),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_SL g2230 ( 
.A(n_1805),
.B(n_1146),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_SL g2231 ( 
.A(n_1856),
.B(n_1149),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_1888),
.B(n_1154),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_1882),
.B(n_1155),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_SL g2234 ( 
.A(n_1668),
.B(n_1156),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_1884),
.B(n_1164),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1734),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_SL g2237 ( 
.A(n_1682),
.B(n_1700),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_1832),
.B(n_1165),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_1716),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2085),
.B(n_2091),
.Y(n_2240)
);

AOI22xp33_ASAP7_75t_SL g2241 ( 
.A1(n_2153),
.A2(n_1880),
.B1(n_1874),
.B2(n_1704),
.Y(n_2241)
);

A2O1A1Ixp33_ASAP7_75t_L g2242 ( 
.A1(n_2090),
.A2(n_1711),
.B(n_1762),
.C(n_1761),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_SL g2243 ( 
.A(n_1926),
.B(n_1839),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_1926),
.B(n_1905),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1952),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_2078),
.B(n_1894),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2078),
.B(n_1891),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_1979),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_1959),
.B(n_1705),
.Y(n_2249)
);

BUFx2_ASAP7_75t_L g2250 ( 
.A(n_1963),
.Y(n_2250)
);

OAI21xp33_ASAP7_75t_L g2251 ( 
.A1(n_2124),
.A2(n_1774),
.B(n_1918),
.Y(n_2251)
);

BUFx6f_ASAP7_75t_L g2252 ( 
.A(n_1924),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_1971),
.B(n_1892),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_1930),
.B(n_1892),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2033),
.B(n_1168),
.Y(n_2255)
);

INVx2_ASAP7_75t_L g2256 ( 
.A(n_1984),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_1932),
.B(n_1874),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1985),
.Y(n_2258)
);

OAI22xp5_ASAP7_75t_L g2259 ( 
.A1(n_1932),
.A2(n_1918),
.B1(n_1897),
.B2(n_1724),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_1938),
.B(n_1939),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_SL g2261 ( 
.A(n_2106),
.B(n_1839),
.Y(n_2261)
);

O2A1O1Ixp33_ASAP7_75t_L g2262 ( 
.A1(n_2062),
.A2(n_2016),
.B(n_2132),
.C(n_2129),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_1989),
.Y(n_2263)
);

AO21x1_ASAP7_75t_L g2264 ( 
.A1(n_2231),
.A2(n_1912),
.B(n_1830),
.Y(n_2264)
);

O2A1O1Ixp33_ASAP7_75t_L g2265 ( 
.A1(n_2082),
.A2(n_994),
.B(n_996),
.C(n_989),
.Y(n_2265)
);

OAI21xp5_ASAP7_75t_L g2266 ( 
.A1(n_2037),
.A2(n_1745),
.B(n_1743),
.Y(n_2266)
);

NOR2xp33_ASAP7_75t_L g2267 ( 
.A(n_1939),
.B(n_1716),
.Y(n_2267)
);

NOR2xp33_ASAP7_75t_L g2268 ( 
.A(n_1955),
.B(n_1169),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_SL g2269 ( 
.A(n_2106),
.B(n_1857),
.Y(n_2269)
);

OAI21xp5_ASAP7_75t_L g2270 ( 
.A1(n_2201),
.A2(n_1748),
.B(n_1756),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1995),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_1955),
.B(n_1173),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_1998),
.Y(n_2273)
);

AO21x1_ASAP7_75t_L g2274 ( 
.A1(n_2133),
.A2(n_1802),
.B(n_1004),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2017),
.B(n_1174),
.Y(n_2275)
);

AOI21xp5_ASAP7_75t_L g2276 ( 
.A1(n_2048),
.A2(n_1791),
.B(n_1790),
.Y(n_2276)
);

AOI21xp5_ASAP7_75t_L g2277 ( 
.A1(n_2123),
.A2(n_1811),
.B(n_1794),
.Y(n_2277)
);

OAI21xp33_ASAP7_75t_L g2278 ( 
.A1(n_1920),
.A2(n_1177),
.B(n_1176),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_SL g2279 ( 
.A(n_2106),
.B(n_1857),
.Y(n_2279)
);

AOI21xp5_ASAP7_75t_L g2280 ( 
.A1(n_2123),
.A2(n_1833),
.B(n_1813),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2014),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_2019),
.Y(n_2282)
);

AOI21xp5_ASAP7_75t_L g2283 ( 
.A1(n_2125),
.A2(n_2126),
.B(n_2077),
.Y(n_2283)
);

AOI21xp5_ASAP7_75t_L g2284 ( 
.A1(n_2125),
.A2(n_1854),
.B(n_1842),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2017),
.B(n_1188),
.Y(n_2285)
);

HB1xp67_ASAP7_75t_L g2286 ( 
.A(n_1970),
.Y(n_2286)
);

AND2x4_ASAP7_75t_L g2287 ( 
.A(n_2074),
.B(n_1862),
.Y(n_2287)
);

BUFx2_ASAP7_75t_L g2288 ( 
.A(n_1988),
.Y(n_2288)
);

OAI22xp5_ASAP7_75t_L g2289 ( 
.A1(n_1928),
.A2(n_1192),
.B1(n_1195),
.B2(n_1189),
.Y(n_2289)
);

AOI21xp5_ASAP7_75t_L g2290 ( 
.A1(n_2206),
.A2(n_2208),
.B(n_2088),
.Y(n_2290)
);

AOI21xp5_ASAP7_75t_L g2291 ( 
.A1(n_2083),
.A2(n_1919),
.B(n_1910),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_SL g2292 ( 
.A(n_2106),
.B(n_1862),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_2084),
.B(n_1208),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2022),
.B(n_1209),
.Y(n_2294)
);

AND2x2_ASAP7_75t_SL g2295 ( 
.A(n_2093),
.B(n_1862),
.Y(n_2295)
);

OAI21xp5_ASAP7_75t_L g2296 ( 
.A1(n_2083),
.A2(n_1908),
.B(n_1899),
.Y(n_2296)
);

OAI21xp5_ASAP7_75t_L g2297 ( 
.A1(n_2088),
.A2(n_1908),
.B(n_1899),
.Y(n_2297)
);

AND2x2_ASAP7_75t_SL g2298 ( 
.A(n_1969),
.B(n_1128),
.Y(n_2298)
);

AND2x2_ASAP7_75t_SL g2299 ( 
.A(n_2015),
.B(n_1162),
.Y(n_2299)
);

NOR2xp33_ASAP7_75t_L g2300 ( 
.A(n_2101),
.B(n_2108),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_2027),
.Y(n_2301)
);

O2A1O1Ixp33_ASAP7_75t_L g2302 ( 
.A1(n_2082),
.A2(n_1005),
.B(n_1013),
.C(n_998),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2022),
.B(n_2031),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2031),
.B(n_1216),
.Y(n_2304)
);

AOI21xp5_ASAP7_75t_L g2305 ( 
.A1(n_2101),
.A2(n_1019),
.B(n_1018),
.Y(n_2305)
);

NAND2xp33_ASAP7_75t_L g2306 ( 
.A(n_2182),
.B(n_1219),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2036),
.B(n_1223),
.Y(n_2307)
);

CKINVDCx8_ASAP7_75t_R g2308 ( 
.A(n_2198),
.Y(n_2308)
);

OAI21xp5_ASAP7_75t_L g2309 ( 
.A1(n_2108),
.A2(n_1031),
.B(n_1025),
.Y(n_2309)
);

AOI21xp5_ASAP7_75t_L g2310 ( 
.A1(n_2222),
.A2(n_1047),
.B(n_1036),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2036),
.B(n_1226),
.Y(n_2311)
);

O2A1O1Ixp5_ASAP7_75t_L g2312 ( 
.A1(n_2009),
.A2(n_1182),
.B(n_1198),
.C(n_1109),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_1922),
.B(n_1263),
.Y(n_2313)
);

NOR3xp33_ASAP7_75t_L g2314 ( 
.A(n_2029),
.B(n_1277),
.C(n_1067),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2189),
.B(n_1065),
.Y(n_2315)
);

OAI22xp5_ASAP7_75t_L g2316 ( 
.A1(n_1942),
.A2(n_2183),
.B1(n_1987),
.B2(n_2164),
.Y(n_2316)
);

AND2x2_ASAP7_75t_L g2317 ( 
.A(n_2096),
.B(n_1076),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2189),
.B(n_1089),
.Y(n_2318)
);

INVx2_ASAP7_75t_SL g2319 ( 
.A(n_1954),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2028),
.Y(n_2320)
);

AOI21xp5_ASAP7_75t_L g2321 ( 
.A1(n_2222),
.A2(n_1106),
.B(n_1090),
.Y(n_2321)
);

AOI21xp5_ASAP7_75t_L g2322 ( 
.A1(n_2195),
.A2(n_2197),
.B(n_2226),
.Y(n_2322)
);

BUFx2_ASAP7_75t_L g2323 ( 
.A(n_2006),
.Y(n_2323)
);

OAI21xp5_ASAP7_75t_L g2324 ( 
.A1(n_2195),
.A2(n_1126),
.B(n_1115),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2095),
.B(n_1129),
.Y(n_2325)
);

BUFx4f_ASAP7_75t_L g2326 ( 
.A(n_2198),
.Y(n_2326)
);

AOI22xp5_ASAP7_75t_L g2327 ( 
.A1(n_2055),
.A2(n_1142),
.B1(n_1145),
.B2(n_1132),
.Y(n_2327)
);

NOR2xp33_ASAP7_75t_L g2328 ( 
.A(n_1961),
.B(n_1148),
.Y(n_2328)
);

A2O1A1Ixp33_ASAP7_75t_L g2329 ( 
.A1(n_2138),
.A2(n_1157),
.B(n_1160),
.C(n_1151),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_1987),
.B(n_1161),
.Y(n_2330)
);

AOI21xp5_ASAP7_75t_L g2331 ( 
.A1(n_2197),
.A2(n_1186),
.B(n_1184),
.Y(n_2331)
);

OAI21xp5_ASAP7_75t_L g2332 ( 
.A1(n_1967),
.A2(n_1203),
.B(n_1199),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_SL g2333 ( 
.A(n_2004),
.B(n_1266),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2034),
.Y(n_2334)
);

NOR2xp33_ASAP7_75t_L g2335 ( 
.A(n_1962),
.B(n_1237),
.Y(n_2335)
);

INVxp67_ASAP7_75t_L g2336 ( 
.A(n_2001),
.Y(n_2336)
);

AOI21xp5_ASAP7_75t_L g2337 ( 
.A1(n_2226),
.A2(n_1247),
.B(n_1243),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2044),
.B(n_1182),
.Y(n_2338)
);

AOI21xp5_ASAP7_75t_L g2339 ( 
.A1(n_2228),
.A2(n_1217),
.B(n_1198),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2053),
.B(n_2073),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2080),
.Y(n_2341)
);

NOR2xp33_ASAP7_75t_L g2342 ( 
.A(n_2228),
.B(n_7),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_1958),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2003),
.B(n_7),
.Y(n_2344)
);

INVx3_ASAP7_75t_L g2345 ( 
.A(n_2182),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2007),
.B(n_8),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_SL g2347 ( 
.A(n_2004),
.B(n_1273),
.Y(n_2347)
);

NOR2x1p5_ASAP7_75t_L g2348 ( 
.A(n_2002),
.B(n_913),
.Y(n_2348)
);

BUFx3_ASAP7_75t_L g2349 ( 
.A(n_1948),
.Y(n_2349)
);

A2O1A1Ixp33_ASAP7_75t_L g2350 ( 
.A1(n_2021),
.A2(n_1273),
.B(n_1071),
.C(n_1079),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_1964),
.Y(n_2351)
);

OAI22xp5_ASAP7_75t_L g2352 ( 
.A1(n_2164),
.A2(n_1273),
.B1(n_933),
.B2(n_941),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_SL g2353 ( 
.A(n_2004),
.B(n_913),
.Y(n_2353)
);

AOI21xp5_ASAP7_75t_L g2354 ( 
.A1(n_2038),
.A2(n_1616),
.B(n_1610),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_1996),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_SL g2356 ( 
.A(n_2004),
.B(n_913),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2046),
.B(n_8),
.Y(n_2357)
);

INVxp67_ASAP7_75t_L g2358 ( 
.A(n_2164),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2162),
.Y(n_2359)
);

NOR2xp33_ASAP7_75t_L g2360 ( 
.A(n_2047),
.B(n_9),
.Y(n_2360)
);

OAI21xp5_ASAP7_75t_L g2361 ( 
.A1(n_2185),
.A2(n_933),
.B(n_913),
.Y(n_2361)
);

OAI21xp5_ASAP7_75t_L g2362 ( 
.A1(n_2185),
.A2(n_933),
.B(n_913),
.Y(n_2362)
);

NOR2xp33_ASAP7_75t_L g2363 ( 
.A(n_2050),
.B(n_9),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2052),
.B(n_10),
.Y(n_2364)
);

NOR2xp33_ASAP7_75t_L g2365 ( 
.A(n_2165),
.B(n_10),
.Y(n_2365)
);

AOI21xp5_ASAP7_75t_L g2366 ( 
.A1(n_2117),
.A2(n_1616),
.B(n_1610),
.Y(n_2366)
);

INVx6_ASAP7_75t_L g2367 ( 
.A(n_1954),
.Y(n_2367)
);

NOR2xp33_ASAP7_75t_L g2368 ( 
.A(n_1968),
.B(n_10),
.Y(n_2368)
);

AND2x2_ASAP7_75t_L g2369 ( 
.A(n_2122),
.B(n_11),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_SL g2370 ( 
.A(n_2042),
.B(n_2079),
.Y(n_2370)
);

OAI21xp5_ASAP7_75t_L g2371 ( 
.A1(n_2233),
.A2(n_941),
.B(n_933),
.Y(n_2371)
);

AND2x2_ASAP7_75t_L g2372 ( 
.A(n_1972),
.B(n_11),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2172),
.Y(n_2373)
);

A2O1A1Ixp33_ASAP7_75t_L g2374 ( 
.A1(n_2113),
.A2(n_2056),
.B(n_1992),
.C(n_1982),
.Y(n_2374)
);

O2A1O1Ixp5_ASAP7_75t_L g2375 ( 
.A1(n_2020),
.A2(n_2237),
.B(n_2178),
.C(n_2214),
.Y(n_2375)
);

AOI21xp5_ASAP7_75t_L g2376 ( 
.A1(n_2235),
.A2(n_1630),
.B(n_1619),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_1973),
.B(n_11),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2173),
.Y(n_2378)
);

BUFx6f_ASAP7_75t_L g2379 ( 
.A(n_1924),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_1975),
.B(n_12),
.Y(n_2380)
);

O2A1O1Ixp33_ASAP7_75t_L g2381 ( 
.A1(n_2129),
.A2(n_14),
.B(n_12),
.C(n_13),
.Y(n_2381)
);

AOI22xp5_ASAP7_75t_L g2382 ( 
.A1(n_2060),
.A2(n_943),
.B1(n_945),
.B2(n_941),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2000),
.B(n_12),
.Y(n_2383)
);

AO21x1_ASAP7_75t_L g2384 ( 
.A1(n_2141),
.A2(n_415),
.B(n_414),
.Y(n_2384)
);

INVx3_ASAP7_75t_L g2385 ( 
.A(n_2182),
.Y(n_2385)
);

AOI21xp5_ASAP7_75t_L g2386 ( 
.A1(n_2097),
.A2(n_2110),
.B(n_2099),
.Y(n_2386)
);

AOI21xp5_ASAP7_75t_L g2387 ( 
.A1(n_2065),
.A2(n_1630),
.B(n_1619),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_2012),
.Y(n_2388)
);

AOI21xp5_ASAP7_75t_L g2389 ( 
.A1(n_2067),
.A2(n_1635),
.B(n_1633),
.Y(n_2389)
);

HB1xp67_ASAP7_75t_L g2390 ( 
.A(n_2074),
.Y(n_2390)
);

INVxp67_ASAP7_75t_L g2391 ( 
.A(n_2042),
.Y(n_2391)
);

O2A1O1Ixp33_ASAP7_75t_L g2392 ( 
.A1(n_2032),
.A2(n_1953),
.B(n_2061),
.C(n_2068),
.Y(n_2392)
);

NOR2xp33_ASAP7_75t_L g2393 ( 
.A(n_2159),
.B(n_15),
.Y(n_2393)
);

BUFx12f_ASAP7_75t_L g2394 ( 
.A(n_2025),
.Y(n_2394)
);

O2A1O1Ixp33_ASAP7_75t_L g2395 ( 
.A1(n_2032),
.A2(n_18),
.B(n_16),
.C(n_17),
.Y(n_2395)
);

INVx2_ASAP7_75t_SL g2396 ( 
.A(n_2198),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_SL g2397 ( 
.A(n_2004),
.B(n_2191),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_1951),
.B(n_17),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_1974),
.B(n_17),
.Y(n_2399)
);

NOR3xp33_ASAP7_75t_L g2400 ( 
.A(n_1949),
.B(n_18),
.C(n_19),
.Y(n_2400)
);

AOI22xp33_ASAP7_75t_L g2401 ( 
.A1(n_1957),
.A2(n_943),
.B1(n_945),
.B2(n_941),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_2018),
.Y(n_2402)
);

AOI21xp5_ASAP7_75t_L g2403 ( 
.A1(n_2105),
.A2(n_945),
.B(n_943),
.Y(n_2403)
);

BUFx2_ASAP7_75t_L g2404 ( 
.A(n_2074),
.Y(n_2404)
);

NOR2xp33_ASAP7_75t_L g2405 ( 
.A(n_2109),
.B(n_18),
.Y(n_2405)
);

INVx11_ASAP7_75t_L g2406 ( 
.A(n_2025),
.Y(n_2406)
);

NOR2xp33_ASAP7_75t_L g2407 ( 
.A(n_2005),
.B(n_19),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_1965),
.B(n_20),
.Y(n_2408)
);

AOI21xp5_ASAP7_75t_L g2409 ( 
.A1(n_2066),
.A2(n_945),
.B(n_943),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_SL g2410 ( 
.A(n_2191),
.B(n_2155),
.Y(n_2410)
);

AND2x2_ASAP7_75t_L g2411 ( 
.A(n_1921),
.B(n_20),
.Y(n_2411)
);

AOI21xp5_ASAP7_75t_L g2412 ( 
.A1(n_2054),
.A2(n_945),
.B(n_943),
.Y(n_2412)
);

INVx3_ASAP7_75t_L g2413 ( 
.A(n_1991),
.Y(n_2413)
);

AOI21xp5_ASAP7_75t_L g2414 ( 
.A1(n_2059),
.A2(n_2039),
.B(n_2174),
.Y(n_2414)
);

NOR2xp33_ASAP7_75t_L g2415 ( 
.A(n_2008),
.B(n_20),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_SL g2416 ( 
.A(n_2191),
.B(n_1058),
.Y(n_2416)
);

INVx3_ASAP7_75t_L g2417 ( 
.A(n_1991),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2064),
.B(n_21),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2100),
.Y(n_2419)
);

NOR2xp33_ASAP7_75t_L g2420 ( 
.A(n_2010),
.B(n_21),
.Y(n_2420)
);

AOI21xp5_ASAP7_75t_L g2421 ( 
.A1(n_1947),
.A2(n_1071),
.B(n_1058),
.Y(n_2421)
);

BUFx3_ASAP7_75t_L g2422 ( 
.A(n_1948),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_2064),
.B(n_1960),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_2030),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2102),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2063),
.B(n_21),
.Y(n_2426)
);

AOI21xp5_ASAP7_75t_L g2427 ( 
.A1(n_1956),
.A2(n_1071),
.B(n_1058),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_1977),
.B(n_22),
.Y(n_2428)
);

NAND3xp33_ASAP7_75t_L g2429 ( 
.A(n_1934),
.B(n_1071),
.C(n_1058),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2040),
.B(n_22),
.Y(n_2430)
);

OAI22xp5_ASAP7_75t_L g2431 ( 
.A1(n_2076),
.A2(n_2112),
.B1(n_2140),
.B2(n_2139),
.Y(n_2431)
);

OAI21xp5_ASAP7_75t_L g2432 ( 
.A1(n_2035),
.A2(n_1071),
.B(n_1058),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2043),
.Y(n_2433)
);

AOI22xp5_ASAP7_75t_L g2434 ( 
.A1(n_2023),
.A2(n_1083),
.B1(n_1288),
.B2(n_1079),
.Y(n_2434)
);

INVx3_ASAP7_75t_L g2435 ( 
.A(n_1991),
.Y(n_2435)
);

BUFx2_ASAP7_75t_L g2436 ( 
.A(n_1997),
.Y(n_2436)
);

AOI21xp5_ASAP7_75t_L g2437 ( 
.A1(n_2194),
.A2(n_1083),
.B(n_1079),
.Y(n_2437)
);

OAI21xp5_ASAP7_75t_L g2438 ( 
.A1(n_2045),
.A2(n_1288),
.B(n_1083),
.Y(n_2438)
);

AOI21xp5_ASAP7_75t_L g2439 ( 
.A1(n_1927),
.A2(n_1288),
.B(n_1083),
.Y(n_2439)
);

OAI22xp5_ASAP7_75t_L g2440 ( 
.A1(n_2076),
.A2(n_1288),
.B1(n_25),
.B2(n_23),
.Y(n_2440)
);

AND2x4_ASAP7_75t_L g2441 ( 
.A(n_2087),
.B(n_23),
.Y(n_2441)
);

AOI21xp5_ASAP7_75t_L g2442 ( 
.A1(n_1931),
.A2(n_24),
.B(n_25),
.Y(n_2442)
);

AND2x2_ASAP7_75t_L g2443 ( 
.A(n_2144),
.B(n_24),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2098),
.B(n_24),
.Y(n_2444)
);

AOI21xp5_ASAP7_75t_L g2445 ( 
.A1(n_1935),
.A2(n_26),
.B(n_27),
.Y(n_2445)
);

AOI21xp5_ASAP7_75t_L g2446 ( 
.A1(n_1937),
.A2(n_26),
.B(n_27),
.Y(n_2446)
);

BUFx3_ASAP7_75t_L g2447 ( 
.A(n_1997),
.Y(n_2447)
);

NOR2xp67_ASAP7_75t_L g2448 ( 
.A(n_2171),
.B(n_26),
.Y(n_2448)
);

AOI21xp33_ASAP7_75t_L g2449 ( 
.A1(n_1999),
.A2(n_29),
.B(n_30),
.Y(n_2449)
);

AOI21xp5_ASAP7_75t_L g2450 ( 
.A1(n_1978),
.A2(n_29),
.B(n_31),
.Y(n_2450)
);

AOI21xp5_ASAP7_75t_L g2451 ( 
.A1(n_1980),
.A2(n_31),
.B(n_32),
.Y(n_2451)
);

A2O1A1Ixp33_ASAP7_75t_L g2452 ( 
.A1(n_2188),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_2452)
);

AOI21xp5_ASAP7_75t_L g2453 ( 
.A1(n_1990),
.A2(n_32),
.B(n_33),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2120),
.B(n_34),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2128),
.B(n_2150),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_1944),
.Y(n_2456)
);

A2O1A1Ixp33_ASAP7_75t_L g2457 ( 
.A1(n_2160),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_2457)
);

BUFx12f_ASAP7_75t_L g2458 ( 
.A(n_2149),
.Y(n_2458)
);

INVx3_ASAP7_75t_L g2459 ( 
.A(n_2169),
.Y(n_2459)
);

NOR3xp33_ASAP7_75t_L g2460 ( 
.A(n_2081),
.B(n_35),
.C(n_36),
.Y(n_2460)
);

OAI22xp5_ASAP7_75t_L g2461 ( 
.A1(n_2076),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_2461)
);

AOI21x1_ASAP7_75t_L g2462 ( 
.A1(n_2236),
.A2(n_38),
.B(n_39),
.Y(n_2462)
);

O2A1O1Ixp33_ASAP7_75t_L g2463 ( 
.A1(n_2224),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_2463)
);

BUFx6f_ASAP7_75t_L g2464 ( 
.A(n_1924),
.Y(n_2464)
);

AOI21xp5_ASAP7_75t_L g2465 ( 
.A1(n_2161),
.A2(n_38),
.B(n_39),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2150),
.B(n_41),
.Y(n_2466)
);

AOI21xp5_ASAP7_75t_L g2467 ( 
.A1(n_2179),
.A2(n_41),
.B(n_42),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_2151),
.B(n_42),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2089),
.B(n_42),
.Y(n_2469)
);

O2A1O1Ixp5_ASAP7_75t_L g2470 ( 
.A1(n_2234),
.A2(n_45),
.B(n_43),
.C(n_44),
.Y(n_2470)
);

OAI22xp5_ASAP7_75t_L g2471 ( 
.A1(n_2112),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2094),
.B(n_46),
.Y(n_2472)
);

A2O1A1Ixp33_ASAP7_75t_L g2473 ( 
.A1(n_2209),
.A2(n_48),
.B(n_46),
.C(n_47),
.Y(n_2473)
);

NAND3xp33_ASAP7_75t_L g2474 ( 
.A(n_2069),
.B(n_47),
.C(n_48),
.Y(n_2474)
);

AOI21x1_ASAP7_75t_L g2475 ( 
.A1(n_1925),
.A2(n_47),
.B(n_49),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2086),
.Y(n_2476)
);

INVx2_ASAP7_75t_L g2477 ( 
.A(n_2092),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2104),
.B(n_50),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2156),
.B(n_50),
.Y(n_2479)
);

INVx3_ASAP7_75t_L g2480 ( 
.A(n_2169),
.Y(n_2480)
);

O2A1O1Ixp33_ASAP7_75t_L g2481 ( 
.A1(n_2224),
.A2(n_52),
.B(n_50),
.C(n_51),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_2156),
.B(n_51),
.Y(n_2482)
);

BUFx4f_ASAP7_75t_L g2483 ( 
.A(n_2112),
.Y(n_2483)
);

NOR3xp33_ASAP7_75t_L g2484 ( 
.A(n_1929),
.B(n_53),
.C(n_54),
.Y(n_2484)
);

NOR2x1p5_ASAP7_75t_L g2485 ( 
.A(n_1983),
.B(n_54),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_2115),
.Y(n_2486)
);

INVx1_ASAP7_75t_SL g2487 ( 
.A(n_1941),
.Y(n_2487)
);

OAI21xp33_ASAP7_75t_SL g2488 ( 
.A1(n_1923),
.A2(n_2147),
.B(n_2207),
.Y(n_2488)
);

AND2x4_ASAP7_75t_L g2489 ( 
.A(n_2026),
.B(n_55),
.Y(n_2489)
);

O2A1O1Ixp33_ASAP7_75t_L g2490 ( 
.A1(n_2225),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_2490)
);

NAND3xp33_ASAP7_75t_L g2491 ( 
.A(n_2146),
.B(n_56),
.C(n_58),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_1950),
.Y(n_2492)
);

OAI21xp5_ASAP7_75t_L g2493 ( 
.A1(n_2127),
.A2(n_58),
.B(n_59),
.Y(n_2493)
);

AOI22xp5_ASAP7_75t_L g2494 ( 
.A1(n_1945),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2180),
.B(n_59),
.Y(n_2495)
);

OAI21xp5_ASAP7_75t_L g2496 ( 
.A1(n_2134),
.A2(n_60),
.B(n_61),
.Y(n_2496)
);

AO21x1_ASAP7_75t_L g2497 ( 
.A1(n_2118),
.A2(n_420),
.B(n_419),
.Y(n_2497)
);

AND2x4_ASAP7_75t_L g2498 ( 
.A(n_2024),
.B(n_60),
.Y(n_2498)
);

A2O1A1Ixp33_ASAP7_75t_L g2499 ( 
.A1(n_1946),
.A2(n_64),
.B(n_62),
.C(n_63),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_2190),
.B(n_62),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2143),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_2225),
.B(n_62),
.Y(n_2502)
);

OAI22xp5_ASAP7_75t_L g2503 ( 
.A1(n_2011),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_2503)
);

NOR2x1_ASAP7_75t_L g2504 ( 
.A(n_2152),
.B(n_63),
.Y(n_2504)
);

AOI21xp5_ASAP7_75t_L g2505 ( 
.A1(n_2154),
.A2(n_2200),
.B(n_2166),
.Y(n_2505)
);

HB1xp67_ASAP7_75t_L g2506 ( 
.A(n_2070),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2158),
.B(n_64),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2103),
.B(n_65),
.Y(n_2508)
);

AOI21xp5_ASAP7_75t_L g2509 ( 
.A1(n_2157),
.A2(n_2176),
.B(n_2170),
.Y(n_2509)
);

AND2x2_ASAP7_75t_L g2510 ( 
.A(n_2168),
.B(n_65),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2107),
.B(n_2111),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_2114),
.B(n_66),
.Y(n_2512)
);

NOR2xp33_ASAP7_75t_L g2513 ( 
.A(n_1993),
.B(n_66),
.Y(n_2513)
);

AND2x4_ASAP7_75t_L g2514 ( 
.A(n_2051),
.B(n_66),
.Y(n_2514)
);

AOI21xp33_ASAP7_75t_L g2515 ( 
.A1(n_2202),
.A2(n_67),
.B(n_68),
.Y(n_2515)
);

A2O1A1Ixp33_ASAP7_75t_L g2516 ( 
.A1(n_1943),
.A2(n_69),
.B(n_67),
.C(n_68),
.Y(n_2516)
);

INVx2_ASAP7_75t_L g2517 ( 
.A(n_2121),
.Y(n_2517)
);

AOI21xp5_ASAP7_75t_L g2518 ( 
.A1(n_2193),
.A2(n_2217),
.B(n_2057),
.Y(n_2518)
);

BUFx3_ASAP7_75t_L g2519 ( 
.A(n_2041),
.Y(n_2519)
);

BUFx6f_ASAP7_75t_L g2520 ( 
.A(n_1976),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_SL g2521 ( 
.A(n_2191),
.B(n_67),
.Y(n_2521)
);

OAI21xp33_ASAP7_75t_L g2522 ( 
.A1(n_1940),
.A2(n_68),
.B(n_69),
.Y(n_2522)
);

NOR2xp33_ASAP7_75t_L g2523 ( 
.A(n_2220),
.B(n_69),
.Y(n_2523)
);

AOI21x1_ASAP7_75t_L g2524 ( 
.A1(n_1933),
.A2(n_70),
.B(n_71),
.Y(n_2524)
);

AOI21xp5_ASAP7_75t_L g2525 ( 
.A1(n_2049),
.A2(n_74),
.B(n_75),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2130),
.B(n_74),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2142),
.B(n_75),
.Y(n_2527)
);

INVx4_ASAP7_75t_L g2528 ( 
.A(n_2216),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_2148),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2135),
.B(n_77),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2136),
.B(n_77),
.Y(n_2531)
);

BUFx6f_ASAP7_75t_L g2532 ( 
.A(n_1976),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2181),
.Y(n_2533)
);

OAI21xp5_ASAP7_75t_L g2534 ( 
.A1(n_2163),
.A2(n_2131),
.B(n_2184),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_2199),
.B(n_77),
.Y(n_2535)
);

AND2x2_ASAP7_75t_L g2536 ( 
.A(n_2013),
.B(n_78),
.Y(n_2536)
);

HB1xp67_ASAP7_75t_L g2537 ( 
.A(n_2071),
.Y(n_2537)
);

INVx3_ASAP7_75t_L g2538 ( 
.A(n_2169),
.Y(n_2538)
);

OR2x2_ASAP7_75t_L g2539 ( 
.A(n_2227),
.B(n_78),
.Y(n_2539)
);

BUFx4f_ASAP7_75t_L g2540 ( 
.A(n_2075),
.Y(n_2540)
);

AOI22xp5_ASAP7_75t_L g2541 ( 
.A1(n_2204),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_2541)
);

AOI21xp5_ASAP7_75t_L g2542 ( 
.A1(n_1981),
.A2(n_2239),
.B(n_2215),
.Y(n_2542)
);

AOI22xp33_ASAP7_75t_L g2543 ( 
.A1(n_2186),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_2543)
);

A2O1A1Ixp33_ASAP7_75t_L g2544 ( 
.A1(n_2167),
.A2(n_82),
.B(n_79),
.C(n_81),
.Y(n_2544)
);

AOI21xp5_ASAP7_75t_L g2545 ( 
.A1(n_2212),
.A2(n_82),
.B(n_83),
.Y(n_2545)
);

NOR2xp33_ASAP7_75t_L g2546 ( 
.A(n_2232),
.B(n_82),
.Y(n_2546)
);

AO21x1_ASAP7_75t_L g2547 ( 
.A1(n_2118),
.A2(n_421),
.B(n_420),
.Y(n_2547)
);

OAI21xp5_ASAP7_75t_L g2548 ( 
.A1(n_2232),
.A2(n_83),
.B(n_84),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2119),
.B(n_2205),
.Y(n_2549)
);

AOI21xp5_ASAP7_75t_L g2550 ( 
.A1(n_2238),
.A2(n_85),
.B(n_86),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_SL g2551 ( 
.A(n_2211),
.B(n_86),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2119),
.B(n_85),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2229),
.B(n_86),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2210),
.B(n_87),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2219),
.B(n_87),
.Y(n_2555)
);

AND2x2_ASAP7_75t_SL g2556 ( 
.A(n_2187),
.B(n_87),
.Y(n_2556)
);

NOR2xp33_ASAP7_75t_SL g2557 ( 
.A(n_2216),
.B(n_88),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2203),
.Y(n_2558)
);

AOI21xp5_ASAP7_75t_L g2559 ( 
.A1(n_2145),
.A2(n_88),
.B(n_89),
.Y(n_2559)
);

OAI21xp5_ASAP7_75t_L g2560 ( 
.A1(n_2192),
.A2(n_88),
.B(n_89),
.Y(n_2560)
);

AOI22xp33_ASAP7_75t_L g2561 ( 
.A1(n_2072),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_1966),
.Y(n_2562)
);

AOI21x1_ASAP7_75t_L g2563 ( 
.A1(n_2213),
.A2(n_92),
.B(n_93),
.Y(n_2563)
);

AOI21x1_ASAP7_75t_L g2564 ( 
.A1(n_2218),
.A2(n_93),
.B(n_94),
.Y(n_2564)
);

AOI21xp5_ASAP7_75t_L g2565 ( 
.A1(n_2071),
.A2(n_94),
.B(n_95),
.Y(n_2565)
);

INVx2_ASAP7_75t_L g2566 ( 
.A(n_1966),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2175),
.B(n_94),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_SL g2568 ( 
.A(n_1976),
.B(n_95),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_1994),
.Y(n_2569)
);

OAI21xp5_ASAP7_75t_L g2570 ( 
.A1(n_2221),
.A2(n_96),
.B(n_97),
.Y(n_2570)
);

NOR2xp33_ASAP7_75t_L g2571 ( 
.A(n_2137),
.B(n_96),
.Y(n_2571)
);

BUFx6f_ASAP7_75t_L g2572 ( 
.A(n_1986),
.Y(n_2572)
);

AOI21xp5_ASAP7_75t_L g2573 ( 
.A1(n_2230),
.A2(n_97),
.B(n_98),
.Y(n_2573)
);

NOR2xp33_ASAP7_75t_L g2574 ( 
.A(n_2223),
.B(n_97),
.Y(n_2574)
);

AND2x4_ASAP7_75t_L g2575 ( 
.A(n_1936),
.B(n_2058),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_SL g2576 ( 
.A(n_1986),
.B(n_98),
.Y(n_2576)
);

AOI21xp5_ASAP7_75t_L g2577 ( 
.A1(n_1994),
.A2(n_1986),
.B(n_2116),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2177),
.Y(n_2578)
);

AOI21xp5_ASAP7_75t_L g2579 ( 
.A1(n_2177),
.A2(n_99),
.B(n_100),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2177),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2196),
.Y(n_2581)
);

AND2x2_ASAP7_75t_L g2582 ( 
.A(n_2196),
.B(n_99),
.Y(n_2582)
);

AOI21xp5_ASAP7_75t_L g2583 ( 
.A1(n_2196),
.A2(n_99),
.B(n_100),
.Y(n_2583)
);

HB1xp67_ASAP7_75t_L g2584 ( 
.A(n_1926),
.Y(n_2584)
);

AOI21xp5_ASAP7_75t_L g2585 ( 
.A1(n_1926),
.A2(n_101),
.B(n_102),
.Y(n_2585)
);

NOR2xp33_ASAP7_75t_L g2586 ( 
.A(n_2090),
.B(n_102),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2085),
.B(n_102),
.Y(n_2587)
);

NOR2xp33_ASAP7_75t_L g2588 ( 
.A(n_2090),
.B(n_103),
.Y(n_2588)
);

BUFx3_ASAP7_75t_L g2589 ( 
.A(n_1948),
.Y(n_2589)
);

BUFx3_ASAP7_75t_L g2590 ( 
.A(n_1948),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2085),
.Y(n_2591)
);

AOI21xp5_ASAP7_75t_L g2592 ( 
.A1(n_1926),
.A2(n_103),
.B(n_104),
.Y(n_2592)
);

OAI21xp5_ASAP7_75t_L g2593 ( 
.A1(n_1971),
.A2(n_103),
.B(n_104),
.Y(n_2593)
);

AOI21xp5_ASAP7_75t_L g2594 ( 
.A1(n_1926),
.A2(n_105),
.B(n_106),
.Y(n_2594)
);

INVx1_ASAP7_75t_SL g2595 ( 
.A(n_1959),
.Y(n_2595)
);

NAND2x1p5_ASAP7_75t_L g2596 ( 
.A(n_2106),
.B(n_105),
.Y(n_2596)
);

AOI21xp5_ASAP7_75t_L g2597 ( 
.A1(n_1926),
.A2(n_106),
.B(n_107),
.Y(n_2597)
);

O2A1O1Ixp33_ASAP7_75t_SL g2598 ( 
.A1(n_1926),
.A2(n_108),
.B(n_106),
.C(n_107),
.Y(n_2598)
);

A2O1A1Ixp33_ASAP7_75t_L g2599 ( 
.A1(n_2090),
.A2(n_109),
.B(n_107),
.C(n_108),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2085),
.B(n_109),
.Y(n_2600)
);

HB1xp67_ASAP7_75t_L g2601 ( 
.A(n_1926),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_L g2602 ( 
.A(n_2085),
.B(n_109),
.Y(n_2602)
);

INVx3_ASAP7_75t_L g2603 ( 
.A(n_2182),
.Y(n_2603)
);

NOR2xp33_ASAP7_75t_L g2604 ( 
.A(n_2090),
.B(n_110),
.Y(n_2604)
);

NOR2xp33_ASAP7_75t_SL g2605 ( 
.A(n_2006),
.B(n_110),
.Y(n_2605)
);

AOI33xp33_ASAP7_75t_L g2606 ( 
.A1(n_1951),
.A2(n_113),
.A3(n_115),
.B1(n_111),
.B2(n_112),
.B3(n_114),
.Y(n_2606)
);

O2A1O1Ixp33_ASAP7_75t_L g2607 ( 
.A1(n_2062),
.A2(n_113),
.B(n_111),
.C(n_112),
.Y(n_2607)
);

OAI22xp5_ASAP7_75t_L g2608 ( 
.A1(n_1926),
.A2(n_115),
.B1(n_112),
.B2(n_113),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2085),
.B(n_115),
.Y(n_2609)
);

OAI22xp5_ASAP7_75t_L g2610 ( 
.A1(n_1926),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.Y(n_2610)
);

O2A1O1Ixp33_ASAP7_75t_L g2611 ( 
.A1(n_2062),
.A2(n_119),
.B(n_117),
.C(n_118),
.Y(n_2611)
);

A2O1A1Ixp33_ASAP7_75t_L g2612 ( 
.A1(n_2090),
.A2(n_120),
.B(n_118),
.C(n_119),
.Y(n_2612)
);

INVx3_ASAP7_75t_L g2613 ( 
.A(n_2182),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_2085),
.B(n_120),
.Y(n_2614)
);

NOR2xp33_ASAP7_75t_L g2615 ( 
.A(n_2090),
.B(n_121),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_2085),
.B(n_122),
.Y(n_2616)
);

NOR2xp33_ASAP7_75t_L g2617 ( 
.A(n_2090),
.B(n_122),
.Y(n_2617)
);

O2A1O1Ixp33_ASAP7_75t_L g2618 ( 
.A1(n_2062),
.A2(n_124),
.B(n_122),
.C(n_123),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_SL g2619 ( 
.A(n_1963),
.B(n_124),
.Y(n_2619)
);

INVx3_ASAP7_75t_L g2620 ( 
.A(n_2182),
.Y(n_2620)
);

AOI22xp5_ASAP7_75t_L g2621 ( 
.A1(n_1926),
.A2(n_126),
.B1(n_123),
.B2(n_125),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_L g2622 ( 
.A(n_2085),
.B(n_126),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_SL g2623 ( 
.A(n_1926),
.B(n_126),
.Y(n_2623)
);

OR2x2_ASAP7_75t_L g2624 ( 
.A(n_1963),
.B(n_127),
.Y(n_2624)
);

AOI22xp33_ASAP7_75t_L g2625 ( 
.A1(n_2033),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_2625)
);

AO21x1_ASAP7_75t_L g2626 ( 
.A1(n_2231),
.A2(n_423),
.B(n_422),
.Y(n_2626)
);

BUFx12f_ASAP7_75t_L g2627 ( 
.A(n_2025),
.Y(n_2627)
);

OAI21xp33_ASAP7_75t_L g2628 ( 
.A1(n_2090),
.A2(n_127),
.B(n_128),
.Y(n_2628)
);

OAI22xp5_ASAP7_75t_L g2629 ( 
.A1(n_1926),
.A2(n_131),
.B1(n_128),
.B2(n_130),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_2085),
.B(n_130),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_L g2631 ( 
.A(n_2085),
.B(n_131),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_L g2632 ( 
.A(n_2085),
.B(n_132),
.Y(n_2632)
);

AOI21xp5_ASAP7_75t_L g2633 ( 
.A1(n_1926),
.A2(n_132),
.B(n_133),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2085),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_1926),
.Y(n_2635)
);

AND2x2_ASAP7_75t_L g2636 ( 
.A(n_1959),
.B(n_132),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2085),
.B(n_133),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_L g2638 ( 
.A(n_2085),
.B(n_134),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2085),
.Y(n_2639)
);

AOI22xp5_ASAP7_75t_L g2640 ( 
.A1(n_1926),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.Y(n_2640)
);

OAI22xp5_ASAP7_75t_L g2641 ( 
.A1(n_1926),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_2641)
);

NOR2xp33_ASAP7_75t_L g2642 ( 
.A(n_2090),
.B(n_135),
.Y(n_2642)
);

INVx3_ASAP7_75t_L g2643 ( 
.A(n_2182),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2085),
.Y(n_2644)
);

OAI22xp5_ASAP7_75t_L g2645 ( 
.A1(n_1926),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.Y(n_2645)
);

INVx2_ASAP7_75t_L g2646 ( 
.A(n_1926),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2085),
.Y(n_2647)
);

NAND2xp5_ASAP7_75t_L g2648 ( 
.A(n_2085),
.B(n_138),
.Y(n_2648)
);

HB1xp67_ASAP7_75t_L g2649 ( 
.A(n_1926),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_2085),
.B(n_139),
.Y(n_2650)
);

OAI21xp5_ASAP7_75t_L g2651 ( 
.A1(n_1971),
.A2(n_140),
.B(n_141),
.Y(n_2651)
);

AOI21x1_ASAP7_75t_L g2652 ( 
.A1(n_2133),
.A2(n_141),
.B(n_142),
.Y(n_2652)
);

AOI21xp5_ASAP7_75t_L g2653 ( 
.A1(n_1926),
.A2(n_142),
.B(n_143),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2085),
.B(n_142),
.Y(n_2654)
);

O2A1O1Ixp33_ASAP7_75t_L g2655 ( 
.A1(n_2062),
.A2(n_145),
.B(n_143),
.C(n_144),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_L g2656 ( 
.A(n_2085),
.B(n_144),
.Y(n_2656)
);

AOI21xp5_ASAP7_75t_L g2657 ( 
.A1(n_1926),
.A2(n_145),
.B(n_146),
.Y(n_2657)
);

AOI21xp5_ASAP7_75t_L g2658 ( 
.A1(n_1926),
.A2(n_145),
.B(n_146),
.Y(n_2658)
);

AOI21xp5_ASAP7_75t_L g2659 ( 
.A1(n_1926),
.A2(n_146),
.B(n_147),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_SL g2660 ( 
.A(n_1926),
.B(n_147),
.Y(n_2660)
);

AOI21xp5_ASAP7_75t_L g2661 ( 
.A1(n_1926),
.A2(n_148),
.B(n_149),
.Y(n_2661)
);

AND2x6_ASAP7_75t_L g2662 ( 
.A(n_1926),
.B(n_149),
.Y(n_2662)
);

AOI22xp5_ASAP7_75t_L g2663 ( 
.A1(n_1926),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_SL g2664 ( 
.A(n_1926),
.B(n_148),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_1926),
.Y(n_2665)
);

AOI21xp5_ASAP7_75t_L g2666 ( 
.A1(n_1926),
.A2(n_150),
.B(n_152),
.Y(n_2666)
);

NOR2xp33_ASAP7_75t_L g2667 ( 
.A(n_2090),
.B(n_150),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2085),
.Y(n_2668)
);

OAI22xp5_ASAP7_75t_L g2669 ( 
.A1(n_1926),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_2669)
);

A2O1A1Ixp33_ASAP7_75t_L g2670 ( 
.A1(n_2090),
.A2(n_155),
.B(n_153),
.C(n_154),
.Y(n_2670)
);

HB1xp67_ASAP7_75t_L g2671 ( 
.A(n_1926),
.Y(n_2671)
);

INVx2_ASAP7_75t_L g2672 ( 
.A(n_1926),
.Y(n_2672)
);

NOR2xp33_ASAP7_75t_L g2673 ( 
.A(n_2090),
.B(n_153),
.Y(n_2673)
);

OAI21xp5_ASAP7_75t_L g2674 ( 
.A1(n_1971),
.A2(n_154),
.B(n_155),
.Y(n_2674)
);

A2O1A1Ixp33_ASAP7_75t_L g2675 ( 
.A1(n_2090),
.A2(n_157),
.B(n_155),
.C(n_156),
.Y(n_2675)
);

NOR2xp33_ASAP7_75t_R g2676 ( 
.A(n_2198),
.B(n_156),
.Y(n_2676)
);

AOI22xp5_ASAP7_75t_L g2677 ( 
.A1(n_1926),
.A2(n_158),
.B1(n_156),
.B2(n_157),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2085),
.B(n_158),
.Y(n_2678)
);

OAI21xp5_ASAP7_75t_L g2679 ( 
.A1(n_1971),
.A2(n_158),
.B(n_159),
.Y(n_2679)
);

AOI21xp5_ASAP7_75t_L g2680 ( 
.A1(n_1926),
.A2(n_159),
.B(n_160),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_SL g2681 ( 
.A(n_1926),
.B(n_160),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_2085),
.B(n_160),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_SL g2683 ( 
.A(n_2483),
.B(n_424),
.Y(n_2683)
);

AND2x2_ASAP7_75t_L g2684 ( 
.A(n_2255),
.B(n_161),
.Y(n_2684)
);

OAI22x1_ASAP7_75t_L g2685 ( 
.A1(n_2485),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.Y(n_2685)
);

AOI21xp33_ASAP7_75t_L g2686 ( 
.A1(n_2392),
.A2(n_162),
.B(n_163),
.Y(n_2686)
);

INVxp67_ASAP7_75t_SL g2687 ( 
.A(n_2584),
.Y(n_2687)
);

INVx1_ASAP7_75t_SL g2688 ( 
.A(n_2595),
.Y(n_2688)
);

INVx2_ASAP7_75t_SL g2689 ( 
.A(n_2326),
.Y(n_2689)
);

NAND2x1p5_ASAP7_75t_L g2690 ( 
.A(n_2326),
.B(n_2483),
.Y(n_2690)
);

A2O1A1Ixp33_ASAP7_75t_L g2691 ( 
.A1(n_2322),
.A2(n_165),
.B(n_163),
.C(n_164),
.Y(n_2691)
);

AOI21xp5_ASAP7_75t_L g2692 ( 
.A1(n_2283),
.A2(n_164),
.B(n_165),
.Y(n_2692)
);

AOI22xp5_ASAP7_75t_L g2693 ( 
.A1(n_2584),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_2693)
);

AOI21xp5_ASAP7_75t_L g2694 ( 
.A1(n_2635),
.A2(n_166),
.B(n_167),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2293),
.B(n_166),
.Y(n_2695)
);

NAND3xp33_ASAP7_75t_SL g2696 ( 
.A(n_2676),
.B(n_167),
.C(n_168),
.Y(n_2696)
);

AOI21xp5_ASAP7_75t_L g2697 ( 
.A1(n_2646),
.A2(n_168),
.B(n_169),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_2665),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2256),
.Y(n_2699)
);

NAND2x1p5_ASAP7_75t_L g2700 ( 
.A(n_2349),
.B(n_168),
.Y(n_2700)
);

INVx4_ASAP7_75t_L g2701 ( 
.A(n_2406),
.Y(n_2701)
);

HB1xp67_ASAP7_75t_L g2702 ( 
.A(n_2288),
.Y(n_2702)
);

NOR2xp33_ASAP7_75t_SL g2703 ( 
.A(n_2308),
.B(n_169),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_SL g2704 ( 
.A(n_2298),
.B(n_425),
.Y(n_2704)
);

AOI21xp5_ASAP7_75t_L g2705 ( 
.A1(n_2672),
.A2(n_170),
.B(n_171),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2240),
.B(n_170),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2258),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2601),
.B(n_171),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2601),
.B(n_171),
.Y(n_2709)
);

A2O1A1Ixp33_ASAP7_75t_L g2710 ( 
.A1(n_2300),
.A2(n_174),
.B(n_172),
.C(n_173),
.Y(n_2710)
);

AOI22xp33_ASAP7_75t_L g2711 ( 
.A1(n_2314),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2263),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2649),
.B(n_174),
.Y(n_2713)
);

A2O1A1Ixp33_ASAP7_75t_L g2714 ( 
.A1(n_2300),
.A2(n_177),
.B(n_175),
.C(n_176),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_SL g2715 ( 
.A(n_2298),
.B(n_426),
.Y(n_2715)
);

AOI21xp5_ASAP7_75t_L g2716 ( 
.A1(n_2649),
.A2(n_175),
.B(n_176),
.Y(n_2716)
);

INVxp67_ASAP7_75t_L g2717 ( 
.A(n_2605),
.Y(n_2717)
);

OAI22x1_ASAP7_75t_L g2718 ( 
.A1(n_2348),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_2718)
);

OAI22xp5_ASAP7_75t_L g2719 ( 
.A1(n_2671),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.Y(n_2719)
);

NOR2xp33_ASAP7_75t_L g2720 ( 
.A(n_2549),
.B(n_178),
.Y(n_2720)
);

AOI21xp5_ASAP7_75t_L g2721 ( 
.A1(n_2671),
.A2(n_178),
.B(n_179),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2282),
.Y(n_2722)
);

NOR2x1_ASAP7_75t_L g2723 ( 
.A(n_2422),
.B(n_180),
.Y(n_2723)
);

OAI21xp5_ASAP7_75t_L g2724 ( 
.A1(n_2260),
.A2(n_180),
.B(n_181),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2591),
.B(n_181),
.Y(n_2725)
);

AOI21xp5_ASAP7_75t_L g2726 ( 
.A1(n_2290),
.A2(n_182),
.B(n_183),
.Y(n_2726)
);

A2O1A1Ixp33_ASAP7_75t_L g2727 ( 
.A1(n_2342),
.A2(n_185),
.B(n_183),
.C(n_184),
.Y(n_2727)
);

NOR2xp33_ASAP7_75t_L g2728 ( 
.A(n_2358),
.B(n_183),
.Y(n_2728)
);

INVx4_ASAP7_75t_L g2729 ( 
.A(n_2394),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_L g2730 ( 
.A(n_2634),
.B(n_184),
.Y(n_2730)
);

BUFx6f_ASAP7_75t_L g2731 ( 
.A(n_2252),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2301),
.Y(n_2732)
);

AOI21xp5_ASAP7_75t_L g2733 ( 
.A1(n_2316),
.A2(n_184),
.B(n_185),
.Y(n_2733)
);

CKINVDCx5p33_ASAP7_75t_R g2734 ( 
.A(n_2627),
.Y(n_2734)
);

CKINVDCx20_ASAP7_75t_R g2735 ( 
.A(n_2676),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2639),
.B(n_186),
.Y(n_2736)
);

AOI22xp5_ASAP7_75t_L g2737 ( 
.A1(n_2556),
.A2(n_188),
.B1(n_186),
.B2(n_187),
.Y(n_2737)
);

AOI21xp5_ASAP7_75t_L g2738 ( 
.A1(n_2387),
.A2(n_187),
.B(n_189),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2341),
.Y(n_2739)
);

A2O1A1Ixp33_ASAP7_75t_L g2740 ( 
.A1(n_2342),
.A2(n_190),
.B(n_187),
.C(n_189),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2245),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2248),
.Y(n_2742)
);

OAI22xp5_ASAP7_75t_L g2743 ( 
.A1(n_2299),
.A2(n_191),
.B1(n_189),
.B2(n_190),
.Y(n_2743)
);

BUFx6f_ASAP7_75t_L g2744 ( 
.A(n_2252),
.Y(n_2744)
);

AOI21xp5_ASAP7_75t_L g2745 ( 
.A1(n_2389),
.A2(n_190),
.B(n_191),
.Y(n_2745)
);

OAI22xp5_ASAP7_75t_L g2746 ( 
.A1(n_2299),
.A2(n_2588),
.B1(n_2604),
.B2(n_2586),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2271),
.Y(n_2747)
);

AOI21xp5_ASAP7_75t_L g2748 ( 
.A1(n_2376),
.A2(n_191),
.B(n_192),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2273),
.Y(n_2749)
);

O2A1O1Ixp33_ASAP7_75t_L g2750 ( 
.A1(n_2449),
.A2(n_194),
.B(n_192),
.C(n_193),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2644),
.B(n_192),
.Y(n_2751)
);

OAI22xp5_ASAP7_75t_SL g2752 ( 
.A1(n_2556),
.A2(n_2436),
.B1(n_2561),
.B2(n_2447),
.Y(n_2752)
);

INVx3_ASAP7_75t_L g2753 ( 
.A(n_2345),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2281),
.Y(n_2754)
);

OR2x2_ASAP7_75t_L g2755 ( 
.A(n_2323),
.B(n_193),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_2647),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2668),
.B(n_193),
.Y(n_2757)
);

BUFx2_ASAP7_75t_L g2758 ( 
.A(n_2336),
.Y(n_2758)
);

AOI21xp5_ASAP7_75t_L g2759 ( 
.A1(n_2303),
.A2(n_194),
.B(n_195),
.Y(n_2759)
);

INVx4_ASAP7_75t_L g2760 ( 
.A(n_2589),
.Y(n_2760)
);

AND2x4_ASAP7_75t_L g2761 ( 
.A(n_2287),
.B(n_196),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2320),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2586),
.B(n_196),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2334),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_2588),
.B(n_196),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2359),
.Y(n_2766)
);

INVx4_ASAP7_75t_L g2767 ( 
.A(n_2590),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2373),
.Y(n_2768)
);

OAI22xp5_ASAP7_75t_R g2769 ( 
.A1(n_2458),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.Y(n_2769)
);

HB1xp67_ASAP7_75t_L g2770 ( 
.A(n_2286),
.Y(n_2770)
);

AND2x4_ASAP7_75t_L g2771 ( 
.A(n_2287),
.B(n_198),
.Y(n_2771)
);

BUFx2_ASAP7_75t_L g2772 ( 
.A(n_2336),
.Y(n_2772)
);

OAI22xp5_ASAP7_75t_L g2773 ( 
.A1(n_2604),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.Y(n_2773)
);

AOI21xp5_ASAP7_75t_L g2774 ( 
.A1(n_2243),
.A2(n_200),
.B(n_201),
.Y(n_2774)
);

AOI21xp5_ASAP7_75t_L g2775 ( 
.A1(n_2243),
.A2(n_201),
.B(n_202),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_L g2776 ( 
.A(n_2615),
.B(n_202),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_SL g2777 ( 
.A(n_2250),
.B(n_427),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2378),
.Y(n_2778)
);

OR2x6_ASAP7_75t_SL g2779 ( 
.A(n_2461),
.B(n_203),
.Y(n_2779)
);

OA21x2_ASAP7_75t_L g2780 ( 
.A1(n_2438),
.A2(n_2362),
.B(n_2361),
.Y(n_2780)
);

A2O1A1Ixp33_ASAP7_75t_L g2781 ( 
.A1(n_2615),
.A2(n_205),
.B(n_203),
.C(n_204),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_L g2782 ( 
.A(n_2617),
.B(n_204),
.Y(n_2782)
);

BUFx2_ASAP7_75t_L g2783 ( 
.A(n_2662),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_L g2784 ( 
.A(n_2642),
.B(n_205),
.Y(n_2784)
);

INVx6_ASAP7_75t_L g2785 ( 
.A(n_2367),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2456),
.Y(n_2786)
);

A2O1A1Ixp33_ASAP7_75t_SL g2787 ( 
.A1(n_2328),
.A2(n_208),
.B(n_206),
.C(n_207),
.Y(n_2787)
);

AND2x4_ASAP7_75t_L g2788 ( 
.A(n_2396),
.B(n_206),
.Y(n_2788)
);

OR2x2_ASAP7_75t_L g2789 ( 
.A(n_2539),
.B(n_206),
.Y(n_2789)
);

BUFx6f_ASAP7_75t_L g2790 ( 
.A(n_2252),
.Y(n_2790)
);

NOR2xp33_ASAP7_75t_R g2791 ( 
.A(n_2557),
.B(n_207),
.Y(n_2791)
);

AOI21xp5_ASAP7_75t_L g2792 ( 
.A1(n_2291),
.A2(n_208),
.B(n_209),
.Y(n_2792)
);

AOI21xp33_ASAP7_75t_L g2793 ( 
.A1(n_2262),
.A2(n_209),
.B(n_210),
.Y(n_2793)
);

AOI21xp5_ASAP7_75t_L g2794 ( 
.A1(n_2277),
.A2(n_209),
.B(n_210),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2492),
.Y(n_2795)
);

INVx2_ASAP7_75t_L g2796 ( 
.A(n_2343),
.Y(n_2796)
);

AND2x4_ASAP7_75t_L g2797 ( 
.A(n_2345),
.B(n_210),
.Y(n_2797)
);

INVx2_ASAP7_75t_SL g2798 ( 
.A(n_2367),
.Y(n_2798)
);

BUFx2_ASAP7_75t_L g2799 ( 
.A(n_2662),
.Y(n_2799)
);

BUFx2_ASAP7_75t_L g2800 ( 
.A(n_2662),
.Y(n_2800)
);

AOI21xp5_ASAP7_75t_L g2801 ( 
.A1(n_2280),
.A2(n_211),
.B(n_212),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_SL g2802 ( 
.A(n_2391),
.B(n_2241),
.Y(n_2802)
);

AND3x1_ASAP7_75t_SL g2803 ( 
.A(n_2504),
.B(n_211),
.C(n_212),
.Y(n_2803)
);

INVx6_ASAP7_75t_L g2804 ( 
.A(n_2367),
.Y(n_2804)
);

AOI21xp5_ASAP7_75t_L g2805 ( 
.A1(n_2284),
.A2(n_211),
.B(n_212),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2642),
.B(n_213),
.Y(n_2806)
);

NOR2xp33_ASAP7_75t_L g2807 ( 
.A(n_2249),
.B(n_213),
.Y(n_2807)
);

A2O1A1Ixp33_ASAP7_75t_L g2808 ( 
.A1(n_2667),
.A2(n_216),
.B(n_214),
.C(n_215),
.Y(n_2808)
);

AOI22x1_ASAP7_75t_L g2809 ( 
.A1(n_2403),
.A2(n_2437),
.B1(n_2421),
.B2(n_2427),
.Y(n_2809)
);

BUFx6f_ASAP7_75t_L g2810 ( 
.A(n_2252),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_SL g2811 ( 
.A(n_2391),
.B(n_428),
.Y(n_2811)
);

INVx4_ASAP7_75t_L g2812 ( 
.A(n_2528),
.Y(n_2812)
);

A2O1A1Ixp33_ASAP7_75t_L g2813 ( 
.A1(n_2667),
.A2(n_216),
.B(n_214),
.C(n_215),
.Y(n_2813)
);

INVx3_ASAP7_75t_L g2814 ( 
.A(n_2385),
.Y(n_2814)
);

NOR2xp33_ASAP7_75t_L g2815 ( 
.A(n_2268),
.B(n_215),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_2673),
.B(n_217),
.Y(n_2816)
);

AOI21xp5_ASAP7_75t_L g2817 ( 
.A1(n_2257),
.A2(n_218),
.B(n_219),
.Y(n_2817)
);

A2O1A1Ixp33_ASAP7_75t_L g2818 ( 
.A1(n_2673),
.A2(n_220),
.B(n_218),
.C(n_219),
.Y(n_2818)
);

AOI22xp5_ASAP7_75t_L g2819 ( 
.A1(n_2662),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.Y(n_2819)
);

AOI21x1_ASAP7_75t_L g2820 ( 
.A1(n_2353),
.A2(n_220),
.B(n_223),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2624),
.Y(n_2821)
);

INVx2_ASAP7_75t_SL g2822 ( 
.A(n_2540),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2419),
.Y(n_2823)
);

O2A1O1Ixp33_ASAP7_75t_L g2824 ( 
.A1(n_2325),
.A2(n_225),
.B(n_223),
.C(n_224),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_SL g2825 ( 
.A(n_2241),
.B(n_428),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_L g2826 ( 
.A(n_2423),
.B(n_223),
.Y(n_2826)
);

OAI22xp5_ASAP7_75t_L g2827 ( 
.A1(n_2244),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.Y(n_2827)
);

O2A1O1Ixp33_ASAP7_75t_L g2828 ( 
.A1(n_2426),
.A2(n_227),
.B(n_225),
.C(n_226),
.Y(n_2828)
);

CKINVDCx5p33_ASAP7_75t_R g2829 ( 
.A(n_2528),
.Y(n_2829)
);

NOR2xp33_ASAP7_75t_L g2830 ( 
.A(n_2390),
.B(n_226),
.Y(n_2830)
);

OAI21xp5_ASAP7_75t_L g2831 ( 
.A1(n_2310),
.A2(n_227),
.B(n_228),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_SL g2832 ( 
.A(n_2286),
.B(n_429),
.Y(n_2832)
);

HB1xp67_ASAP7_75t_L g2833 ( 
.A(n_2489),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_SL g2834 ( 
.A(n_2488),
.B(n_429),
.Y(n_2834)
);

NOR2xp33_ASAP7_75t_L g2835 ( 
.A(n_2390),
.B(n_227),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_L g2836 ( 
.A(n_2317),
.B(n_228),
.Y(n_2836)
);

AOI21xp5_ASAP7_75t_L g2837 ( 
.A1(n_2371),
.A2(n_229),
.B(n_230),
.Y(n_2837)
);

AOI21xp5_ASAP7_75t_L g2838 ( 
.A1(n_2242),
.A2(n_229),
.B(n_230),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2314),
.B(n_231),
.Y(n_2839)
);

INVx2_ASAP7_75t_L g2840 ( 
.A(n_2351),
.Y(n_2840)
);

AOI21xp5_ASAP7_75t_L g2841 ( 
.A1(n_2505),
.A2(n_231),
.B(n_232),
.Y(n_2841)
);

O2A1O1Ixp33_ASAP7_75t_L g2842 ( 
.A1(n_2515),
.A2(n_2484),
.B(n_2516),
.C(n_2455),
.Y(n_2842)
);

INVx3_ASAP7_75t_L g2843 ( 
.A(n_2385),
.Y(n_2843)
);

AND2x4_ASAP7_75t_SL g2844 ( 
.A(n_2575),
.B(n_232),
.Y(n_2844)
);

A2O1A1Ixp33_ASAP7_75t_L g2845 ( 
.A1(n_2405),
.A2(n_235),
.B(n_233),
.C(n_234),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2425),
.Y(n_2846)
);

A2O1A1Ixp33_ASAP7_75t_L g2847 ( 
.A1(n_2405),
.A2(n_235),
.B(n_233),
.C(n_234),
.Y(n_2847)
);

BUFx2_ASAP7_75t_L g2848 ( 
.A(n_2662),
.Y(n_2848)
);

OAI22xp5_ASAP7_75t_L g2849 ( 
.A1(n_2407),
.A2(n_2420),
.B1(n_2415),
.B2(n_2365),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2340),
.Y(n_2850)
);

HB1xp67_ASAP7_75t_L g2851 ( 
.A(n_2489),
.Y(n_2851)
);

CKINVDCx10_ASAP7_75t_R g2852 ( 
.A(n_2540),
.Y(n_2852)
);

AOI21xp5_ASAP7_75t_L g2853 ( 
.A1(n_2246),
.A2(n_236),
.B(n_237),
.Y(n_2853)
);

A2O1A1Ixp33_ASAP7_75t_L g2854 ( 
.A1(n_2368),
.A2(n_238),
.B(n_236),
.C(n_237),
.Y(n_2854)
);

O2A1O1Ixp33_ASAP7_75t_L g2855 ( 
.A1(n_2484),
.A2(n_240),
.B(n_238),
.C(n_239),
.Y(n_2855)
);

HB1xp67_ASAP7_75t_L g2856 ( 
.A(n_2441),
.Y(n_2856)
);

O2A1O1Ixp5_ASAP7_75t_L g2857 ( 
.A1(n_2353),
.A2(n_2416),
.B(n_2356),
.C(n_2333),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_L g2858 ( 
.A(n_2365),
.B(n_239),
.Y(n_2858)
);

AOI21xp5_ASAP7_75t_L g2859 ( 
.A1(n_2315),
.A2(n_239),
.B(n_240),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2393),
.B(n_241),
.Y(n_2860)
);

BUFx6f_ASAP7_75t_L g2861 ( 
.A(n_2379),
.Y(n_2861)
);

O2A1O1Ixp33_ASAP7_75t_L g2862 ( 
.A1(n_2329),
.A2(n_244),
.B(n_242),
.C(n_243),
.Y(n_2862)
);

CKINVDCx20_ASAP7_75t_R g2863 ( 
.A(n_2519),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_2393),
.B(n_243),
.Y(n_2864)
);

NOR2xp33_ASAP7_75t_L g2865 ( 
.A(n_2404),
.B(n_243),
.Y(n_2865)
);

CKINVDCx5p33_ASAP7_75t_R g2866 ( 
.A(n_2536),
.Y(n_2866)
);

AOI21xp5_ASAP7_75t_L g2867 ( 
.A1(n_2318),
.A2(n_244),
.B(n_245),
.Y(n_2867)
);

INVx3_ASAP7_75t_L g2868 ( 
.A(n_2603),
.Y(n_2868)
);

CKINVDCx5p33_ASAP7_75t_R g2869 ( 
.A(n_2575),
.Y(n_2869)
);

OAI22xp5_ASAP7_75t_L g2870 ( 
.A1(n_2407),
.A2(n_246),
.B1(n_244),
.B2(n_245),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_L g2871 ( 
.A(n_2309),
.B(n_245),
.Y(n_2871)
);

AOI21xp5_ASAP7_75t_L g2872 ( 
.A1(n_2397),
.A2(n_247),
.B(n_248),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2355),
.Y(n_2873)
);

AOI21xp5_ASAP7_75t_L g2874 ( 
.A1(n_2276),
.A2(n_247),
.B(n_249),
.Y(n_2874)
);

NAND2x1p5_ASAP7_75t_L g2875 ( 
.A(n_2319),
.B(n_247),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2487),
.B(n_2328),
.Y(n_2876)
);

INVx3_ASAP7_75t_L g2877 ( 
.A(n_2603),
.Y(n_2877)
);

AOI21xp5_ASAP7_75t_L g2878 ( 
.A1(n_2354),
.A2(n_250),
.B(n_252),
.Y(n_2878)
);

OAI22x1_ASAP7_75t_L g2879 ( 
.A1(n_2441),
.A2(n_253),
.B1(n_250),
.B2(n_252),
.Y(n_2879)
);

BUFx4f_ASAP7_75t_L g2880 ( 
.A(n_2596),
.Y(n_2880)
);

BUFx6f_ASAP7_75t_L g2881 ( 
.A(n_2379),
.Y(n_2881)
);

BUFx2_ASAP7_75t_L g2882 ( 
.A(n_2506),
.Y(n_2882)
);

OAI22xp5_ASAP7_75t_L g2883 ( 
.A1(n_2415),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_2883)
);

OAI22xp5_ASAP7_75t_L g2884 ( 
.A1(n_2420),
.A2(n_256),
.B1(n_254),
.B2(n_255),
.Y(n_2884)
);

CKINVDCx10_ASAP7_75t_R g2885 ( 
.A(n_2460),
.Y(n_2885)
);

OAI22xp5_ASAP7_75t_SL g2886 ( 
.A1(n_2561),
.A2(n_257),
.B1(n_255),
.B2(n_256),
.Y(n_2886)
);

A2O1A1Ixp33_ASAP7_75t_L g2887 ( 
.A1(n_2368),
.A2(n_258),
.B(n_256),
.C(n_257),
.Y(n_2887)
);

AOI21xp5_ASAP7_75t_L g2888 ( 
.A1(n_2366),
.A2(n_257),
.B(n_258),
.Y(n_2888)
);

INVx2_ASAP7_75t_L g2889 ( 
.A(n_2388),
.Y(n_2889)
);

NOR2xp67_ASAP7_75t_L g2890 ( 
.A(n_2413),
.B(n_260),
.Y(n_2890)
);

OAI22xp5_ASAP7_75t_L g2891 ( 
.A1(n_2625),
.A2(n_261),
.B1(n_259),
.B2(n_260),
.Y(n_2891)
);

BUFx2_ASAP7_75t_L g2892 ( 
.A(n_2506),
.Y(n_2892)
);

A2O1A1Ixp33_ASAP7_75t_L g2893 ( 
.A1(n_2360),
.A2(n_262),
.B(n_259),
.C(n_261),
.Y(n_2893)
);

NOR2xp33_ASAP7_75t_R g2894 ( 
.A(n_2306),
.B(n_2613),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_SL g2895 ( 
.A(n_2431),
.B(n_430),
.Y(n_2895)
);

OAI22xp5_ASAP7_75t_L g2896 ( 
.A1(n_2625),
.A2(n_262),
.B1(n_259),
.B2(n_261),
.Y(n_2896)
);

BUFx2_ASAP7_75t_L g2897 ( 
.A(n_2596),
.Y(n_2897)
);

A2O1A1Ixp33_ASAP7_75t_L g2898 ( 
.A1(n_2360),
.A2(n_264),
.B(n_262),
.C(n_263),
.Y(n_2898)
);

INVx3_ASAP7_75t_L g2899 ( 
.A(n_2613),
.Y(n_2899)
);

INVxp67_ASAP7_75t_L g2900 ( 
.A(n_2372),
.Y(n_2900)
);

AND3x1_ASAP7_75t_SL g2901 ( 
.A(n_2558),
.B(n_263),
.C(n_264),
.Y(n_2901)
);

OAI22xp5_ASAP7_75t_L g2902 ( 
.A1(n_2682),
.A2(n_266),
.B1(n_264),
.B2(n_265),
.Y(n_2902)
);

INVx1_ASAP7_75t_SL g2903 ( 
.A(n_2636),
.Y(n_2903)
);

BUFx6f_ASAP7_75t_L g2904 ( 
.A(n_2379),
.Y(n_2904)
);

HB1xp67_ASAP7_75t_L g2905 ( 
.A(n_2498),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2587),
.Y(n_2906)
);

OAI22xp5_ASAP7_75t_SL g2907 ( 
.A1(n_2327),
.A2(n_2523),
.B1(n_2418),
.B2(n_2543),
.Y(n_2907)
);

AOI21xp5_ASAP7_75t_L g2908 ( 
.A1(n_2330),
.A2(n_266),
.B(n_268),
.Y(n_2908)
);

OR2x6_ASAP7_75t_SL g2909 ( 
.A(n_2471),
.B(n_269),
.Y(n_2909)
);

AOI21xp5_ASAP7_75t_L g2910 ( 
.A1(n_2270),
.A2(n_269),
.B(n_270),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2600),
.Y(n_2911)
);

AND2x2_ASAP7_75t_L g2912 ( 
.A(n_2510),
.B(n_270),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_SL g2913 ( 
.A(n_2370),
.B(n_431),
.Y(n_2913)
);

INVx2_ASAP7_75t_L g2914 ( 
.A(n_2402),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2335),
.B(n_271),
.Y(n_2915)
);

CKINVDCx5p33_ASAP7_75t_R g2916 ( 
.A(n_2369),
.Y(n_2916)
);

INVx3_ASAP7_75t_L g2917 ( 
.A(n_2620),
.Y(n_2917)
);

AOI21xp5_ASAP7_75t_L g2918 ( 
.A1(n_2251),
.A2(n_271),
.B(n_272),
.Y(n_2918)
);

AOI22xp5_ASAP7_75t_L g2919 ( 
.A1(n_2523),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_SL g2920 ( 
.A(n_2498),
.B(n_431),
.Y(n_2920)
);

AOI21xp5_ASAP7_75t_L g2921 ( 
.A1(n_2509),
.A2(n_272),
.B(n_273),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_SL g2922 ( 
.A(n_2514),
.B(n_432),
.Y(n_2922)
);

A2O1A1Ixp33_ASAP7_75t_L g2923 ( 
.A1(n_2363),
.A2(n_276),
.B(n_274),
.C(n_275),
.Y(n_2923)
);

HB1xp67_ASAP7_75t_L g2924 ( 
.A(n_2514),
.Y(n_2924)
);

A2O1A1Ixp33_ASAP7_75t_L g2925 ( 
.A1(n_2363),
.A2(n_276),
.B(n_274),
.C(n_275),
.Y(n_2925)
);

OAI22xp5_ASAP7_75t_L g2926 ( 
.A1(n_2602),
.A2(n_277),
.B1(n_275),
.B2(n_276),
.Y(n_2926)
);

O2A1O1Ixp5_ASAP7_75t_L g2927 ( 
.A1(n_2416),
.A2(n_279),
.B(n_277),
.C(n_278),
.Y(n_2927)
);

INVx3_ASAP7_75t_L g2928 ( 
.A(n_2620),
.Y(n_2928)
);

BUFx6f_ASAP7_75t_L g2929 ( 
.A(n_2379),
.Y(n_2929)
);

OAI22xp5_ASAP7_75t_L g2930 ( 
.A1(n_2609),
.A2(n_280),
.B1(n_278),
.B2(n_279),
.Y(n_2930)
);

NOR2xp33_ASAP7_75t_L g2931 ( 
.A(n_2272),
.B(n_278),
.Y(n_2931)
);

A2O1A1Ixp33_ASAP7_75t_L g2932 ( 
.A1(n_2267),
.A2(n_281),
.B(n_279),
.C(n_280),
.Y(n_2932)
);

AOI21xp5_ASAP7_75t_L g2933 ( 
.A1(n_2296),
.A2(n_280),
.B(n_281),
.Y(n_2933)
);

INVx3_ASAP7_75t_SL g2934 ( 
.A(n_2582),
.Y(n_2934)
);

INVx8_ASAP7_75t_L g2935 ( 
.A(n_2643),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_2335),
.B(n_281),
.Y(n_2936)
);

NAND3xp33_ASAP7_75t_SL g2937 ( 
.A(n_2460),
.B(n_282),
.C(n_283),
.Y(n_2937)
);

OAI21xp33_ASAP7_75t_L g2938 ( 
.A1(n_2628),
.A2(n_284),
.B(n_285),
.Y(n_2938)
);

BUFx6f_ASAP7_75t_SL g2939 ( 
.A(n_2295),
.Y(n_2939)
);

AOI21xp5_ASAP7_75t_L g2940 ( 
.A1(n_2297),
.A2(n_284),
.B(n_285),
.Y(n_2940)
);

OAI22xp5_ASAP7_75t_L g2941 ( 
.A1(n_2614),
.A2(n_288),
.B1(n_286),
.B2(n_287),
.Y(n_2941)
);

BUFx8_ASAP7_75t_SL g2942 ( 
.A(n_2552),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2324),
.B(n_286),
.Y(n_2943)
);

AOI21xp5_ASAP7_75t_L g2944 ( 
.A1(n_2254),
.A2(n_286),
.B(n_287),
.Y(n_2944)
);

NOR2xp33_ASAP7_75t_L g2945 ( 
.A(n_2275),
.B(n_287),
.Y(n_2945)
);

AND2x2_ASAP7_75t_L g2946 ( 
.A(n_2443),
.B(n_288),
.Y(n_2946)
);

CKINVDCx5p33_ASAP7_75t_R g2947 ( 
.A(n_2513),
.Y(n_2947)
);

BUFx6f_ASAP7_75t_L g2948 ( 
.A(n_2464),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_L g2949 ( 
.A(n_2265),
.B(n_288),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_L g2950 ( 
.A(n_2302),
.B(n_289),
.Y(n_2950)
);

AOI22xp33_ASAP7_75t_L g2951 ( 
.A1(n_2400),
.A2(n_2546),
.B1(n_2513),
.B2(n_2574),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_L g2952 ( 
.A(n_2546),
.B(n_289),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_L g2953 ( 
.A(n_2305),
.B(n_289),
.Y(n_2953)
);

AND2x4_ASAP7_75t_L g2954 ( 
.A(n_2643),
.B(n_290),
.Y(n_2954)
);

OR2x2_ASAP7_75t_L g2955 ( 
.A(n_2289),
.B(n_290),
.Y(n_2955)
);

INVx3_ASAP7_75t_L g2956 ( 
.A(n_2413),
.Y(n_2956)
);

AOI21x1_ASAP7_75t_L g2957 ( 
.A1(n_2333),
.A2(n_290),
.B(n_291),
.Y(n_2957)
);

NOR2xp33_ASAP7_75t_L g2958 ( 
.A(n_2285),
.B(n_291),
.Y(n_2958)
);

O2A1O1Ixp33_ASAP7_75t_L g2959 ( 
.A1(n_2530),
.A2(n_294),
.B(n_292),
.C(n_293),
.Y(n_2959)
);

BUFx6f_ASAP7_75t_L g2960 ( 
.A(n_2464),
.Y(n_2960)
);

AOI21xp5_ASAP7_75t_L g2961 ( 
.A1(n_2542),
.A2(n_292),
.B(n_293),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_SL g2962 ( 
.A(n_2593),
.B(n_433),
.Y(n_2962)
);

INVx3_ASAP7_75t_L g2963 ( 
.A(n_2417),
.Y(n_2963)
);

NOR2xp33_ASAP7_75t_L g2964 ( 
.A(n_2294),
.B(n_292),
.Y(n_2964)
);

AOI22xp33_ASAP7_75t_L g2965 ( 
.A1(n_2400),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_2965)
);

INVx3_ASAP7_75t_L g2966 ( 
.A(n_2417),
.Y(n_2966)
);

OR2x6_ASAP7_75t_L g2967 ( 
.A(n_2253),
.B(n_2381),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_SL g2968 ( 
.A(n_2651),
.B(n_2674),
.Y(n_2968)
);

NOR3xp33_ASAP7_75t_L g2969 ( 
.A(n_2551),
.B(n_295),
.C(n_296),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2321),
.B(n_295),
.Y(n_2970)
);

AO22x1_ASAP7_75t_L g2971 ( 
.A1(n_2679),
.A2(n_299),
.B1(n_297),
.B2(n_298),
.Y(n_2971)
);

O2A1O1Ixp5_ASAP7_75t_L g2972 ( 
.A1(n_2347),
.A2(n_2623),
.B(n_2664),
.C(n_2660),
.Y(n_2972)
);

AND2x2_ASAP7_75t_L g2973 ( 
.A(n_2411),
.B(n_297),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_SL g2974 ( 
.A(n_2247),
.B(n_433),
.Y(n_2974)
);

BUFx6f_ASAP7_75t_L g2975 ( 
.A(n_2464),
.Y(n_2975)
);

A2O1A1Ixp33_ASAP7_75t_L g2976 ( 
.A1(n_2267),
.A2(n_299),
.B(n_297),
.C(n_298),
.Y(n_2976)
);

AOI21xp5_ASAP7_75t_L g2977 ( 
.A1(n_2259),
.A2(n_300),
.B(n_301),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_L g2978 ( 
.A(n_2337),
.B(n_300),
.Y(n_2978)
);

INVx5_ASAP7_75t_L g2979 ( 
.A(n_2464),
.Y(n_2979)
);

BUFx8_ASAP7_75t_L g2980 ( 
.A(n_2424),
.Y(n_2980)
);

CKINVDCx16_ASAP7_75t_R g2981 ( 
.A(n_2440),
.Y(n_2981)
);

A2O1A1Ixp33_ASAP7_75t_L g2982 ( 
.A1(n_2463),
.A2(n_302),
.B(n_300),
.C(n_301),
.Y(n_2982)
);

AOI21xp5_ASAP7_75t_L g2983 ( 
.A1(n_2518),
.A2(n_301),
.B(n_303),
.Y(n_2983)
);

AOI22xp5_ASAP7_75t_L g2984 ( 
.A1(n_2571),
.A2(n_305),
.B1(n_303),
.B2(n_304),
.Y(n_2984)
);

NOR2xp33_ASAP7_75t_L g2985 ( 
.A(n_2304),
.B(n_303),
.Y(n_2985)
);

A2O1A1Ixp33_ASAP7_75t_SL g2986 ( 
.A1(n_2548),
.A2(n_307),
.B(n_304),
.C(n_306),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_2313),
.B(n_304),
.Y(n_2987)
);

OAI22xp5_ASAP7_75t_L g2988 ( 
.A1(n_2616),
.A2(n_308),
.B1(n_306),
.B2(n_307),
.Y(n_2988)
);

AOI21xp5_ASAP7_75t_L g2989 ( 
.A1(n_2347),
.A2(n_308),
.B(n_309),
.Y(n_2989)
);

O2A1O1Ixp33_ASAP7_75t_SL g2990 ( 
.A1(n_2521),
.A2(n_310),
.B(n_308),
.C(n_309),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_SL g2991 ( 
.A(n_2448),
.B(n_434),
.Y(n_2991)
);

A2O1A1Ixp33_ASAP7_75t_L g2992 ( 
.A1(n_2481),
.A2(n_311),
.B(n_309),
.C(n_310),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_2331),
.B(n_310),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2468),
.B(n_311),
.Y(n_2994)
);

HB1xp67_ASAP7_75t_L g2995 ( 
.A(n_2537),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2433),
.Y(n_2996)
);

INVx2_ASAP7_75t_L g2997 ( 
.A(n_2476),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_SL g2998 ( 
.A(n_2520),
.B(n_434),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2408),
.B(n_311),
.Y(n_2999)
);

BUFx6f_ASAP7_75t_L g3000 ( 
.A(n_2520),
.Y(n_3000)
);

NOR2xp33_ASAP7_75t_L g3001 ( 
.A(n_2307),
.B(n_312),
.Y(n_3001)
);

NAND2x1_ASAP7_75t_SL g3002 ( 
.A(n_2621),
.B(n_312),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2311),
.B(n_312),
.Y(n_3003)
);

OAI22xp5_ASAP7_75t_SL g3004 ( 
.A1(n_2543),
.A2(n_315),
.B1(n_313),
.B2(n_314),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_2502),
.B(n_315),
.Y(n_3005)
);

INVx4_ASAP7_75t_L g3006 ( 
.A(n_2435),
.Y(n_3006)
);

AND2x4_ASAP7_75t_L g3007 ( 
.A(n_2517),
.B(n_316),
.Y(n_3007)
);

AND2x4_ASAP7_75t_L g3008 ( 
.A(n_2529),
.B(n_2533),
.Y(n_3008)
);

NOR2xp33_ASAP7_75t_L g3009 ( 
.A(n_2278),
.B(n_316),
.Y(n_3009)
);

AOI22xp33_ASAP7_75t_L g3010 ( 
.A1(n_2574),
.A2(n_2398),
.B1(n_2571),
.B2(n_2507),
.Y(n_3010)
);

OAI22xp5_ASAP7_75t_L g3011 ( 
.A1(n_2622),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2630),
.Y(n_3012)
);

OAI22xp5_ASAP7_75t_L g3013 ( 
.A1(n_2631),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.Y(n_3013)
);

A2O1A1Ixp33_ASAP7_75t_L g3014 ( 
.A1(n_2490),
.A2(n_320),
.B(n_318),
.C(n_319),
.Y(n_3014)
);

AOI21x1_ASAP7_75t_L g3015 ( 
.A1(n_2410),
.A2(n_320),
.B(n_321),
.Y(n_3015)
);

INVx2_ASAP7_75t_L g3016 ( 
.A(n_2477),
.Y(n_3016)
);

AOI21xp5_ASAP7_75t_L g3017 ( 
.A1(n_2375),
.A2(n_321),
.B(n_323),
.Y(n_3017)
);

OAI22xp5_ASAP7_75t_L g3018 ( 
.A1(n_2632),
.A2(n_325),
.B1(n_323),
.B2(n_324),
.Y(n_3018)
);

OAI22xp5_ASAP7_75t_L g3019 ( 
.A1(n_2637),
.A2(n_325),
.B1(n_323),
.B2(n_324),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2638),
.Y(n_3020)
);

NOR2xp33_ASAP7_75t_R g3021 ( 
.A(n_2295),
.B(n_324),
.Y(n_3021)
);

O2A1O1Ixp33_ASAP7_75t_SL g3022 ( 
.A1(n_2623),
.A2(n_327),
.B(n_325),
.C(n_326),
.Y(n_3022)
);

INVx2_ASAP7_75t_L g3023 ( 
.A(n_2486),
.Y(n_3023)
);

NOR2xp33_ASAP7_75t_L g3024 ( 
.A(n_2531),
.B(n_326),
.Y(n_3024)
);

A2O1A1Ixp33_ASAP7_75t_L g3025 ( 
.A1(n_2607),
.A2(n_328),
.B(n_326),
.C(n_327),
.Y(n_3025)
);

INVx2_ASAP7_75t_L g3026 ( 
.A(n_2501),
.Y(n_3026)
);

BUFx10_ASAP7_75t_L g3027 ( 
.A(n_2537),
.Y(n_3027)
);

O2A1O1Ixp33_ASAP7_75t_L g3028 ( 
.A1(n_2473),
.A2(n_330),
.B(n_328),
.C(n_329),
.Y(n_3028)
);

AOI22xp5_ASAP7_75t_L g3029 ( 
.A1(n_2619),
.A2(n_331),
.B1(n_329),
.B2(n_330),
.Y(n_3029)
);

AOI22xp5_ASAP7_75t_L g3030 ( 
.A1(n_2660),
.A2(n_332),
.B1(n_329),
.B2(n_331),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2648),
.Y(n_3031)
);

NAND2x1p5_ASAP7_75t_L g3032 ( 
.A(n_2435),
.B(n_331),
.Y(n_3032)
);

O2A1O1Ixp33_ASAP7_75t_SL g3033 ( 
.A1(n_2664),
.A2(n_334),
.B(n_332),
.C(n_333),
.Y(n_3033)
);

OAI22xp5_ASAP7_75t_L g3034 ( 
.A1(n_2650),
.A2(n_337),
.B1(n_335),
.B2(n_336),
.Y(n_3034)
);

OAI22xp5_ASAP7_75t_L g3035 ( 
.A1(n_2654),
.A2(n_337),
.B1(n_335),
.B2(n_336),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_SL g3036 ( 
.A(n_2520),
.B(n_435),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2656),
.B(n_336),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2678),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2567),
.B(n_337),
.Y(n_3039)
);

AOI21xp5_ASAP7_75t_L g3040 ( 
.A1(n_2375),
.A2(n_338),
.B(n_339),
.Y(n_3040)
);

AND2x2_ASAP7_75t_L g3041 ( 
.A(n_2479),
.B(n_338),
.Y(n_3041)
);

INVx5_ASAP7_75t_L g3042 ( 
.A(n_2520),
.Y(n_3042)
);

AOI21xp5_ASAP7_75t_L g3043 ( 
.A1(n_2534),
.A2(n_339),
.B(n_340),
.Y(n_3043)
);

NOR3xp33_ASAP7_75t_SL g3044 ( 
.A(n_2499),
.B(n_340),
.C(n_341),
.Y(n_3044)
);

AND2x2_ASAP7_75t_L g3045 ( 
.A(n_2482),
.B(n_341),
.Y(n_3045)
);

A2O1A1Ixp33_ASAP7_75t_L g3046 ( 
.A1(n_2611),
.A2(n_344),
.B(n_342),
.C(n_343),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2606),
.Y(n_3047)
);

AOI21xp5_ASAP7_75t_L g3048 ( 
.A1(n_2377),
.A2(n_342),
.B(n_343),
.Y(n_3048)
);

OR2x6_ASAP7_75t_L g3049 ( 
.A(n_2395),
.B(n_2414),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_L g3050 ( 
.A(n_2344),
.B(n_344),
.Y(n_3050)
);

AOI21xp5_ASAP7_75t_L g3051 ( 
.A1(n_2380),
.A2(n_344),
.B(n_345),
.Y(n_3051)
);

NAND2xp5_ASAP7_75t_SL g3052 ( 
.A(n_2532),
.B(n_436),
.Y(n_3052)
);

O2A1O1Ixp33_ASAP7_75t_L g3053 ( 
.A1(n_2544),
.A2(n_347),
.B(n_345),
.C(n_346),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_L g3054 ( 
.A(n_2346),
.B(n_345),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2399),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_2357),
.B(n_347),
.Y(n_3056)
);

INVx5_ASAP7_75t_L g3057 ( 
.A(n_2532),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2508),
.Y(n_3058)
);

INVx2_ASAP7_75t_L g3059 ( 
.A(n_2475),
.Y(n_3059)
);

INVxp67_ASAP7_75t_L g3060 ( 
.A(n_2681),
.Y(n_3060)
);

BUFx3_ASAP7_75t_L g3061 ( 
.A(n_2459),
.Y(n_3061)
);

INVx1_ASAP7_75t_SL g3062 ( 
.A(n_2469),
.Y(n_3062)
);

AOI22xp33_ASAP7_75t_L g3063 ( 
.A1(n_2430),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.Y(n_3063)
);

O2A1O1Ixp5_ASAP7_75t_L g3064 ( 
.A1(n_2274),
.A2(n_350),
.B(n_348),
.C(n_349),
.Y(n_3064)
);

O2A1O1Ixp5_ASAP7_75t_SL g3065 ( 
.A1(n_2568),
.A2(n_438),
.B(n_439),
.C(n_436),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_2364),
.B(n_349),
.Y(n_3066)
);

INVxp67_ASAP7_75t_L g3067 ( 
.A(n_2500),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2512),
.Y(n_3068)
);

AO32x2_ASAP7_75t_L g3069 ( 
.A1(n_2886),
.A2(n_2503),
.A3(n_2608),
.B1(n_2629),
.B2(n_2610),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2786),
.Y(n_3070)
);

HB1xp67_ASAP7_75t_L g3071 ( 
.A(n_2702),
.Y(n_3071)
);

O2A1O1Ixp33_ASAP7_75t_L g3072 ( 
.A1(n_2849),
.A2(n_2374),
.B(n_2675),
.C(n_2670),
.Y(n_3072)
);

AO31x2_ASAP7_75t_L g3073 ( 
.A1(n_3059),
.A2(n_2547),
.A3(n_2497),
.B(n_2384),
.Y(n_3073)
);

AO31x2_ASAP7_75t_L g3074 ( 
.A1(n_2746),
.A2(n_2350),
.A3(n_2626),
.B(n_2264),
.Y(n_3074)
);

NOR2xp33_ASAP7_75t_L g3075 ( 
.A(n_2752),
.B(n_2947),
.Y(n_3075)
);

AOI21xp5_ASAP7_75t_L g3076 ( 
.A1(n_2968),
.A2(n_2269),
.B(n_2261),
.Y(n_3076)
);

INVx2_ASAP7_75t_L g3077 ( 
.A(n_2698),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2795),
.Y(n_3078)
);

OAI21x1_ASAP7_75t_L g3079 ( 
.A1(n_2857),
.A2(n_2652),
.B(n_2269),
.Y(n_3079)
);

INVx2_ASAP7_75t_L g3080 ( 
.A(n_2756),
.Y(n_3080)
);

AO22x2_ASAP7_75t_L g3081 ( 
.A1(n_2743),
.A2(n_2669),
.B1(n_2645),
.B2(n_2641),
.Y(n_3081)
);

OAI22xp5_ASAP7_75t_L g3082 ( 
.A1(n_2880),
.A2(n_2541),
.B1(n_2663),
.B2(n_2640),
.Y(n_3082)
);

O2A1O1Ixp33_ASAP7_75t_L g3083 ( 
.A1(n_2787),
.A2(n_2612),
.B(n_2599),
.C(n_2457),
.Y(n_3083)
);

OAI21x1_ASAP7_75t_L g3084 ( 
.A1(n_2809),
.A2(n_2279),
.B(n_2261),
.Y(n_3084)
);

NOR2xp33_ASAP7_75t_SL g3085 ( 
.A(n_2735),
.B(n_2522),
.Y(n_3085)
);

INVx2_ASAP7_75t_L g3086 ( 
.A(n_2699),
.Y(n_3086)
);

BUFx6f_ASAP7_75t_L g3087 ( 
.A(n_2701),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_SL g3088 ( 
.A(n_2880),
.B(n_2493),
.Y(n_3088)
);

AO31x2_ASAP7_75t_L g3089 ( 
.A1(n_2783),
.A2(n_2352),
.A3(n_2452),
.B(n_2633),
.Y(n_3089)
);

AOI21xp5_ASAP7_75t_L g3090 ( 
.A1(n_2780),
.A2(n_2279),
.B(n_2576),
.Y(n_3090)
);

A2O1A1Ixp33_ASAP7_75t_L g3091 ( 
.A1(n_2842),
.A2(n_2655),
.B(n_2618),
.C(n_2559),
.Y(n_3091)
);

AOI21xp5_ASAP7_75t_L g3092 ( 
.A1(n_2780),
.A2(n_2568),
.B(n_2576),
.Y(n_3092)
);

AO31x2_ASAP7_75t_L g3093 ( 
.A1(n_2799),
.A2(n_2666),
.A3(n_2680),
.B(n_2661),
.Y(n_3093)
);

NOR2xp67_ASAP7_75t_L g3094 ( 
.A(n_2701),
.B(n_2677),
.Y(n_3094)
);

AOI21x1_ASAP7_75t_L g3095 ( 
.A1(n_2802),
.A2(n_2524),
.B(n_2462),
.Y(n_3095)
);

BUFx2_ASAP7_75t_L g3096 ( 
.A(n_2980),
.Y(n_3096)
);

OAI21xp5_ASAP7_75t_SL g3097 ( 
.A1(n_2737),
.A2(n_2494),
.B(n_2496),
.Y(n_3097)
);

AO31x2_ASAP7_75t_L g3098 ( 
.A1(n_2800),
.A2(n_2592),
.A3(n_2597),
.B(n_2594),
.Y(n_3098)
);

AO21x1_ASAP7_75t_L g3099 ( 
.A1(n_2704),
.A2(n_2565),
.B(n_2585),
.Y(n_3099)
);

AOI21xp5_ASAP7_75t_L g3100 ( 
.A1(n_2972),
.A2(n_2687),
.B(n_2715),
.Y(n_3100)
);

OAI21xp5_ASAP7_75t_L g3101 ( 
.A1(n_2733),
.A2(n_2312),
.B(n_2491),
.Y(n_3101)
);

AO31x2_ASAP7_75t_L g3102 ( 
.A1(n_2848),
.A2(n_2691),
.A3(n_2838),
.B(n_2692),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2850),
.B(n_2466),
.Y(n_3103)
);

AOI21xp5_ASAP7_75t_L g3104 ( 
.A1(n_2962),
.A2(n_2572),
.B(n_2532),
.Y(n_3104)
);

NOR2xp33_ASAP7_75t_L g3105 ( 
.A(n_2885),
.B(n_2472),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_SL g3106 ( 
.A(n_3021),
.B(n_2532),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2741),
.Y(n_3107)
);

OAI21xp5_ASAP7_75t_L g3108 ( 
.A1(n_2951),
.A2(n_2312),
.B(n_2442),
.Y(n_3108)
);

OAI21xp5_ASAP7_75t_L g3109 ( 
.A1(n_2815),
.A2(n_2446),
.B(n_2445),
.Y(n_3109)
);

AOI21xp5_ASAP7_75t_L g3110 ( 
.A1(n_3049),
.A2(n_2572),
.B(n_2432),
.Y(n_3110)
);

OAI21x1_ASAP7_75t_L g3111 ( 
.A1(n_3015),
.A2(n_2577),
.B(n_2292),
.Y(n_3111)
);

AOI21xp5_ASAP7_75t_L g3112 ( 
.A1(n_3049),
.A2(n_2826),
.B(n_2834),
.Y(n_3112)
);

BUFx4f_ASAP7_75t_L g3113 ( 
.A(n_2690),
.Y(n_3113)
);

O2A1O1Ixp33_ASAP7_75t_L g3114 ( 
.A1(n_3067),
.A2(n_2915),
.B(n_2936),
.C(n_2937),
.Y(n_3114)
);

OAI21xp5_ASAP7_75t_L g3115 ( 
.A1(n_3060),
.A2(n_2474),
.B(n_2553),
.Y(n_3115)
);

AOI221xp5_ASAP7_75t_L g3116 ( 
.A1(n_2686),
.A2(n_2339),
.B1(n_2598),
.B2(n_2467),
.C(n_2465),
.Y(n_3116)
);

OR2x2_ASAP7_75t_L g3117 ( 
.A(n_2688),
.B(n_2478),
.Y(n_3117)
);

BUFx6f_ASAP7_75t_L g3118 ( 
.A(n_2785),
.Y(n_3118)
);

AOI21x1_ASAP7_75t_L g3119 ( 
.A1(n_2897),
.A2(n_2292),
.B(n_2563),
.Y(n_3119)
);

AND2x4_ASAP7_75t_L g3120 ( 
.A(n_2761),
.B(n_2459),
.Y(n_3120)
);

O2A1O1Ixp33_ASAP7_75t_L g3121 ( 
.A1(n_2696),
.A2(n_2555),
.B(n_2554),
.C(n_2383),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_3047),
.B(n_2444),
.Y(n_3122)
);

AOI21xp5_ASAP7_75t_L g3123 ( 
.A1(n_3049),
.A2(n_2967),
.B(n_2793),
.Y(n_3123)
);

NAND2x1p5_ASAP7_75t_L g3124 ( 
.A(n_2760),
.B(n_2480),
.Y(n_3124)
);

AOI21xp5_ASAP7_75t_L g3125 ( 
.A1(n_2967),
.A2(n_2572),
.B(n_2428),
.Y(n_3125)
);

AOI21xp5_ASAP7_75t_L g3126 ( 
.A1(n_2967),
.A2(n_2572),
.B(n_2495),
.Y(n_3126)
);

AOI21x1_ASAP7_75t_L g3127 ( 
.A1(n_2825),
.A2(n_2564),
.B(n_2338),
.Y(n_3127)
);

AND2x2_ASAP7_75t_L g3128 ( 
.A(n_2973),
.B(n_2454),
.Y(n_3128)
);

AO31x2_ASAP7_75t_L g3129 ( 
.A1(n_3043),
.A2(n_2657),
.A3(n_2658),
.B(n_2653),
.Y(n_3129)
);

NOR3xp33_ASAP7_75t_L g3130 ( 
.A(n_2717),
.B(n_2855),
.C(n_2723),
.Y(n_3130)
);

OAI22x1_ASAP7_75t_L g3131 ( 
.A1(n_2819),
.A2(n_2382),
.B1(n_2434),
.B2(n_2578),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_L g3132 ( 
.A(n_2876),
.B(n_2720),
.Y(n_3132)
);

OAI21xp5_ASAP7_75t_L g3133 ( 
.A1(n_2931),
.A2(n_2470),
.B(n_2659),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2903),
.B(n_2545),
.Y(n_3134)
);

OR2x2_ASAP7_75t_L g3135 ( 
.A(n_2789),
.B(n_2526),
.Y(n_3135)
);

OR2x6_ASAP7_75t_L g3136 ( 
.A(n_2729),
.B(n_2450),
.Y(n_3136)
);

NOR2xp33_ASAP7_75t_L g3137 ( 
.A(n_2885),
.B(n_2386),
.Y(n_3137)
);

NOR2xp33_ASAP7_75t_L g3138 ( 
.A(n_2916),
.B(n_2562),
.Y(n_3138)
);

AOI21xp5_ASAP7_75t_L g3139 ( 
.A1(n_2906),
.A2(n_2535),
.B(n_2527),
.Y(n_3139)
);

BUFx3_ASAP7_75t_L g3140 ( 
.A(n_2980),
.Y(n_3140)
);

CKINVDCx5p33_ASAP7_75t_R g3141 ( 
.A(n_2734),
.Y(n_3141)
);

NAND3xp33_ASAP7_75t_SL g3142 ( 
.A(n_2791),
.B(n_2470),
.C(n_2550),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2742),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2747),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_2749),
.B(n_2451),
.Y(n_3145)
);

OAI22xp5_ASAP7_75t_L g3146 ( 
.A1(n_2981),
.A2(n_2570),
.B1(n_2560),
.B2(n_2401),
.Y(n_3146)
);

NOR2xp33_ASAP7_75t_L g3147 ( 
.A(n_2866),
.B(n_2566),
.Y(n_3147)
);

O2A1O1Ixp33_ASAP7_75t_SL g3148 ( 
.A1(n_2781),
.A2(n_2579),
.B(n_2583),
.C(n_2525),
.Y(n_3148)
);

O2A1O1Ixp5_ASAP7_75t_L g3149 ( 
.A1(n_2895),
.A2(n_2971),
.B(n_2974),
.C(n_2913),
.Y(n_3149)
);

AOI22xp5_ASAP7_75t_L g3150 ( 
.A1(n_2907),
.A2(n_2453),
.B1(n_2429),
.B2(n_2511),
.Y(n_3150)
);

AOI21xp5_ASAP7_75t_SL g3151 ( 
.A1(n_2939),
.A2(n_2332),
.B(n_2580),
.Y(n_3151)
);

INVx4_ASAP7_75t_L g3152 ( 
.A(n_2760),
.Y(n_3152)
);

HB1xp67_ASAP7_75t_L g3153 ( 
.A(n_2758),
.Y(n_3153)
);

OAI21x1_ASAP7_75t_L g3154 ( 
.A1(n_2820),
.A2(n_2439),
.B(n_2480),
.Y(n_3154)
);

BUFx3_ASAP7_75t_L g3155 ( 
.A(n_2863),
.Y(n_3155)
);

AOI22xp33_ASAP7_75t_L g3156 ( 
.A1(n_2969),
.A2(n_2573),
.B1(n_2412),
.B2(n_2409),
.Y(n_3156)
);

AOI21xp5_ASAP7_75t_L g3157 ( 
.A1(n_2911),
.A2(n_2581),
.B(n_2266),
.Y(n_3157)
);

NAND2xp5_ASAP7_75t_L g3158 ( 
.A(n_2754),
.B(n_2569),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2762),
.B(n_2401),
.Y(n_3159)
);

OAI21x1_ASAP7_75t_L g3160 ( 
.A1(n_2957),
.A2(n_2538),
.B(n_350),
.Y(n_3160)
);

INVx3_ASAP7_75t_L g3161 ( 
.A(n_2767),
.Y(n_3161)
);

OAI22xp5_ASAP7_75t_L g3162 ( 
.A1(n_2819),
.A2(n_353),
.B1(n_351),
.B2(n_352),
.Y(n_3162)
);

AO31x2_ASAP7_75t_L g3163 ( 
.A1(n_2837),
.A2(n_353),
.A3(n_351),
.B(n_352),
.Y(n_3163)
);

AOI21xp5_ASAP7_75t_L g3164 ( 
.A1(n_3012),
.A2(n_351),
.B(n_353),
.Y(n_3164)
);

INVx2_ASAP7_75t_L g3165 ( 
.A(n_2707),
.Y(n_3165)
);

A2O1A1Ixp33_ASAP7_75t_L g3166 ( 
.A1(n_3053),
.A2(n_356),
.B(n_354),
.C(n_355),
.Y(n_3166)
);

O2A1O1Ixp33_ASAP7_75t_SL g3167 ( 
.A1(n_2808),
.A2(n_356),
.B(n_354),
.C(n_355),
.Y(n_3167)
);

AOI21xp5_ASAP7_75t_L g3168 ( 
.A1(n_3020),
.A2(n_358),
.B(n_359),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2764),
.Y(n_3169)
);

AOI21xp5_ASAP7_75t_L g3170 ( 
.A1(n_3031),
.A2(n_358),
.B(n_359),
.Y(n_3170)
);

NOR2xp33_ASAP7_75t_L g3171 ( 
.A(n_2833),
.B(n_360),
.Y(n_3171)
);

A2O1A1Ixp33_ASAP7_75t_L g3172 ( 
.A1(n_3028),
.A2(n_362),
.B(n_360),
.C(n_361),
.Y(n_3172)
);

AO31x2_ASAP7_75t_L g3173 ( 
.A1(n_2918),
.A2(n_364),
.A3(n_361),
.B(n_363),
.Y(n_3173)
);

AOI21xp5_ASAP7_75t_L g3174 ( 
.A1(n_3038),
.A2(n_363),
.B(n_364),
.Y(n_3174)
);

AO32x2_ASAP7_75t_L g3175 ( 
.A1(n_3004),
.A2(n_2719),
.A3(n_2773),
.B1(n_2883),
.B2(n_2870),
.Y(n_3175)
);

INVx2_ASAP7_75t_L g3176 ( 
.A(n_2712),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_2766),
.B(n_364),
.Y(n_3177)
);

AOI22xp5_ASAP7_75t_L g3178 ( 
.A1(n_2703),
.A2(n_368),
.B1(n_366),
.B2(n_367),
.Y(n_3178)
);

AND2x2_ASAP7_75t_L g3179 ( 
.A(n_2912),
.B(n_366),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_L g3180 ( 
.A(n_2768),
.B(n_367),
.Y(n_3180)
);

AOI21xp5_ASAP7_75t_L g3181 ( 
.A1(n_2986),
.A2(n_368),
.B(n_369),
.Y(n_3181)
);

OAI21xp33_ASAP7_75t_L g3182 ( 
.A1(n_3024),
.A2(n_368),
.B(n_369),
.Y(n_3182)
);

OAI21xp5_ASAP7_75t_L g3183 ( 
.A1(n_2945),
.A2(n_369),
.B(n_370),
.Y(n_3183)
);

AOI21xp33_ASAP7_75t_L g3184 ( 
.A1(n_3050),
.A2(n_370),
.B(n_371),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_L g3185 ( 
.A(n_2778),
.B(n_371),
.Y(n_3185)
);

BUFx2_ASAP7_75t_L g3186 ( 
.A(n_2894),
.Y(n_3186)
);

O2A1O1Ixp33_ASAP7_75t_SL g3187 ( 
.A1(n_2813),
.A2(n_373),
.B(n_371),
.C(n_372),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2823),
.Y(n_3188)
);

NAND2xp33_ASAP7_75t_L g3189 ( 
.A(n_2869),
.B(n_372),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_2846),
.Y(n_3190)
);

NAND2xp5_ASAP7_75t_L g3191 ( 
.A(n_2958),
.B(n_372),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_2722),
.Y(n_3192)
);

AOI21xp5_ASAP7_75t_L g3193 ( 
.A1(n_3058),
.A2(n_373),
.B(n_374),
.Y(n_3193)
);

BUFx3_ASAP7_75t_L g3194 ( 
.A(n_2767),
.Y(n_3194)
);

BUFx2_ASAP7_75t_L g3195 ( 
.A(n_2772),
.Y(n_3195)
);

OAI21xp5_ASAP7_75t_SL g3196 ( 
.A1(n_2700),
.A2(n_373),
.B(n_374),
.Y(n_3196)
);

OAI21x1_ASAP7_75t_L g3197 ( 
.A1(n_3065),
.A2(n_374),
.B(n_375),
.Y(n_3197)
);

A2O1A1Ixp33_ASAP7_75t_L g3198 ( 
.A1(n_2724),
.A2(n_377),
.B(n_375),
.C(n_376),
.Y(n_3198)
);

A2O1A1Ixp33_ASAP7_75t_L g3199 ( 
.A1(n_2862),
.A2(n_378),
.B(n_376),
.C(n_377),
.Y(n_3199)
);

NOR2xp33_ASAP7_75t_L g3200 ( 
.A(n_2851),
.B(n_376),
.Y(n_3200)
);

INVx2_ASAP7_75t_L g3201 ( 
.A(n_2732),
.Y(n_3201)
);

HB1xp67_ASAP7_75t_L g3202 ( 
.A(n_2770),
.Y(n_3202)
);

BUFx10_ASAP7_75t_L g3203 ( 
.A(n_2844),
.Y(n_3203)
);

AO31x2_ASAP7_75t_L g3204 ( 
.A1(n_3017),
.A2(n_3040),
.A3(n_2940),
.B(n_2933),
.Y(n_3204)
);

O2A1O1Ixp33_ASAP7_75t_L g3205 ( 
.A1(n_3025),
.A2(n_379),
.B(n_377),
.C(n_378),
.Y(n_3205)
);

HB1xp67_ASAP7_75t_L g3206 ( 
.A(n_2856),
.Y(n_3206)
);

AND2x4_ASAP7_75t_L g3207 ( 
.A(n_2761),
.B(n_379),
.Y(n_3207)
);

AO31x2_ASAP7_75t_L g3208 ( 
.A1(n_2910),
.A2(n_3046),
.A3(n_2841),
.B(n_2992),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_2739),
.Y(n_3209)
);

OAI21xp5_ASAP7_75t_L g3210 ( 
.A1(n_2964),
.A2(n_379),
.B(n_380),
.Y(n_3210)
);

AOI21xp33_ASAP7_75t_L g3211 ( 
.A1(n_3054),
.A2(n_380),
.B(n_381),
.Y(n_3211)
);

CKINVDCx20_ASAP7_75t_R g3212 ( 
.A(n_2729),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_3007),
.Y(n_3213)
);

A2O1A1Ixp33_ASAP7_75t_L g3214 ( 
.A1(n_3002),
.A2(n_383),
.B(n_381),
.C(n_382),
.Y(n_3214)
);

AND2x4_ASAP7_75t_L g3215 ( 
.A(n_2771),
.B(n_382),
.Y(n_3215)
);

INVx4_ASAP7_75t_L g3216 ( 
.A(n_2812),
.Y(n_3216)
);

NAND3xp33_ASAP7_75t_SL g3217 ( 
.A(n_2875),
.B(n_382),
.C(n_383),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_2985),
.B(n_383),
.Y(n_3218)
);

AOI21xp5_ASAP7_75t_L g3219 ( 
.A1(n_3068),
.A2(n_384),
.B(n_385),
.Y(n_3219)
);

OAI22xp5_ASAP7_75t_L g3220 ( 
.A1(n_2779),
.A2(n_387),
.B1(n_384),
.B2(n_386),
.Y(n_3220)
);

NAND3xp33_ASAP7_75t_L g3221 ( 
.A(n_3001),
.B(n_384),
.C(n_386),
.Y(n_3221)
);

AOI21xp5_ASAP7_75t_L g3222 ( 
.A1(n_3055),
.A2(n_386),
.B(n_387),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_3007),
.Y(n_3223)
);

OAI21x1_ASAP7_75t_L g3224 ( 
.A1(n_2961),
.A2(n_388),
.B(n_389),
.Y(n_3224)
);

AO31x2_ASAP7_75t_L g3225 ( 
.A1(n_2982),
.A2(n_390),
.A3(n_388),
.B(n_389),
.Y(n_3225)
);

AOI21xp5_ASAP7_75t_L g3226 ( 
.A1(n_2990),
.A2(n_390),
.B(n_391),
.Y(n_3226)
);

O2A1O1Ixp33_ASAP7_75t_SL g3227 ( 
.A1(n_2818),
.A2(n_393),
.B(n_391),
.C(n_392),
.Y(n_3227)
);

CKINVDCx20_ASAP7_75t_R g3228 ( 
.A(n_2829),
.Y(n_3228)
);

BUFx4f_ASAP7_75t_SL g3229 ( 
.A(n_2812),
.Y(n_3229)
);

OAI21x1_ASAP7_75t_L g3230 ( 
.A1(n_2748),
.A2(n_392),
.B(n_393),
.Y(n_3230)
);

OAI21x1_ASAP7_75t_L g3231 ( 
.A1(n_2738),
.A2(n_394),
.B(n_395),
.Y(n_3231)
);

OAI21x1_ASAP7_75t_L g3232 ( 
.A1(n_2745),
.A2(n_394),
.B(n_395),
.Y(n_3232)
);

BUFx2_ASAP7_75t_R g3233 ( 
.A(n_2909),
.Y(n_3233)
);

OAI22x1_ASAP7_75t_L g3234 ( 
.A1(n_2771),
.A2(n_396),
.B1(n_394),
.B2(n_395),
.Y(n_3234)
);

BUFx3_ASAP7_75t_L g3235 ( 
.A(n_2785),
.Y(n_3235)
);

BUFx6f_ASAP7_75t_L g3236 ( 
.A(n_2804),
.Y(n_3236)
);

CKINVDCx8_ASAP7_75t_R g3237 ( 
.A(n_2852),
.Y(n_3237)
);

NOR2xp33_ASAP7_75t_L g3238 ( 
.A(n_2934),
.B(n_2942),
.Y(n_3238)
);

AO31x2_ASAP7_75t_L g3239 ( 
.A1(n_3014),
.A2(n_398),
.A3(n_396),
.B(n_397),
.Y(n_3239)
);

AOI22xp5_ASAP7_75t_L g3240 ( 
.A1(n_2807),
.A2(n_399),
.B1(n_396),
.B2(n_398),
.Y(n_3240)
);

AOI21xp5_ASAP7_75t_L g3241 ( 
.A1(n_2708),
.A2(n_399),
.B(n_400),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_SL g3242 ( 
.A(n_2890),
.B(n_400),
.Y(n_3242)
);

AOI21xp5_ASAP7_75t_L g3243 ( 
.A1(n_2709),
.A2(n_400),
.B(n_401),
.Y(n_3243)
);

AOI21xp5_ASAP7_75t_L g3244 ( 
.A1(n_2713),
.A2(n_401),
.B(n_402),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_2796),
.Y(n_3245)
);

AOI21xp5_ASAP7_75t_L g3246 ( 
.A1(n_3022),
.A2(n_401),
.B(n_403),
.Y(n_3246)
);

HB1xp67_ASAP7_75t_L g3247 ( 
.A(n_2995),
.Y(n_3247)
);

O2A1O1Ixp5_ASAP7_75t_L g3248 ( 
.A1(n_2991),
.A2(n_405),
.B(n_403),
.C(n_404),
.Y(n_3248)
);

AOI21xp5_ASAP7_75t_L g3249 ( 
.A1(n_3033),
.A2(n_403),
.B(n_404),
.Y(n_3249)
);

AND2x4_ASAP7_75t_L g3250 ( 
.A(n_3008),
.B(n_404),
.Y(n_3250)
);

AOI21xp5_ASAP7_75t_L g3251 ( 
.A1(n_3056),
.A2(n_405),
.B(n_406),
.Y(n_3251)
);

OA21x2_ASAP7_75t_L g3252 ( 
.A1(n_2938),
.A2(n_405),
.B(n_406),
.Y(n_3252)
);

BUFx2_ASAP7_75t_L g3253 ( 
.A(n_2804),
.Y(n_3253)
);

AO32x2_ASAP7_75t_L g3254 ( 
.A1(n_2884),
.A2(n_409),
.A3(n_407),
.B1(n_408),
.B2(n_410),
.Y(n_3254)
);

OAI21x1_ASAP7_75t_L g3255 ( 
.A1(n_2956),
.A2(n_407),
.B(n_408),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_2840),
.Y(n_3256)
);

AOI21xp5_ASAP7_75t_L g3257 ( 
.A1(n_3066),
.A2(n_407),
.B(n_408),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_2873),
.Y(n_3258)
);

AOI21xp5_ASAP7_75t_L g3259 ( 
.A1(n_3037),
.A2(n_409),
.B(n_410),
.Y(n_3259)
);

NOR2xp67_ASAP7_75t_L g3260 ( 
.A(n_2689),
.B(n_409),
.Y(n_3260)
);

OAI21x1_ASAP7_75t_L g3261 ( 
.A1(n_2956),
.A2(n_411),
.B(n_412),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_2889),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_2914),
.Y(n_3263)
);

A2O1A1Ixp33_ASAP7_75t_L g3264 ( 
.A1(n_2831),
.A2(n_413),
.B(n_411),
.C(n_412),
.Y(n_3264)
);

A2O1A1Ixp33_ASAP7_75t_L g3265 ( 
.A1(n_3044),
.A2(n_411),
.B(n_413),
.C(n_441),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_L g3266 ( 
.A(n_2821),
.B(n_413),
.Y(n_3266)
);

AND2x2_ASAP7_75t_L g3267 ( 
.A(n_2684),
.B(n_441),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_2996),
.Y(n_3268)
);

INVx2_ASAP7_75t_L g3269 ( 
.A(n_2997),
.Y(n_3269)
);

CKINVDCx11_ASAP7_75t_R g3270 ( 
.A(n_3027),
.Y(n_3270)
);

OA21x2_ASAP7_75t_L g3271 ( 
.A1(n_3064),
.A2(n_442),
.B(n_444),
.Y(n_3271)
);

AO31x2_ASAP7_75t_L g3272 ( 
.A1(n_2792),
.A2(n_2801),
.A3(n_2805),
.B(n_2794),
.Y(n_3272)
);

INVx1_ASAP7_75t_SL g3273 ( 
.A(n_2852),
.Y(n_3273)
);

INVx2_ASAP7_75t_L g3274 ( 
.A(n_3016),
.Y(n_3274)
);

AOI21xp5_ASAP7_75t_L g3275 ( 
.A1(n_3005),
.A2(n_442),
.B(n_445),
.Y(n_3275)
);

INVxp67_ASAP7_75t_SL g3276 ( 
.A(n_2905),
.Y(n_3276)
);

AOI21xp5_ASAP7_75t_L g3277 ( 
.A1(n_2731),
.A2(n_445),
.B(n_446),
.Y(n_3277)
);

AO21x2_ASAP7_75t_L g3278 ( 
.A1(n_2998),
.A2(n_447),
.B(n_449),
.Y(n_3278)
);

AOI21xp5_ASAP7_75t_L g3279 ( 
.A1(n_2731),
.A2(n_450),
.B(n_451),
.Y(n_3279)
);

OAI21x1_ASAP7_75t_L g3280 ( 
.A1(n_2963),
.A2(n_450),
.B(n_451),
.Y(n_3280)
);

AOI21xp5_ASAP7_75t_L g3281 ( 
.A1(n_2731),
.A2(n_452),
.B(n_453),
.Y(n_3281)
);

AO21x1_ASAP7_75t_L g3282 ( 
.A1(n_2811),
.A2(n_452),
.B(n_455),
.Y(n_3282)
);

OAI21x1_ASAP7_75t_L g3283 ( 
.A1(n_2966),
.A2(n_455),
.B(n_457),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_3010),
.B(n_813),
.Y(n_3284)
);

AOI21xp5_ASAP7_75t_L g3285 ( 
.A1(n_2744),
.A2(n_457),
.B(n_459),
.Y(n_3285)
);

INVx6_ASAP7_75t_SL g3286 ( 
.A(n_2788),
.Y(n_3286)
);

NOR2xp33_ASAP7_75t_SL g3287 ( 
.A(n_2939),
.B(n_459),
.Y(n_3287)
);

AOI21xp5_ASAP7_75t_L g3288 ( 
.A1(n_2744),
.A2(n_460),
.B(n_461),
.Y(n_3288)
);

BUFx6f_ASAP7_75t_L g3289 ( 
.A(n_2979),
.Y(n_3289)
);

OAI22xp5_ASAP7_75t_L g3290 ( 
.A1(n_2965),
.A2(n_462),
.B1(n_460),
.B2(n_461),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_2725),
.Y(n_3291)
);

OAI21xp5_ASAP7_75t_L g3292 ( 
.A1(n_2927),
.A2(n_462),
.B(n_463),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_SL g3293 ( 
.A(n_3027),
.B(n_463),
.Y(n_3293)
);

NOR2xp33_ASAP7_75t_SL g3294 ( 
.A(n_2822),
.B(n_464),
.Y(n_3294)
);

OAI21x1_ASAP7_75t_L g3295 ( 
.A1(n_2966),
.A2(n_464),
.B(n_465),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_SL g3296 ( 
.A(n_2718),
.B(n_465),
.Y(n_3296)
);

AO31x2_ASAP7_75t_L g3297 ( 
.A1(n_2977),
.A2(n_468),
.A3(n_466),
.B(n_467),
.Y(n_3297)
);

AOI21xp5_ASAP7_75t_L g3298 ( 
.A1(n_2744),
.A2(n_466),
.B(n_468),
.Y(n_3298)
);

NAND2x1_ASAP7_75t_L g3299 ( 
.A(n_3006),
.B(n_2790),
.Y(n_3299)
);

AOI21xp5_ASAP7_75t_L g3300 ( 
.A1(n_2790),
.A2(n_469),
.B(n_470),
.Y(n_3300)
);

INVx2_ASAP7_75t_SL g3301 ( 
.A(n_2935),
.Y(n_3301)
);

CKINVDCx5p33_ASAP7_75t_R g3302 ( 
.A(n_2769),
.Y(n_3302)
);

INVx3_ASAP7_75t_L g3303 ( 
.A(n_2935),
.Y(n_3303)
);

A2O1A1Ixp33_ASAP7_75t_L g3304 ( 
.A1(n_2828),
.A2(n_471),
.B(n_469),
.C(n_470),
.Y(n_3304)
);

AO32x2_ASAP7_75t_L g3305 ( 
.A1(n_2891),
.A2(n_474),
.A3(n_472),
.B1(n_473),
.B2(n_475),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_2763),
.B(n_813),
.Y(n_3306)
);

AOI21xp5_ASAP7_75t_L g3307 ( 
.A1(n_2790),
.A2(n_474),
.B(n_475),
.Y(n_3307)
);

OAI21xp5_ASAP7_75t_L g3308 ( 
.A1(n_2765),
.A2(n_476),
.B(n_477),
.Y(n_3308)
);

A2O1A1Ixp33_ASAP7_75t_L g3309 ( 
.A1(n_2959),
.A2(n_480),
.B(n_478),
.C(n_479),
.Y(n_3309)
);

AOI22xp5_ASAP7_75t_L g3310 ( 
.A1(n_2788),
.A2(n_2865),
.B1(n_2839),
.B2(n_2920),
.Y(n_3310)
);

OAI21x1_ASAP7_75t_L g3311 ( 
.A1(n_2878),
.A2(n_479),
.B(n_480),
.Y(n_3311)
);

INVx3_ASAP7_75t_SL g3312 ( 
.A(n_2798),
.Y(n_3312)
);

OAI21x1_ASAP7_75t_L g3313 ( 
.A1(n_2888),
.A2(n_481),
.B(n_482),
.Y(n_3313)
);

OAI21x1_ASAP7_75t_L g3314 ( 
.A1(n_2774),
.A2(n_481),
.B(n_483),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_2730),
.Y(n_3315)
);

OA21x2_ASAP7_75t_L g3316 ( 
.A1(n_2726),
.A2(n_484),
.B(n_485),
.Y(n_3316)
);

OAI22xp5_ASAP7_75t_L g3317 ( 
.A1(n_2776),
.A2(n_487),
.B1(n_485),
.B2(n_486),
.Y(n_3317)
);

BUFx2_ASAP7_75t_L g3318 ( 
.A(n_2882),
.Y(n_3318)
);

AO32x2_ASAP7_75t_L g3319 ( 
.A1(n_2896),
.A2(n_488),
.A3(n_486),
.B1(n_487),
.B2(n_489),
.Y(n_3319)
);

OAI21x1_ASAP7_75t_L g3320 ( 
.A1(n_2775),
.A2(n_488),
.B(n_489),
.Y(n_3320)
);

BUFx8_ASAP7_75t_SL g3321 ( 
.A(n_2892),
.Y(n_3321)
);

O2A1O1Ixp33_ASAP7_75t_SL g3322 ( 
.A1(n_2710),
.A2(n_492),
.B(n_490),
.C(n_491),
.Y(n_3322)
);

AO31x2_ASAP7_75t_L g3323 ( 
.A1(n_2874),
.A2(n_493),
.A3(n_490),
.B(n_491),
.Y(n_3323)
);

NAND3xp33_ASAP7_75t_L g3324 ( 
.A(n_3009),
.B(n_493),
.C(n_494),
.Y(n_3324)
);

BUFx3_ASAP7_75t_L g3325 ( 
.A(n_2935),
.Y(n_3325)
);

AO31x2_ASAP7_75t_L g3326 ( 
.A1(n_2983),
.A2(n_497),
.A3(n_495),
.B(n_496),
.Y(n_3326)
);

OR2x2_ASAP7_75t_L g3327 ( 
.A(n_2755),
.B(n_496),
.Y(n_3327)
);

OAI221xp5_ASAP7_75t_L g3328 ( 
.A1(n_2919),
.A2(n_499),
.B1(n_497),
.B2(n_498),
.C(n_500),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_2736),
.Y(n_3329)
);

AOI221x1_ASAP7_75t_L g3330 ( 
.A1(n_2685),
.A2(n_501),
.B1(n_498),
.B2(n_499),
.C(n_502),
.Y(n_3330)
);

AOI31xp67_ASAP7_75t_L g3331 ( 
.A1(n_3036),
.A2(n_503),
.A3(n_501),
.B(n_502),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_2782),
.B(n_504),
.Y(n_3332)
);

AND2x2_ASAP7_75t_L g3333 ( 
.A(n_2946),
.B(n_505),
.Y(n_3333)
);

AOI22xp5_ASAP7_75t_L g3334 ( 
.A1(n_2922),
.A2(n_507),
.B1(n_505),
.B2(n_506),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_2751),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_2784),
.B(n_2806),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_L g3337 ( 
.A(n_2816),
.B(n_812),
.Y(n_3337)
);

BUFx10_ASAP7_75t_L g3338 ( 
.A(n_2797),
.Y(n_3338)
);

OR2x6_ASAP7_75t_L g3339 ( 
.A(n_2797),
.B(n_506),
.Y(n_3339)
);

OR2x2_ASAP7_75t_L g3340 ( 
.A(n_3008),
.B(n_508),
.Y(n_3340)
);

AOI21xp5_ASAP7_75t_L g3341 ( 
.A1(n_2810),
.A2(n_508),
.B(n_509),
.Y(n_3341)
);

O2A1O1Ixp33_ASAP7_75t_L g3342 ( 
.A1(n_2893),
.A2(n_511),
.B(n_509),
.C(n_510),
.Y(n_3342)
);

OAI22xp5_ASAP7_75t_L g3343 ( 
.A1(n_2924),
.A2(n_514),
.B1(n_512),
.B2(n_513),
.Y(n_3343)
);

AO21x1_ASAP7_75t_L g3344 ( 
.A1(n_3052),
.A2(n_513),
.B(n_514),
.Y(n_3344)
);

INVx2_ASAP7_75t_L g3345 ( 
.A(n_3023),
.Y(n_3345)
);

AOI22xp33_ASAP7_75t_L g3346 ( 
.A1(n_2695),
.A2(n_517),
.B1(n_515),
.B2(n_516),
.Y(n_3346)
);

OAI21xp5_ASAP7_75t_L g3347 ( 
.A1(n_2859),
.A2(n_2867),
.B(n_2952),
.Y(n_3347)
);

AOI21xp5_ASAP7_75t_L g3348 ( 
.A1(n_2810),
.A2(n_516),
.B(n_517),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_2858),
.B(n_811),
.Y(n_3349)
);

AOI221x1_ASAP7_75t_L g3350 ( 
.A1(n_2879),
.A2(n_520),
.B1(n_518),
.B2(n_519),
.C(n_522),
.Y(n_3350)
);

INVx2_ASAP7_75t_L g3351 ( 
.A(n_3026),
.Y(n_3351)
);

OAI21xp5_ASAP7_75t_L g3352 ( 
.A1(n_2987),
.A2(n_518),
.B(n_520),
.Y(n_3352)
);

NAND3xp33_ASAP7_75t_L g3353 ( 
.A(n_2845),
.B(n_522),
.C(n_524),
.Y(n_3353)
);

INVx2_ASAP7_75t_L g3354 ( 
.A(n_2979),
.Y(n_3354)
);

OA21x2_ASAP7_75t_L g3355 ( 
.A1(n_2921),
.A2(n_525),
.B(n_527),
.Y(n_3355)
);

O2A1O1Ixp33_ASAP7_75t_L g3356 ( 
.A1(n_2898),
.A2(n_528),
.B(n_525),
.C(n_527),
.Y(n_3356)
);

CKINVDCx16_ASAP7_75t_R g3357 ( 
.A(n_2954),
.Y(n_3357)
);

AO32x2_ASAP7_75t_L g3358 ( 
.A1(n_2902),
.A2(n_530),
.A3(n_528),
.B1(n_529),
.B2(n_531),
.Y(n_3358)
);

AOI21xp5_ASAP7_75t_L g3359 ( 
.A1(n_2810),
.A2(n_529),
.B(n_531),
.Y(n_3359)
);

AOI21xp5_ASAP7_75t_L g3360 ( 
.A1(n_2861),
.A2(n_532),
.B(n_533),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_2757),
.Y(n_3361)
);

OAI22x1_ASAP7_75t_L g3362 ( 
.A1(n_2954),
.A2(n_535),
.B1(n_532),
.B2(n_534),
.Y(n_3362)
);

AOI22xp33_ASAP7_75t_L g3363 ( 
.A1(n_2949),
.A2(n_536),
.B1(n_534),
.B2(n_535),
.Y(n_3363)
);

AO22x2_ASAP7_75t_L g3364 ( 
.A1(n_2955),
.A2(n_540),
.B1(n_536),
.B2(n_539),
.Y(n_3364)
);

OA21x2_ASAP7_75t_L g3365 ( 
.A1(n_2817),
.A2(n_2872),
.B(n_2989),
.Y(n_3365)
);

NOR2x1_ASAP7_75t_L g3366 ( 
.A(n_2683),
.B(n_2777),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_2706),
.Y(n_3367)
);

OA21x2_ASAP7_75t_L g3368 ( 
.A1(n_2853),
.A2(n_539),
.B(n_540),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_2943),
.B(n_811),
.Y(n_3369)
);

AOI21xp5_ASAP7_75t_L g3370 ( 
.A1(n_2861),
.A2(n_541),
.B(n_542),
.Y(n_3370)
);

NOR2xp33_ASAP7_75t_L g3371 ( 
.A(n_2900),
.B(n_544),
.Y(n_3371)
);

BUFx8_ASAP7_75t_L g3372 ( 
.A(n_3041),
.Y(n_3372)
);

OR2x2_ASAP7_75t_L g3373 ( 
.A(n_3318),
.B(n_2836),
.Y(n_3373)
);

CKINVDCx20_ASAP7_75t_R g3374 ( 
.A(n_3212),
.Y(n_3374)
);

HB1xp67_ASAP7_75t_L g3375 ( 
.A(n_3202),
.Y(n_3375)
);

AOI22xp33_ASAP7_75t_SL g3376 ( 
.A1(n_3357),
.A2(n_3032),
.B1(n_2835),
.B2(n_2830),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_L g3377 ( 
.A(n_3367),
.B(n_2728),
.Y(n_3377)
);

CKINVDCx11_ASAP7_75t_R g3378 ( 
.A(n_3237),
.Y(n_3378)
);

BUFx2_ASAP7_75t_L g3379 ( 
.A(n_3286),
.Y(n_3379)
);

INVx2_ASAP7_75t_L g3380 ( 
.A(n_3269),
.Y(n_3380)
);

AOI21xp5_ASAP7_75t_SL g3381 ( 
.A1(n_3339),
.A2(n_2714),
.B(n_2727),
.Y(n_3381)
);

INVx8_ASAP7_75t_L g3382 ( 
.A(n_3087),
.Y(n_3382)
);

HB1xp67_ASAP7_75t_L g3383 ( 
.A(n_3071),
.Y(n_3383)
);

INVx6_ASAP7_75t_L g3384 ( 
.A(n_3152),
.Y(n_3384)
);

BUFx12f_ASAP7_75t_L g3385 ( 
.A(n_3141),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_3070),
.Y(n_3386)
);

BUFx6f_ASAP7_75t_SL g3387 ( 
.A(n_3140),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_3078),
.Y(n_3388)
);

OAI22xp5_ASAP7_75t_L g3389 ( 
.A1(n_3339),
.A2(n_2711),
.B1(n_2693),
.B2(n_3030),
.Y(n_3389)
);

OAI22xp33_ASAP7_75t_L g3390 ( 
.A1(n_3196),
.A2(n_2984),
.B1(n_2871),
.B2(n_3029),
.Y(n_3390)
);

AOI22xp33_ASAP7_75t_L g3391 ( 
.A1(n_3130),
.A2(n_2950),
.B1(n_2864),
.B2(n_2860),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3107),
.Y(n_3392)
);

CKINVDCx11_ASAP7_75t_R g3393 ( 
.A(n_3273),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3143),
.Y(n_3394)
);

OAI22xp33_ASAP7_75t_L g3395 ( 
.A1(n_3287),
.A2(n_2827),
.B1(n_2721),
.B2(n_2716),
.Y(n_3395)
);

OR2x2_ASAP7_75t_L g3396 ( 
.A(n_3247),
.B(n_3062),
.Y(n_3396)
);

BUFx10_ASAP7_75t_L g3397 ( 
.A(n_3087),
.Y(n_3397)
);

AOI22xp33_ASAP7_75t_L g3398 ( 
.A1(n_3082),
.A2(n_2930),
.B1(n_2941),
.B2(n_2926),
.Y(n_3398)
);

INVx1_ASAP7_75t_SL g3399 ( 
.A(n_3286),
.Y(n_3399)
);

INVx1_ASAP7_75t_L g3400 ( 
.A(n_3144),
.Y(n_3400)
);

CKINVDCx11_ASAP7_75t_R g3401 ( 
.A(n_3228),
.Y(n_3401)
);

CKINVDCx11_ASAP7_75t_R g3402 ( 
.A(n_3096),
.Y(n_3402)
);

INVx6_ASAP7_75t_L g3403 ( 
.A(n_3216),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_3169),
.Y(n_3404)
);

CKINVDCx20_ASAP7_75t_R g3405 ( 
.A(n_3229),
.Y(n_3405)
);

AOI22xp33_ASAP7_75t_L g3406 ( 
.A1(n_3217),
.A2(n_3011),
.B1(n_3013),
.B2(n_2988),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_3188),
.Y(n_3407)
);

AOI22xp5_ASAP7_75t_L g3408 ( 
.A1(n_3189),
.A2(n_2901),
.B1(n_2803),
.B2(n_3018),
.Y(n_3408)
);

INVx1_ASAP7_75t_L g3409 ( 
.A(n_3190),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3192),
.Y(n_3410)
);

CKINVDCx20_ASAP7_75t_R g3411 ( 
.A(n_3270),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_3274),
.Y(n_3412)
);

BUFx12f_ASAP7_75t_L g3413 ( 
.A(n_3203),
.Y(n_3413)
);

INVx6_ASAP7_75t_L g3414 ( 
.A(n_3325),
.Y(n_3414)
);

BUFx6f_ASAP7_75t_SL g3415 ( 
.A(n_3194),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_3209),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_L g3417 ( 
.A(n_3132),
.B(n_3045),
.Y(n_3417)
);

OAI21xp33_ASAP7_75t_L g3418 ( 
.A1(n_3233),
.A2(n_2740),
.B(n_2847),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_3086),
.Y(n_3419)
);

INVx6_ASAP7_75t_L g3420 ( 
.A(n_3338),
.Y(n_3420)
);

AOI22xp33_ASAP7_75t_L g3421 ( 
.A1(n_3146),
.A2(n_3034),
.B1(n_3035),
.B2(n_3019),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_3165),
.Y(n_3422)
);

BUFx6f_ASAP7_75t_L g3423 ( 
.A(n_3289),
.Y(n_3423)
);

CKINVDCx11_ASAP7_75t_R g3424 ( 
.A(n_3155),
.Y(n_3424)
);

AOI22xp33_ASAP7_75t_L g3425 ( 
.A1(n_3081),
.A2(n_2832),
.B1(n_2953),
.B2(n_2970),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_L g3426 ( 
.A(n_3128),
.B(n_3291),
.Y(n_3426)
);

INVx2_ASAP7_75t_L g3427 ( 
.A(n_3345),
.Y(n_3427)
);

INVx6_ASAP7_75t_L g3428 ( 
.A(n_3372),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_3176),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_L g3430 ( 
.A(n_3315),
.B(n_2923),
.Y(n_3430)
);

CKINVDCx20_ASAP7_75t_R g3431 ( 
.A(n_3321),
.Y(n_3431)
);

NAND2x1p5_ASAP7_75t_L g3432 ( 
.A(n_3113),
.B(n_2979),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_3201),
.Y(n_3433)
);

INVx6_ASAP7_75t_L g3434 ( 
.A(n_3118),
.Y(n_3434)
);

AOI22xp33_ASAP7_75t_L g3435 ( 
.A1(n_3081),
.A2(n_2993),
.B1(n_2978),
.B2(n_3039),
.Y(n_3435)
);

AOI22xp5_ASAP7_75t_L g3436 ( 
.A1(n_3097),
.A2(n_3003),
.B1(n_2999),
.B2(n_3063),
.Y(n_3436)
);

INVx6_ASAP7_75t_L g3437 ( 
.A(n_3118),
.Y(n_3437)
);

INVx1_ASAP7_75t_L g3438 ( 
.A(n_3080),
.Y(n_3438)
);

AOI22xp33_ASAP7_75t_L g3439 ( 
.A1(n_3296),
.A2(n_2908),
.B1(n_2759),
.B2(n_3048),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3245),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_3256),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_3258),
.Y(n_3442)
);

AND2x2_ASAP7_75t_L g3443 ( 
.A(n_3179),
.B(n_544),
.Y(n_3443)
);

INVx2_ASAP7_75t_L g3444 ( 
.A(n_3351),
.Y(n_3444)
);

BUFx4f_ASAP7_75t_SL g3445 ( 
.A(n_3161),
.Y(n_3445)
);

CKINVDCx14_ASAP7_75t_R g3446 ( 
.A(n_3238),
.Y(n_3446)
);

CKINVDCx11_ASAP7_75t_R g3447 ( 
.A(n_3312),
.Y(n_3447)
);

AOI22xp33_ASAP7_75t_L g3448 ( 
.A1(n_3094),
.A2(n_3051),
.B1(n_2944),
.B2(n_2994),
.Y(n_3448)
);

CKINVDCx11_ASAP7_75t_R g3449 ( 
.A(n_3186),
.Y(n_3449)
);

BUFx3_ASAP7_75t_L g3450 ( 
.A(n_3235),
.Y(n_3450)
);

AOI22xp33_ASAP7_75t_SL g3451 ( 
.A1(n_3220),
.A2(n_3207),
.B1(n_3215),
.B2(n_3085),
.Y(n_3451)
);

OAI22xp5_ASAP7_75t_L g3452 ( 
.A1(n_3310),
.A2(n_2925),
.B1(n_2887),
.B2(n_2854),
.Y(n_3452)
);

INVx2_ASAP7_75t_L g3453 ( 
.A(n_3077),
.Y(n_3453)
);

INVx2_ASAP7_75t_L g3454 ( 
.A(n_3262),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_3263),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3268),
.Y(n_3456)
);

OAI22xp5_ASAP7_75t_L g3457 ( 
.A1(n_3207),
.A2(n_2976),
.B1(n_2932),
.B2(n_2824),
.Y(n_3457)
);

INVx3_ASAP7_75t_L g3458 ( 
.A(n_3289),
.Y(n_3458)
);

AOI22xp5_ASAP7_75t_L g3459 ( 
.A1(n_3162),
.A2(n_2697),
.B1(n_2705),
.B2(n_2694),
.Y(n_3459)
);

AOI22xp33_ASAP7_75t_L g3460 ( 
.A1(n_3215),
.A2(n_3250),
.B1(n_3137),
.B2(n_3182),
.Y(n_3460)
);

OAI22xp33_ASAP7_75t_R g3461 ( 
.A1(n_3075),
.A2(n_548),
.B1(n_545),
.B2(n_546),
.Y(n_3461)
);

OAI22xp5_ASAP7_75t_L g3462 ( 
.A1(n_3265),
.A2(n_2750),
.B1(n_3006),
.B2(n_3061),
.Y(n_3462)
);

INVx6_ASAP7_75t_L g3463 ( 
.A(n_3236),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3158),
.Y(n_3464)
);

AOI22xp33_ASAP7_75t_SL g3465 ( 
.A1(n_3294),
.A2(n_3057),
.B1(n_3042),
.B2(n_2814),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_3340),
.Y(n_3466)
);

INVxp67_ASAP7_75t_L g3467 ( 
.A(n_3195),
.Y(n_3467)
);

AOI22xp33_ASAP7_75t_L g3468 ( 
.A1(n_3250),
.A2(n_2814),
.B1(n_2843),
.B2(n_2753),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3177),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3180),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3185),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3266),
.Y(n_3472)
);

AOI22xp33_ASAP7_75t_L g3473 ( 
.A1(n_3364),
.A2(n_2843),
.B1(n_2868),
.B2(n_2753),
.Y(n_3473)
);

AOI22xp33_ASAP7_75t_SL g3474 ( 
.A1(n_3364),
.A2(n_3057),
.B1(n_3042),
.B2(n_2868),
.Y(n_3474)
);

AOI22xp33_ASAP7_75t_SL g3475 ( 
.A1(n_3153),
.A2(n_3057),
.B1(n_3042),
.B2(n_2877),
.Y(n_3475)
);

AOI22xp33_ASAP7_75t_L g3476 ( 
.A1(n_3328),
.A2(n_2877),
.B1(n_2917),
.B2(n_2899),
.Y(n_3476)
);

BUFx6f_ASAP7_75t_L g3477 ( 
.A(n_3301),
.Y(n_3477)
);

BUFx12f_ASAP7_75t_L g3478 ( 
.A(n_3236),
.Y(n_3478)
);

NAND2xp5_ASAP7_75t_L g3479 ( 
.A(n_3329),
.B(n_3335),
.Y(n_3479)
);

AOI22xp5_ASAP7_75t_L g3480 ( 
.A1(n_3240),
.A2(n_2917),
.B1(n_2928),
.B2(n_2899),
.Y(n_3480)
);

AOI22xp33_ASAP7_75t_L g3481 ( 
.A1(n_3142),
.A2(n_2928),
.B1(n_2881),
.B2(n_2904),
.Y(n_3481)
);

AOI22xp33_ASAP7_75t_SL g3482 ( 
.A1(n_3183),
.A2(n_3210),
.B1(n_3302),
.B2(n_3276),
.Y(n_3482)
);

AOI22xp33_ASAP7_75t_L g3483 ( 
.A1(n_3088),
.A2(n_2881),
.B1(n_2904),
.B2(n_2861),
.Y(n_3483)
);

INVx2_ASAP7_75t_L g3484 ( 
.A(n_3255),
.Y(n_3484)
);

AOI22xp33_ASAP7_75t_L g3485 ( 
.A1(n_3221),
.A2(n_3123),
.B1(n_3347),
.B2(n_3136),
.Y(n_3485)
);

CKINVDCx5p33_ASAP7_75t_R g3486 ( 
.A(n_3138),
.Y(n_3486)
);

BUFx4_ASAP7_75t_SL g3487 ( 
.A(n_3136),
.Y(n_3487)
);

AOI22xp33_ASAP7_75t_L g3488 ( 
.A1(n_3105),
.A2(n_3366),
.B1(n_3290),
.B2(n_3336),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3163),
.Y(n_3489)
);

BUFx12f_ASAP7_75t_L g3490 ( 
.A(n_3253),
.Y(n_3490)
);

AOI22xp33_ASAP7_75t_L g3491 ( 
.A1(n_3284),
.A2(n_2904),
.B1(n_2929),
.B2(n_2881),
.Y(n_3491)
);

INVx2_ASAP7_75t_L g3492 ( 
.A(n_3261),
.Y(n_3492)
);

OAI21xp33_ASAP7_75t_L g3493 ( 
.A1(n_3234),
.A2(n_2948),
.B(n_2929),
.Y(n_3493)
);

AOI22xp33_ASAP7_75t_SL g3494 ( 
.A1(n_3308),
.A2(n_2948),
.B1(n_2960),
.B2(n_2929),
.Y(n_3494)
);

INVx2_ASAP7_75t_L g3495 ( 
.A(n_3280),
.Y(n_3495)
);

AOI22xp5_ASAP7_75t_L g3496 ( 
.A1(n_3260),
.A2(n_2960),
.B1(n_2975),
.B2(n_2948),
.Y(n_3496)
);

AOI22xp33_ASAP7_75t_L g3497 ( 
.A1(n_3353),
.A2(n_3191),
.B1(n_3218),
.B2(n_3361),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_3163),
.Y(n_3498)
);

INVx2_ASAP7_75t_L g3499 ( 
.A(n_3283),
.Y(n_3499)
);

INVx2_ASAP7_75t_L g3500 ( 
.A(n_3295),
.Y(n_3500)
);

AOI22xp33_ASAP7_75t_L g3501 ( 
.A1(n_3134),
.A2(n_2975),
.B1(n_3000),
.B2(n_2960),
.Y(n_3501)
);

AOI22xp33_ASAP7_75t_SL g3502 ( 
.A1(n_3333),
.A2(n_3000),
.B1(n_2975),
.B2(n_549),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_3103),
.B(n_3000),
.Y(n_3503)
);

BUFx12f_ASAP7_75t_L g3504 ( 
.A(n_3124),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_3163),
.Y(n_3505)
);

AOI22xp33_ASAP7_75t_L g3506 ( 
.A1(n_3184),
.A2(n_550),
.B1(n_546),
.B2(n_548),
.Y(n_3506)
);

OAI22xp33_ASAP7_75t_L g3507 ( 
.A1(n_3178),
.A2(n_3362),
.B1(n_3106),
.B2(n_3334),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_L g3508 ( 
.A(n_3135),
.B(n_3206),
.Y(n_3508)
);

CKINVDCx11_ASAP7_75t_R g3509 ( 
.A(n_3354),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_3326),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_3326),
.Y(n_3511)
);

BUFx2_ASAP7_75t_L g3512 ( 
.A(n_3120),
.Y(n_3512)
);

CKINVDCx11_ASAP7_75t_R g3513 ( 
.A(n_3120),
.Y(n_3513)
);

OAI22xp5_ASAP7_75t_L g3514 ( 
.A1(n_3264),
.A2(n_553),
.B1(n_551),
.B2(n_552),
.Y(n_3514)
);

BUFx2_ASAP7_75t_L g3515 ( 
.A(n_3303),
.Y(n_3515)
);

INVx1_ASAP7_75t_SL g3516 ( 
.A(n_3147),
.Y(n_3516)
);

INVx1_ASAP7_75t_L g3517 ( 
.A(n_3213),
.Y(n_3517)
);

AND2x2_ASAP7_75t_L g3518 ( 
.A(n_3267),
.B(n_810),
.Y(n_3518)
);

OR2x2_ASAP7_75t_L g3519 ( 
.A(n_3327),
.B(n_552),
.Y(n_3519)
);

AOI22xp5_ASAP7_75t_L g3520 ( 
.A1(n_3317),
.A2(n_555),
.B1(n_553),
.B2(n_554),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_3223),
.Y(n_3521)
);

CKINVDCx20_ASAP7_75t_R g3522 ( 
.A(n_3117),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3297),
.Y(n_3523)
);

AOI22xp33_ASAP7_75t_SL g3524 ( 
.A1(n_3352),
.A2(n_556),
.B1(n_554),
.B2(n_555),
.Y(n_3524)
);

CKINVDCx5p33_ASAP7_75t_R g3525 ( 
.A(n_3371),
.Y(n_3525)
);

AOI22xp33_ASAP7_75t_L g3526 ( 
.A1(n_3211),
.A2(n_558),
.B1(n_556),
.B2(n_557),
.Y(n_3526)
);

OAI22xp5_ASAP7_75t_L g3527 ( 
.A1(n_3198),
.A2(n_559),
.B1(n_557),
.B2(n_558),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_3122),
.B(n_559),
.Y(n_3528)
);

AOI22xp33_ASAP7_75t_L g3529 ( 
.A1(n_3109),
.A2(n_564),
.B1(n_560),
.B2(n_561),
.Y(n_3529)
);

CKINVDCx20_ASAP7_75t_R g3530 ( 
.A(n_3171),
.Y(n_3530)
);

AOI22xp33_ASAP7_75t_L g3531 ( 
.A1(n_3133),
.A2(n_567),
.B1(n_560),
.B2(n_565),
.Y(n_3531)
);

INVx6_ASAP7_75t_L g3532 ( 
.A(n_3299),
.Y(n_3532)
);

INVx11_ASAP7_75t_L g3533 ( 
.A(n_3151),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3297),
.Y(n_3534)
);

AOI22xp33_ASAP7_75t_L g3535 ( 
.A1(n_3200),
.A2(n_569),
.B1(n_565),
.B2(n_567),
.Y(n_3535)
);

OAI22xp33_ASAP7_75t_L g3536 ( 
.A1(n_3330),
.A2(n_571),
.B1(n_569),
.B2(n_570),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3297),
.Y(n_3537)
);

AOI22xp33_ASAP7_75t_L g3538 ( 
.A1(n_3131),
.A2(n_573),
.B1(n_570),
.B2(n_572),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_3323),
.Y(n_3539)
);

HB1xp67_ASAP7_75t_L g3540 ( 
.A(n_3159),
.Y(n_3540)
);

AOI22xp33_ASAP7_75t_L g3541 ( 
.A1(n_3343),
.A2(n_574),
.B1(n_572),
.B2(n_573),
.Y(n_3541)
);

OAI22xp5_ASAP7_75t_L g3542 ( 
.A1(n_3346),
.A2(n_577),
.B1(n_575),
.B2(n_576),
.Y(n_3542)
);

BUFx12f_ASAP7_75t_L g3543 ( 
.A(n_3350),
.Y(n_3543)
);

BUFx2_ASAP7_75t_SL g3544 ( 
.A(n_3293),
.Y(n_3544)
);

AOI22xp5_ASAP7_75t_L g3545 ( 
.A1(n_3369),
.A2(n_579),
.B1(n_575),
.B2(n_577),
.Y(n_3545)
);

NAND2x1p5_ASAP7_75t_L g3546 ( 
.A(n_3242),
.B(n_580),
.Y(n_3546)
);

INVx6_ASAP7_75t_L g3547 ( 
.A(n_3214),
.Y(n_3547)
);

NAND2xp5_ASAP7_75t_L g3548 ( 
.A(n_3114),
.B(n_580),
.Y(n_3548)
);

AOI22xp33_ASAP7_75t_SL g3549 ( 
.A1(n_3252),
.A2(n_583),
.B1(n_581),
.B2(n_582),
.Y(n_3549)
);

INVx8_ASAP7_75t_L g3550 ( 
.A(n_3167),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_L g3551 ( 
.A(n_3139),
.B(n_581),
.Y(n_3551)
);

AND2x2_ASAP7_75t_L g3552 ( 
.A(n_3175),
.B(n_582),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_3323),
.Y(n_3553)
);

AOI22xp33_ASAP7_75t_SL g3554 ( 
.A1(n_3252),
.A2(n_585),
.B1(n_583),
.B2(n_584),
.Y(n_3554)
);

OAI22xp5_ASAP7_75t_L g3555 ( 
.A1(n_3166),
.A2(n_586),
.B1(n_584),
.B2(n_585),
.Y(n_3555)
);

BUFx2_ASAP7_75t_L g3556 ( 
.A(n_3305),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3145),
.Y(n_3557)
);

AOI22xp33_ASAP7_75t_L g3558 ( 
.A1(n_3112),
.A2(n_588),
.B1(n_586),
.B2(n_587),
.Y(n_3558)
);

AOI22xp33_ASAP7_75t_SL g3559 ( 
.A1(n_3316),
.A2(n_591),
.B1(n_589),
.B2(n_590),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_L g3560 ( 
.A(n_3349),
.B(n_590),
.Y(n_3560)
);

BUFx6f_ASAP7_75t_L g3561 ( 
.A(n_3084),
.Y(n_3561)
);

INVx1_ASAP7_75t_L g3562 ( 
.A(n_3173),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3173),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3254),
.Y(n_3564)
);

AOI22xp33_ASAP7_75t_L g3565 ( 
.A1(n_3363),
.A2(n_593),
.B1(n_591),
.B2(n_592),
.Y(n_3565)
);

AOI22xp33_ASAP7_75t_L g3566 ( 
.A1(n_3251),
.A2(n_596),
.B1(n_594),
.B2(n_595),
.Y(n_3566)
);

AOI22xp33_ASAP7_75t_SL g3567 ( 
.A1(n_3316),
.A2(n_598),
.B1(n_594),
.B2(n_597),
.Y(n_3567)
);

AOI22xp33_ASAP7_75t_SL g3568 ( 
.A1(n_3368),
.A2(n_599),
.B1(n_597),
.B2(n_598),
.Y(n_3568)
);

CKINVDCx6p67_ASAP7_75t_R g3569 ( 
.A(n_3306),
.Y(n_3569)
);

AND2x2_ASAP7_75t_L g3570 ( 
.A(n_3175),
.B(n_600),
.Y(n_3570)
);

BUFx3_ASAP7_75t_L g3571 ( 
.A(n_3314),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3254),
.Y(n_3572)
);

INVx1_ASAP7_75t_SL g3573 ( 
.A(n_3110),
.Y(n_3573)
);

BUFx8_ASAP7_75t_L g3574 ( 
.A(n_3254),
.Y(n_3574)
);

AOI22xp33_ASAP7_75t_L g3575 ( 
.A1(n_3257),
.A2(n_603),
.B1(n_601),
.B2(n_602),
.Y(n_3575)
);

AND2x2_ASAP7_75t_L g3576 ( 
.A(n_3175),
.B(n_604),
.Y(n_3576)
);

AOI22xp33_ASAP7_75t_SL g3577 ( 
.A1(n_3368),
.A2(n_606),
.B1(n_604),
.B2(n_605),
.Y(n_3577)
);

CKINVDCx5p33_ASAP7_75t_R g3578 ( 
.A(n_3332),
.Y(n_3578)
);

OAI22xp5_ASAP7_75t_L g3579 ( 
.A1(n_3172),
.A2(n_608),
.B1(n_605),
.B2(n_606),
.Y(n_3579)
);

AOI22xp33_ASAP7_75t_L g3580 ( 
.A1(n_3282),
.A2(n_611),
.B1(n_609),
.B2(n_610),
.Y(n_3580)
);

BUFx3_ASAP7_75t_L g3581 ( 
.A(n_3320),
.Y(n_3581)
);

CKINVDCx8_ASAP7_75t_R g3582 ( 
.A(n_3355),
.Y(n_3582)
);

CKINVDCx5p33_ASAP7_75t_R g3583 ( 
.A(n_3337),
.Y(n_3583)
);

AOI22xp33_ASAP7_75t_SL g3584 ( 
.A1(n_3355),
.A2(n_612),
.B1(n_609),
.B2(n_610),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3225),
.Y(n_3585)
);

BUFx2_ASAP7_75t_L g3586 ( 
.A(n_3305),
.Y(n_3586)
);

AOI22xp5_ASAP7_75t_L g3587 ( 
.A1(n_3150),
.A2(n_615),
.B1(n_612),
.B2(n_614),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3225),
.Y(n_3588)
);

OR2x2_ASAP7_75t_L g3589 ( 
.A(n_3225),
.B(n_614),
.Y(n_3589)
);

CKINVDCx11_ASAP7_75t_R g3590 ( 
.A(n_3305),
.Y(n_3590)
);

BUFx3_ASAP7_75t_L g3591 ( 
.A(n_3230),
.Y(n_3591)
);

INVx4_ASAP7_75t_L g3592 ( 
.A(n_3278),
.Y(n_3592)
);

AOI22xp33_ASAP7_75t_L g3593 ( 
.A1(n_3259),
.A2(n_618),
.B1(n_615),
.B2(n_617),
.Y(n_3593)
);

AOI22xp33_ASAP7_75t_L g3594 ( 
.A1(n_3108),
.A2(n_621),
.B1(n_619),
.B2(n_620),
.Y(n_3594)
);

BUFx10_ASAP7_75t_L g3595 ( 
.A(n_3319),
.Y(n_3595)
);

AOI22xp33_ASAP7_75t_L g3596 ( 
.A1(n_3241),
.A2(n_622),
.B1(n_620),
.B2(n_621),
.Y(n_3596)
);

AOI22xp33_ASAP7_75t_SL g3597 ( 
.A1(n_3292),
.A2(n_624),
.B1(n_622),
.B2(n_623),
.Y(n_3597)
);

OAI22xp5_ASAP7_75t_L g3598 ( 
.A1(n_3199),
.A2(n_626),
.B1(n_623),
.B2(n_625),
.Y(n_3598)
);

AND2x2_ASAP7_75t_L g3599 ( 
.A(n_3319),
.B(n_810),
.Y(n_3599)
);

AOI22xp33_ASAP7_75t_L g3600 ( 
.A1(n_3243),
.A2(n_628),
.B1(n_625),
.B2(n_627),
.Y(n_3600)
);

CKINVDCx20_ASAP7_75t_R g3601 ( 
.A(n_3344),
.Y(n_3601)
);

AOI21xp5_ASAP7_75t_L g3602 ( 
.A1(n_3092),
.A2(n_3126),
.B(n_3090),
.Y(n_3602)
);

INVxp67_ASAP7_75t_SL g3603 ( 
.A(n_3100),
.Y(n_3603)
);

BUFx3_ASAP7_75t_L g3604 ( 
.A(n_3231),
.Y(n_3604)
);

AND2x2_ASAP7_75t_L g3605 ( 
.A(n_3319),
.B(n_809),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_L g3606 ( 
.A(n_3244),
.B(n_627),
.Y(n_3606)
);

INVx2_ASAP7_75t_SL g3607 ( 
.A(n_3232),
.Y(n_3607)
);

AOI22xp33_ASAP7_75t_L g3608 ( 
.A1(n_3324),
.A2(n_631),
.B1(n_628),
.B2(n_630),
.Y(n_3608)
);

INVx1_ASAP7_75t_SL g3609 ( 
.A(n_3365),
.Y(n_3609)
);

OAI22xp5_ASAP7_75t_SL g3610 ( 
.A1(n_3271),
.A2(n_634),
.B1(n_631),
.B2(n_633),
.Y(n_3610)
);

AOI22xp33_ASAP7_75t_L g3611 ( 
.A1(n_3099),
.A2(n_637),
.B1(n_635),
.B2(n_636),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_L g3612 ( 
.A(n_3239),
.B(n_3072),
.Y(n_3612)
);

CKINVDCx20_ASAP7_75t_R g3613 ( 
.A(n_3275),
.Y(n_3613)
);

CKINVDCx8_ASAP7_75t_R g3614 ( 
.A(n_3271),
.Y(n_3614)
);

AOI22xp33_ASAP7_75t_L g3615 ( 
.A1(n_3116),
.A2(n_638),
.B1(n_635),
.B2(n_637),
.Y(n_3615)
);

BUFx12f_ASAP7_75t_L g3616 ( 
.A(n_3358),
.Y(n_3616)
);

INVx4_ASAP7_75t_L g3617 ( 
.A(n_3365),
.Y(n_3617)
);

INVx2_ASAP7_75t_SL g3618 ( 
.A(n_3224),
.Y(n_3618)
);

INVxp67_ASAP7_75t_SL g3619 ( 
.A(n_3076),
.Y(n_3619)
);

OAI21xp33_ASAP7_75t_L g3620 ( 
.A1(n_3091),
.A2(n_638),
.B(n_639),
.Y(n_3620)
);

AOI22xp5_ASAP7_75t_L g3621 ( 
.A1(n_3222),
.A2(n_642),
.B1(n_640),
.B2(n_641),
.Y(n_3621)
);

CKINVDCx11_ASAP7_75t_R g3622 ( 
.A(n_3331),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_3358),
.Y(n_3623)
);

CKINVDCx20_ASAP7_75t_R g3624 ( 
.A(n_3181),
.Y(n_3624)
);

NAND2x1p5_ASAP7_75t_L g3625 ( 
.A(n_3311),
.B(n_640),
.Y(n_3625)
);

INVx4_ASAP7_75t_SL g3626 ( 
.A(n_3403),
.Y(n_3626)
);

AND2x2_ASAP7_75t_L g3627 ( 
.A(n_3426),
.B(n_3358),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_3386),
.Y(n_3628)
);

NOR2xp67_ASAP7_75t_L g3629 ( 
.A(n_3616),
.B(n_3226),
.Y(n_3629)
);

INVx1_ASAP7_75t_L g3630 ( 
.A(n_3388),
.Y(n_3630)
);

HB1xp67_ASAP7_75t_L g3631 ( 
.A(n_3375),
.Y(n_3631)
);

AND2x4_ASAP7_75t_L g3632 ( 
.A(n_3489),
.B(n_3079),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3392),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3394),
.Y(n_3634)
);

OR2x2_ASAP7_75t_L g3635 ( 
.A(n_3383),
.B(n_3073),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_3400),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3404),
.Y(n_3637)
);

AND2x2_ASAP7_75t_L g3638 ( 
.A(n_3466),
.B(n_3073),
.Y(n_3638)
);

OAI21xp5_ASAP7_75t_L g3639 ( 
.A1(n_3548),
.A2(n_3482),
.B(n_3620),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3407),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3409),
.Y(n_3641)
);

INVx2_ASAP7_75t_L g3642 ( 
.A(n_3557),
.Y(n_3642)
);

BUFx2_ASAP7_75t_SL g3643 ( 
.A(n_3405),
.Y(n_3643)
);

BUFx12f_ASAP7_75t_L g3644 ( 
.A(n_3447),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3410),
.Y(n_3645)
);

AO21x2_ASAP7_75t_L g3646 ( 
.A1(n_3602),
.A2(n_3095),
.B(n_3125),
.Y(n_3646)
);

AND2x4_ASAP7_75t_L g3647 ( 
.A(n_3498),
.B(n_3073),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3416),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_3419),
.Y(n_3649)
);

INVx2_ASAP7_75t_L g3650 ( 
.A(n_3617),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_3422),
.Y(n_3651)
);

BUFx6f_ASAP7_75t_L g3652 ( 
.A(n_3423),
.Y(n_3652)
);

INVx2_ASAP7_75t_L g3653 ( 
.A(n_3609),
.Y(n_3653)
);

OA21x2_ASAP7_75t_L g3654 ( 
.A1(n_3603),
.A2(n_3111),
.B(n_3160),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3429),
.Y(n_3655)
);

INVx1_ASAP7_75t_L g3656 ( 
.A(n_3433),
.Y(n_3656)
);

BUFx3_ASAP7_75t_L g3657 ( 
.A(n_3384),
.Y(n_3657)
);

OA21x2_ASAP7_75t_L g3658 ( 
.A1(n_3612),
.A2(n_3197),
.B(n_3154),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_3440),
.Y(n_3659)
);

OAI21x1_ASAP7_75t_L g3660 ( 
.A1(n_3495),
.A2(n_3119),
.B(n_3104),
.Y(n_3660)
);

INVx1_ASAP7_75t_L g3661 ( 
.A(n_3441),
.Y(n_3661)
);

INVx3_ASAP7_75t_L g3662 ( 
.A(n_3532),
.Y(n_3662)
);

AND2x4_ASAP7_75t_L g3663 ( 
.A(n_3505),
.B(n_3074),
.Y(n_3663)
);

NOR2xp33_ASAP7_75t_L g3664 ( 
.A(n_3418),
.B(n_3121),
.Y(n_3664)
);

INVx2_ASAP7_75t_L g3665 ( 
.A(n_3562),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3442),
.Y(n_3666)
);

INVx4_ASAP7_75t_L g3667 ( 
.A(n_3403),
.Y(n_3667)
);

BUFx2_ASAP7_75t_L g3668 ( 
.A(n_3384),
.Y(n_3668)
);

AOI22xp5_ASAP7_75t_L g3669 ( 
.A1(n_3418),
.A2(n_3164),
.B1(n_3170),
.B2(n_3168),
.Y(n_3669)
);

AO21x1_ASAP7_75t_L g3670 ( 
.A1(n_3552),
.A2(n_3249),
.B(n_3246),
.Y(n_3670)
);

INVx2_ASAP7_75t_L g3671 ( 
.A(n_3563),
.Y(n_3671)
);

INVx2_ASAP7_75t_L g3672 ( 
.A(n_3510),
.Y(n_3672)
);

NAND2xp5_ASAP7_75t_L g3673 ( 
.A(n_3464),
.B(n_3157),
.Y(n_3673)
);

OR2x2_ASAP7_75t_L g3674 ( 
.A(n_3508),
.B(n_3093),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_L g3675 ( 
.A(n_3438),
.B(n_3174),
.Y(n_3675)
);

INVx1_ASAP7_75t_L g3676 ( 
.A(n_3455),
.Y(n_3676)
);

NAND2x1p5_ASAP7_75t_L g3677 ( 
.A(n_3399),
.B(n_3313),
.Y(n_3677)
);

INVx2_ASAP7_75t_L g3678 ( 
.A(n_3511),
.Y(n_3678)
);

INVx2_ASAP7_75t_L g3679 ( 
.A(n_3380),
.Y(n_3679)
);

AND2x2_ASAP7_75t_L g3680 ( 
.A(n_3443),
.B(n_3102),
.Y(n_3680)
);

INVx1_ASAP7_75t_L g3681 ( 
.A(n_3456),
.Y(n_3681)
);

AND2x2_ASAP7_75t_L g3682 ( 
.A(n_3467),
.B(n_3102),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3454),
.Y(n_3683)
);

INVx2_ASAP7_75t_L g3684 ( 
.A(n_3412),
.Y(n_3684)
);

AND2x2_ASAP7_75t_L g3685 ( 
.A(n_3518),
.B(n_3093),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3396),
.Y(n_3686)
);

OAI21x1_ASAP7_75t_L g3687 ( 
.A1(n_3499),
.A2(n_3127),
.B(n_3101),
.Y(n_3687)
);

BUFx3_ASAP7_75t_L g3688 ( 
.A(n_3504),
.Y(n_3688)
);

BUFx8_ASAP7_75t_SL g3689 ( 
.A(n_3374),
.Y(n_3689)
);

INVx3_ASAP7_75t_L g3690 ( 
.A(n_3532),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3479),
.Y(n_3691)
);

BUFx6f_ASAP7_75t_L g3692 ( 
.A(n_3423),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3517),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3521),
.Y(n_3694)
);

INVx2_ASAP7_75t_L g3695 ( 
.A(n_3427),
.Y(n_3695)
);

INVx3_ASAP7_75t_L g3696 ( 
.A(n_3423),
.Y(n_3696)
);

INVx2_ASAP7_75t_L g3697 ( 
.A(n_3444),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_3453),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3540),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3503),
.Y(n_3700)
);

INVx2_ASAP7_75t_L g3701 ( 
.A(n_3523),
.Y(n_3701)
);

INVx2_ASAP7_75t_L g3702 ( 
.A(n_3534),
.Y(n_3702)
);

INVx3_ASAP7_75t_L g3703 ( 
.A(n_3533),
.Y(n_3703)
);

INVx2_ASAP7_75t_L g3704 ( 
.A(n_3537),
.Y(n_3704)
);

OAI21x1_ASAP7_75t_L g3705 ( 
.A1(n_3500),
.A2(n_3149),
.B(n_3115),
.Y(n_3705)
);

INVx2_ASAP7_75t_L g3706 ( 
.A(n_3585),
.Y(n_3706)
);

INVx2_ASAP7_75t_L g3707 ( 
.A(n_3588),
.Y(n_3707)
);

OA21x2_ASAP7_75t_L g3708 ( 
.A1(n_3485),
.A2(n_3309),
.B(n_3304),
.Y(n_3708)
);

OAI21x1_ASAP7_75t_L g3709 ( 
.A1(n_3484),
.A2(n_3279),
.B(n_3277),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3570),
.Y(n_3710)
);

OAI21x1_ASAP7_75t_L g3711 ( 
.A1(n_3492),
.A2(n_3083),
.B(n_3281),
.Y(n_3711)
);

HB1xp67_ASAP7_75t_SL g3712 ( 
.A(n_3574),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3576),
.Y(n_3713)
);

OR2x2_ASAP7_75t_L g3714 ( 
.A(n_3373),
.B(n_3098),
.Y(n_3714)
);

INVx2_ASAP7_75t_SL g3715 ( 
.A(n_3397),
.Y(n_3715)
);

BUFx8_ASAP7_75t_L g3716 ( 
.A(n_3387),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3564),
.Y(n_3717)
);

INVx2_ASAP7_75t_L g3718 ( 
.A(n_3539),
.Y(n_3718)
);

AND2x2_ASAP7_75t_L g3719 ( 
.A(n_3512),
.B(n_3098),
.Y(n_3719)
);

OAI22xp5_ASAP7_75t_L g3720 ( 
.A1(n_3451),
.A2(n_3219),
.B1(n_3193),
.B2(n_3342),
.Y(n_3720)
);

INVx2_ASAP7_75t_L g3721 ( 
.A(n_3553),
.Y(n_3721)
);

BUFx3_ASAP7_75t_L g3722 ( 
.A(n_3445),
.Y(n_3722)
);

AO21x2_ASAP7_75t_L g3723 ( 
.A1(n_3620),
.A2(n_3288),
.B(n_3285),
.Y(n_3723)
);

AND2x2_ASAP7_75t_L g3724 ( 
.A(n_3472),
.B(n_3074),
.Y(n_3724)
);

INVxp67_ASAP7_75t_L g3725 ( 
.A(n_3556),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3572),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_3469),
.Y(n_3727)
);

OAI21x1_ASAP7_75t_L g3728 ( 
.A1(n_3481),
.A2(n_3300),
.B(n_3298),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_3470),
.Y(n_3729)
);

INVx1_ASAP7_75t_SL g3730 ( 
.A(n_3509),
.Y(n_3730)
);

NOR2xp33_ASAP7_75t_L g3731 ( 
.A(n_3507),
.B(n_3187),
.Y(n_3731)
);

HB1xp67_ASAP7_75t_L g3732 ( 
.A(n_3586),
.Y(n_3732)
);

OAI21x1_ASAP7_75t_L g3733 ( 
.A1(n_3501),
.A2(n_3341),
.B(n_3307),
.Y(n_3733)
);

AND2x4_ASAP7_75t_L g3734 ( 
.A(n_3573),
.B(n_3074),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_3471),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3589),
.Y(n_3736)
);

INVx3_ASAP7_75t_L g3737 ( 
.A(n_3477),
.Y(n_3737)
);

AND2x2_ASAP7_75t_L g3738 ( 
.A(n_3516),
.B(n_3069),
.Y(n_3738)
);

INVx2_ASAP7_75t_L g3739 ( 
.A(n_3561),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3623),
.Y(n_3740)
);

INVx2_ASAP7_75t_L g3741 ( 
.A(n_3561),
.Y(n_3741)
);

HB1xp67_ASAP7_75t_L g3742 ( 
.A(n_3607),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3595),
.Y(n_3743)
);

AND2x2_ASAP7_75t_L g3744 ( 
.A(n_3522),
.B(n_3069),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3595),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3487),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3599),
.Y(n_3747)
);

AND2x2_ASAP7_75t_L g3748 ( 
.A(n_3515),
.B(n_3069),
.Y(n_3748)
);

INVx2_ASAP7_75t_L g3749 ( 
.A(n_3561),
.Y(n_3749)
);

INVx2_ASAP7_75t_L g3750 ( 
.A(n_3618),
.Y(n_3750)
);

INVx1_ASAP7_75t_L g3751 ( 
.A(n_3605),
.Y(n_3751)
);

INVx2_ASAP7_75t_SL g3752 ( 
.A(n_3397),
.Y(n_3752)
);

OAI21x1_ASAP7_75t_L g3753 ( 
.A1(n_3491),
.A2(n_3359),
.B(n_3348),
.Y(n_3753)
);

OAI21x1_ASAP7_75t_L g3754 ( 
.A1(n_3619),
.A2(n_3370),
.B(n_3360),
.Y(n_3754)
);

INVx2_ASAP7_75t_L g3755 ( 
.A(n_3573),
.Y(n_3755)
);

INVx2_ASAP7_75t_L g3756 ( 
.A(n_3591),
.Y(n_3756)
);

INVx2_ASAP7_75t_L g3757 ( 
.A(n_3604),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_3415),
.Y(n_3758)
);

INVx2_ASAP7_75t_L g3759 ( 
.A(n_3582),
.Y(n_3759)
);

INVx2_ASAP7_75t_L g3760 ( 
.A(n_3571),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3415),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3574),
.Y(n_3762)
);

OAI22xp5_ASAP7_75t_L g3763 ( 
.A1(n_3408),
.A2(n_3356),
.B1(n_3205),
.B2(n_3156),
.Y(n_3763)
);

INVx2_ASAP7_75t_L g3764 ( 
.A(n_3581),
.Y(n_3764)
);

AO21x2_ASAP7_75t_L g3765 ( 
.A1(n_3493),
.A2(n_3322),
.B(n_3227),
.Y(n_3765)
);

INVx2_ASAP7_75t_L g3766 ( 
.A(n_3614),
.Y(n_3766)
);

INVx2_ASAP7_75t_L g3767 ( 
.A(n_3592),
.Y(n_3767)
);

BUFx2_ASAP7_75t_L g3768 ( 
.A(n_3382),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_3377),
.Y(n_3769)
);

INVx2_ASAP7_75t_SL g3770 ( 
.A(n_3382),
.Y(n_3770)
);

HB1xp67_ASAP7_75t_L g3771 ( 
.A(n_3592),
.Y(n_3771)
);

OAI21x1_ASAP7_75t_L g3772 ( 
.A1(n_3483),
.A2(n_3625),
.B(n_3493),
.Y(n_3772)
);

AND2x2_ASAP7_75t_L g3773 ( 
.A(n_3435),
.B(n_3089),
.Y(n_3773)
);

INVx2_ASAP7_75t_L g3774 ( 
.A(n_3551),
.Y(n_3774)
);

OAI21x1_ASAP7_75t_L g3775 ( 
.A1(n_3425),
.A2(n_3248),
.B(n_3204),
.Y(n_3775)
);

INVx2_ASAP7_75t_L g3776 ( 
.A(n_3590),
.Y(n_3776)
);

INVx2_ASAP7_75t_L g3777 ( 
.A(n_3430),
.Y(n_3777)
);

OR2x2_ASAP7_75t_L g3778 ( 
.A(n_3417),
.B(n_641),
.Y(n_3778)
);

INVx1_ASAP7_75t_L g3779 ( 
.A(n_3519),
.Y(n_3779)
);

INVx1_ASAP7_75t_L g3780 ( 
.A(n_3528),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3399),
.Y(n_3781)
);

INVx1_ASAP7_75t_L g3782 ( 
.A(n_3379),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3543),
.Y(n_3783)
);

NAND2x1p5_ASAP7_75t_L g3784 ( 
.A(n_3496),
.B(n_3148),
.Y(n_3784)
);

AND2x2_ASAP7_75t_L g3785 ( 
.A(n_3477),
.B(n_643),
.Y(n_3785)
);

INVx2_ASAP7_75t_L g3786 ( 
.A(n_3550),
.Y(n_3786)
);

INVx2_ASAP7_75t_L g3787 ( 
.A(n_3550),
.Y(n_3787)
);

NOR2xp33_ASAP7_75t_L g3788 ( 
.A(n_3569),
.B(n_3613),
.Y(n_3788)
);

HB1xp67_ASAP7_75t_L g3789 ( 
.A(n_3458),
.Y(n_3789)
);

INVx2_ASAP7_75t_L g3790 ( 
.A(n_3550),
.Y(n_3790)
);

AND2x2_ASAP7_75t_L g3791 ( 
.A(n_3477),
.B(n_643),
.Y(n_3791)
);

INVx1_ASAP7_75t_L g3792 ( 
.A(n_3601),
.Y(n_3792)
);

INVx3_ASAP7_75t_L g3793 ( 
.A(n_3458),
.Y(n_3793)
);

NAND2x1p5_ASAP7_75t_L g3794 ( 
.A(n_3496),
.B(n_3129),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3587),
.Y(n_3795)
);

INVx2_ASAP7_75t_L g3796 ( 
.A(n_3610),
.Y(n_3796)
);

NOR2xp33_ASAP7_75t_L g3797 ( 
.A(n_3408),
.B(n_645),
.Y(n_3797)
);

AND2x4_ASAP7_75t_L g3798 ( 
.A(n_3743),
.B(n_3450),
.Y(n_3798)
);

NOR2x1p5_ASAP7_75t_L g3799 ( 
.A(n_3703),
.B(n_3413),
.Y(n_3799)
);

AND2x2_ASAP7_75t_L g3800 ( 
.A(n_3776),
.B(n_3460),
.Y(n_3800)
);

AND2x2_ASAP7_75t_L g3801 ( 
.A(n_3776),
.B(n_3473),
.Y(n_3801)
);

AND2x2_ASAP7_75t_L g3802 ( 
.A(n_3686),
.B(n_3474),
.Y(n_3802)
);

BUFx3_ASAP7_75t_L g3803 ( 
.A(n_3688),
.Y(n_3803)
);

AOI22xp5_ASAP7_75t_L g3804 ( 
.A1(n_3731),
.A2(n_3461),
.B1(n_3389),
.B2(n_3488),
.Y(n_3804)
);

AOI221xp5_ASAP7_75t_L g3805 ( 
.A1(n_3664),
.A2(n_3381),
.B1(n_3391),
.B2(n_3497),
.C(n_3390),
.Y(n_3805)
);

AND2x2_ASAP7_75t_L g3806 ( 
.A(n_3762),
.B(n_3513),
.Y(n_3806)
);

OAI21xp5_ASAP7_75t_L g3807 ( 
.A1(n_3664),
.A2(n_3524),
.B(n_3502),
.Y(n_3807)
);

OA21x2_ASAP7_75t_L g3808 ( 
.A1(n_3772),
.A2(n_3611),
.B(n_3538),
.Y(n_3808)
);

AND2x2_ASAP7_75t_L g3809 ( 
.A(n_3781),
.B(n_3578),
.Y(n_3809)
);

AND2x2_ASAP7_75t_L g3810 ( 
.A(n_3631),
.B(n_3583),
.Y(n_3810)
);

AND2x6_ASAP7_75t_L g3811 ( 
.A(n_3703),
.B(n_3480),
.Y(n_3811)
);

A2O1A1Ixp33_ASAP7_75t_L g3812 ( 
.A1(n_3731),
.A2(n_3544),
.B(n_3545),
.C(n_3465),
.Y(n_3812)
);

AND2x2_ASAP7_75t_L g3813 ( 
.A(n_3631),
.B(n_3468),
.Y(n_3813)
);

AND2x6_ASAP7_75t_L g3814 ( 
.A(n_3786),
.B(n_3480),
.Y(n_3814)
);

OAI21xp5_ASAP7_75t_L g3815 ( 
.A1(n_3797),
.A2(n_3577),
.B(n_3568),
.Y(n_3815)
);

AO32x2_ASAP7_75t_L g3816 ( 
.A1(n_3763),
.A2(n_3610),
.A3(n_3452),
.B1(n_3457),
.B2(n_3462),
.Y(n_3816)
);

OAI21xp5_ASAP7_75t_L g3817 ( 
.A1(n_3797),
.A2(n_3545),
.B(n_3559),
.Y(n_3817)
);

NOR2xp33_ASAP7_75t_L g3818 ( 
.A(n_3758),
.B(n_3393),
.Y(n_3818)
);

OR2x6_ASAP7_75t_L g3819 ( 
.A(n_3667),
.B(n_3428),
.Y(n_3819)
);

AND2x2_ASAP7_75t_L g3820 ( 
.A(n_3744),
.B(n_3486),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3706),
.Y(n_3821)
);

AND2x2_ASAP7_75t_L g3822 ( 
.A(n_3699),
.B(n_3449),
.Y(n_3822)
);

AND2x2_ASAP7_75t_L g3823 ( 
.A(n_3782),
.B(n_3475),
.Y(n_3823)
);

AND2x2_ASAP7_75t_L g3824 ( 
.A(n_3738),
.B(n_3494),
.Y(n_3824)
);

OA21x2_ASAP7_75t_L g3825 ( 
.A1(n_3705),
.A2(n_3587),
.B(n_3448),
.Y(n_3825)
);

INVx2_ASAP7_75t_L g3826 ( 
.A(n_3679),
.Y(n_3826)
);

BUFx4f_ASAP7_75t_SL g3827 ( 
.A(n_3688),
.Y(n_3827)
);

AOI221xp5_ASAP7_75t_L g3828 ( 
.A1(n_3639),
.A2(n_3560),
.B1(n_3535),
.B2(n_3536),
.C(n_3398),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_3627),
.B(n_3436),
.Y(n_3829)
);

NOR2x1_ASAP7_75t_SL g3830 ( 
.A(n_3667),
.B(n_3490),
.Y(n_3830)
);

INVx1_ASAP7_75t_L g3831 ( 
.A(n_3628),
.Y(n_3831)
);

BUFx6f_ASAP7_75t_L g3832 ( 
.A(n_3652),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_L g3833 ( 
.A(n_3691),
.B(n_3436),
.Y(n_3833)
);

AND2x4_ASAP7_75t_L g3834 ( 
.A(n_3745),
.B(n_3624),
.Y(n_3834)
);

AOI21xp5_ASAP7_75t_SL g3835 ( 
.A1(n_3786),
.A2(n_3790),
.B(n_3787),
.Y(n_3835)
);

A2O1A1Ixp33_ASAP7_75t_L g3836 ( 
.A1(n_3788),
.A2(n_3376),
.B(n_3382),
.C(n_3520),
.Y(n_3836)
);

NOR2x1_ASAP7_75t_SL g3837 ( 
.A(n_3787),
.B(n_3478),
.Y(n_3837)
);

INVx2_ASAP7_75t_L g3838 ( 
.A(n_3679),
.Y(n_3838)
);

AND2x2_ASAP7_75t_L g3839 ( 
.A(n_3685),
.B(n_3414),
.Y(n_3839)
);

AND2x2_ASAP7_75t_L g3840 ( 
.A(n_3700),
.B(n_3414),
.Y(n_3840)
);

AO32x2_ASAP7_75t_L g3841 ( 
.A1(n_3720),
.A2(n_3514),
.A3(n_3555),
.B1(n_3598),
.B2(n_3579),
.Y(n_3841)
);

INVx2_ASAP7_75t_L g3842 ( 
.A(n_3684),
.Y(n_3842)
);

OAI22xp5_ASAP7_75t_L g3843 ( 
.A1(n_3712),
.A2(n_3421),
.B1(n_3547),
.B2(n_3520),
.Y(n_3843)
);

OAI21xp5_ASAP7_75t_L g3844 ( 
.A1(n_3783),
.A2(n_3584),
.B(n_3567),
.Y(n_3844)
);

INVx2_ASAP7_75t_L g3845 ( 
.A(n_3684),
.Y(n_3845)
);

OAI211xp5_ASAP7_75t_L g3846 ( 
.A1(n_3792),
.A2(n_3402),
.B(n_3424),
.C(n_3378),
.Y(n_3846)
);

NOR2xp33_ASAP7_75t_L g3847 ( 
.A(n_3761),
.B(n_3387),
.Y(n_3847)
);

INVx2_ASAP7_75t_L g3848 ( 
.A(n_3695),
.Y(n_3848)
);

AND2x4_ASAP7_75t_L g3849 ( 
.A(n_3759),
.B(n_3411),
.Y(n_3849)
);

AND2x4_ASAP7_75t_L g3850 ( 
.A(n_3759),
.B(n_3431),
.Y(n_3850)
);

AND2x2_ASAP7_75t_L g3851 ( 
.A(n_3769),
.B(n_3434),
.Y(n_3851)
);

AND2x2_ASAP7_75t_L g3852 ( 
.A(n_3779),
.B(n_3434),
.Y(n_3852)
);

AO32x2_ASAP7_75t_L g3853 ( 
.A1(n_3715),
.A2(n_3527),
.A3(n_3542),
.B1(n_3622),
.B2(n_3549),
.Y(n_3853)
);

INVx2_ASAP7_75t_SL g3854 ( 
.A(n_3716),
.Y(n_3854)
);

AOI221x1_ASAP7_75t_L g3855 ( 
.A1(n_3746),
.A2(n_3606),
.B1(n_3446),
.B2(n_3554),
.C(n_3547),
.Y(n_3855)
);

AO21x2_ASAP7_75t_L g3856 ( 
.A1(n_3767),
.A2(n_3621),
.B(n_3395),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_L g3857 ( 
.A(n_3748),
.B(n_3476),
.Y(n_3857)
);

NOR2xp33_ASAP7_75t_L g3858 ( 
.A(n_3657),
.B(n_3437),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_3706),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_3707),
.Y(n_3860)
);

AND2x2_ASAP7_75t_L g3861 ( 
.A(n_3727),
.B(n_3437),
.Y(n_3861)
);

AOI221xp5_ASAP7_75t_L g3862 ( 
.A1(n_3780),
.A2(n_3526),
.B1(n_3506),
.B2(n_3439),
.C(n_3566),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3707),
.Y(n_3863)
);

AND2x2_ASAP7_75t_L g3864 ( 
.A(n_3729),
.B(n_3463),
.Y(n_3864)
);

OAI22xp5_ASAP7_75t_L g3865 ( 
.A1(n_3712),
.A2(n_3546),
.B1(n_3621),
.B2(n_3597),
.Y(n_3865)
);

AO32x2_ASAP7_75t_L g3866 ( 
.A1(n_3752),
.A2(n_3204),
.A3(n_3558),
.B1(n_3615),
.B2(n_3580),
.Y(n_3866)
);

AND2x4_ASAP7_75t_L g3867 ( 
.A(n_3766),
.B(n_3459),
.Y(n_3867)
);

AND2x2_ASAP7_75t_L g3868 ( 
.A(n_3735),
.B(n_3463),
.Y(n_3868)
);

INVx1_ASAP7_75t_SL g3869 ( 
.A(n_3768),
.Y(n_3869)
);

AO21x2_ASAP7_75t_L g3870 ( 
.A1(n_3767),
.A2(n_3459),
.B(n_3420),
.Y(n_3870)
);

AOI221xp5_ASAP7_75t_L g3871 ( 
.A1(n_3724),
.A2(n_3593),
.B1(n_3575),
.B2(n_3596),
.C(n_3600),
.Y(n_3871)
);

AND2x2_ASAP7_75t_L g3872 ( 
.A(n_3777),
.B(n_3420),
.Y(n_3872)
);

BUFx12f_ASAP7_75t_L g3873 ( 
.A(n_3716),
.Y(n_3873)
);

INVx3_ASAP7_75t_L g3874 ( 
.A(n_3650),
.Y(n_3874)
);

A2O1A1Ixp33_ASAP7_75t_L g3875 ( 
.A1(n_3788),
.A2(n_3406),
.B(n_3525),
.C(n_3530),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_L g3876 ( 
.A(n_3777),
.B(n_3529),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_L g3877 ( 
.A(n_3638),
.B(n_3710),
.Y(n_3877)
);

OR2x6_ASAP7_75t_L g3878 ( 
.A(n_3644),
.B(n_3668),
.Y(n_3878)
);

A2O1A1Ixp33_ASAP7_75t_L g3879 ( 
.A1(n_3657),
.A2(n_3722),
.B(n_3790),
.C(n_3796),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_SL g3880 ( 
.A(n_3626),
.B(n_3432),
.Y(n_3880)
);

AND2x2_ASAP7_75t_L g3881 ( 
.A(n_3680),
.B(n_3428),
.Y(n_3881)
);

OR2x2_ASAP7_75t_L g3882 ( 
.A(n_3674),
.B(n_3129),
.Y(n_3882)
);

OAI21xp5_ASAP7_75t_L g3883 ( 
.A1(n_3796),
.A2(n_3608),
.B(n_3531),
.Y(n_3883)
);

OR2x2_ASAP7_75t_L g3884 ( 
.A(n_3714),
.B(n_646),
.Y(n_3884)
);

A2O1A1Ixp33_ASAP7_75t_L g3885 ( 
.A1(n_3722),
.A2(n_3541),
.B(n_3594),
.C(n_3565),
.Y(n_3885)
);

BUFx3_ASAP7_75t_L g3886 ( 
.A(n_3716),
.Y(n_3886)
);

OAI21x1_ASAP7_75t_L g3887 ( 
.A1(n_3660),
.A2(n_3208),
.B(n_3272),
.Y(n_3887)
);

AND2x6_ASAP7_75t_L g3888 ( 
.A(n_3766),
.B(n_3208),
.Y(n_3888)
);

INVx2_ASAP7_75t_L g3889 ( 
.A(n_3821),
.Y(n_3889)
);

OR2x2_ASAP7_75t_L g3890 ( 
.A(n_3877),
.B(n_3829),
.Y(n_3890)
);

INVx1_ASAP7_75t_L g3891 ( 
.A(n_3831),
.Y(n_3891)
);

AND2x2_ASAP7_75t_L g3892 ( 
.A(n_3839),
.B(n_3682),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_L g3893 ( 
.A(n_3833),
.B(n_3713),
.Y(n_3893)
);

BUFx6f_ASAP7_75t_L g3894 ( 
.A(n_3886),
.Y(n_3894)
);

OR2x2_ASAP7_75t_L g3895 ( 
.A(n_3882),
.B(n_3725),
.Y(n_3895)
);

HB1xp67_ASAP7_75t_L g3896 ( 
.A(n_3874),
.Y(n_3896)
);

BUFx6f_ASAP7_75t_L g3897 ( 
.A(n_3832),
.Y(n_3897)
);

INVx2_ASAP7_75t_L g3898 ( 
.A(n_3821),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_3872),
.Y(n_3899)
);

AND2x2_ASAP7_75t_L g3900 ( 
.A(n_3881),
.B(n_3719),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_3859),
.Y(n_3901)
);

INVx2_ASAP7_75t_L g3902 ( 
.A(n_3859),
.Y(n_3902)
);

AND2x2_ASAP7_75t_L g3903 ( 
.A(n_3820),
.B(n_3800),
.Y(n_3903)
);

AND2x2_ASAP7_75t_L g3904 ( 
.A(n_3834),
.B(n_3725),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3860),
.Y(n_3905)
);

INVx1_ASAP7_75t_L g3906 ( 
.A(n_3860),
.Y(n_3906)
);

CKINVDCx20_ASAP7_75t_R g3907 ( 
.A(n_3827),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3863),
.Y(n_3908)
);

INVx2_ASAP7_75t_L g3909 ( 
.A(n_3863),
.Y(n_3909)
);

OAI22xp5_ASAP7_75t_L g3910 ( 
.A1(n_3836),
.A2(n_3730),
.B1(n_3629),
.B2(n_3669),
.Y(n_3910)
);

INVx1_ASAP7_75t_L g3911 ( 
.A(n_3861),
.Y(n_3911)
);

OR2x2_ASAP7_75t_L g3912 ( 
.A(n_3826),
.B(n_3732),
.Y(n_3912)
);

INVx2_ASAP7_75t_L g3913 ( 
.A(n_3838),
.Y(n_3913)
);

INVx2_ASAP7_75t_L g3914 ( 
.A(n_3842),
.Y(n_3914)
);

AOI22xp33_ASAP7_75t_L g3915 ( 
.A1(n_3805),
.A2(n_3795),
.B1(n_3708),
.B2(n_3773),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3864),
.Y(n_3916)
);

AOI22xp33_ASAP7_75t_L g3917 ( 
.A1(n_3804),
.A2(n_3708),
.B1(n_3774),
.B2(n_3736),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3868),
.Y(n_3918)
);

AOI22xp33_ASAP7_75t_L g3919 ( 
.A1(n_3843),
.A2(n_3708),
.B1(n_3774),
.B2(n_3778),
.Y(n_3919)
);

AND2x2_ASAP7_75t_L g3920 ( 
.A(n_3834),
.B(n_3732),
.Y(n_3920)
);

NAND2xp5_ASAP7_75t_L g3921 ( 
.A(n_3802),
.B(n_3747),
.Y(n_3921)
);

AND2x2_ASAP7_75t_L g3922 ( 
.A(n_3810),
.B(n_3751),
.Y(n_3922)
);

AOI22xp5_ASAP7_75t_L g3923 ( 
.A1(n_3865),
.A2(n_3791),
.B1(n_3785),
.B2(n_3626),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3845),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3848),
.Y(n_3925)
);

AND2x2_ASAP7_75t_L g3926 ( 
.A(n_3801),
.B(n_3771),
.Y(n_3926)
);

INVxp67_ASAP7_75t_SL g3927 ( 
.A(n_3874),
.Y(n_3927)
);

AND2x4_ASAP7_75t_L g3928 ( 
.A(n_3867),
.B(n_3771),
.Y(n_3928)
);

AND2x4_ASAP7_75t_L g3929 ( 
.A(n_3867),
.B(n_3663),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3852),
.Y(n_3930)
);

AND2x4_ASAP7_75t_L g3931 ( 
.A(n_3870),
.B(n_3663),
.Y(n_3931)
);

AOI22xp33_ASAP7_75t_L g3932 ( 
.A1(n_3817),
.A2(n_3670),
.B1(n_3644),
.B2(n_3647),
.Y(n_3932)
);

HB1xp67_ASAP7_75t_L g3933 ( 
.A(n_3869),
.Y(n_3933)
);

HB1xp67_ASAP7_75t_L g3934 ( 
.A(n_3887),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3840),
.Y(n_3935)
);

OAI21xp33_ASAP7_75t_L g3936 ( 
.A1(n_3812),
.A2(n_3635),
.B(n_3663),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3851),
.Y(n_3937)
);

AND2x2_ASAP7_75t_L g3938 ( 
.A(n_3798),
.B(n_3813),
.Y(n_3938)
);

AOI22xp33_ASAP7_75t_SL g3939 ( 
.A1(n_3830),
.A2(n_3789),
.B1(n_3793),
.B2(n_3737),
.Y(n_3939)
);

HB1xp67_ASAP7_75t_L g3940 ( 
.A(n_3798),
.Y(n_3940)
);

INVx3_ASAP7_75t_L g3941 ( 
.A(n_3832),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3823),
.Y(n_3942)
);

AOI22xp33_ASAP7_75t_SL g3943 ( 
.A1(n_3830),
.A2(n_3789),
.B1(n_3793),
.B2(n_3737),
.Y(n_3943)
);

HB1xp67_ASAP7_75t_L g3944 ( 
.A(n_3824),
.Y(n_3944)
);

INVxp67_ASAP7_75t_SL g3945 ( 
.A(n_3884),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3822),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_3879),
.Y(n_3947)
);

AOI22xp33_ASAP7_75t_L g3948 ( 
.A1(n_3828),
.A2(n_3647),
.B1(n_3765),
.B2(n_3633),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_3857),
.B(n_3642),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3876),
.Y(n_3950)
);

NOR2xp33_ASAP7_75t_L g3951 ( 
.A(n_3875),
.B(n_3662),
.Y(n_3951)
);

AND2x2_ASAP7_75t_L g3952 ( 
.A(n_3809),
.B(n_3630),
.Y(n_3952)
);

INVx1_ASAP7_75t_L g3953 ( 
.A(n_3849),
.Y(n_3953)
);

INVx2_ASAP7_75t_L g3954 ( 
.A(n_3832),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3849),
.Y(n_3955)
);

INVx1_ASAP7_75t_L g3956 ( 
.A(n_3850),
.Y(n_3956)
);

OR2x2_ASAP7_75t_SL g3957 ( 
.A(n_3873),
.B(n_3808),
.Y(n_3957)
);

INVxp67_ASAP7_75t_L g3958 ( 
.A(n_3803),
.Y(n_3958)
);

AND2x4_ASAP7_75t_L g3959 ( 
.A(n_3929),
.B(n_3850),
.Y(n_3959)
);

NOR2xp33_ASAP7_75t_L g3960 ( 
.A(n_3894),
.B(n_3846),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3891),
.Y(n_3961)
);

INVx1_ASAP7_75t_L g3962 ( 
.A(n_3901),
.Y(n_3962)
);

OAI31xp33_ASAP7_75t_L g3963 ( 
.A1(n_3910),
.A2(n_3936),
.A3(n_3932),
.B(n_3951),
.Y(n_3963)
);

NOR2x1p5_ASAP7_75t_L g3964 ( 
.A(n_3894),
.B(n_3837),
.Y(n_3964)
);

AND2x4_ASAP7_75t_L g3965 ( 
.A(n_3929),
.B(n_3837),
.Y(n_3965)
);

AOI211xp5_ASAP7_75t_L g3966 ( 
.A1(n_3951),
.A2(n_3835),
.B(n_3807),
.C(n_3880),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_3905),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_3906),
.Y(n_3968)
);

AOI221xp5_ASAP7_75t_L g3969 ( 
.A1(n_3948),
.A2(n_3815),
.B1(n_3844),
.B2(n_3883),
.C(n_3862),
.Y(n_3969)
);

AND2x2_ASAP7_75t_L g3970 ( 
.A(n_3938),
.B(n_3806),
.Y(n_3970)
);

INVx2_ASAP7_75t_L g3971 ( 
.A(n_3896),
.Y(n_3971)
);

AND2x4_ASAP7_75t_L g3972 ( 
.A(n_3929),
.B(n_3940),
.Y(n_3972)
);

INVx1_ASAP7_75t_L g3973 ( 
.A(n_3908),
.Y(n_3973)
);

INVx1_ASAP7_75t_L g3974 ( 
.A(n_3949),
.Y(n_3974)
);

INVx1_ASAP7_75t_SL g3975 ( 
.A(n_3933),
.Y(n_3975)
);

NAND4xp25_ASAP7_75t_L g3976 ( 
.A(n_3932),
.B(n_3855),
.C(n_3885),
.D(n_3818),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_L g3977 ( 
.A(n_3950),
.B(n_3740),
.Y(n_3977)
);

INVxp67_ASAP7_75t_L g3978 ( 
.A(n_3933),
.Y(n_3978)
);

INVxp67_ASAP7_75t_SL g3979 ( 
.A(n_3896),
.Y(n_3979)
);

AND2x2_ASAP7_75t_L g3980 ( 
.A(n_3940),
.B(n_3878),
.Y(n_3980)
);

AOI21x1_ASAP7_75t_L g3981 ( 
.A1(n_3947),
.A2(n_3819),
.B(n_3878),
.Y(n_3981)
);

AND2x2_ASAP7_75t_L g3982 ( 
.A(n_3926),
.B(n_3742),
.Y(n_3982)
);

INVx2_ASAP7_75t_L g3983 ( 
.A(n_3912),
.Y(n_3983)
);

CKINVDCx20_ASAP7_75t_R g3984 ( 
.A(n_3907),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3895),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_L g3986 ( 
.A(n_3944),
.B(n_3717),
.Y(n_3986)
);

INVx1_ASAP7_75t_SL g3987 ( 
.A(n_3907),
.Y(n_3987)
);

AND2x2_ASAP7_75t_L g3988 ( 
.A(n_3903),
.B(n_3742),
.Y(n_3988)
);

INVx1_ASAP7_75t_L g3989 ( 
.A(n_3889),
.Y(n_3989)
);

AND2x4_ASAP7_75t_L g3990 ( 
.A(n_3928),
.B(n_3904),
.Y(n_3990)
);

AOI221xp5_ASAP7_75t_SL g3991 ( 
.A1(n_3957),
.A2(n_3847),
.B1(n_3643),
.B2(n_3637),
.C(n_3640),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3889),
.Y(n_3992)
);

AND2x2_ASAP7_75t_L g3993 ( 
.A(n_3920),
.B(n_3650),
.Y(n_3993)
);

OR2x2_ASAP7_75t_L g3994 ( 
.A(n_3890),
.B(n_3755),
.Y(n_3994)
);

INVx5_ASAP7_75t_L g3995 ( 
.A(n_3894),
.Y(n_3995)
);

INVx2_ASAP7_75t_L g3996 ( 
.A(n_3928),
.Y(n_3996)
);

AND2x4_ASAP7_75t_L g3997 ( 
.A(n_3928),
.B(n_3931),
.Y(n_3997)
);

INVx1_ASAP7_75t_L g3998 ( 
.A(n_3898),
.Y(n_3998)
);

OR2x2_ASAP7_75t_L g3999 ( 
.A(n_3944),
.B(n_3755),
.Y(n_3999)
);

INVx2_ASAP7_75t_L g4000 ( 
.A(n_3898),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_3902),
.Y(n_4001)
);

INVx2_ASAP7_75t_L g4002 ( 
.A(n_3902),
.Y(n_4002)
);

NOR2xp33_ASAP7_75t_L g4003 ( 
.A(n_3894),
.B(n_3854),
.Y(n_4003)
);

INVx1_ASAP7_75t_L g4004 ( 
.A(n_3909),
.Y(n_4004)
);

INVx1_ASAP7_75t_L g4005 ( 
.A(n_3909),
.Y(n_4005)
);

AND2x2_ASAP7_75t_L g4006 ( 
.A(n_3900),
.B(n_3756),
.Y(n_4006)
);

AND2x2_ASAP7_75t_L g4007 ( 
.A(n_3892),
.B(n_3756),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_3924),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_L g4009 ( 
.A(n_3925),
.B(n_3726),
.Y(n_4009)
);

OAI221xp5_ASAP7_75t_L g4010 ( 
.A1(n_3948),
.A2(n_3819),
.B1(n_3871),
.B2(n_3808),
.C(n_3858),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3913),
.Y(n_4011)
);

AND2x2_ASAP7_75t_L g4012 ( 
.A(n_3956),
.B(n_3757),
.Y(n_4012)
);

NAND3xp33_ASAP7_75t_L g4013 ( 
.A(n_3917),
.B(n_3825),
.C(n_3683),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_L g4014 ( 
.A(n_3917),
.B(n_3642),
.Y(n_4014)
);

INVx3_ASAP7_75t_L g4015 ( 
.A(n_3931),
.Y(n_4015)
);

INVx2_ASAP7_75t_L g4016 ( 
.A(n_3913),
.Y(n_4016)
);

OAI221xp5_ASAP7_75t_L g4017 ( 
.A1(n_3923),
.A2(n_3919),
.B1(n_3915),
.B2(n_3943),
.C(n_3939),
.Y(n_4017)
);

AOI221xp5_ASAP7_75t_L g4018 ( 
.A1(n_3915),
.A2(n_3636),
.B1(n_3645),
.B2(n_3641),
.C(n_3634),
.Y(n_4018)
);

INVx1_ASAP7_75t_L g4019 ( 
.A(n_3914),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_3914),
.Y(n_4020)
);

OR2x2_ASAP7_75t_L g4021 ( 
.A(n_3986),
.B(n_3942),
.Y(n_4021)
);

INVx1_ASAP7_75t_L g4022 ( 
.A(n_4009),
.Y(n_4022)
);

AND2x4_ASAP7_75t_SL g4023 ( 
.A(n_3965),
.B(n_3953),
.Y(n_4023)
);

AND2x2_ASAP7_75t_L g4024 ( 
.A(n_3988),
.B(n_3955),
.Y(n_4024)
);

OR2x2_ASAP7_75t_L g4025 ( 
.A(n_3986),
.B(n_3893),
.Y(n_4025)
);

INVx1_ASAP7_75t_L g4026 ( 
.A(n_3989),
.Y(n_4026)
);

AND2x4_ASAP7_75t_L g4027 ( 
.A(n_3964),
.B(n_3931),
.Y(n_4027)
);

INVx1_ASAP7_75t_L g4028 ( 
.A(n_4009),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_3962),
.Y(n_4029)
);

NAND4xp25_ASAP7_75t_L g4030 ( 
.A(n_3969),
.B(n_3919),
.C(n_3958),
.D(n_3946),
.Y(n_4030)
);

AND2x2_ASAP7_75t_L g4031 ( 
.A(n_3996),
.B(n_3952),
.Y(n_4031)
);

NOR3xp33_ASAP7_75t_L g4032 ( 
.A(n_3976),
.B(n_3934),
.C(n_3690),
.Y(n_4032)
);

INVx2_ASAP7_75t_L g4033 ( 
.A(n_4000),
.Y(n_4033)
);

OR2x2_ASAP7_75t_L g4034 ( 
.A(n_3975),
.B(n_3921),
.Y(n_4034)
);

AND2x2_ASAP7_75t_L g4035 ( 
.A(n_3997),
.B(n_3922),
.Y(n_4035)
);

INVx2_ASAP7_75t_L g4036 ( 
.A(n_4002),
.Y(n_4036)
);

INVx1_ASAP7_75t_L g4037 ( 
.A(n_3992),
.Y(n_4037)
);

NAND2xp5_ASAP7_75t_L g4038 ( 
.A(n_4018),
.B(n_3945),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3998),
.Y(n_4039)
);

INVx3_ASAP7_75t_L g4040 ( 
.A(n_3965),
.Y(n_4040)
);

INVx1_ASAP7_75t_L g4041 ( 
.A(n_3967),
.Y(n_4041)
);

AND2x4_ASAP7_75t_L g4042 ( 
.A(n_3981),
.B(n_3934),
.Y(n_4042)
);

INVx2_ASAP7_75t_L g4043 ( 
.A(n_4016),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_3968),
.Y(n_4044)
);

AND2x2_ASAP7_75t_L g4045 ( 
.A(n_3997),
.B(n_3935),
.Y(n_4045)
);

AND2x2_ASAP7_75t_L g4046 ( 
.A(n_3975),
.B(n_3899),
.Y(n_4046)
);

INVx2_ASAP7_75t_L g4047 ( 
.A(n_3999),
.Y(n_4047)
);

AND2x2_ASAP7_75t_L g4048 ( 
.A(n_3972),
.B(n_3930),
.Y(n_4048)
);

AND2x2_ASAP7_75t_L g4049 ( 
.A(n_3972),
.B(n_3937),
.Y(n_4049)
);

AND2x2_ASAP7_75t_L g4050 ( 
.A(n_4015),
.B(n_3911),
.Y(n_4050)
);

AND2x2_ASAP7_75t_L g4051 ( 
.A(n_4015),
.B(n_3916),
.Y(n_4051)
);

AND2x2_ASAP7_75t_L g4052 ( 
.A(n_3982),
.B(n_3918),
.Y(n_4052)
);

AOI22xp5_ASAP7_75t_L g4053 ( 
.A1(n_3976),
.A2(n_3811),
.B1(n_3856),
.B2(n_3814),
.Y(n_4053)
);

OR2x2_ASAP7_75t_L g4054 ( 
.A(n_3974),
.B(n_3927),
.Y(n_4054)
);

NAND2xp5_ASAP7_75t_L g4055 ( 
.A(n_4014),
.B(n_3888),
.Y(n_4055)
);

AND2x2_ASAP7_75t_L g4056 ( 
.A(n_3980),
.B(n_3954),
.Y(n_4056)
);

AND2x4_ASAP7_75t_L g4057 ( 
.A(n_3959),
.B(n_3941),
.Y(n_4057)
);

NAND2xp5_ASAP7_75t_L g4058 ( 
.A(n_4014),
.B(n_3888),
.Y(n_4058)
);

INVx2_ASAP7_75t_L g4059 ( 
.A(n_3971),
.Y(n_4059)
);

INVx1_ASAP7_75t_L g4060 ( 
.A(n_3973),
.Y(n_4060)
);

AND2x2_ASAP7_75t_L g4061 ( 
.A(n_3979),
.B(n_3954),
.Y(n_4061)
);

AOI21xp33_ASAP7_75t_L g4062 ( 
.A1(n_4038),
.A2(n_4010),
.B(n_3963),
.Y(n_4062)
);

AND2x2_ASAP7_75t_L g4063 ( 
.A(n_4040),
.B(n_3959),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_4021),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_4021),
.Y(n_4065)
);

INVx2_ASAP7_75t_SL g4066 ( 
.A(n_4023),
.Y(n_4066)
);

INVx1_ASAP7_75t_L g4067 ( 
.A(n_4022),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_4028),
.Y(n_4068)
);

NAND2xp5_ASAP7_75t_L g4069 ( 
.A(n_4025),
.B(n_3978),
.Y(n_4069)
);

NAND2xp5_ASAP7_75t_L g4070 ( 
.A(n_4025),
.B(n_3963),
.Y(n_4070)
);

INVx2_ASAP7_75t_L g4071 ( 
.A(n_4054),
.Y(n_4071)
);

INVx1_ASAP7_75t_L g4072 ( 
.A(n_4029),
.Y(n_4072)
);

AND2x2_ASAP7_75t_L g4073 ( 
.A(n_4040),
.B(n_3990),
.Y(n_4073)
);

NAND2xp5_ASAP7_75t_L g4074 ( 
.A(n_4030),
.B(n_3985),
.Y(n_4074)
);

INVx1_ASAP7_75t_L g4075 ( 
.A(n_4041),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_4044),
.Y(n_4076)
);

AND2x2_ASAP7_75t_L g4077 ( 
.A(n_4040),
.B(n_3990),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_4060),
.Y(n_4078)
);

OR2x2_ASAP7_75t_L g4079 ( 
.A(n_4034),
.B(n_3994),
.Y(n_4079)
);

NAND2xp5_ASAP7_75t_L g4080 ( 
.A(n_4026),
.B(n_3961),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_4034),
.Y(n_4081)
);

INVx1_ASAP7_75t_L g4082 ( 
.A(n_4046),
.Y(n_4082)
);

NAND2xp5_ASAP7_75t_L g4083 ( 
.A(n_4026),
.B(n_4037),
.Y(n_4083)
);

NOR2x1_ASAP7_75t_L g4084 ( 
.A(n_4027),
.B(n_3799),
.Y(n_4084)
);

AND2x2_ASAP7_75t_L g4085 ( 
.A(n_4023),
.B(n_3970),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_L g4086 ( 
.A(n_4037),
.B(n_3977),
.Y(n_4086)
);

INVxp67_ASAP7_75t_L g4087 ( 
.A(n_4032),
.Y(n_4087)
);

INVx2_ASAP7_75t_L g4088 ( 
.A(n_4054),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_4046),
.Y(n_4089)
);

NOR2xp67_ASAP7_75t_L g4090 ( 
.A(n_4027),
.B(n_3995),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_4039),
.Y(n_4091)
);

NOR2xp33_ASAP7_75t_SL g4092 ( 
.A(n_4027),
.B(n_3995),
.Y(n_4092)
);

NAND2xp5_ASAP7_75t_L g4093 ( 
.A(n_4053),
.B(n_3966),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_4039),
.Y(n_4094)
);

INVx1_ASAP7_75t_L g4095 ( 
.A(n_4052),
.Y(n_4095)
);

INVx2_ASAP7_75t_L g4096 ( 
.A(n_4061),
.Y(n_4096)
);

CKINVDCx16_ASAP7_75t_R g4097 ( 
.A(n_4035),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_L g4098 ( 
.A(n_4033),
.B(n_3977),
.Y(n_4098)
);

NAND2xp5_ASAP7_75t_L g4099 ( 
.A(n_4033),
.B(n_4008),
.Y(n_4099)
);

OR2x6_ASAP7_75t_L g4100 ( 
.A(n_4042),
.B(n_3960),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_4052),
.Y(n_4101)
);

AND2x2_ASAP7_75t_L g4102 ( 
.A(n_4097),
.B(n_4050),
.Y(n_4102)
);

NAND2xp5_ASAP7_75t_L g4103 ( 
.A(n_4070),
.B(n_3966),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_4086),
.Y(n_4104)
);

INVx2_ASAP7_75t_L g4105 ( 
.A(n_4071),
.Y(n_4105)
);

AOI22xp33_ASAP7_75t_L g4106 ( 
.A1(n_4062),
.A2(n_4017),
.B1(n_4042),
.B2(n_4013),
.Y(n_4106)
);

NAND2xp5_ASAP7_75t_L g4107 ( 
.A(n_4074),
.B(n_4013),
.Y(n_4107)
);

AND2x2_ASAP7_75t_L g4108 ( 
.A(n_4087),
.B(n_4050),
.Y(n_4108)
);

NOR2xp33_ASAP7_75t_L g4109 ( 
.A(n_4066),
.B(n_3987),
.Y(n_4109)
);

AND2x2_ASAP7_75t_L g4110 ( 
.A(n_4088),
.B(n_4051),
.Y(n_4110)
);

INVx2_ASAP7_75t_L g4111 ( 
.A(n_4096),
.Y(n_4111)
);

OR2x2_ASAP7_75t_L g4112 ( 
.A(n_4086),
.B(n_4036),
.Y(n_4112)
);

INVx3_ASAP7_75t_L g4113 ( 
.A(n_4100),
.Y(n_4113)
);

INVxp67_ASAP7_75t_SL g4114 ( 
.A(n_4093),
.Y(n_4114)
);

AND2x2_ASAP7_75t_L g4115 ( 
.A(n_4063),
.B(n_4051),
.Y(n_4115)
);

AND2x2_ASAP7_75t_SL g4116 ( 
.A(n_4092),
.B(n_4042),
.Y(n_4116)
);

INVxp67_ASAP7_75t_L g4117 ( 
.A(n_4100),
.Y(n_4117)
);

OR2x2_ASAP7_75t_L g4118 ( 
.A(n_4067),
.B(n_4036),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_4098),
.Y(n_4119)
);

INVx2_ASAP7_75t_L g4120 ( 
.A(n_4081),
.Y(n_4120)
);

NAND2xp5_ASAP7_75t_L g4121 ( 
.A(n_4062),
.B(n_4045),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_4098),
.Y(n_4122)
);

NAND2xp5_ASAP7_75t_L g4123 ( 
.A(n_4095),
.B(n_4045),
.Y(n_4123)
);

AND2x2_ASAP7_75t_L g4124 ( 
.A(n_4073),
.B(n_4056),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_4083),
.Y(n_4125)
);

INVx2_ASAP7_75t_L g4126 ( 
.A(n_4082),
.Y(n_4126)
);

INVx1_ASAP7_75t_L g4127 ( 
.A(n_4083),
.Y(n_4127)
);

INVx1_ASAP7_75t_L g4128 ( 
.A(n_4080),
.Y(n_4128)
);

NAND2xp5_ASAP7_75t_L g4129 ( 
.A(n_4128),
.B(n_4064),
.Y(n_4129)
);

INVx2_ASAP7_75t_L g4130 ( 
.A(n_4110),
.Y(n_4130)
);

AOI21xp33_ASAP7_75t_L g4131 ( 
.A1(n_4114),
.A2(n_4100),
.B(n_3987),
.Y(n_4131)
);

INVxp67_ASAP7_75t_L g4132 ( 
.A(n_4109),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_4108),
.Y(n_4133)
);

NOR2xp33_ASAP7_75t_L g4134 ( 
.A(n_4117),
.B(n_3984),
.Y(n_4134)
);

INVx2_ASAP7_75t_L g4135 ( 
.A(n_4110),
.Y(n_4135)
);

CKINVDCx14_ASAP7_75t_R g4136 ( 
.A(n_4113),
.Y(n_4136)
);

NAND3xp33_ASAP7_75t_L g4137 ( 
.A(n_4106),
.B(n_4092),
.C(n_4084),
.Y(n_4137)
);

AND2x2_ASAP7_75t_L g4138 ( 
.A(n_4102),
.B(n_4077),
.Y(n_4138)
);

NAND2x1p5_ASAP7_75t_L g4139 ( 
.A(n_4113),
.B(n_3995),
.Y(n_4139)
);

OAI21xp33_ASAP7_75t_L g4140 ( 
.A1(n_4103),
.A2(n_4069),
.B(n_4065),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_4108),
.Y(n_4141)
);

INVx1_ASAP7_75t_L g4142 ( 
.A(n_4120),
.Y(n_4142)
);

OR2x2_ASAP7_75t_L g4143 ( 
.A(n_4105),
.B(n_4089),
.Y(n_4143)
);

NAND2xp5_ASAP7_75t_SL g4144 ( 
.A(n_4116),
.B(n_4090),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_4120),
.Y(n_4145)
);

INVx2_ASAP7_75t_SL g4146 ( 
.A(n_4113),
.Y(n_4146)
);

INVx2_ASAP7_75t_L g4147 ( 
.A(n_4105),
.Y(n_4147)
);

NAND2xp5_ASAP7_75t_L g4148 ( 
.A(n_4128),
.B(n_4119),
.Y(n_4148)
);

INVxp67_ASAP7_75t_L g4149 ( 
.A(n_4121),
.Y(n_4149)
);

AOI21xp33_ASAP7_75t_SL g4150 ( 
.A1(n_4116),
.A2(n_4003),
.B(n_4068),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_L g4151 ( 
.A(n_4146),
.B(n_4102),
.Y(n_4151)
);

AOI21xp33_ASAP7_75t_L g4152 ( 
.A1(n_4136),
.A2(n_4107),
.B(n_4125),
.Y(n_4152)
);

NAND2xp5_ASAP7_75t_SL g4153 ( 
.A(n_4137),
.B(n_4111),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_4147),
.Y(n_4154)
);

INVxp67_ASAP7_75t_SL g4155 ( 
.A(n_4134),
.Y(n_4155)
);

AOI22xp5_ASAP7_75t_L g4156 ( 
.A1(n_4132),
.A2(n_4126),
.B1(n_4122),
.B2(n_4119),
.Y(n_4156)
);

AOI22xp5_ASAP7_75t_L g4157 ( 
.A1(n_4140),
.A2(n_4126),
.B1(n_4122),
.B2(n_4104),
.Y(n_4157)
);

OAI21xp5_ASAP7_75t_SL g4158 ( 
.A1(n_4131),
.A2(n_4127),
.B(n_4125),
.Y(n_4158)
);

AOI22xp5_ASAP7_75t_L g4159 ( 
.A1(n_4149),
.A2(n_4115),
.B1(n_4127),
.B2(n_4111),
.Y(n_4159)
);

NOR2x1_ASAP7_75t_L g4160 ( 
.A(n_4144),
.B(n_4118),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_SL g4161 ( 
.A(n_4131),
.B(n_4118),
.Y(n_4161)
);

O2A1O1Ixp33_ASAP7_75t_SL g4162 ( 
.A1(n_4150),
.A2(n_4133),
.B(n_4141),
.C(n_4129),
.Y(n_4162)
);

OAI221xp5_ASAP7_75t_L g4163 ( 
.A1(n_4139),
.A2(n_3991),
.B1(n_4112),
.B2(n_4123),
.C(n_4115),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_4142),
.Y(n_4164)
);

OAI22xp5_ASAP7_75t_L g4165 ( 
.A1(n_4130),
.A2(n_4112),
.B1(n_4124),
.B2(n_4101),
.Y(n_4165)
);

AOI222xp33_ASAP7_75t_L g4166 ( 
.A1(n_4148),
.A2(n_4075),
.B1(n_4076),
.B2(n_4078),
.C1(n_4072),
.C2(n_4091),
.Y(n_4166)
);

OAI21xp5_ASAP7_75t_L g4167 ( 
.A1(n_4148),
.A2(n_4124),
.B(n_3991),
.Y(n_4167)
);

AO21x1_ASAP7_75t_L g4168 ( 
.A1(n_4139),
.A2(n_4094),
.B(n_4080),
.Y(n_4168)
);

AND4x1_ASAP7_75t_L g4169 ( 
.A(n_4138),
.B(n_4085),
.C(n_3401),
.D(n_3385),
.Y(n_4169)
);

OAI21xp5_ASAP7_75t_SL g4170 ( 
.A1(n_4129),
.A2(n_4058),
.B(n_4055),
.Y(n_4170)
);

OAI21xp5_ASAP7_75t_SL g4171 ( 
.A1(n_4145),
.A2(n_4057),
.B(n_3770),
.Y(n_4171)
);

AOI22xp33_ASAP7_75t_L g4172 ( 
.A1(n_4135),
.A2(n_3811),
.B1(n_3814),
.B2(n_4057),
.Y(n_4172)
);

AOI22xp5_ASAP7_75t_L g4173 ( 
.A1(n_4143),
.A2(n_4057),
.B1(n_4056),
.B2(n_4061),
.Y(n_4173)
);

AND2x2_ASAP7_75t_L g4174 ( 
.A(n_4138),
.B(n_4035),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_4151),
.Y(n_4175)
);

INVx1_ASAP7_75t_SL g4176 ( 
.A(n_4154),
.Y(n_4176)
);

AOI22xp5_ASAP7_75t_L g4177 ( 
.A1(n_4155),
.A2(n_4165),
.B1(n_4153),
.B2(n_4161),
.Y(n_4177)
);

AOI211xp5_ASAP7_75t_SL g4178 ( 
.A1(n_4152),
.A2(n_3689),
.B(n_4099),
.C(n_3690),
.Y(n_4178)
);

OAI331xp33_ASAP7_75t_L g4179 ( 
.A1(n_4164),
.A2(n_3853),
.A3(n_3689),
.B1(n_3626),
.B2(n_4099),
.B3(n_3816),
.C1(n_4059),
.Y(n_4179)
);

AOI31xp33_ASAP7_75t_SL g4180 ( 
.A1(n_4166),
.A2(n_4079),
.A3(n_4059),
.B(n_4047),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_4159),
.Y(n_4181)
);

NAND2xp5_ASAP7_75t_L g4182 ( 
.A(n_4174),
.B(n_4048),
.Y(n_4182)
);

OAI22xp33_ASAP7_75t_SL g4183 ( 
.A1(n_4163),
.A2(n_3995),
.B1(n_4043),
.B2(n_4047),
.Y(n_4183)
);

OAI222xp33_ASAP7_75t_L g4184 ( 
.A1(n_4160),
.A2(n_4156),
.B1(n_4157),
.B2(n_4172),
.C1(n_4173),
.C2(n_4162),
.Y(n_4184)
);

OAI22xp33_ASAP7_75t_SL g4185 ( 
.A1(n_4167),
.A2(n_4043),
.B1(n_3662),
.B2(n_3677),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_4168),
.Y(n_4186)
);

INVx2_ASAP7_75t_SL g4187 ( 
.A(n_4169),
.Y(n_4187)
);

OAI21xp33_ASAP7_75t_L g4188 ( 
.A1(n_4158),
.A2(n_4049),
.B(n_4048),
.Y(n_4188)
);

OR2x2_ASAP7_75t_L g4189 ( 
.A(n_4167),
.B(n_3983),
.Y(n_4189)
);

NOR2xp33_ASAP7_75t_L g4190 ( 
.A(n_4171),
.B(n_4049),
.Y(n_4190)
);

INVx3_ASAP7_75t_L g4191 ( 
.A(n_4170),
.Y(n_4191)
);

O2A1O1Ixp5_ASAP7_75t_L g4192 ( 
.A1(n_4153),
.A2(n_4024),
.B(n_4031),
.C(n_3941),
.Y(n_4192)
);

AOI22xp5_ASAP7_75t_L g4193 ( 
.A1(n_4155),
.A2(n_3811),
.B1(n_4024),
.B2(n_4031),
.Y(n_4193)
);

OR2x2_ASAP7_75t_L g4194 ( 
.A(n_4151),
.B(n_3993),
.Y(n_4194)
);

INVx1_ASAP7_75t_L g4195 ( 
.A(n_4151),
.Y(n_4195)
);

HB1xp67_ASAP7_75t_L g4196 ( 
.A(n_4154),
.Y(n_4196)
);

NAND2xp33_ASAP7_75t_L g4197 ( 
.A(n_4151),
.B(n_3811),
.Y(n_4197)
);

AND2x2_ASAP7_75t_L g4198 ( 
.A(n_4174),
.B(n_4007),
.Y(n_4198)
);

NAND3x2_ASAP7_75t_L g4199 ( 
.A(n_4154),
.B(n_3853),
.C(n_4012),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_4151),
.Y(n_4200)
);

NAND2xp5_ASAP7_75t_L g4201 ( 
.A(n_4177),
.B(n_4001),
.Y(n_4201)
);

AOI22xp5_ASAP7_75t_L g4202 ( 
.A1(n_4179),
.A2(n_3814),
.B1(n_3825),
.B2(n_3888),
.Y(n_4202)
);

OAI22xp5_ASAP7_75t_L g4203 ( 
.A1(n_4187),
.A2(n_3941),
.B1(n_4019),
.B2(n_4011),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_4196),
.Y(n_4204)
);

NAND2xp5_ASAP7_75t_L g4205 ( 
.A(n_4176),
.B(n_4004),
.Y(n_4205)
);

NAND3xp33_ASAP7_75t_L g4206 ( 
.A(n_4181),
.B(n_4005),
.C(n_3648),
.Y(n_4206)
);

NAND2xp5_ASAP7_75t_L g4207 ( 
.A(n_4188),
.B(n_4020),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_SL g4208 ( 
.A(n_4183),
.B(n_4191),
.Y(n_4208)
);

NAND4xp25_ASAP7_75t_L g4209 ( 
.A(n_4178),
.B(n_3853),
.C(n_3696),
.D(n_3816),
.Y(n_4209)
);

INVx1_ASAP7_75t_SL g4210 ( 
.A(n_4175),
.Y(n_4210)
);

BUFx4f_ASAP7_75t_SL g4211 ( 
.A(n_4195),
.Y(n_4211)
);

NOR3xp33_ASAP7_75t_L g4212 ( 
.A(n_4184),
.B(n_646),
.C(n_647),
.Y(n_4212)
);

NOR2x1_ASAP7_75t_L g4213 ( 
.A(n_4186),
.B(n_3765),
.Y(n_4213)
);

AND2x2_ASAP7_75t_L g4214 ( 
.A(n_4198),
.B(n_4006),
.Y(n_4214)
);

NAND2xp5_ASAP7_75t_SL g4215 ( 
.A(n_4191),
.B(n_3897),
.Y(n_4215)
);

AOI21xp5_ASAP7_75t_L g4216 ( 
.A1(n_4200),
.A2(n_3673),
.B(n_3661),
.Y(n_4216)
);

NOR3xp33_ASAP7_75t_SL g4217 ( 
.A(n_4188),
.B(n_647),
.C(n_648),
.Y(n_4217)
);

INVx1_ASAP7_75t_L g4218 ( 
.A(n_4189),
.Y(n_4218)
);

NOR2xp33_ASAP7_75t_L g4219 ( 
.A(n_4194),
.B(n_3659),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_L g4220 ( 
.A(n_4182),
.B(n_3666),
.Y(n_4220)
);

NOR2x1_ASAP7_75t_L g4221 ( 
.A(n_4180),
.B(n_3723),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_L g4222 ( 
.A(n_4190),
.B(n_3676),
.Y(n_4222)
);

NOR2xp33_ASAP7_75t_SL g4223 ( 
.A(n_4185),
.B(n_4197),
.Y(n_4223)
);

NAND5xp2_ASAP7_75t_L g4224 ( 
.A(n_4193),
.B(n_3677),
.C(n_3784),
.D(n_3794),
.E(n_3816),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_4192),
.Y(n_4225)
);

NAND2xp33_ASAP7_75t_L g4226 ( 
.A(n_4199),
.B(n_3652),
.Y(n_4226)
);

AOI211xp5_ASAP7_75t_SL g4227 ( 
.A1(n_4184),
.A2(n_3696),
.B(n_3681),
.C(n_3675),
.Y(n_4227)
);

NAND2xp5_ASAP7_75t_L g4228 ( 
.A(n_4177),
.B(n_3649),
.Y(n_4228)
);

OAI221xp5_ASAP7_75t_L g4229 ( 
.A1(n_4187),
.A2(n_3784),
.B1(n_3794),
.B2(n_3897),
.C(n_3655),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_4196),
.Y(n_4230)
);

NAND3xp33_ASAP7_75t_L g4231 ( 
.A(n_4177),
.B(n_3656),
.C(n_3651),
.Y(n_4231)
);

AOI31xp33_ASAP7_75t_L g4232 ( 
.A1(n_4210),
.A2(n_651),
.A3(n_649),
.B(n_650),
.Y(n_4232)
);

AOI21xp5_ASAP7_75t_L g4233 ( 
.A1(n_4208),
.A2(n_3723),
.B(n_3775),
.Y(n_4233)
);

INVx1_ASAP7_75t_SL g4234 ( 
.A(n_4211),
.Y(n_4234)
);

O2A1O1Ixp33_ASAP7_75t_L g4235 ( 
.A1(n_4212),
.A2(n_652),
.B(n_650),
.C(n_651),
.Y(n_4235)
);

AOI221x1_ASAP7_75t_L g4236 ( 
.A1(n_4204),
.A2(n_3897),
.B1(n_653),
.B2(n_654),
.C(n_655),
.Y(n_4236)
);

INVx1_ASAP7_75t_L g4237 ( 
.A(n_4218),
.Y(n_4237)
);

NOR2xp33_ASAP7_75t_R g4238 ( 
.A(n_4230),
.B(n_652),
.Y(n_4238)
);

NAND4xp25_ASAP7_75t_L g4239 ( 
.A(n_4227),
.B(n_657),
.C(n_653),
.D(n_656),
.Y(n_4239)
);

AOI221xp5_ASAP7_75t_L g4240 ( 
.A1(n_4225),
.A2(n_3693),
.B1(n_3694),
.B2(n_3647),
.C(n_3734),
.Y(n_4240)
);

NAND2xp5_ASAP7_75t_L g4241 ( 
.A(n_4217),
.B(n_3888),
.Y(n_4241)
);

O2A1O1Ixp33_ASAP7_75t_L g4242 ( 
.A1(n_4215),
.A2(n_658),
.B(n_656),
.C(n_657),
.Y(n_4242)
);

NAND2x1_ASAP7_75t_L g4243 ( 
.A(n_4205),
.B(n_4201),
.Y(n_4243)
);

OAI22xp33_ASAP7_75t_L g4244 ( 
.A1(n_4209),
.A2(n_3897),
.B1(n_3692),
.B2(n_3652),
.Y(n_4244)
);

NAND4xp25_ASAP7_75t_L g4245 ( 
.A(n_4223),
.B(n_660),
.C(n_658),
.D(n_659),
.Y(n_4245)
);

NOR3xp33_ASAP7_75t_SL g4246 ( 
.A(n_4229),
.B(n_660),
.C(n_661),
.Y(n_4246)
);

AOI221xp5_ASAP7_75t_L g4247 ( 
.A1(n_4228),
.A2(n_4203),
.B1(n_4207),
.B2(n_4231),
.C(n_4224),
.Y(n_4247)
);

A2O1A1Ixp33_ASAP7_75t_L g4248 ( 
.A1(n_4219),
.A2(n_3775),
.B(n_3754),
.C(n_3728),
.Y(n_4248)
);

AOI221xp5_ASAP7_75t_L g4249 ( 
.A1(n_4226),
.A2(n_3734),
.B1(n_3698),
.B2(n_3764),
.C(n_3760),
.Y(n_4249)
);

NAND2x1_ASAP7_75t_SL g4250 ( 
.A(n_4213),
.B(n_662),
.Y(n_4250)
);

OAI21xp33_ASAP7_75t_SL g4251 ( 
.A1(n_4221),
.A2(n_3753),
.B(n_3754),
.Y(n_4251)
);

A2O1A1Ixp33_ASAP7_75t_SL g4252 ( 
.A1(n_4222),
.A2(n_666),
.B(n_663),
.C(n_664),
.Y(n_4252)
);

NOR2xp33_ASAP7_75t_L g4253 ( 
.A(n_4206),
.B(n_4220),
.Y(n_4253)
);

OAI22xp5_ASAP7_75t_L g4254 ( 
.A1(n_4202),
.A2(n_4216),
.B1(n_4214),
.B2(n_3652),
.Y(n_4254)
);

AOI21x1_ASAP7_75t_L g4255 ( 
.A1(n_4216),
.A2(n_663),
.B(n_664),
.Y(n_4255)
);

AOI21xp5_ASAP7_75t_L g4256 ( 
.A1(n_4208),
.A2(n_3711),
.B(n_3709),
.Y(n_4256)
);

NOR2x1p5_ASAP7_75t_L g4257 ( 
.A(n_4218),
.B(n_3692),
.Y(n_4257)
);

AOI211xp5_ASAP7_75t_L g4258 ( 
.A1(n_4212),
.A2(n_3692),
.B(n_669),
.C(n_666),
.Y(n_4258)
);

OAI21xp5_ASAP7_75t_L g4259 ( 
.A1(n_4234),
.A2(n_3711),
.B(n_3733),
.Y(n_4259)
);

AOI21xp5_ASAP7_75t_SL g4260 ( 
.A1(n_4236),
.A2(n_668),
.B(n_669),
.Y(n_4260)
);

OAI221xp5_ASAP7_75t_L g4261 ( 
.A1(n_4245),
.A2(n_3692),
.B1(n_3757),
.B2(n_3760),
.C(n_3764),
.Y(n_4261)
);

AOI221xp5_ASAP7_75t_SL g4262 ( 
.A1(n_4237),
.A2(n_3841),
.B1(n_3866),
.B2(n_671),
.C(n_673),
.Y(n_4262)
);

OAI221xp5_ASAP7_75t_L g4263 ( 
.A1(n_4239),
.A2(n_3841),
.B1(n_3750),
.B2(n_671),
.C(n_673),
.Y(n_4263)
);

XNOR2xp5_ASAP7_75t_L g4264 ( 
.A(n_4258),
.B(n_668),
.Y(n_4264)
);

AOI321xp33_ASAP7_75t_L g4265 ( 
.A1(n_4247),
.A2(n_3841),
.A3(n_3734),
.B1(n_3866),
.B2(n_3632),
.C(n_680),
.Y(n_4265)
);

OAI221xp5_ASAP7_75t_L g4266 ( 
.A1(n_4252),
.A2(n_3750),
.B1(n_674),
.B2(n_678),
.C(n_679),
.Y(n_4266)
);

NAND2xp5_ASAP7_75t_L g4267 ( 
.A(n_4232),
.B(n_670),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_4242),
.Y(n_4268)
);

XNOR2x1_ASAP7_75t_L g4269 ( 
.A(n_4243),
.B(n_681),
.Y(n_4269)
);

O2A1O1Ixp33_ASAP7_75t_L g4270 ( 
.A1(n_4235),
.A2(n_683),
.B(n_681),
.C(n_682),
.Y(n_4270)
);

XNOR2x1_ASAP7_75t_L g4271 ( 
.A(n_4257),
.B(n_682),
.Y(n_4271)
);

A2O1A1Ixp33_ASAP7_75t_L g4272 ( 
.A1(n_4246),
.A2(n_4253),
.B(n_4250),
.C(n_4241),
.Y(n_4272)
);

AOI221x1_ASAP7_75t_L g4273 ( 
.A1(n_4254),
.A2(n_4233),
.B1(n_4256),
.B2(n_4238),
.C(n_4255),
.Y(n_4273)
);

INVx1_ASAP7_75t_SL g4274 ( 
.A(n_4244),
.Y(n_4274)
);

NOR2xp33_ASAP7_75t_L g4275 ( 
.A(n_4251),
.B(n_683),
.Y(n_4275)
);

HB1xp67_ASAP7_75t_L g4276 ( 
.A(n_4240),
.Y(n_4276)
);

OAI211xp5_ASAP7_75t_L g4277 ( 
.A1(n_4249),
.A2(n_687),
.B(n_684),
.C(n_685),
.Y(n_4277)
);

AOI21xp33_ASAP7_75t_L g4278 ( 
.A1(n_4248),
.A2(n_684),
.B(n_685),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_4232),
.Y(n_4279)
);

O2A1O1Ixp33_ASAP7_75t_L g4280 ( 
.A1(n_4232),
.A2(n_689),
.B(n_687),
.C(n_688),
.Y(n_4280)
);

OAI322xp33_ASAP7_75t_SL g4281 ( 
.A1(n_4237),
.A2(n_3866),
.A3(n_3739),
.B1(n_3749),
.B2(n_3741),
.C1(n_3653),
.C2(n_3814),
.Y(n_4281)
);

NAND5xp2_ASAP7_75t_SL g4282 ( 
.A(n_4247),
.B(n_688),
.C(n_690),
.D(n_691),
.E(n_692),
.Y(n_4282)
);

AOI221xp5_ASAP7_75t_L g4283 ( 
.A1(n_4234),
.A2(n_3632),
.B1(n_3741),
.B2(n_3739),
.C(n_3749),
.Y(n_4283)
);

NAND4xp75_ASAP7_75t_L g4284 ( 
.A(n_4268),
.B(n_694),
.C(n_692),
.D(n_693),
.Y(n_4284)
);

AOI22xp5_ASAP7_75t_L g4285 ( 
.A1(n_4274),
.A2(n_3646),
.B1(n_3733),
.B2(n_3632),
.Y(n_4285)
);

AND2x2_ASAP7_75t_L g4286 ( 
.A(n_4279),
.B(n_693),
.Y(n_4286)
);

XNOR2xp5_ASAP7_75t_L g4287 ( 
.A(n_4264),
.B(n_694),
.Y(n_4287)
);

HB1xp67_ASAP7_75t_L g4288 ( 
.A(n_4271),
.Y(n_4288)
);

XOR2xp5_ASAP7_75t_L g4289 ( 
.A(n_4282),
.B(n_695),
.Y(n_4289)
);

NOR2x1_ASAP7_75t_L g4290 ( 
.A(n_4269),
.B(n_695),
.Y(n_4290)
);

NAND2xp5_ASAP7_75t_L g4291 ( 
.A(n_4275),
.B(n_696),
.Y(n_4291)
);

INVx2_ASAP7_75t_L g4292 ( 
.A(n_4267),
.Y(n_4292)
);

NAND4xp75_ASAP7_75t_L g4293 ( 
.A(n_4273),
.B(n_696),
.C(n_698),
.D(n_699),
.Y(n_4293)
);

NOR2xp67_ASAP7_75t_L g4294 ( 
.A(n_4277),
.B(n_698),
.Y(n_4294)
);

INVx2_ASAP7_75t_L g4295 ( 
.A(n_4260),
.Y(n_4295)
);

NAND2xp5_ASAP7_75t_L g4296 ( 
.A(n_4262),
.B(n_701),
.Y(n_4296)
);

NAND4xp75_ASAP7_75t_L g4297 ( 
.A(n_4262),
.B(n_701),
.C(n_702),
.D(n_704),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_4280),
.Y(n_4298)
);

AND2x2_ASAP7_75t_SL g4299 ( 
.A(n_4276),
.B(n_702),
.Y(n_4299)
);

AOI22xp5_ASAP7_75t_L g4300 ( 
.A1(n_4263),
.A2(n_3646),
.B1(n_3658),
.B2(n_3654),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_4270),
.Y(n_4301)
);

AND2x4_ASAP7_75t_L g4302 ( 
.A(n_4272),
.B(n_3695),
.Y(n_4302)
);

NAND2x1p5_ASAP7_75t_L g4303 ( 
.A(n_4266),
.B(n_705),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_4265),
.Y(n_4304)
);

NOR2xp67_ASAP7_75t_L g4305 ( 
.A(n_4261),
.B(n_705),
.Y(n_4305)
);

NAND4xp75_ASAP7_75t_L g4306 ( 
.A(n_4278),
.B(n_706),
.C(n_707),
.D(n_708),
.Y(n_4306)
);

INVx1_ASAP7_75t_L g4307 ( 
.A(n_4259),
.Y(n_4307)
);

INVxp67_ASAP7_75t_L g4308 ( 
.A(n_4283),
.Y(n_4308)
);

OR3x1_ASAP7_75t_L g4309 ( 
.A(n_4304),
.B(n_4281),
.C(n_706),
.Y(n_4309)
);

NAND3xp33_ASAP7_75t_L g4310 ( 
.A(n_4301),
.B(n_707),
.C(n_708),
.Y(n_4310)
);

NAND3xp33_ASAP7_75t_L g4311 ( 
.A(n_4301),
.B(n_709),
.C(n_710),
.Y(n_4311)
);

AND4x1_ASAP7_75t_L g4312 ( 
.A(n_4290),
.B(n_709),
.C(n_711),
.D(n_712),
.Y(n_4312)
);

NOR2xp67_ASAP7_75t_SL g4313 ( 
.A(n_4284),
.B(n_711),
.Y(n_4313)
);

NOR2x1p5_ASAP7_75t_L g4314 ( 
.A(n_4293),
.B(n_713),
.Y(n_4314)
);

NOR2x1_ASAP7_75t_L g4315 ( 
.A(n_4295),
.B(n_715),
.Y(n_4315)
);

OR4x1_ASAP7_75t_L g4316 ( 
.A(n_4298),
.B(n_715),
.C(n_717),
.D(n_718),
.Y(n_4316)
);

AOI221xp5_ASAP7_75t_L g4317 ( 
.A1(n_4289),
.A2(n_717),
.B1(n_718),
.B2(n_719),
.C(n_720),
.Y(n_4317)
);

AND4x1_ASAP7_75t_L g4318 ( 
.A(n_4286),
.B(n_719),
.C(n_720),
.D(n_721),
.Y(n_4318)
);

INVx2_ASAP7_75t_L g4319 ( 
.A(n_4302),
.Y(n_4319)
);

XOR2xp5_ASAP7_75t_L g4320 ( 
.A(n_4287),
.B(n_4297),
.Y(n_4320)
);

INVxp67_ASAP7_75t_L g4321 ( 
.A(n_4306),
.Y(n_4321)
);

NAND4xp25_ASAP7_75t_L g4322 ( 
.A(n_4294),
.B(n_721),
.C(n_722),
.D(n_723),
.Y(n_4322)
);

NOR3xp33_ASAP7_75t_SL g4323 ( 
.A(n_4291),
.B(n_722),
.C(n_723),
.Y(n_4323)
);

AND2x2_ASAP7_75t_L g4324 ( 
.A(n_4303),
.B(n_724),
.Y(n_4324)
);

OAI21xp5_ASAP7_75t_L g4325 ( 
.A1(n_4296),
.A2(n_3687),
.B(n_726),
.Y(n_4325)
);

NOR2x1p5_ASAP7_75t_L g4326 ( 
.A(n_4292),
.B(n_726),
.Y(n_4326)
);

NAND3xp33_ASAP7_75t_SL g4327 ( 
.A(n_4288),
.B(n_727),
.C(n_728),
.Y(n_4327)
);

NAND2xp5_ASAP7_75t_L g4328 ( 
.A(n_4305),
.B(n_729),
.Y(n_4328)
);

AND2x2_ASAP7_75t_L g4329 ( 
.A(n_4308),
.B(n_730),
.Y(n_4329)
);

OAI211xp5_ASAP7_75t_L g4330 ( 
.A1(n_4307),
.A2(n_730),
.B(n_731),
.C(n_733),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_4329),
.Y(n_4331)
);

INVx1_ASAP7_75t_L g4332 ( 
.A(n_4328),
.Y(n_4332)
);

NAND2xp5_ASAP7_75t_L g4333 ( 
.A(n_4319),
.B(n_4299),
.Y(n_4333)
);

AO221x1_ASAP7_75t_L g4334 ( 
.A1(n_4321),
.A2(n_4302),
.B1(n_4285),
.B2(n_4300),
.C(n_737),
.Y(n_4334)
);

AND2x4_ASAP7_75t_L g4335 ( 
.A(n_4324),
.B(n_733),
.Y(n_4335)
);

INVx2_ASAP7_75t_SL g4336 ( 
.A(n_4315),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_4310),
.Y(n_4337)
);

OAI211xp5_ASAP7_75t_SL g4338 ( 
.A1(n_4317),
.A2(n_734),
.B(n_736),
.C(n_737),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_4311),
.Y(n_4339)
);

INVx2_ASAP7_75t_L g4340 ( 
.A(n_4316),
.Y(n_4340)
);

OAI22xp5_ASAP7_75t_L g4341 ( 
.A1(n_4309),
.A2(n_4320),
.B1(n_4314),
.B2(n_4323),
.Y(n_4341)
);

INVx2_ASAP7_75t_L g4342 ( 
.A(n_4326),
.Y(n_4342)
);

NAND2xp5_ASAP7_75t_L g4343 ( 
.A(n_4313),
.B(n_736),
.Y(n_4343)
);

NAND2xp5_ASAP7_75t_L g4344 ( 
.A(n_4318),
.B(n_738),
.Y(n_4344)
);

INVx1_ASAP7_75t_L g4345 ( 
.A(n_4330),
.Y(n_4345)
);

NAND5xp2_ASAP7_75t_L g4346 ( 
.A(n_4325),
.B(n_4327),
.C(n_4312),
.D(n_4322),
.E(n_741),
.Y(n_4346)
);

AOI22xp33_ASAP7_75t_L g4347 ( 
.A1(n_4329),
.A2(n_3658),
.B1(n_3665),
.B2(n_3671),
.Y(n_4347)
);

NAND2xp5_ASAP7_75t_L g4348 ( 
.A(n_4329),
.B(n_738),
.Y(n_4348)
);

INVx1_ASAP7_75t_L g4349 ( 
.A(n_4348),
.Y(n_4349)
);

AOI31xp33_ASAP7_75t_L g4350 ( 
.A1(n_4340),
.A2(n_739),
.A3(n_740),
.B(n_741),
.Y(n_4350)
);

OAI22x1_ASAP7_75t_L g4351 ( 
.A1(n_4345),
.A2(n_3658),
.B1(n_3653),
.B2(n_3654),
.Y(n_4351)
);

INVx2_ASAP7_75t_L g4352 ( 
.A(n_4335),
.Y(n_4352)
);

OA22x2_ASAP7_75t_L g4353 ( 
.A1(n_4334),
.A2(n_4343),
.B1(n_4339),
.B2(n_4337),
.Y(n_4353)
);

OAI22x1_ASAP7_75t_L g4354 ( 
.A1(n_4335),
.A2(n_4331),
.B1(n_4336),
.B2(n_4344),
.Y(n_4354)
);

OAI22x1_ASAP7_75t_L g4355 ( 
.A1(n_4342),
.A2(n_3654),
.B1(n_742),
.B2(n_743),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_4333),
.Y(n_4356)
);

OAI22x1_ASAP7_75t_L g4357 ( 
.A1(n_4332),
.A2(n_739),
.B1(n_742),
.B2(n_743),
.Y(n_4357)
);

AO22x2_ASAP7_75t_L g4358 ( 
.A1(n_4341),
.A2(n_744),
.B1(n_745),
.B2(n_746),
.Y(n_4358)
);

AOI22xp5_ASAP7_75t_L g4359 ( 
.A1(n_4338),
.A2(n_3671),
.B1(n_3665),
.B2(n_3721),
.Y(n_4359)
);

OAI22xp5_ASAP7_75t_L g4360 ( 
.A1(n_4347),
.A2(n_3721),
.B1(n_3718),
.B2(n_3702),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_4346),
.Y(n_4361)
);

AOI22xp5_ASAP7_75t_L g4362 ( 
.A1(n_4345),
.A2(n_3718),
.B1(n_3672),
.B2(n_3702),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_4348),
.Y(n_4363)
);

AOI21xp5_ASAP7_75t_L g4364 ( 
.A1(n_4358),
.A2(n_744),
.B(n_748),
.Y(n_4364)
);

INVx1_ASAP7_75t_L g4365 ( 
.A(n_4358),
.Y(n_4365)
);

HB1xp67_ASAP7_75t_L g4366 ( 
.A(n_4357),
.Y(n_4366)
);

OAI22x1_ASAP7_75t_L g4367 ( 
.A1(n_4356),
.A2(n_748),
.B1(n_749),
.B2(n_751),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_4353),
.Y(n_4368)
);

OAI22x1_ASAP7_75t_L g4369 ( 
.A1(n_4361),
.A2(n_749),
.B1(n_751),
.B2(n_752),
.Y(n_4369)
);

HB1xp67_ASAP7_75t_L g4370 ( 
.A(n_4352),
.Y(n_4370)
);

INVx1_ASAP7_75t_L g4371 ( 
.A(n_4350),
.Y(n_4371)
);

OA21x2_ASAP7_75t_L g4372 ( 
.A1(n_4349),
.A2(n_752),
.B(n_753),
.Y(n_4372)
);

AO22x2_ASAP7_75t_L g4373 ( 
.A1(n_4363),
.A2(n_3697),
.B1(n_754),
.B2(n_755),
.Y(n_4373)
);

XOR2x1_ASAP7_75t_L g4374 ( 
.A(n_4354),
.B(n_753),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_4355),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4368),
.Y(n_4376)
);

HB1xp67_ASAP7_75t_L g4377 ( 
.A(n_4370),
.Y(n_4377)
);

BUFx2_ASAP7_75t_L g4378 ( 
.A(n_4372),
.Y(n_4378)
);

NAND3xp33_ASAP7_75t_L g4379 ( 
.A(n_4375),
.B(n_4362),
.C(n_4360),
.Y(n_4379)
);

BUFx2_ASAP7_75t_L g4380 ( 
.A(n_4366),
.Y(n_4380)
);

CKINVDCx20_ASAP7_75t_R g4381 ( 
.A(n_4371),
.Y(n_4381)
);

BUFx2_ASAP7_75t_L g4382 ( 
.A(n_4365),
.Y(n_4382)
);

AND3x1_ASAP7_75t_L g4383 ( 
.A(n_4364),
.B(n_4359),
.C(n_4351),
.Y(n_4383)
);

HB1xp67_ASAP7_75t_L g4384 ( 
.A(n_4369),
.Y(n_4384)
);

AOI22xp33_ASAP7_75t_R g4385 ( 
.A1(n_4377),
.A2(n_4374),
.B1(n_4367),
.B2(n_4373),
.Y(n_4385)
);

INVx1_ASAP7_75t_L g4386 ( 
.A(n_4376),
.Y(n_4386)
);

AND2x2_ASAP7_75t_L g4387 ( 
.A(n_4380),
.B(n_754),
.Y(n_4387)
);

OAI21xp5_ASAP7_75t_L g4388 ( 
.A1(n_4379),
.A2(n_755),
.B(n_756),
.Y(n_4388)
);

OAI22xp5_ASAP7_75t_L g4389 ( 
.A1(n_4381),
.A2(n_3697),
.B1(n_3672),
.B2(n_3704),
.Y(n_4389)
);

XOR2x2_ASAP7_75t_L g4390 ( 
.A(n_4383),
.B(n_756),
.Y(n_4390)
);

NAND2xp5_ASAP7_75t_L g4391 ( 
.A(n_4386),
.B(n_4378),
.Y(n_4391)
);

AOI21xp5_ASAP7_75t_L g4392 ( 
.A1(n_4388),
.A2(n_4384),
.B(n_4382),
.Y(n_4392)
);

OAI21x1_ASAP7_75t_SL g4393 ( 
.A1(n_4385),
.A2(n_3704),
.B(n_3701),
.Y(n_4393)
);

OAI21x1_ASAP7_75t_L g4394 ( 
.A1(n_4391),
.A2(n_4387),
.B(n_4390),
.Y(n_4394)
);

XNOR2xp5_ASAP7_75t_L g4395 ( 
.A(n_4392),
.B(n_4389),
.Y(n_4395)
);

AOI22xp5_ASAP7_75t_L g4396 ( 
.A1(n_4395),
.A2(n_4393),
.B1(n_3678),
.B2(n_3701),
.Y(n_4396)
);

OAI221xp5_ASAP7_75t_R g4397 ( 
.A1(n_4396),
.A2(n_4394),
.B1(n_759),
.B2(n_760),
.C(n_761),
.Y(n_4397)
);

AOI211xp5_ASAP7_75t_L g4398 ( 
.A1(n_4397),
.A2(n_758),
.B(n_760),
.C(n_761),
.Y(n_4398)
);


endmodule