module fake_jpeg_11968_n_474 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_474);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_474;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_9),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_0),
.B(n_16),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_3),
.B(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_16),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_5),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_57),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_58),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_59),
.B(n_90),
.Y(n_139)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_60),
.Y(n_167)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_61),
.Y(n_151)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_62),
.Y(n_172)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_64),
.Y(n_164)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_67),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_70),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_71),
.Y(n_169)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_35),
.Y(n_72)
);

INVx6_ASAP7_75t_SL g133 ( 
.A(n_72),
.Y(n_133)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx11_ASAP7_75t_L g162 ( 
.A(n_73),
.Y(n_162)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_75),
.Y(n_185)
);

BUFx10_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_76),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_14),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_107),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_79),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_80),
.Y(n_182)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_81),
.Y(n_163)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_82),
.Y(n_175)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_83),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

INVx4_ASAP7_75t_SL g85 ( 
.A(n_35),
.Y(n_85)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_46),
.B(n_14),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_86),
.B(n_104),
.Y(n_141)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_87),
.Y(n_190)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_89),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_14),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_92),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_93),
.Y(n_186)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_40),
.B(n_0),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_94),
.B(n_95),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_30),
.B(n_13),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_96),
.Y(n_177)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_97),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_99),
.Y(n_178)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_100),
.Y(n_181)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_101),
.Y(n_183)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_102),
.Y(n_184)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_103),
.B(n_105),
.Y(n_118)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_20),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_19),
.B(n_12),
.Y(n_105)
);

BUFx24_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_106),
.Y(n_179)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_22),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_112),
.Y(n_146)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_34),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_110),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_23),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_23),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_26),
.Y(n_153)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_28),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_42),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_115),
.Y(n_142)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_28),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_114),
.B(n_41),
.Y(n_170)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_34),
.Y(n_115)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_42),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_116),
.B(n_52),
.Y(n_132)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

BUFx16f_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_33),
.C(n_42),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_120),
.B(n_137),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_95),
.A2(n_51),
.B1(n_28),
.B2(n_53),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_122),
.B(n_129),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_91),
.A2(n_51),
.B1(n_53),
.B2(n_19),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_59),
.A2(n_51),
.B1(n_24),
.B2(n_39),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_131),
.A2(n_144),
.B1(n_161),
.B2(n_26),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_132),
.B(n_170),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_105),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_135),
.B(n_149),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_106),
.A2(n_52),
.B1(n_48),
.B2(n_47),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_136),
.A2(n_138),
.B(n_180),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_90),
.B(n_56),
.C(n_48),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_78),
.A2(n_47),
.B1(n_43),
.B2(n_56),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_110),
.A2(n_24),
.B1(n_49),
.B2(n_18),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_76),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_153),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_76),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_157),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_43),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_113),
.A2(n_71),
.B1(n_58),
.B2(n_67),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_159),
.A2(n_26),
.B1(n_2),
.B2(n_5),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_57),
.A2(n_49),
.B1(n_41),
.B2(n_39),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_98),
.B(n_37),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_173),
.B(n_176),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_92),
.B(n_37),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_85),
.A2(n_25),
.B(n_18),
.C(n_10),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_80),
.B(n_25),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_187),
.B(n_174),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_84),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_9),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_93),
.A2(n_26),
.B(n_9),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_189),
.Y(n_194)
);

AO22x1_ASAP7_75t_L g193 ( 
.A1(n_184),
.A2(n_75),
.B1(n_70),
.B2(n_4),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_193),
.A2(n_213),
.B(n_251),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_197),
.B(n_209),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_199),
.A2(n_207),
.B1(n_211),
.B2(n_216),
.Y(n_257)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_201),
.Y(n_253)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_202),
.Y(n_258)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_124),
.Y(n_203)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_203),
.Y(n_259)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_142),
.Y(n_204)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_204),
.Y(n_261)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_134),
.Y(n_205)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_205),
.Y(n_288)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_157),
.A2(n_153),
.B1(n_120),
.B2(n_180),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_206),
.A2(n_235),
.B1(n_236),
.B2(n_193),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_119),
.B(n_171),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_208),
.B(n_210),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_146),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_1),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_154),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_133),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_212),
.B(n_214),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_137),
.A2(n_2),
.B1(n_6),
.B2(n_8),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_136),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_127),
.Y(n_215)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_215),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_179),
.A2(n_8),
.B1(n_190),
.B2(n_163),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_138),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_217),
.B(n_220),
.Y(n_267)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_151),
.Y(n_219)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_219),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_164),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_159),
.A2(n_8),
.B1(n_118),
.B2(n_139),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_221),
.A2(n_222),
.B1(n_224),
.B2(n_238),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_143),
.A2(n_148),
.B1(n_169),
.B2(n_156),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_141),
.B(n_140),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_223),
.B(n_228),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_178),
.A2(n_156),
.B1(n_185),
.B2(n_148),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_177),
.Y(n_225)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_225),
.Y(n_263)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_125),
.Y(n_226)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_226),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_121),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_227),
.B(n_229),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_140),
.B(n_168),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_121),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_179),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_230),
.B(n_244),
.Y(n_290)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_167),
.Y(n_231)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_231),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_123),
.B(n_160),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_232),
.B(n_245),
.Y(n_293)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_177),
.Y(n_233)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_233),
.Y(n_299)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_125),
.Y(n_234)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_234),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_179),
.A2(n_190),
.B1(n_165),
.B2(n_163),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_165),
.A2(n_166),
.B1(n_186),
.B2(n_134),
.Y(n_236)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_182),
.Y(n_237)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_237),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_143),
.A2(n_185),
.B1(n_169),
.B2(n_147),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_147),
.A2(n_150),
.B1(n_128),
.B2(n_130),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_240),
.A2(n_229),
.B1(n_244),
.B2(n_200),
.Y(n_279)
);

AOI32xp33_ASAP7_75t_L g241 ( 
.A1(n_162),
.A2(n_158),
.A3(n_175),
.B1(n_128),
.B2(n_130),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_241),
.B(n_250),
.Y(n_286)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_182),
.Y(n_242)
);

BUFx2_ASAP7_75t_SL g260 ( 
.A(n_242),
.Y(n_260)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_167),
.Y(n_243)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_243),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_186),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_123),
.B(n_160),
.Y(n_245)
);

NAND2x1_ASAP7_75t_SL g246 ( 
.A(n_172),
.B(n_152),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_246),
.A2(n_196),
.B(n_227),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_247),
.B(n_252),
.Y(n_295)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_172),
.Y(n_248)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_248),
.Y(n_282)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_158),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_249),
.Y(n_278)
);

AOI32xp33_ASAP7_75t_L g250 ( 
.A1(n_162),
.A2(n_158),
.A3(n_126),
.B1(n_145),
.B2(n_152),
.Y(n_250)
);

BUFx10_ASAP7_75t_L g251 ( 
.A(n_174),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_251),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_126),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_214),
.A2(n_145),
.B(n_217),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_264),
.A2(n_297),
.B(n_279),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_207),
.A2(n_239),
.B1(n_204),
.B2(n_203),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_268),
.A2(n_271),
.B1(n_279),
.B2(n_281),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_239),
.A2(n_191),
.B1(n_194),
.B2(n_208),
.Y(n_271)
);

O2A1O1Ixp33_ASAP7_75t_SL g273 ( 
.A1(n_221),
.A2(n_191),
.B(n_199),
.C(n_250),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_273),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_276),
.A2(n_267),
.B(n_255),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_198),
.B(n_210),
.C(n_218),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_291),
.C(n_292),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_200),
.A2(n_192),
.B1(n_213),
.B2(n_198),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_294),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_284),
.A2(n_238),
.B1(n_226),
.B2(n_242),
.Y(n_309)
);

O2A1O1Ixp33_ASAP7_75t_L g289 ( 
.A1(n_218),
.A2(n_193),
.B(n_195),
.C(n_246),
.Y(n_289)
);

O2A1O1Ixp33_ASAP7_75t_L g327 ( 
.A1(n_289),
.A2(n_264),
.B(n_276),
.C(n_258),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_218),
.B(n_219),
.C(n_201),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_209),
.B(n_202),
.C(n_215),
.Y(n_292)
);

AND2x2_ASAP7_75t_SL g294 ( 
.A(n_246),
.B(n_231),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_220),
.B(n_252),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_251),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_248),
.B(n_240),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_249),
.C(n_224),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_212),
.B(n_243),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_298),
.B(n_237),
.Y(n_310)
);

NAND2x1_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_225),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_301),
.A2(n_320),
.B(n_303),
.Y(n_357)
);

INVx8_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_302),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_233),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_304),
.B(n_317),
.C(n_318),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_305),
.B(n_300),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_269),
.B(n_205),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_307),
.B(n_308),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_269),
.B(n_234),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_309),
.A2(n_326),
.B(n_278),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_310),
.B(n_311),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_251),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_266),
.Y(n_312)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_312),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_296),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_313),
.B(n_321),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_314),
.B(n_319),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_268),
.A2(n_272),
.B1(n_271),
.B2(n_286),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_315),
.A2(n_323),
.B1(n_332),
.B2(n_290),
.Y(n_336)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_253),
.Y(n_316)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_316),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_281),
.B(n_256),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_292),
.B(n_259),
.C(n_261),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_273),
.A2(n_259),
.B1(n_261),
.B2(n_286),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_254),
.B(n_295),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_293),
.B(n_285),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_322),
.B(n_328),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_272),
.A2(n_257),
.B1(n_273),
.B2(n_289),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_256),
.B(n_293),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_324),
.B(n_325),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_283),
.B(n_294),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_330),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_253),
.B(n_265),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_265),
.Y(n_329)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_329),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_258),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_287),
.A2(n_262),
.B1(n_280),
.B2(n_288),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_331),
.B(n_335),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_262),
.A2(n_282),
.B1(n_266),
.B2(n_274),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_282),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_333),
.Y(n_345)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_275),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_336),
.A2(n_346),
.B1(n_305),
.B2(n_313),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_304),
.B(n_275),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_337),
.B(n_359),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_338),
.B(n_354),
.Y(n_376)
);

AND2x6_ASAP7_75t_L g343 ( 
.A(n_315),
.B(n_278),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_343),
.B(n_356),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_323),
.A2(n_280),
.B1(n_288),
.B2(n_278),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_326),
.A2(n_270),
.B(n_274),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_347),
.A2(n_348),
.B(n_351),
.Y(n_382)
);

OA21x2_ASAP7_75t_L g348 ( 
.A1(n_334),
.A2(n_270),
.B(n_263),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_325),
.A2(n_263),
.B(n_299),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_327),
.A2(n_299),
.B(n_260),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_332),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_357),
.A2(n_360),
.B(n_301),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_320),
.A2(n_303),
.B(n_319),
.Y(n_360)
);

CKINVDCx12_ASAP7_75t_R g362 ( 
.A(n_318),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_362),
.Y(n_366)
);

INVx4_ASAP7_75t_SL g364 ( 
.A(n_302),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_364),
.Y(n_367)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_363),
.Y(n_365)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_365),
.Y(n_395)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_363),
.Y(n_368)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_368),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_369),
.A2(n_348),
.B1(n_346),
.B2(n_345),
.Y(n_406)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_350),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_370),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_339),
.A2(n_334),
.B1(n_306),
.B2(n_309),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_L g408 ( 
.A1(n_371),
.A2(n_372),
.B1(n_375),
.B2(n_385),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_339),
.A2(n_306),
.B1(n_360),
.B2(n_356),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_342),
.B(n_302),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_373),
.B(n_378),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_349),
.A2(n_324),
.B1(n_314),
.B2(n_310),
.Y(n_375)
);

OAI21xp33_ASAP7_75t_SL g377 ( 
.A1(n_348),
.A2(n_301),
.B(n_303),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_377),
.B(n_382),
.Y(n_409)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_350),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_358),
.B(n_316),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_379),
.B(n_381),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_355),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_380),
.B(n_388),
.Y(n_398)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_352),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_336),
.A2(n_317),
.B1(n_300),
.B2(n_330),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_384),
.A2(n_353),
.B1(n_354),
.B2(n_338),
.Y(n_402)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_352),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_358),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_386),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_387),
.A2(n_355),
.B(n_353),
.Y(n_404)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_341),
.Y(n_388)
);

OAI32xp33_ASAP7_75t_L g389 ( 
.A1(n_365),
.A2(n_361),
.A3(n_348),
.B1(n_343),
.B2(n_340),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_389),
.B(n_374),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_383),
.B(n_359),
.C(n_344),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_391),
.B(n_394),
.C(n_396),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_376),
.A2(n_355),
.B(n_357),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_392),
.B(n_393),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_373),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_383),
.B(n_344),
.C(n_337),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_384),
.B(n_366),
.C(n_387),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_372),
.B(n_361),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_397),
.B(n_404),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_369),
.B(n_347),
.C(n_351),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_401),
.B(n_405),
.C(n_379),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_402),
.B(n_382),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_371),
.B(n_368),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_406),
.A2(n_395),
.B1(n_399),
.B2(n_401),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_409),
.B(n_385),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_410),
.B(n_413),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_411),
.B(n_416),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_402),
.A2(n_376),
.B1(n_380),
.B2(n_367),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_408),
.A2(n_376),
.B1(n_378),
.B2(n_370),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_414),
.A2(n_406),
.B1(n_399),
.B2(n_400),
.Y(n_429)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_403),
.Y(n_415)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_415),
.Y(n_433)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_403),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_417),
.B(n_419),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_391),
.B(n_328),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_418),
.B(n_396),
.Y(n_428)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_398),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_400),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_420),
.B(n_425),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_423),
.B(n_424),
.C(n_394),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_395),
.A2(n_367),
.B1(n_381),
.B2(n_345),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_426),
.B(n_422),
.C(n_424),
.Y(n_442)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_428),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_429),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_414),
.A2(n_409),
.B1(n_404),
.B2(n_405),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_430),
.B(n_435),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_415),
.A2(n_407),
.B1(n_389),
.B2(n_397),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_412),
.B(n_392),
.C(n_407),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_436),
.B(n_390),
.C(n_341),
.Y(n_447)
);

INVx11_ASAP7_75t_L g437 ( 
.A(n_421),
.Y(n_437)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_437),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_413),
.A2(n_388),
.B(n_364),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_438),
.B(n_416),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_432),
.A2(n_411),
.B1(n_423),
.B2(n_412),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_440),
.B(n_442),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g456 ( 
.A(n_443),
.B(n_430),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_434),
.B(n_437),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_444),
.B(n_427),
.Y(n_451)
);

OAI21xp33_ASAP7_75t_L g445 ( 
.A1(n_432),
.A2(n_410),
.B(n_422),
.Y(n_445)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_445),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_447),
.B(n_431),
.C(n_426),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_439),
.A2(n_436),
.B(n_438),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_450),
.A2(n_456),
.B(n_443),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_451),
.B(n_453),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_441),
.B(n_431),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_452),
.B(n_455),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_446),
.A2(n_435),
.B1(n_429),
.B2(n_433),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_449),
.A2(n_433),
.B1(n_454),
.B2(n_456),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_458),
.B(n_455),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_453),
.B(n_441),
.Y(n_459)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_459),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_461),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_452),
.A2(n_447),
.B(n_448),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_462),
.B(n_364),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_465),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_466),
.Y(n_467)
);

OAI211xp5_ASAP7_75t_L g469 ( 
.A1(n_464),
.A2(n_460),
.B(n_457),
.C(n_445),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_469),
.B(n_329),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_468),
.B(n_463),
.C(n_331),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_470),
.A2(n_471),
.B(n_467),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_472),
.A2(n_335),
.B(n_333),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_473),
.B(n_312),
.Y(n_474)
);


endmodule