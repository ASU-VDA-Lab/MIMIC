module real_aes_5416_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_959, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_957, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_960, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_958, n_154, n_127, n_199, n_245, n_161, n_189, n_961, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_959;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_957;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_960;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_958;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_961;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_919;
wire n_857;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_260;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_889;
wire n_955;
wire n_696;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_932;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_925;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_261;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_954;
wire n_702;
wire n_296;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_915;
wire n_470;
wire n_851;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_928;
wire n_637;
wire n_899;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_922;
wire n_679;
wire n_926;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_949;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_911;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_500;
wire n_601;
wire n_307;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_259;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_0), .A2(n_510), .B(n_513), .Y(n_509) );
INVx1_ASAP7_75t_L g533 ( .A(n_1), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_2), .A2(n_5), .B1(n_406), .B2(n_553), .Y(n_552) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_3), .Y(n_662) );
AND2x4_ASAP7_75t_L g674 ( .A(n_3), .B(n_242), .Y(n_674) );
AND2x4_ASAP7_75t_L g679 ( .A(n_3), .B(n_680), .Y(n_679) );
AOI22xp33_ASAP7_75t_SL g709 ( .A1(n_4), .A2(n_46), .B1(n_702), .B2(n_703), .Y(n_709) );
INVx1_ASAP7_75t_L g938 ( .A(n_6), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_7), .A2(n_204), .B1(n_458), .B2(n_459), .Y(n_457) );
INVx1_ASAP7_75t_L g568 ( .A(n_8), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_9), .A2(n_218), .B1(n_443), .B2(n_456), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_10), .A2(n_94), .B1(n_913), .B2(n_934), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_11), .A2(n_104), .B1(n_671), .B2(n_675), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_12), .A2(n_22), .B1(n_453), .B2(n_459), .Y(n_627) );
INVx1_ASAP7_75t_L g329 ( .A(n_13), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_14), .A2(n_77), .B1(n_440), .B2(n_458), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_15), .A2(n_236), .B1(n_447), .B2(n_638), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_16), .A2(n_73), .B1(n_500), .B2(n_550), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g301 ( .A1(n_17), .A2(n_76), .B1(n_302), .B2(n_309), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_18), .A2(n_142), .B1(n_388), .B2(n_476), .Y(n_516) );
INVx1_ASAP7_75t_L g611 ( .A(n_19), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_20), .A2(n_107), .B1(n_606), .B2(n_908), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_21), .B(n_580), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_23), .A2(n_96), .B1(n_356), .B2(n_416), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_24), .A2(n_64), .B1(n_577), .B2(n_578), .Y(n_576) );
INVx1_ASAP7_75t_SL g362 ( .A(n_25), .Y(n_362) );
INVx1_ASAP7_75t_L g785 ( .A(n_26), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_27), .A2(n_157), .B1(n_580), .B2(n_581), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_28), .A2(n_93), .B1(n_698), .B2(n_700), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_29), .A2(n_153), .B1(n_282), .B2(n_547), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_30), .A2(n_75), .B1(n_406), .B2(n_599), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_31), .A2(n_247), .B1(n_356), .B2(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g279 ( .A(n_32), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_32), .B(n_182), .Y(n_336) );
INVxp67_ASAP7_75t_L g355 ( .A(n_32), .Y(n_355) );
AOI221xp5_ASAP7_75t_L g565 ( .A1(n_33), .A2(n_35), .B1(n_378), .B2(n_566), .C(n_567), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_34), .A2(n_203), .B1(n_643), .B2(n_644), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_36), .A2(n_141), .B1(n_452), .B2(n_453), .Y(n_451) );
CKINVDCx5p33_ASAP7_75t_R g892 ( .A(n_37), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_38), .A2(n_79), .B1(n_343), .B2(n_915), .Y(n_914) );
INVx1_ASAP7_75t_L g536 ( .A(n_39), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_40), .A2(n_170), .B1(n_702), .B2(n_703), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_41), .A2(n_44), .B1(n_409), .B2(n_411), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_42), .A2(n_229), .B1(n_691), .B2(n_694), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_43), .B(n_476), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_45), .A2(n_197), .B1(n_371), .B2(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_47), .B(n_264), .Y(n_274) );
INVx1_ASAP7_75t_L g524 ( .A(n_48), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_49), .A2(n_160), .B1(n_526), .B2(n_634), .Y(n_633) );
AOI21xp33_ASAP7_75t_L g422 ( .A1(n_50), .A2(n_341), .B(n_423), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_51), .A2(n_227), .B1(n_395), .B2(n_449), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_52), .A2(n_117), .B1(n_671), .B2(n_675), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_53), .A2(n_245), .B1(n_282), .B2(n_373), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_54), .A2(n_146), .B1(n_309), .B2(n_371), .Y(n_582) );
INVx2_ASAP7_75t_L g660 ( .A(n_55), .Y(n_660) );
INVx1_ASAP7_75t_L g673 ( .A(n_56), .Y(n_673) );
AND2x4_ASAP7_75t_L g676 ( .A(n_56), .B(n_660), .Y(n_676) );
INVx1_ASAP7_75t_SL g699 ( .A(n_56), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_57), .A2(n_172), .B1(n_416), .B2(n_421), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g258 ( .A1(n_58), .A2(n_177), .B1(n_259), .B2(n_282), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_59), .A2(n_235), .B1(n_413), .B2(n_545), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_60), .A2(n_120), .B1(n_461), .B2(n_462), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_61), .A2(n_185), .B1(n_369), .B2(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g530 ( .A(n_62), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g313 ( .A1(n_63), .A2(n_210), .B1(n_314), .B2(n_316), .Y(n_313) );
INVx1_ASAP7_75t_L g479 ( .A(n_65), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_66), .A2(n_206), .B1(n_368), .B2(n_369), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_67), .A2(n_187), .B1(n_297), .B2(n_366), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_68), .A2(n_119), .B1(n_282), .B2(n_368), .Y(n_583) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_69), .Y(n_264) );
INVx1_ASAP7_75t_L g517 ( .A(n_70), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_71), .A2(n_154), .B1(n_702), .B2(n_703), .Y(n_712) );
INVx1_ASAP7_75t_L g688 ( .A(n_72), .Y(n_688) );
XOR2x2_ASAP7_75t_L g630 ( .A(n_74), .B(n_631), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_78), .A2(n_243), .B1(n_698), .B2(n_700), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g340 ( .A1(n_80), .A2(n_166), .B1(n_341), .B2(n_343), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_81), .A2(n_189), .B1(n_461), .B2(n_462), .Y(n_460) );
INVx1_ASAP7_75t_L g265 ( .A(n_82), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_82), .B(n_181), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_83), .A2(n_224), .B1(n_394), .B2(n_395), .Y(n_393) );
AOI33xp33_ASAP7_75t_R g649 ( .A1(n_84), .A2(n_212), .A3(n_261), .B1(n_285), .B2(n_650), .B3(n_959), .Y(n_649) );
INVx1_ASAP7_75t_L g527 ( .A(n_85), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_86), .A2(n_90), .B1(n_698), .B2(n_700), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g947 ( .A1(n_87), .A2(n_208), .B1(n_948), .B2(n_949), .Y(n_947) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_88), .A2(n_173), .B1(n_302), .B2(n_404), .Y(n_602) );
AOI21xp5_ASAP7_75t_SL g323 ( .A1(n_89), .A2(n_324), .B(n_328), .Y(n_323) );
INVx1_ASAP7_75t_L g563 ( .A(n_90), .Y(n_563) );
OAI222xp33_ASAP7_75t_L g574 ( .A1(n_90), .A2(n_575), .B1(n_582), .B2(n_583), .C1(n_957), .C2(n_958), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_90), .B(n_583), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_91), .A2(n_222), .B1(n_302), .B2(n_646), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_92), .A2(n_99), .B1(n_443), .B2(n_444), .Y(n_442) );
INVx1_ASAP7_75t_L g436 ( .A(n_93), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g358 ( .A(n_95), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_97), .A2(n_180), .B1(n_455), .B2(n_456), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_98), .A2(n_237), .B1(n_316), .B2(n_368), .Y(n_502) );
INVx1_ASAP7_75t_L g400 ( .A(n_100), .Y(n_400) );
INVx1_ASAP7_75t_L g384 ( .A(n_101), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_102), .A2(n_192), .B1(n_413), .B2(n_545), .Y(n_603) );
AOI21xp33_ASAP7_75t_L g609 ( .A1(n_103), .A2(n_449), .B(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g482 ( .A(n_105), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_106), .A2(n_195), .B1(n_371), .B2(n_404), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_108), .A2(n_136), .B1(n_297), .B2(n_406), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_109), .A2(n_131), .B1(n_373), .B2(n_411), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_110), .A2(n_221), .B1(n_259), .B2(n_282), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_111), .A2(n_188), .B1(n_694), .B2(n_702), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_112), .A2(n_144), .B1(n_440), .B2(n_441), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g904 ( .A(n_113), .Y(n_904) );
AOI22x1_ASAP7_75t_L g466 ( .A1(n_114), .A2(n_467), .B1(n_468), .B2(n_491), .Y(n_466) );
INVx1_ASAP7_75t_L g491 ( .A(n_114), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_115), .A2(n_214), .B1(n_297), .B2(n_366), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_116), .A2(n_184), .B1(n_347), .B2(n_421), .Y(n_420) );
INVxp33_ASAP7_75t_SL g695 ( .A(n_118), .Y(n_695) );
AO22x1_ASAP7_75t_L g573 ( .A1(n_121), .A2(n_122), .B1(n_366), .B2(n_373), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_123), .A2(n_130), .B1(n_901), .B2(n_902), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_124), .A2(n_129), .B1(n_309), .B2(n_371), .Y(n_370) );
OAI22xp5_ASAP7_75t_L g927 ( .A1(n_125), .A2(n_928), .B1(n_929), .B2(n_953), .Y(n_927) );
CKINVDCx20_ASAP7_75t_R g928 ( .A(n_125), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_126), .A2(n_159), .B1(n_678), .B2(n_681), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_127), .B(n_580), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_128), .A2(n_133), .B1(n_888), .B2(n_889), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_132), .A2(n_143), .B1(n_888), .B2(n_889), .Y(n_887) );
INVx1_ASAP7_75t_L g514 ( .A(n_134), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_135), .A2(n_320), .B(n_472), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_137), .A2(n_156), .B1(n_547), .B2(n_601), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_138), .A2(n_246), .B1(n_911), .B2(n_913), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_139), .A2(n_230), .B1(n_452), .B2(n_455), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_140), .A2(n_213), .B1(n_944), .B2(n_946), .Y(n_943) );
XOR2xp5_ASAP7_75t_L g616 ( .A(n_145), .B(n_617), .Y(n_616) );
XOR2xp5_ASAP7_75t_L g653 ( .A(n_145), .B(n_617), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_147), .A2(n_244), .B1(n_293), .B2(n_297), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g895 ( .A(n_148), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_149), .B(n_485), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_150), .A2(n_176), .B1(n_314), .B2(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g692 ( .A(n_151), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_152), .B(n_941), .Y(n_940) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_155), .A2(n_196), .B1(n_441), .B2(n_540), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_158), .A2(n_161), .B1(n_441), .B2(n_444), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_162), .A2(n_186), .B1(n_356), .B2(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_163), .B(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_164), .B(n_447), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_165), .A2(n_248), .B1(n_373), .B2(n_505), .Y(n_504) );
OA22x2_ASAP7_75t_L g269 ( .A1(n_167), .A2(n_182), .B1(n_264), .B2(n_268), .Y(n_269) );
INVx1_ASAP7_75t_L g289 ( .A(n_167), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_168), .A2(n_219), .B1(n_282), .B2(n_373), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_169), .A2(n_233), .B1(n_446), .B2(n_447), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_171), .A2(n_239), .B1(n_678), .B2(n_681), .Y(n_725) );
AO22x2_ASAP7_75t_L g518 ( .A1(n_174), .A2(n_519), .B1(n_520), .B2(n_521), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_174), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_175), .A2(n_191), .B1(n_368), .B2(n_369), .Y(n_367) );
INVx1_ASAP7_75t_L g386 ( .A(n_178), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_179), .A2(n_223), .B1(n_343), .B2(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g281 ( .A(n_181), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_181), .B(n_287), .Y(n_339) );
OAI21xp33_ASAP7_75t_L g290 ( .A1(n_182), .A2(n_200), .B(n_291), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_183), .A2(n_199), .B1(n_297), .B2(n_406), .Y(n_487) );
INVx1_ASAP7_75t_L g595 ( .A(n_190), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_190), .A2(n_207), .B1(n_698), .B2(n_700), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_193), .B(n_532), .Y(n_619) );
INVx1_ASAP7_75t_L g784 ( .A(n_194), .Y(n_784) );
INVx1_ASAP7_75t_L g376 ( .A(n_198), .Y(n_376) );
INVx1_ASAP7_75t_L g267 ( .A(n_200), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_200), .B(n_234), .Y(n_337) );
INVx1_ASAP7_75t_L g379 ( .A(n_201), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_202), .B(n_449), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_205), .A2(n_228), .B1(n_545), .B2(n_648), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g935 ( .A1(n_209), .A2(n_936), .B(n_937), .Y(n_935) );
INVx1_ASAP7_75t_L g390 ( .A(n_211), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_215), .A2(n_231), .B1(n_302), .B2(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_216), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g480 ( .A(n_217), .Y(n_480) );
INVx1_ASAP7_75t_L g473 ( .A(n_220), .Y(n_473) );
INVx1_ASAP7_75t_L g424 ( .A(n_225), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_226), .A2(n_238), .B1(n_378), .B2(n_508), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g916 ( .A(n_229), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_229), .A2(n_925), .B1(n_927), .B2(n_954), .Y(n_924) );
AOI22x1_ASAP7_75t_L g346 ( .A1(n_232), .A2(n_241), .B1(n_347), .B2(n_356), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_234), .B(n_273), .Y(n_272) );
INVxp33_ASAP7_75t_L g686 ( .A(n_240), .Y(n_686) );
INVx1_ASAP7_75t_L g680 ( .A(n_242), .Y(n_680) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_557), .B(n_654), .C(n_663), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g654 ( .A1(n_250), .A2(n_557), .B(n_655), .Y(n_654) );
XNOR2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_429), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_397), .B1(n_427), .B2(n_428), .Y(n_251) );
INVx1_ASAP7_75t_L g427 ( .A(n_252), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_359), .B1(n_360), .B2(n_396), .Y(n_252) );
INVx1_ASAP7_75t_L g396 ( .A(n_253), .Y(n_396) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
XNOR2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_358), .Y(n_255) );
NOR3xp33_ASAP7_75t_SL g256 ( .A(n_257), .B(n_300), .C(n_318), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_292), .Y(n_257) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
BUFx8_ASAP7_75t_L g373 ( .A(n_260), .Y(n_373) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_270), .Y(n_260) );
AND2x4_ASAP7_75t_L g294 ( .A(n_261), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g322 ( .A(n_261), .B(n_311), .Y(n_322) );
AND2x2_ASAP7_75t_L g357 ( .A(n_261), .B(n_307), .Y(n_357) );
AND2x2_ASAP7_75t_L g410 ( .A(n_261), .B(n_270), .Y(n_410) );
AND2x4_ASAP7_75t_L g443 ( .A(n_261), .B(n_307), .Y(n_443) );
AND2x2_ASAP7_75t_L g449 ( .A(n_261), .B(n_311), .Y(n_449) );
AND2x4_ASAP7_75t_L g452 ( .A(n_261), .B(n_299), .Y(n_452) );
AND2x4_ASAP7_75t_L g458 ( .A(n_261), .B(n_270), .Y(n_458) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_269), .Y(n_261) );
INVx1_ASAP7_75t_L g305 ( .A(n_262), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_266), .Y(n_262) );
NAND2xp33_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx2_ASAP7_75t_L g268 ( .A(n_264), .Y(n_268) );
INVx3_ASAP7_75t_L g273 ( .A(n_264), .Y(n_273) );
NAND2xp33_ASAP7_75t_L g280 ( .A(n_264), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g291 ( .A(n_264), .Y(n_291) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_264), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_265), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
OAI21xp5_ASAP7_75t_L g354 ( .A1(n_267), .A2(n_291), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g306 ( .A(n_269), .Y(n_306) );
AND2x2_ASAP7_75t_L g327 ( .A(n_269), .B(n_305), .Y(n_327) );
AND2x2_ASAP7_75t_L g353 ( .A(n_269), .B(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g284 ( .A(n_270), .B(n_285), .Y(n_284) );
AND2x4_ASAP7_75t_L g315 ( .A(n_270), .B(n_304), .Y(n_315) );
AND2x4_ASAP7_75t_L g455 ( .A(n_270), .B(n_304), .Y(n_455) );
AND2x4_ASAP7_75t_L g459 ( .A(n_270), .B(n_285), .Y(n_459) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_270), .Y(n_650) );
AND2x4_ASAP7_75t_L g270 ( .A(n_271), .B(n_275), .Y(n_270) );
OR2x2_ASAP7_75t_L g296 ( .A(n_271), .B(n_276), .Y(n_296) );
AND2x4_ASAP7_75t_L g307 ( .A(n_271), .B(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g312 ( .A(n_271), .Y(n_312) );
AND2x2_ASAP7_75t_L g350 ( .A(n_271), .B(n_351), .Y(n_350) );
AND2x4_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_273), .B(n_279), .Y(n_278) );
INVxp67_ASAP7_75t_L g287 ( .A(n_273), .Y(n_287) );
NAND3xp33_ASAP7_75t_L g338 ( .A(n_274), .B(n_286), .C(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g308 ( .A(n_277), .Y(n_308) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
INVx4_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx4_ASAP7_75t_L g411 ( .A(n_283), .Y(n_411) );
INVx4_ASAP7_75t_L g505 ( .A(n_283), .Y(n_505) );
INVx2_ASAP7_75t_SL g601 ( .A(n_283), .Y(n_601) );
INVx8_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g298 ( .A(n_285), .B(n_299), .Y(n_298) );
AND2x4_ASAP7_75t_L g345 ( .A(n_285), .B(n_311), .Y(n_345) );
AND2x4_ASAP7_75t_L g444 ( .A(n_285), .B(n_311), .Y(n_444) );
AND2x4_ASAP7_75t_L g453 ( .A(n_285), .B(n_299), .Y(n_453) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_290), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
BUFx12f_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_294), .Y(n_366) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_294), .Y(n_406) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_294), .Y(n_644) );
BUFx3_ASAP7_75t_L g948 ( .A(n_294), .Y(n_948) );
AND2x4_ASAP7_75t_L g456 ( .A(n_295), .B(n_304), .Y(n_456) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g299 ( .A(n_296), .Y(n_299) );
BUFx12f_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx6_ASAP7_75t_L g554 ( .A(n_298), .Y(n_554) );
AND2x4_ASAP7_75t_L g317 ( .A(n_299), .B(n_304), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_313), .Y(n_300) );
BUFx12f_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_303), .Y(n_371) );
INVx3_ASAP7_75t_L g551 ( .A(n_303), .Y(n_551) );
AND2x4_ASAP7_75t_L g303 ( .A(n_304), .B(n_307), .Y(n_303) );
AND2x2_ASAP7_75t_L g310 ( .A(n_304), .B(n_311), .Y(n_310) );
AND2x4_ASAP7_75t_L g461 ( .A(n_304), .B(n_307), .Y(n_461) );
AND2x4_ASAP7_75t_L g462 ( .A(n_304), .B(n_311), .Y(n_462) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
AND2x4_ASAP7_75t_L g326 ( .A(n_307), .B(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g440 ( .A(n_307), .B(n_327), .Y(n_440) );
AND2x4_ASAP7_75t_L g311 ( .A(n_308), .B(n_312), .Y(n_311) );
BUFx5_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_310), .Y(n_404) );
INVx1_ASAP7_75t_L g501 ( .A(n_310), .Y(n_501) );
BUFx3_ASAP7_75t_L g646 ( .A(n_310), .Y(n_646) );
AND2x4_ASAP7_75t_L g342 ( .A(n_311), .B(n_327), .Y(n_342) );
AND2x2_ASAP7_75t_L g446 ( .A(n_311), .B(n_327), .Y(n_446) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx6f_ASAP7_75t_L g368 ( .A(n_315), .Y(n_368) );
BUFx12f_ASAP7_75t_L g545 ( .A(n_315), .Y(n_545) );
HB1xp67_ASAP7_75t_L g894 ( .A(n_316), .Y(n_894) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_317), .Y(n_369) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_317), .Y(n_413) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_317), .Y(n_648) );
NAND4xp25_ASAP7_75t_L g318 ( .A(n_319), .B(n_323), .C(n_340), .D(n_346), .Y(n_318) );
INVx3_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g392 ( .A(n_321), .Y(n_392) );
INVx2_ASAP7_75t_L g418 ( .A(n_321), .Y(n_418) );
INVx2_ASAP7_75t_L g512 ( .A(n_321), .Y(n_512) );
INVx3_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx3_ASAP7_75t_L g538 ( .A(n_322), .Y(n_538) );
INVx2_ASAP7_75t_L g639 ( .A(n_322), .Y(n_639) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_326), .Y(n_378) );
BUFx3_ASAP7_75t_L g421 ( .A(n_326), .Y(n_421) );
BUFx3_ASAP7_75t_L g526 ( .A(n_326), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_330), .B(n_611), .Y(n_610) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_SL g395 ( .A(n_331), .Y(n_395) );
INVx2_ASAP7_75t_L g447 ( .A(n_331), .Y(n_447) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_331), .Y(n_541) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx3_ASAP7_75t_L g426 ( .A(n_332), .Y(n_426) );
AO21x2_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_335), .B(n_338), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_334), .B(n_352), .Y(n_351) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_335), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
BUFx6f_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g385 ( .A(n_342), .Y(n_385) );
INVx2_ASAP7_75t_L g477 ( .A(n_342), .Y(n_477) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_342), .Y(n_532) );
BUFx3_ASAP7_75t_L g580 ( .A(n_342), .Y(n_580) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx3_ASAP7_75t_L g388 ( .A(n_344), .Y(n_388) );
INVx2_ASAP7_75t_L g634 ( .A(n_344), .Y(n_634) );
INVx3_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_345), .Y(n_416) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_345), .Y(n_581) );
INVx4_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g394 ( .A(n_348), .Y(n_394) );
INVx3_ASAP7_75t_L g485 ( .A(n_348), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g513 ( .A1(n_348), .A2(n_514), .B(n_515), .Y(n_513) );
INVx2_ASAP7_75t_L g578 ( .A(n_348), .Y(n_578) );
INVx5_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx4f_ASAP7_75t_L g606 ( .A(n_349), .Y(n_606) );
BUFx2_ASAP7_75t_L g636 ( .A(n_349), .Y(n_636) );
AND2x4_ASAP7_75t_L g349 ( .A(n_350), .B(n_353), .Y(n_349) );
AND2x2_ASAP7_75t_L g441 ( .A(n_350), .B(n_353), .Y(n_441) );
INVx3_ASAP7_75t_L g528 ( .A(n_356), .Y(n_528) );
BUFx3_ASAP7_75t_L g913 ( .A(n_356), .Y(n_913) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g382 ( .A(n_357), .Y(n_382) );
BUFx3_ASAP7_75t_L g577 ( .A(n_357), .Y(n_577) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
XNOR2x1_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_374), .Y(n_363) );
AND4x1_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .C(n_370), .D(n_372), .Y(n_364) );
NOR3xp33_ASAP7_75t_L g374 ( .A(n_375), .B(n_383), .C(n_389), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_377), .B1(n_379), .B2(n_380), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_377), .A2(n_387), .B1(n_479), .B2(n_480), .Y(n_478) );
INVx4_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_382), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B1(n_386), .B2(n_387), .Y(n_383) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI21xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B(n_393), .Y(n_389) );
INVx1_ASAP7_75t_L g936 ( .A(n_391), .Y(n_936) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g428 ( .A(n_397), .Y(n_428) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx3_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
XNOR2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
NOR4xp75_ASAP7_75t_L g401 ( .A(n_402), .B(n_407), .C(n_414), .D(n_419), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_405), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_408), .B(n_412), .Y(n_407) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx4f_ASAP7_75t_L g547 ( .A(n_410), .Y(n_547) );
BUFx3_ASAP7_75t_L g946 ( .A(n_413), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_417), .Y(n_414) );
INVx3_ASAP7_75t_L g534 ( .A(n_416), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_420), .B(n_422), .Y(n_419) );
INVx2_ASAP7_75t_L g912 ( .A(n_421), .Y(n_912) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_425), .B(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g908 ( .A(n_425), .Y(n_908) );
INVx1_ASAP7_75t_L g941 ( .A(n_425), .Y(n_941) );
INVx4_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_431), .B1(n_492), .B2(n_493), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B1(n_463), .B2(n_464), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
XNOR2x1_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
OR2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_450), .Y(n_437) );
NAND4xp25_ASAP7_75t_L g438 ( .A(n_439), .B(n_442), .C(n_445), .D(n_448), .Y(n_438) );
INVx3_ASAP7_75t_L g474 ( .A(n_447), .Y(n_474) );
NAND4xp25_ASAP7_75t_L g450 ( .A(n_451), .B(n_454), .C(n_457), .D(n_460), .Y(n_450) );
INVx2_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_486), .Y(n_468) );
NOR3xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_478), .C(n_481), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_471), .B(n_475), .Y(n_470) );
NOR2xp33_ASAP7_75t_SL g472 ( .A(n_473), .B(n_474), .Y(n_472) );
INVx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g915 ( .A(n_477), .Y(n_915) );
OAI21xp33_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .B(n_484), .Y(n_481) );
INVx2_ASAP7_75t_L g508 ( .A(n_483), .Y(n_508) );
AND4x1_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .C(n_489), .D(n_490), .Y(n_486) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx2_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
AO22x2_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_518), .B1(n_555), .B2(n_556), .Y(n_494) );
INVx1_ASAP7_75t_L g555 ( .A(n_495), .Y(n_555) );
XOR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_517), .Y(n_495) );
NOR2x1_ASAP7_75t_L g496 ( .A(n_497), .B(n_506), .Y(n_496) );
NAND4xp25_ASAP7_75t_L g497 ( .A(n_498), .B(n_502), .C(n_503), .D(n_504), .Y(n_497) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NAND3xp33_ASAP7_75t_L g506 ( .A(n_507), .B(n_509), .C(n_516), .Y(n_506) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g556 ( .A(n_518), .Y(n_556) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_542), .Y(n_521) );
NOR3xp33_ASAP7_75t_SL g522 ( .A(n_523), .B(n_529), .C(n_535), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B1(n_527), .B2(n_528), .Y(n_523) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx2_ASAP7_75t_L g934 ( .A(n_526), .Y(n_934) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B1(n_533), .B2(n_534), .Y(n_529) );
INVx1_ASAP7_75t_L g932 ( .A(n_531), .Y(n_932) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
OAI21xp33_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_537), .B(n_539), .Y(n_535) );
INVx2_ASAP7_75t_L g566 ( .A(n_537), .Y(n_566) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx3_ASAP7_75t_L g906 ( .A(n_538), .Y(n_906) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_548), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_546), .Y(n_543) );
BUFx6f_ASAP7_75t_L g897 ( .A(n_545), .Y(n_897) );
INVx1_ASAP7_75t_L g945 ( .A(n_545), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_552), .Y(n_548) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g888 ( .A(n_551), .Y(n_888) );
INVx3_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g572 ( .A(n_554), .Y(n_572) );
INVx2_ASAP7_75t_L g599 ( .A(n_554), .Y(n_599) );
INVx5_ASAP7_75t_L g643 ( .A(n_554), .Y(n_643) );
INVx2_ASAP7_75t_L g950 ( .A(n_554), .Y(n_950) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .B1(n_613), .B2(n_614), .Y(n_557) );
INVx2_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
OA22x2_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B1(n_591), .B2(n_612), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x4_ASAP7_75t_L g561 ( .A(n_562), .B(n_584), .Y(n_561) );
AOI21x1_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_564), .B(n_574), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_569), .Y(n_564) );
BUFx2_ASAP7_75t_L g585 ( .A(n_565), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_573), .Y(n_569) );
INVxp67_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g589 ( .A(n_571), .B(n_582), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_573), .Y(n_590) );
INVx1_ASAP7_75t_L g588 ( .A(n_575), .Y(n_588) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_579), .Y(n_575) );
NAND4xp75_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .C(n_589), .D(n_590), .Y(n_584) );
NOR2x1_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g612 ( .A(n_591), .Y(n_612) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
BUFx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
XNOR2x1_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g594 ( .A(n_595), .Y(n_594) );
NOR2x1_ASAP7_75t_L g596 ( .A(n_597), .B(n_604), .Y(n_596) );
NAND4xp25_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .C(n_602), .D(n_603), .Y(n_597) );
HB1xp67_ASAP7_75t_L g902 ( .A(n_599), .Y(n_902) );
NAND4xp25_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .C(n_608), .D(n_609), .Y(n_604) );
INVx2_ASAP7_75t_SL g939 ( .A(n_606), .Y(n_939) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AO22x1_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_628), .B1(n_629), .B2(n_651), .Y(n_614) );
INVxp67_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OR2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_623), .Y(n_617) );
NAND4xp25_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .C(n_621), .D(n_622), .Y(n_618) );
NAND4xp25_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .C(n_626), .D(n_627), .Y(n_623) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NOR2x1_ASAP7_75t_L g631 ( .A(n_632), .B(n_641), .Y(n_631) );
NAND4xp25_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .C(n_637), .D(n_640), .Y(n_632) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND4xp25_ASAP7_75t_L g641 ( .A(n_642), .B(n_645), .C(n_647), .D(n_649), .Y(n_641) );
BUFx3_ASAP7_75t_L g901 ( .A(n_644), .Y(n_901) );
BUFx2_ASAP7_75t_L g889 ( .A(n_646), .Y(n_889) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
BUFx3_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NAND3xp33_ASAP7_75t_L g657 ( .A(n_658), .B(n_661), .C(n_662), .Y(n_657) );
AND2x2_ASAP7_75t_L g921 ( .A(n_658), .B(n_922), .Y(n_921) );
AND2x2_ASAP7_75t_L g926 ( .A(n_658), .B(n_923), .Y(n_926) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OA21x2_ASAP7_75t_L g954 ( .A1(n_659), .A2(n_699), .B(n_955), .Y(n_954) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g672 ( .A(n_660), .B(n_673), .Y(n_672) );
AND3x4_ASAP7_75t_L g698 ( .A(n_660), .B(n_679), .C(n_699), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g922 ( .A(n_661), .B(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_662), .Y(n_923) );
OAI221xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_881), .B1(n_883), .B2(n_919), .C(n_924), .Y(n_663) );
AOI211x1_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_781), .B(n_787), .C(n_862), .Y(n_664) );
NAND5xp2_ASAP7_75t_L g665 ( .A(n_666), .B(n_739), .C(n_757), .D(n_767), .E(n_772), .Y(n_665) );
AOI332xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_704), .A3(n_714), .B1(n_715), .B2(n_719), .B3(n_728), .C1(n_729), .C2(n_733), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_668), .B(n_682), .Y(n_667) );
INVx2_ASAP7_75t_L g727 ( .A(n_668), .Y(n_727) );
BUFx3_ASAP7_75t_L g800 ( .A(n_668), .Y(n_800) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_668), .B(n_723), .Y(n_807) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g737 ( .A(n_669), .Y(n_737) );
OR2x2_ASAP7_75t_L g834 ( .A(n_669), .B(n_696), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_677), .Y(n_669) );
AND2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_674), .Y(n_671) );
AND2x4_ASAP7_75t_L g678 ( .A(n_672), .B(n_679), .Y(n_678) );
AND2x4_ASAP7_75t_L g691 ( .A(n_672), .B(n_674), .Y(n_691) );
AND2x2_ASAP7_75t_L g702 ( .A(n_672), .B(n_674), .Y(n_702) );
AND2x2_ASAP7_75t_L g675 ( .A(n_674), .B(n_676), .Y(n_675) );
AND2x4_ASAP7_75t_L g694 ( .A(n_674), .B(n_676), .Y(n_694) );
AND2x2_ASAP7_75t_L g703 ( .A(n_674), .B(n_676), .Y(n_703) );
CKINVDCx5p33_ASAP7_75t_R g955 ( .A(n_674), .Y(n_955) );
AND2x4_ASAP7_75t_L g681 ( .A(n_676), .B(n_679), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_676), .B(n_679), .Y(n_687) );
AND2x4_ASAP7_75t_L g700 ( .A(n_676), .B(n_679), .Y(n_700) );
INVx3_ASAP7_75t_L g685 ( .A(n_678), .Y(n_685) );
INVx1_ASAP7_75t_L g797 ( .A(n_682), .Y(n_797) );
NOR2xp33_ASAP7_75t_L g846 ( .A(n_682), .B(n_847), .Y(n_846) );
OR2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_696), .Y(n_682) );
INVx1_ASAP7_75t_L g722 ( .A(n_683), .Y(n_722) );
INVx2_ASAP7_75t_L g760 ( .A(n_683), .Y(n_760) );
AND2x2_ASAP7_75t_L g768 ( .A(n_683), .B(n_769), .Y(n_768) );
AND2x2_ASAP7_75t_L g776 ( .A(n_683), .B(n_696), .Y(n_776) );
AND2x2_ASAP7_75t_L g779 ( .A(n_683), .B(n_723), .Y(n_779) );
AND2x2_ASAP7_75t_L g829 ( .A(n_683), .B(n_724), .Y(n_829) );
OR2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_689), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_686), .B1(n_687), .B2(n_688), .Y(n_684) );
OAI221xp5_ASAP7_75t_L g783 ( .A1(n_685), .A2(n_687), .B1(n_784), .B2(n_785), .C(n_786), .Y(n_783) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_692), .B1(n_693), .B2(n_695), .Y(n_689) );
INVx3_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
BUFx2_ASAP7_75t_L g882 ( .A(n_694), .Y(n_882) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_696), .Y(n_728) );
INVx2_ASAP7_75t_L g747 ( .A(n_696), .Y(n_747) );
OR2x2_ASAP7_75t_L g756 ( .A(n_696), .B(n_737), .Y(n_756) );
AND2x2_ASAP7_75t_L g769 ( .A(n_696), .B(n_737), .Y(n_769) );
AND2x2_ASAP7_75t_L g789 ( .A(n_696), .B(n_736), .Y(n_789) );
OR2x2_ASAP7_75t_L g818 ( .A(n_696), .B(n_760), .Y(n_818) );
AND2x2_ASAP7_75t_L g852 ( .A(n_696), .B(n_760), .Y(n_852) );
AND2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_701), .Y(n_696) );
INVxp67_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_713), .Y(n_705) );
INVx1_ASAP7_75t_L g732 ( .A(n_706), .Y(n_732) );
OR2x2_ASAP7_75t_L g766 ( .A(n_706), .B(n_716), .Y(n_766) );
OAI32xp33_ASAP7_75t_L g871 ( .A1(n_706), .A2(n_771), .A3(n_788), .B1(n_847), .B2(n_867), .Y(n_871) );
NOR2xp33_ASAP7_75t_L g880 ( .A(n_706), .B(n_764), .Y(n_880) );
OR2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_710), .Y(n_706) );
AND2x2_ASAP7_75t_L g714 ( .A(n_707), .B(n_710), .Y(n_714) );
INVx1_ASAP7_75t_L g744 ( .A(n_707), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_707), .B(n_715), .Y(n_755) );
AND2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
OR2x2_ASAP7_75t_L g743 ( .A(n_710), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g762 ( .A(n_710), .Y(n_762) );
AND2x2_ASAP7_75t_L g780 ( .A(n_710), .B(n_730), .Y(n_780) );
AND2x2_ASAP7_75t_L g795 ( .A(n_710), .B(n_744), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_710), .B(n_715), .Y(n_806) );
AOI211xp5_ASAP7_75t_SL g874 ( .A1(n_710), .A2(n_875), .B(n_876), .C(n_877), .Y(n_874) );
AND2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g750 ( .A(n_714), .B(n_730), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_714), .B(n_815), .Y(n_814) );
AND2x2_ASAP7_75t_L g840 ( .A(n_714), .B(n_715), .Y(n_840) );
NOR2x1_ASAP7_75t_R g740 ( .A(n_715), .B(n_741), .Y(n_740) );
AND2x2_ASAP7_75t_L g761 ( .A(n_715), .B(n_762), .Y(n_761) );
AND2x2_ASAP7_75t_L g803 ( .A(n_715), .B(n_795), .Y(n_803) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g731 ( .A(n_716), .Y(n_731) );
OR2x2_ASAP7_75t_L g771 ( .A(n_716), .B(n_743), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_716), .B(n_742), .Y(n_812) );
AND2x2_ASAP7_75t_L g836 ( .A(n_716), .B(n_762), .Y(n_836) );
AND2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_727), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g790 ( .A1(n_721), .A2(n_729), .B1(n_758), .B2(n_765), .C(n_791), .Y(n_790) );
AND2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
INVx2_ASAP7_75t_L g738 ( .A(n_722), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_722), .B(n_861), .Y(n_860) );
NAND2xp5_ASAP7_75t_SL g741 ( .A(n_723), .B(n_742), .Y(n_741) );
BUFx6f_ASAP7_75t_L g753 ( .A(n_723), .Y(n_753) );
INVx2_ASAP7_75t_L g764 ( .A(n_723), .Y(n_764) );
INVx2_ASAP7_75t_L g775 ( .A(n_723), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_723), .B(n_761), .Y(n_824) );
AND2x2_ASAP7_75t_L g835 ( .A(n_723), .B(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g847 ( .A(n_723), .Y(n_847) );
NAND2xp5_ASAP7_75t_SL g878 ( .A(n_723), .B(n_754), .Y(n_878) );
INVx4_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_724), .B(n_760), .Y(n_759) );
OR2x2_ASAP7_75t_L g816 ( .A(n_724), .B(n_730), .Y(n_816) );
AND2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
A2O1A1Ixp33_ASAP7_75t_L g757 ( .A1(n_727), .A2(n_758), .B(n_761), .C(n_763), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_727), .B(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g810 ( .A(n_727), .Y(n_810) );
NOR2xp33_ASAP7_75t_L g873 ( .A(n_727), .B(n_863), .Y(n_873) );
OAI221xp5_ASAP7_75t_L g877 ( .A1(n_728), .A2(n_743), .B1(n_818), .B2(n_878), .C(n_879), .Y(n_877) );
OAI21xp33_ASAP7_75t_L g804 ( .A1(n_729), .A2(n_805), .B(n_807), .Y(n_804) );
AND2x2_ASAP7_75t_L g861 ( .A(n_729), .B(n_764), .Y(n_861) );
A2O1A1O1Ixp25_ASAP7_75t_L g864 ( .A1(n_729), .A2(n_803), .B(n_852), .C(n_865), .D(n_866), .Y(n_864) );
INVx2_ASAP7_75t_SL g870 ( .A(n_729), .Y(n_870) );
AND2x4_ASAP7_75t_L g729 ( .A(n_730), .B(n_732), .Y(n_729) );
AND2x2_ASAP7_75t_L g794 ( .A(n_730), .B(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
AOI221xp5_ASAP7_75t_L g822 ( .A1(n_733), .A2(n_776), .B1(n_823), .B2(n_825), .C(n_827), .Y(n_822) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_738), .Y(n_734) );
INVx1_ASAP7_75t_SL g865 ( .A(n_735), .Y(n_865) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_738), .B(n_789), .Y(n_841) );
NOR2xp33_ASAP7_75t_L g876 ( .A(n_738), .B(n_856), .Y(n_876) );
AOI21xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_745), .B(n_748), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_742), .B(n_815), .Y(n_826) );
INVx3_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_744), .B(n_829), .Y(n_828) );
AOI221xp5_ASAP7_75t_L g879 ( .A1(n_744), .A2(n_765), .B1(n_779), .B2(n_792), .C(n_880), .Y(n_879) );
CKINVDCx14_ASAP7_75t_R g745 ( .A(n_746), .Y(n_745) );
CKINVDCx14_ASAP7_75t_R g746 ( .A(n_747), .Y(n_746) );
AND2x2_ASAP7_75t_L g844 ( .A(n_747), .B(n_829), .Y(n_844) );
AOI21xp33_ASAP7_75t_SL g748 ( .A1(n_749), .A2(n_751), .B(n_756), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g842 ( .A(n_750), .B(n_765), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_750), .B(n_857), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_754), .Y(n_751) );
AND2x2_ASAP7_75t_L g839 ( .A(n_752), .B(n_840), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_752), .B(n_852), .Y(n_851) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_753), .B(n_762), .Y(n_854) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
A2O1A1Ixp33_ASAP7_75t_L g866 ( .A1(n_755), .A2(n_841), .B(n_867), .C(n_868), .Y(n_866) );
INVx1_ASAP7_75t_L g831 ( .A(n_756), .Y(n_831) );
NOR2xp33_ASAP7_75t_L g855 ( .A(n_756), .B(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g792 ( .A(n_760), .Y(n_792) );
AND2x2_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_764), .B(n_803), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_764), .B(n_766), .Y(n_821) );
INVx1_ASAP7_75t_L g857 ( .A(n_764), .Y(n_857) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_770), .Y(n_767) );
OAI21xp5_ASAP7_75t_L g819 ( .A1(n_769), .A2(n_820), .B(n_821), .Y(n_819) );
INVx1_ASAP7_75t_L g859 ( .A(n_769), .Y(n_859) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
OAI21xp33_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_777), .B(n_780), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
NAND2xp67_ASAP7_75t_L g793 ( .A(n_775), .B(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g853 ( .A(n_776), .Y(n_853) );
INVxp67_ASAP7_75t_SL g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g867 ( .A(n_779), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_780), .B(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g850 ( .A(n_780), .Y(n_850) );
INVx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
AOI211xp5_ASAP7_75t_SL g848 ( .A1(n_782), .A2(n_849), .B(n_855), .C(n_858), .Y(n_848) );
HB1xp67_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_783), .B(n_831), .Y(n_830) );
INVx2_ASAP7_75t_L g863 ( .A(n_783), .Y(n_863) );
OAI211xp5_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_790), .B(n_796), .C(n_848), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
NOR2xp67_ASAP7_75t_SL g791 ( .A(n_792), .B(n_793), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g869 ( .A(n_792), .B(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g801 ( .A(n_794), .Y(n_801) );
AOI211xp5_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_798), .B(n_808), .C(n_837), .Y(n_796) );
OAI211xp5_ASAP7_75t_SL g798 ( .A1(n_799), .A2(n_801), .B(n_802), .C(n_804), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g820 ( .A(n_802), .Y(n_820) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
NAND3xp33_ASAP7_75t_SL g808 ( .A(n_809), .B(n_819), .C(n_822), .Y(n_808) );
A2O1A1Ixp33_ASAP7_75t_SL g809 ( .A1(n_810), .A2(n_811), .B(n_813), .C(n_817), .Y(n_809) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
OAI21xp33_ASAP7_75t_L g827 ( .A1(n_828), .A2(n_830), .B(n_832), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_833), .B(n_835), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
OAI221xp5_ASAP7_75t_L g837 ( .A1(n_838), .A2(n_841), .B1(n_842), .B2(n_843), .C(n_845), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g849 ( .A1(n_850), .A2(n_851), .B1(n_853), .B2(n_854), .Y(n_849) );
INVx1_ASAP7_75t_L g875 ( .A(n_851), .Y(n_875) );
NOR2xp33_ASAP7_75t_L g858 ( .A(n_859), .B(n_860), .Y(n_858) );
OAI22xp33_ASAP7_75t_L g862 ( .A1(n_863), .A2(n_864), .B1(n_872), .B2(n_874), .Y(n_862) );
NOR2xp33_ASAP7_75t_SL g868 ( .A(n_869), .B(n_871), .Y(n_868) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
CKINVDCx5p33_ASAP7_75t_R g881 ( .A(n_882), .Y(n_881) );
INVx2_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
AO211x2_ASAP7_75t_L g884 ( .A1(n_885), .A2(n_898), .B(n_917), .C(n_918), .Y(n_884) );
NOR2xp33_ASAP7_75t_L g885 ( .A(n_886), .B(n_891), .Y(n_885) );
AO22x2_ASAP7_75t_L g918 ( .A1(n_886), .A2(n_899), .B1(n_916), .B2(n_961), .Y(n_918) );
NAND2xp5_ASAP7_75t_SL g886 ( .A(n_887), .B(n_890), .Y(n_886) );
AO22x1_ASAP7_75t_L g917 ( .A1(n_891), .A2(n_909), .B1(n_916), .B2(n_960), .Y(n_917) );
OAI22xp5_ASAP7_75t_L g891 ( .A1(n_892), .A2(n_893), .B1(n_895), .B2(n_896), .Y(n_891) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
NOR3xp33_ASAP7_75t_L g898 ( .A(n_899), .B(n_909), .C(n_916), .Y(n_898) );
NAND2x1_ASAP7_75t_L g899 ( .A(n_900), .B(n_903), .Y(n_899) );
OA21x2_ASAP7_75t_L g903 ( .A1(n_904), .A2(n_905), .B(n_907), .Y(n_903) );
INVx1_ASAP7_75t_SL g905 ( .A(n_906), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_910), .B(n_914), .Y(n_909) );
INVx2_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
HB1xp67_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
BUFx2_ASAP7_75t_SL g925 ( .A(n_926), .Y(n_925) );
INVxp67_ASAP7_75t_SL g953 ( .A(n_929), .Y(n_953) );
OR2x2_ASAP7_75t_L g929 ( .A(n_930), .B(n_942), .Y(n_929) );
NAND3xp33_ASAP7_75t_SL g930 ( .A(n_931), .B(n_933), .C(n_935), .Y(n_930) );
OAI21xp33_ASAP7_75t_L g937 ( .A1(n_938), .A2(n_939), .B(n_940), .Y(n_937) );
NAND4xp25_ASAP7_75t_L g942 ( .A(n_943), .B(n_947), .C(n_951), .D(n_952), .Y(n_942) );
INVx1_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
BUFx2_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
endmodule