module fake_jpeg_31665_n_88 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_88);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_88;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_0),
.B(n_19),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_42),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_44),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_3),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_47),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_3),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_57),
.Y(n_59)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_31),
.B1(n_32),
.B2(n_6),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_4),
.B1(n_5),
.B2(n_10),
.Y(n_61)
);

AOI32xp33_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_34),
.A3(n_39),
.B1(n_7),
.B2(n_9),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_60),
.B(n_66),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_67),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_48),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_62),
.B(n_63),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_29),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_56),
.Y(n_64)
);

INVxp33_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_11),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_50),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_68),
.B(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_20),
.Y(n_69)
);

NOR2x1_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_21),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_22),
.Y(n_77)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_23),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_75),
.A2(n_63),
.B1(n_59),
.B2(n_53),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_79),
.C(n_74),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_78),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_73),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_80),
.C(n_72),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_76),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_70),
.B(n_27),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_86),
.A2(n_26),
.B(n_28),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_68),
.Y(n_88)
);


endmodule