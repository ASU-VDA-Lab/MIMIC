module real_aes_7785_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_679;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g110 ( .A(n_0), .Y(n_110) );
INVx1_ASAP7_75t_L g494 ( .A(n_1), .Y(n_494) );
INVx1_ASAP7_75t_L g203 ( .A(n_2), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_3), .A2(n_38), .B1(n_164), .B2(n_524), .Y(n_539) );
AOI21xp33_ASAP7_75t_L g171 ( .A1(n_4), .A2(n_145), .B(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_5), .B(n_138), .Y(n_507) );
AND2x6_ASAP7_75t_L g150 ( .A(n_6), .B(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_7), .A2(n_253), .B(n_254), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_8), .B(n_116), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_8), .B(n_39), .Y(n_461) );
INVx1_ASAP7_75t_L g178 ( .A(n_9), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_10), .B(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g143 ( .A(n_11), .Y(n_143) );
INVx1_ASAP7_75t_L g488 ( .A(n_12), .Y(n_488) );
INVx1_ASAP7_75t_L g259 ( .A(n_13), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_14), .B(n_186), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_15), .B(n_139), .Y(n_565) );
AO32x2_ASAP7_75t_L g537 ( .A1(n_16), .A2(n_138), .A3(n_183), .B1(n_516), .B2(n_538), .Y(n_537) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_17), .A2(n_63), .B1(n_127), .B2(n_128), .Y(n_126) );
INVx1_ASAP7_75t_L g128 ( .A(n_17), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_18), .B(n_164), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_19), .B(n_159), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_20), .B(n_139), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_21), .A2(n_51), .B1(n_164), .B2(n_524), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_22), .B(n_145), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_23), .A2(n_104), .B1(n_117), .B2(n_781), .Y(n_103) );
AOI22xp33_ASAP7_75t_SL g525 ( .A1(n_24), .A2(n_78), .B1(n_164), .B2(n_186), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_25), .B(n_164), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_26), .B(n_167), .Y(n_166) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_27), .A2(n_257), .B(n_258), .C(n_260), .Y(n_256) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_28), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_29), .B(n_180), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_30), .B(n_176), .Y(n_205) );
INVx1_ASAP7_75t_L g192 ( .A(n_31), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g122 ( .A1(n_32), .A2(n_123), .B1(n_124), .B2(n_455), .Y(n_122) );
INVx1_ASAP7_75t_L g455 ( .A(n_32), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_33), .B(n_180), .Y(n_554) );
INVx2_ASAP7_75t_L g148 ( .A(n_34), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_35), .B(n_164), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_36), .B(n_180), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_37), .A2(n_150), .B(n_154), .C(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g116 ( .A(n_39), .Y(n_116) );
INVx1_ASAP7_75t_L g190 ( .A(n_40), .Y(n_190) );
OAI22xp5_ASAP7_75t_SL g768 ( .A1(n_41), .A2(n_769), .B1(n_772), .B2(n_773), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_41), .Y(n_773) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_42), .B(n_176), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_43), .B(n_164), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_44), .A2(n_89), .B1(n_222), .B2(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_45), .B(n_164), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_46), .B(n_164), .Y(n_489) );
CKINVDCx16_ASAP7_75t_R g193 ( .A(n_47), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_48), .A2(n_71), .B1(n_770), .B2(n_771), .Y(n_769) );
CKINVDCx16_ASAP7_75t_R g771 ( .A(n_48), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_49), .B(n_493), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_50), .B(n_145), .Y(n_247) );
AOI22xp33_ASAP7_75t_SL g563 ( .A1(n_52), .A2(n_61), .B1(n_164), .B2(n_186), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_53), .A2(n_154), .B1(n_186), .B2(n_188), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_54), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_55), .B(n_164), .Y(n_515) );
CKINVDCx16_ASAP7_75t_R g200 ( .A(n_56), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_57), .B(n_164), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g174 ( .A1(n_58), .A2(n_163), .B(n_175), .C(n_177), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_59), .Y(n_235) );
INVx1_ASAP7_75t_L g173 ( .A(n_60), .Y(n_173) );
INVx1_ASAP7_75t_L g151 ( .A(n_62), .Y(n_151) );
INVx1_ASAP7_75t_L g127 ( .A(n_63), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_64), .B(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_65), .B(n_164), .Y(n_495) );
INVx1_ASAP7_75t_L g142 ( .A(n_66), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_67), .Y(n_120) );
AO32x2_ASAP7_75t_L g521 ( .A1(n_68), .A2(n_138), .A3(n_239), .B1(n_516), .B2(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g514 ( .A(n_69), .Y(n_514) );
INVx1_ASAP7_75t_L g549 ( .A(n_70), .Y(n_549) );
INVx1_ASAP7_75t_L g770 ( .A(n_71), .Y(n_770) );
A2O1A1Ixp33_ASAP7_75t_SL g158 ( .A1(n_72), .A2(n_159), .B(n_160), .C(n_163), .Y(n_158) );
INVxp67_ASAP7_75t_L g161 ( .A(n_73), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_74), .B(n_186), .Y(n_550) );
INVx1_ASAP7_75t_L g113 ( .A(n_75), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_76), .Y(n_196) );
INVx1_ASAP7_75t_L g228 ( .A(n_77), .Y(n_228) );
AOI222xp33_ASAP7_75t_L g465 ( .A1(n_79), .A2(n_466), .B1(n_767), .B2(n_768), .C1(n_774), .C2(n_775), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_80), .A2(n_150), .B(n_154), .C(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_81), .B(n_524), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_82), .B(n_186), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_83), .B(n_204), .Y(n_218) );
INVx2_ASAP7_75t_L g140 ( .A(n_84), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_85), .B(n_159), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_86), .B(n_186), .Y(n_503) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_87), .A2(n_150), .B(n_154), .C(n_202), .Y(n_201) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_88), .B(n_110), .C(n_111), .Y(n_109) );
OR2x2_ASAP7_75t_L g458 ( .A(n_88), .B(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g471 ( .A(n_88), .B(n_460), .Y(n_471) );
INVx2_ASAP7_75t_L g474 ( .A(n_88), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_90), .A2(n_102), .B1(n_186), .B2(n_187), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_91), .B(n_180), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_92), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g241 ( .A1(n_93), .A2(n_150), .B(n_154), .C(n_242), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_94), .Y(n_249) );
INVx1_ASAP7_75t_L g157 ( .A(n_95), .Y(n_157) );
CKINVDCx16_ASAP7_75t_R g255 ( .A(n_96), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_97), .B(n_204), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_98), .B(n_186), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_99), .B(n_138), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_100), .B(n_113), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_101), .A2(n_145), .B(n_152), .Y(n_144) );
BUFx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_SL g781 ( .A(n_107), .Y(n_781) );
AND2x2_ASAP7_75t_SL g107 ( .A(n_108), .B(n_114), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g460 ( .A(n_110), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
INVxp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AO21x1_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_121), .B(n_464), .Y(n_117) );
INVx2_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g780 ( .A(n_119), .Y(n_780) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_456), .B(n_462), .Y(n_121) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI22xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_126), .B1(n_129), .B2(n_454), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g454 ( .A(n_129), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_129), .A2(n_468), .B1(n_472), .B2(n_475), .Y(n_467) );
INVx1_ASAP7_75t_SL g777 ( .A(n_129), .Y(n_777) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND4x1_ASAP7_75t_L g130 ( .A(n_131), .B(n_372), .C(n_419), .D(n_439), .Y(n_130) );
NOR3xp33_ASAP7_75t_SL g131 ( .A(n_132), .B(n_302), .C(n_327), .Y(n_131) );
OAI211xp5_ASAP7_75t_SL g132 ( .A1(n_133), .A2(n_210), .B(n_262), .C(n_292), .Y(n_132) );
INVxp67_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_135), .B(n_181), .Y(n_134) );
INVx3_ASAP7_75t_SL g344 ( .A(n_135), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_135), .B(n_275), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_135), .B(n_197), .Y(n_425) );
AND2x2_ASAP7_75t_L g448 ( .A(n_135), .B(n_314), .Y(n_448) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_169), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g266 ( .A(n_137), .B(n_170), .Y(n_266) );
INVx3_ASAP7_75t_L g279 ( .A(n_137), .Y(n_279) );
AND2x2_ASAP7_75t_L g284 ( .A(n_137), .B(n_169), .Y(n_284) );
OR2x2_ASAP7_75t_L g335 ( .A(n_137), .B(n_276), .Y(n_335) );
BUFx2_ASAP7_75t_L g355 ( .A(n_137), .Y(n_355) );
AND2x2_ASAP7_75t_L g365 ( .A(n_137), .B(n_276), .Y(n_365) );
AND2x2_ASAP7_75t_L g371 ( .A(n_137), .B(n_182), .Y(n_371) );
OA21x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_144), .B(n_166), .Y(n_137) );
INVx4_ASAP7_75t_L g168 ( .A(n_138), .Y(n_168) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_138), .A2(n_500), .B(n_507), .Y(n_499) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g183 ( .A(n_139), .Y(n_183) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x2_ASAP7_75t_SL g180 ( .A(n_140), .B(n_141), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
BUFx2_ASAP7_75t_L g253 ( .A(n_145), .Y(n_253) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_150), .Y(n_145) );
NAND2x1p5_ASAP7_75t_L g194 ( .A(n_146), .B(n_150), .Y(n_194) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
INVx1_ASAP7_75t_L g493 ( .A(n_147), .Y(n_493) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g155 ( .A(n_148), .Y(n_155) );
INVx1_ASAP7_75t_L g187 ( .A(n_148), .Y(n_187) );
INVx1_ASAP7_75t_L g156 ( .A(n_149), .Y(n_156) );
INVx1_ASAP7_75t_L g159 ( .A(n_149), .Y(n_159) );
INVx3_ASAP7_75t_L g162 ( .A(n_149), .Y(n_162) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_149), .Y(n_176) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_149), .Y(n_189) );
INVx4_ASAP7_75t_SL g165 ( .A(n_150), .Y(n_165) );
OAI21xp5_ASAP7_75t_L g486 ( .A1(n_150), .A2(n_487), .B(n_491), .Y(n_486) );
OAI21xp5_ASAP7_75t_L g500 ( .A1(n_150), .A2(n_501), .B(n_504), .Y(n_500) );
BUFx3_ASAP7_75t_L g516 ( .A(n_150), .Y(n_516) );
OAI21xp5_ASAP7_75t_L g528 ( .A1(n_150), .A2(n_529), .B(n_533), .Y(n_528) );
OAI21xp5_ASAP7_75t_L g547 ( .A1(n_150), .A2(n_548), .B(n_551), .Y(n_547) );
O2A1O1Ixp33_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_157), .B(n_158), .C(n_165), .Y(n_152) );
O2A1O1Ixp33_ASAP7_75t_L g172 ( .A1(n_153), .A2(n_165), .B(n_173), .C(n_174), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_153), .A2(n_165), .B(n_255), .C(n_256), .Y(n_254) );
INVx5_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x6_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_155), .Y(n_164) );
BUFx3_ASAP7_75t_L g222 ( .A(n_155), .Y(n_222) );
INVx1_ASAP7_75t_L g524 ( .A(n_155), .Y(n_524) );
INVx1_ASAP7_75t_L g532 ( .A(n_159), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_162), .B(n_178), .Y(n_177) );
INVx5_ASAP7_75t_L g204 ( .A(n_162), .Y(n_204) );
OAI22xp5_ASAP7_75t_SL g522 ( .A1(n_162), .A2(n_176), .B1(n_523), .B2(n_525), .Y(n_522) );
O2A1O1Ixp5_ASAP7_75t_SL g548 ( .A1(n_163), .A2(n_204), .B(n_549), .C(n_550), .Y(n_548) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_164), .Y(n_246) );
OAI22xp33_ASAP7_75t_L g184 ( .A1(n_165), .A2(n_185), .B1(n_193), .B2(n_194), .Y(n_184) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_167), .A2(n_171), .B(n_179), .Y(n_170) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_SL g224 ( .A(n_168), .B(n_225), .Y(n_224) );
AO21x1_ASAP7_75t_L g560 ( .A1(n_168), .A2(n_561), .B(n_564), .Y(n_560) );
NAND3xp33_ASAP7_75t_L g579 ( .A(n_168), .B(n_516), .C(n_561), .Y(n_579) );
INVx1_ASAP7_75t_SL g169 ( .A(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_170), .B(n_276), .Y(n_290) );
INVx2_ASAP7_75t_L g300 ( .A(n_170), .Y(n_300) );
AND2x2_ASAP7_75t_L g313 ( .A(n_170), .B(n_279), .Y(n_313) );
OR2x2_ASAP7_75t_L g324 ( .A(n_170), .B(n_276), .Y(n_324) );
AND2x2_ASAP7_75t_SL g370 ( .A(n_170), .B(n_371), .Y(n_370) );
BUFx2_ASAP7_75t_L g382 ( .A(n_170), .Y(n_382) );
AND2x2_ASAP7_75t_L g428 ( .A(n_170), .B(n_182), .Y(n_428) );
O2A1O1Ixp5_ASAP7_75t_L g513 ( .A1(n_175), .A2(n_492), .B(n_514), .C(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_175), .A2(n_534), .B(n_535), .Y(n_533) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx4_ASAP7_75t_L g245 ( .A(n_176), .Y(n_245) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_176), .A2(n_496), .B1(n_539), .B2(n_540), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_176), .A2(n_496), .B1(n_562), .B2(n_563), .Y(n_561) );
INVx1_ASAP7_75t_L g209 ( .A(n_180), .Y(n_209) );
INVx2_ASAP7_75t_L g239 ( .A(n_180), .Y(n_239) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_180), .A2(n_252), .B(n_261), .Y(n_251) );
OA21x2_ASAP7_75t_L g527 ( .A1(n_180), .A2(n_528), .B(n_536), .Y(n_527) );
OA21x2_ASAP7_75t_L g546 ( .A1(n_180), .A2(n_547), .B(n_554), .Y(n_546) );
INVx3_ASAP7_75t_SL g301 ( .A(n_181), .Y(n_301) );
OR2x2_ASAP7_75t_L g354 ( .A(n_181), .B(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_197), .Y(n_181) );
INVx3_ASAP7_75t_L g276 ( .A(n_182), .Y(n_276) );
AND2x2_ASAP7_75t_L g343 ( .A(n_182), .B(n_198), .Y(n_343) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_182), .Y(n_411) );
AOI33xp33_ASAP7_75t_L g415 ( .A1(n_182), .A2(n_344), .A3(n_351), .B1(n_360), .B2(n_416), .B3(n_417), .Y(n_415) );
AO21x2_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_195), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_183), .B(n_196), .Y(n_195) );
AO21x2_ASAP7_75t_L g198 ( .A1(n_183), .A2(n_199), .B(n_207), .Y(n_198) );
INVx2_ASAP7_75t_L g223 ( .A(n_183), .Y(n_223) );
INVx2_ASAP7_75t_L g206 ( .A(n_186), .Y(n_206) );
INVx3_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
OAI22xp5_ASAP7_75t_SL g188 ( .A1(n_189), .A2(n_190), .B1(n_191), .B2(n_192), .Y(n_188) );
INVx2_ASAP7_75t_L g191 ( .A(n_189), .Y(n_191) );
INVx4_ASAP7_75t_L g257 ( .A(n_189), .Y(n_257) );
OAI21xp5_ASAP7_75t_L g199 ( .A1(n_194), .A2(n_200), .B(n_201), .Y(n_199) );
OAI21xp5_ASAP7_75t_L g227 ( .A1(n_194), .A2(n_228), .B(n_229), .Y(n_227) );
INVx1_ASAP7_75t_L g264 ( .A(n_197), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_197), .B(n_279), .Y(n_278) );
NOR3xp33_ASAP7_75t_L g338 ( .A(n_197), .B(n_339), .C(n_341), .Y(n_338) );
AND2x2_ASAP7_75t_L g364 ( .A(n_197), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_197), .B(n_371), .Y(n_374) );
AND2x2_ASAP7_75t_L g427 ( .A(n_197), .B(n_428), .Y(n_427) );
INVx3_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx3_ASAP7_75t_L g283 ( .A(n_198), .Y(n_283) );
OR2x2_ASAP7_75t_L g377 ( .A(n_198), .B(n_276), .Y(n_377) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_205), .C(n_206), .Y(n_202) );
INVx2_ASAP7_75t_L g496 ( .A(n_204), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_204), .A2(n_502), .B(n_503), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_204), .A2(n_511), .B(n_512), .Y(n_510) );
O2A1O1Ixp33_ASAP7_75t_L g487 ( .A1(n_206), .A2(n_488), .B(n_489), .C(n_490), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_209), .B(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_209), .B(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_236), .Y(n_210) );
AOI32xp33_ASAP7_75t_L g328 ( .A1(n_211), .A2(n_329), .A3(n_331), .B1(n_333), .B2(n_336), .Y(n_328) );
NOR2xp67_ASAP7_75t_L g401 ( .A(n_211), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g431 ( .A(n_211), .Y(n_431) );
INVx4_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g363 ( .A(n_212), .B(n_347), .Y(n_363) );
AND2x2_ASAP7_75t_L g383 ( .A(n_212), .B(n_309), .Y(n_383) );
AND2x2_ASAP7_75t_L g451 ( .A(n_212), .B(n_369), .Y(n_451) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_226), .Y(n_212) );
INVx3_ASAP7_75t_L g272 ( .A(n_213), .Y(n_272) );
AND2x2_ASAP7_75t_L g286 ( .A(n_213), .B(n_270), .Y(n_286) );
OR2x2_ASAP7_75t_L g291 ( .A(n_213), .B(n_269), .Y(n_291) );
INVx1_ASAP7_75t_L g298 ( .A(n_213), .Y(n_298) );
AND2x2_ASAP7_75t_L g306 ( .A(n_213), .B(n_280), .Y(n_306) );
AND2x2_ASAP7_75t_L g308 ( .A(n_213), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_213), .B(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g361 ( .A(n_213), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_213), .B(n_446), .Y(n_445) );
OR2x6_ASAP7_75t_L g213 ( .A(n_214), .B(n_224), .Y(n_213) );
AOI21xp5_ASAP7_75t_SL g214 ( .A1(n_215), .A2(n_216), .B(n_223), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_220), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_220), .A2(n_231), .B(n_232), .Y(n_230) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g260 ( .A(n_222), .Y(n_260) );
INVx1_ASAP7_75t_L g233 ( .A(n_223), .Y(n_233) );
OA21x2_ASAP7_75t_L g485 ( .A1(n_223), .A2(n_486), .B(n_497), .Y(n_485) );
OA21x2_ASAP7_75t_L g508 ( .A1(n_223), .A2(n_509), .B(n_517), .Y(n_508) );
INVx2_ASAP7_75t_L g270 ( .A(n_226), .Y(n_270) );
AND2x2_ASAP7_75t_L g316 ( .A(n_226), .B(n_237), .Y(n_316) );
AND2x2_ASAP7_75t_L g326 ( .A(n_226), .B(n_251), .Y(n_326) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_233), .B(n_234), .Y(n_226) );
INVx2_ASAP7_75t_L g446 ( .A(n_236), .Y(n_446) );
OR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_250), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_237), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g287 ( .A(n_237), .Y(n_287) );
AND2x2_ASAP7_75t_L g331 ( .A(n_237), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g347 ( .A(n_237), .B(n_310), .Y(n_347) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g295 ( .A(n_238), .Y(n_295) );
AND2x2_ASAP7_75t_L g309 ( .A(n_238), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g360 ( .A(n_238), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_238), .B(n_270), .Y(n_392) );
AO21x2_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_248), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_241), .B(n_247), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_246), .Y(n_242) );
AND2x2_ASAP7_75t_L g271 ( .A(n_250), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g332 ( .A(n_250), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_250), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g369 ( .A(n_250), .Y(n_369) );
INVx1_ASAP7_75t_L g402 ( .A(n_250), .Y(n_402) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g280 ( .A(n_251), .B(n_270), .Y(n_280) );
INVx1_ASAP7_75t_L g310 ( .A(n_251), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_257), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g490 ( .A(n_257), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_257), .A2(n_552), .B(n_553), .Y(n_551) );
AOI221xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_267), .B1(n_273), .B2(n_280), .C(n_281), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_264), .B(n_284), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_264), .B(n_347), .Y(n_424) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_266), .B(n_314), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_266), .B(n_275), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_266), .B(n_289), .Y(n_418) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_271), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g340 ( .A(n_270), .Y(n_340) );
AND2x2_ASAP7_75t_L g315 ( .A(n_271), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g393 ( .A(n_271), .Y(n_393) );
AND2x2_ASAP7_75t_L g325 ( .A(n_272), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_272), .B(n_295), .Y(n_341) );
AND2x2_ASAP7_75t_L g405 ( .A(n_272), .B(n_331), .Y(n_405) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
BUFx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g314 ( .A(n_276), .B(n_283), .Y(n_314) );
AND2x2_ASAP7_75t_L g410 ( .A(n_277), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_279), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_280), .B(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_280), .B(n_287), .Y(n_375) );
AND2x2_ASAP7_75t_L g395 ( .A(n_280), .B(n_295), .Y(n_395) );
AND2x2_ASAP7_75t_L g416 ( .A(n_280), .B(n_360), .Y(n_416) );
OAI32xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_285), .A3(n_287), .B1(n_288), .B2(n_291), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx1_ASAP7_75t_SL g289 ( .A(n_283), .Y(n_289) );
NAND2x1_ASAP7_75t_L g330 ( .A(n_283), .B(n_313), .Y(n_330) );
OR2x2_ASAP7_75t_L g334 ( .A(n_283), .B(n_335), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_283), .B(n_382), .Y(n_435) );
INVx1_ASAP7_75t_L g303 ( .A(n_284), .Y(n_303) );
OAI221xp5_ASAP7_75t_SL g421 ( .A1(n_285), .A2(n_376), .B1(n_422), .B2(n_425), .C(n_426), .Y(n_421) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g293 ( .A(n_286), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g336 ( .A(n_286), .B(n_309), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_286), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g414 ( .A(n_286), .B(n_347), .Y(n_414) );
INVxp67_ASAP7_75t_L g350 ( .A(n_287), .Y(n_350) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
AND2x2_ASAP7_75t_L g420 ( .A(n_289), .B(n_407), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_289), .B(n_370), .Y(n_443) );
INVx1_ASAP7_75t_L g318 ( .A(n_291), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_291), .B(n_400), .Y(n_399) );
OR2x2_ASAP7_75t_L g436 ( .A(n_291), .B(n_437), .Y(n_436) );
OAI21xp5_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_296), .B(n_299), .Y(n_292) );
AND2x2_ASAP7_75t_L g305 ( .A(n_294), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g389 ( .A(n_298), .B(n_309), .Y(n_389) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
AND2x2_ASAP7_75t_L g407 ( .A(n_300), .B(n_365), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_300), .B(n_364), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_301), .B(n_313), .Y(n_387) );
OAI211xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B(n_307), .C(n_317), .Y(n_302) );
AOI221xp5_ASAP7_75t_L g337 ( .A1(n_303), .A2(n_338), .B1(n_342), .B2(n_345), .C(n_348), .Y(n_337) );
AOI31xp33_ASAP7_75t_L g432 ( .A1(n_303), .A2(n_433), .A3(n_434), .B(n_436), .Y(n_432) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_311), .B1(n_313), .B2(n_315), .Y(n_307) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx1_ASAP7_75t_L g433 ( .A(n_313), .Y(n_433) );
INVx1_ASAP7_75t_L g396 ( .A(n_314), .Y(n_396) );
O2A1O1Ixp33_ASAP7_75t_L g439 ( .A1(n_316), .A2(n_440), .B(n_442), .C(n_444), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_319), .B1(n_321), .B2(n_325), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_322), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI221xp5_ASAP7_75t_SL g412 ( .A1(n_324), .A2(n_358), .B1(n_377), .B2(n_413), .C(n_415), .Y(n_412) );
INVx1_ASAP7_75t_L g408 ( .A(n_325), .Y(n_408) );
INVx1_ASAP7_75t_L g362 ( .A(n_326), .Y(n_362) );
NAND3xp33_ASAP7_75t_SL g327 ( .A(n_328), .B(n_337), .C(n_352), .Y(n_327) );
OAI21xp33_ASAP7_75t_L g378 ( .A1(n_329), .A2(n_379), .B(n_383), .Y(n_378) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_331), .B(n_431), .Y(n_430) );
INVxp67_ASAP7_75t_L g438 ( .A(n_332), .Y(n_438) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g376 ( .A(n_339), .B(n_359), .Y(n_376) );
INVx1_ASAP7_75t_L g351 ( .A(n_340), .Y(n_351) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g349 ( .A(n_343), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_343), .B(n_381), .Y(n_380) );
NOR4xp25_ASAP7_75t_L g348 ( .A(n_344), .B(n_349), .C(n_350), .D(n_351), .Y(n_348) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AOI222xp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_357), .B1(n_363), .B2(n_364), .C1(n_366), .C2(n_370), .Y(n_352) );
NAND2xp5_ASAP7_75t_SL g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g450 ( .A(n_354), .Y(n_450) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_362), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_366), .B(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OAI21xp5_ASAP7_75t_SL g426 ( .A1(n_371), .A2(n_427), .B(n_429), .Y(n_426) );
NOR4xp25_ASAP7_75t_L g372 ( .A(n_373), .B(n_384), .C(n_397), .D(n_412), .Y(n_372) );
OAI221xp5_ASAP7_75t_SL g373 ( .A1(n_374), .A2(n_375), .B1(n_376), .B2(n_377), .C(n_378), .Y(n_373) );
INVx1_ASAP7_75t_L g453 ( .A(n_374), .Y(n_453) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_381), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
OAI222xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_388), .B1(n_390), .B2(n_391), .C1(n_394), .C2(n_396), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI211xp5_ASAP7_75t_L g419 ( .A1(n_389), .A2(n_420), .B(n_421), .C(n_432), .Y(n_419) );
OR2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
OAI222xp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_403), .B1(n_404), .B2(n_406), .C1(n_408), .C2(n_409), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVxp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_414), .A2(n_417), .B1(n_450), .B2(n_451), .Y(n_449) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OAI211xp5_ASAP7_75t_SL g444 ( .A1(n_445), .A2(n_447), .B(n_449), .C(n_452), .Y(n_444) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g463 ( .A(n_457), .Y(n_463) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NOR2x2_ASAP7_75t_L g774 ( .A(n_459), .B(n_474), .Y(n_774) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OR2x2_ASAP7_75t_L g473 ( .A(n_460), .B(n_474), .Y(n_473) );
AOI21xp33_ASAP7_75t_L g464 ( .A1(n_462), .A2(n_465), .B(n_779), .Y(n_464) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_470), .A2(n_476), .B1(n_777), .B2(n_778), .Y(n_776) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx6_ASAP7_75t_L g778 ( .A(n_473), .Y(n_778) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_SL g476 ( .A(n_477), .B(n_733), .Y(n_476) );
NOR3xp33_ASAP7_75t_L g477 ( .A(n_478), .B(n_637), .C(n_721), .Y(n_477) );
NAND4xp25_ASAP7_75t_L g478 ( .A(n_479), .B(n_580), .C(n_602), .D(n_618), .Y(n_478) );
AOI221xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_518), .B1(n_541), .B2(n_559), .C(n_566), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_498), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_482), .B(n_559), .Y(n_592) );
NAND4xp25_ASAP7_75t_L g632 ( .A(n_482), .B(n_620), .C(n_633), .D(n_635), .Y(n_632) );
INVxp67_ASAP7_75t_L g749 ( .A(n_482), .Y(n_749) );
INVx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OR2x2_ASAP7_75t_L g631 ( .A(n_483), .B(n_569), .Y(n_631) );
AND2x2_ASAP7_75t_L g655 ( .A(n_483), .B(n_498), .Y(n_655) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g622 ( .A(n_484), .B(n_558), .Y(n_622) );
AND2x2_ASAP7_75t_L g662 ( .A(n_484), .B(n_643), .Y(n_662) );
AND2x2_ASAP7_75t_L g679 ( .A(n_484), .B(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_484), .B(n_499), .Y(n_703) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g557 ( .A(n_485), .B(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g574 ( .A(n_485), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g586 ( .A(n_485), .B(n_499), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_485), .B(n_508), .Y(n_608) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_494), .B(n_495), .C(n_496), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_496), .A2(n_505), .B(n_506), .Y(n_504) );
AND2x2_ASAP7_75t_L g589 ( .A(n_498), .B(n_590), .Y(n_589) );
AOI221xp5_ASAP7_75t_L g638 ( .A1(n_498), .A2(n_639), .B1(n_642), .B2(n_644), .C(n_648), .Y(n_638) );
AND2x2_ASAP7_75t_L g697 ( .A(n_498), .B(n_662), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_498), .B(n_679), .Y(n_731) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_508), .Y(n_498) );
INVx3_ASAP7_75t_L g558 ( .A(n_499), .Y(n_558) );
AND2x2_ASAP7_75t_L g606 ( .A(n_499), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g660 ( .A(n_499), .B(n_575), .Y(n_660) );
AND2x2_ASAP7_75t_L g718 ( .A(n_499), .B(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g559 ( .A(n_508), .B(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g575 ( .A(n_508), .Y(n_575) );
INVx1_ASAP7_75t_L g630 ( .A(n_508), .Y(n_630) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_508), .Y(n_636) );
AND2x2_ASAP7_75t_L g681 ( .A(n_508), .B(n_558), .Y(n_681) );
OR2x2_ASAP7_75t_L g720 ( .A(n_508), .B(n_560), .Y(n_720) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_513), .B(n_516), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_518), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_526), .Y(n_518) );
AND2x2_ASAP7_75t_L g716 ( .A(n_519), .B(n_713), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_519), .B(n_698), .Y(n_748) );
BUFx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g647 ( .A(n_520), .B(n_571), .Y(n_647) );
AND2x2_ASAP7_75t_L g696 ( .A(n_520), .B(n_544), .Y(n_696) );
INVx1_ASAP7_75t_L g742 ( .A(n_520), .Y(n_742) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_521), .Y(n_556) );
AND2x2_ASAP7_75t_L g597 ( .A(n_521), .B(n_571), .Y(n_597) );
INVx1_ASAP7_75t_L g614 ( .A(n_521), .Y(n_614) );
AND2x2_ASAP7_75t_L g620 ( .A(n_521), .B(n_537), .Y(n_620) );
AND2x2_ASAP7_75t_L g688 ( .A(n_526), .B(n_596), .Y(n_688) );
INVx2_ASAP7_75t_L g753 ( .A(n_526), .Y(n_753) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_537), .Y(n_526) );
AND2x2_ASAP7_75t_L g570 ( .A(n_527), .B(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g583 ( .A(n_527), .B(n_545), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_527), .B(n_544), .Y(n_611) );
INVx1_ASAP7_75t_L g617 ( .A(n_527), .Y(n_617) );
INVx1_ASAP7_75t_L g634 ( .A(n_527), .Y(n_634) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_527), .Y(n_646) );
INVx2_ASAP7_75t_L g714 ( .A(n_527), .Y(n_714) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B(n_532), .Y(n_529) );
INVx2_ASAP7_75t_L g571 ( .A(n_537), .Y(n_571) );
BUFx2_ASAP7_75t_L g668 ( .A(n_537), .Y(n_668) );
AND2x2_ASAP7_75t_L g713 ( .A(n_537), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_555), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_543), .B(n_650), .Y(n_649) );
AOI21xp5_ASAP7_75t_L g736 ( .A1(n_543), .A2(n_712), .B(n_726), .Y(n_736) );
AND2x2_ASAP7_75t_L g761 ( .A(n_543), .B(n_647), .Y(n_761) );
BUFx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g683 ( .A(n_545), .Y(n_683) );
AND2x2_ASAP7_75t_L g712 ( .A(n_545), .B(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_546), .Y(n_596) );
INVx2_ASAP7_75t_L g615 ( .A(n_546), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_546), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
INVx2_ASAP7_75t_L g569 ( .A(n_556), .Y(n_569) );
OR2x2_ASAP7_75t_L g582 ( .A(n_556), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g650 ( .A(n_556), .B(n_646), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_556), .B(n_746), .Y(n_745) );
OR2x2_ASAP7_75t_L g751 ( .A(n_556), .B(n_752), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_556), .B(n_688), .Y(n_763) );
AND2x2_ASAP7_75t_L g642 ( .A(n_557), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g665 ( .A(n_557), .B(n_559), .Y(n_665) );
INVx2_ASAP7_75t_L g577 ( .A(n_558), .Y(n_577) );
AND2x2_ASAP7_75t_L g605 ( .A(n_558), .B(n_578), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_558), .B(n_630), .Y(n_686) );
AND2x2_ASAP7_75t_L g600 ( .A(n_559), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g747 ( .A(n_559), .Y(n_747) );
AND2x2_ASAP7_75t_L g759 ( .A(n_559), .B(n_622), .Y(n_759) );
AND2x2_ASAP7_75t_L g585 ( .A(n_560), .B(n_575), .Y(n_585) );
INVx1_ASAP7_75t_L g680 ( .A(n_560), .Y(n_680) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x4_ASAP7_75t_L g578 ( .A(n_565), .B(n_579), .Y(n_578) );
INVxp67_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_572), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_569), .B(n_616), .Y(n_625) );
OR2x2_ASAP7_75t_L g757 ( .A(n_569), .B(n_758), .Y(n_757) );
AND2x2_ASAP7_75t_L g674 ( .A(n_570), .B(n_615), .Y(n_674) );
AND2x2_ASAP7_75t_L g682 ( .A(n_570), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g741 ( .A(n_570), .B(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g765 ( .A(n_570), .B(n_612), .Y(n_765) );
NOR2xp67_ASAP7_75t_L g723 ( .A(n_571), .B(n_724), .Y(n_723) );
OR2x2_ASAP7_75t_L g752 ( .A(n_571), .B(n_615), .Y(n_752) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2x1p5_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
AND2x2_ASAP7_75t_L g604 ( .A(n_574), .B(n_605), .Y(n_604) );
INVxp67_ASAP7_75t_L g766 ( .A(n_574), .Y(n_766) );
NOR2x1_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
INVx1_ASAP7_75t_L g601 ( .A(n_577), .Y(n_601) );
AND2x2_ASAP7_75t_L g652 ( .A(n_577), .B(n_585), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_577), .B(n_720), .Y(n_746) );
INVx2_ASAP7_75t_L g591 ( .A(n_578), .Y(n_591) );
INVx3_ASAP7_75t_L g643 ( .A(n_578), .Y(n_643) );
OR2x2_ASAP7_75t_L g671 ( .A(n_578), .B(n_672), .Y(n_671) );
AOI311xp33_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_584), .A3(n_586), .B(n_587), .C(n_598), .Y(n_580) );
O2A1O1Ixp33_ASAP7_75t_L g618 ( .A1(n_581), .A2(n_619), .B(n_621), .C(n_623), .Y(n_618) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_SL g603 ( .A(n_583), .Y(n_603) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g621 ( .A(n_585), .B(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_585), .B(n_601), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_585), .B(n_586), .Y(n_754) );
AND2x2_ASAP7_75t_L g676 ( .A(n_586), .B(n_590), .Y(n_676) );
AOI21xp33_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_592), .B(n_593), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g734 ( .A(n_590), .B(n_622), .Y(n_734) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_591), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g628 ( .A(n_591), .Y(n_628) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .Y(n_594) );
AND2x2_ASAP7_75t_L g619 ( .A(n_595), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g664 ( .A(n_597), .Y(n_664) );
AND2x4_ASAP7_75t_L g726 ( .A(n_597), .B(n_695), .Y(n_726) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AOI222xp33_ASAP7_75t_L g677 ( .A1(n_600), .A2(n_666), .B1(n_678), .B2(n_682), .C1(n_684), .C2(n_688), .Y(n_677) );
A2O1A1Ixp33_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .B(n_606), .C(n_609), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_603), .B(n_647), .Y(n_670) );
INVx1_ASAP7_75t_L g692 ( .A(n_605), .Y(n_692) );
INVx1_ASAP7_75t_L g626 ( .A(n_607), .Y(n_626) );
OR2x2_ASAP7_75t_L g691 ( .A(n_608), .B(n_692), .Y(n_691) );
OAI21xp33_ASAP7_75t_SL g609 ( .A1(n_610), .A2(n_612), .B(n_616), .Y(n_609) );
NAND3xp33_ASAP7_75t_L g627 ( .A(n_610), .B(n_628), .C(n_629), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g725 ( .A1(n_610), .A2(n_647), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_614), .Y(n_667) );
AND2x2_ASAP7_75t_SL g633 ( .A(n_615), .B(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g724 ( .A(n_615), .Y(n_724) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_615), .Y(n_740) );
INVx2_ASAP7_75t_L g698 ( .A(n_616), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_620), .B(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g672 ( .A(n_622), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_626), .B1(n_627), .B2(n_631), .C(n_632), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_626), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_SL g760 ( .A(n_626), .Y(n_760) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g641 ( .A(n_633), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_633), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g699 ( .A(n_633), .B(n_647), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_633), .B(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g732 ( .A(n_633), .B(n_667), .Y(n_732) );
BUFx3_ASAP7_75t_L g695 ( .A(n_634), .Y(n_695) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND5xp2_ASAP7_75t_L g637 ( .A(n_638), .B(n_656), .C(n_677), .D(n_689), .E(n_704), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AOI32xp33_ASAP7_75t_L g729 ( .A1(n_641), .A2(n_668), .A3(n_684), .B1(n_730), .B2(n_732), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_643), .B(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_SL g653 ( .A(n_647), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_651), .B1(n_653), .B2(n_654), .Y(n_648) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
AOI221xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_663), .B1(n_665), .B2(n_666), .C(n_669), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
OR2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_661), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g728 ( .A(n_660), .B(n_679), .Y(n_728) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g743 ( .A1(n_665), .A2(n_726), .B1(n_744), .B2(n_749), .C(n_750), .Y(n_743) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
INVx2_ASAP7_75t_L g709 ( .A(n_668), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_671), .B1(n_673), .B2(n_675), .Y(n_669) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_681), .Y(n_678) );
INVx1_ASAP7_75t_L g687 ( .A(n_679), .Y(n_687) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
OR2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
AOI222xp33_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_693), .B1(n_697), .B2(n_698), .C1(n_699), .C2(n_700), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .Y(n_693) );
INVxp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OAI22xp33_ASAP7_75t_L g744 ( .A1(n_698), .A2(n_745), .B1(n_747), .B2(n_748), .Y(n_744) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
AOI21xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_707), .B(n_710), .Y(n_704) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AOI21xp33_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_715), .B(n_717), .Y(n_710) );
INVx2_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g758 ( .A(n_713), .Y(n_758) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
A2O1A1Ixp33_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_725), .B(n_727), .C(n_729), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
AOI211xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_735), .B(n_737), .C(n_762), .Y(n_733) );
CKINVDCx16_ASAP7_75t_R g738 ( .A(n_734), .Y(n_738) );
INVxp67_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
OAI211xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_739), .B(n_743), .C(n_755), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
AOI21xp33_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_753), .B(n_754), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_759), .B1(n_760), .B2(n_761), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
AOI21xp33_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_764), .B(n_766), .Y(n_762) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g772 ( .A(n_769), .Y(n_772) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx2_ASAP7_75t_SL g779 ( .A(n_780), .Y(n_779) );
endmodule