module fake_jpeg_22504_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_32),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_36),
.Y(n_51)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_1),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_41),
.A2(n_30),
.B(n_28),
.C(n_21),
.Y(n_42)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_42),
.A2(n_48),
.B(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_22),
.B1(n_25),
.B2(n_18),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_47),
.A2(n_49),
.B1(n_61),
.B2(n_15),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_21),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_34),
.A2(n_22),
.B1(n_25),
.B2(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_18),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_30),
.B(n_19),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_24),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_16),
.Y(n_59)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_15),
.Y(n_60)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_37),
.A2(n_25),
.B1(n_22),
.B2(n_21),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_63),
.A2(n_44),
.B1(n_57),
.B2(n_56),
.Y(n_96)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_68),
.Y(n_95)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_75),
.Y(n_97)
);

BUFx24_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_27),
.B1(n_17),
.B2(n_29),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_74),
.B1(n_50),
.B2(n_46),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_77),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_53),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_37),
.B1(n_39),
.B2(n_30),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_48),
.B1(n_58),
.B2(n_51),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_80),
.A2(n_86),
.B1(n_88),
.B2(n_96),
.Y(n_118)
);

NAND2xp33_ASAP7_75t_SL g81 ( 
.A(n_70),
.B(n_30),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_87),
.B(n_99),
.Y(n_103)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_83),
.Y(n_101)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_90),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_47),
.B1(n_49),
.B2(n_51),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_1),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_91),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_45),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_79),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_78),
.A2(n_44),
.B1(n_57),
.B2(n_56),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_92),
.A2(n_44),
.B1(n_66),
.B2(n_74),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_67),
.B(n_59),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_60),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_76),
.A2(n_52),
.B(n_43),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_66),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_102),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_105),
.Y(n_131)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_SL g106 ( 
.A1(n_93),
.A2(n_74),
.B(n_77),
.C(n_30),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_106),
.A2(n_117),
.B(n_100),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_109),
.A2(n_110),
.B1(n_119),
.B2(n_92),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_74),
.B1(n_57),
.B2(n_67),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_43),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_87),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_64),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_112),
.Y(n_126)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_115),
.B1(n_89),
.B2(n_91),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_81),
.Y(n_115)
);

NOR3xp33_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_16),
.C(n_26),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_116),
.B(n_54),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_2),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_85),
.A2(n_26),
.B1(n_39),
.B2(n_17),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_101),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_120),
.B(n_121),
.Y(n_147)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_123),
.Y(n_139)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_124),
.A2(n_128),
.B(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_136),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_127),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_119),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_106),
.A2(n_91),
.B1(n_90),
.B2(n_84),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_130),
.A2(n_134),
.B1(n_19),
.B2(n_4),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_132),
.B(n_103),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_108),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_88),
.B1(n_84),
.B2(n_89),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_106),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_135)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_103),
.C(n_115),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_143),
.C(n_148),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_141),
.B(n_132),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_108),
.C(n_134),
.Y(n_143)
);

OAI32xp33_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_106),
.A3(n_108),
.B1(n_111),
.B2(n_117),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_130),
.Y(n_157)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_126),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_104),
.C(n_30),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_19),
.C(n_4),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_151),
.A2(n_129),
.B1(n_123),
.B2(n_142),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_120),
.Y(n_152)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_152),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_153),
.A2(n_160),
.B(n_164),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_154),
.Y(n_174)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_165),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_124),
.Y(n_158)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_150),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_150),
.A2(n_128),
.B1(n_137),
.B2(n_5),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_151),
.B1(n_140),
.B2(n_149),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_138),
.C(n_146),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_3),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_143),
.A2(n_3),
.B(n_4),
.Y(n_165)
);

XOR2x2_ASAP7_75t_SL g168 ( 
.A(n_157),
.B(n_146),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_168),
.A2(n_6),
.B(n_8),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_148),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_159),
.C(n_158),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_170),
.A2(n_155),
.B1(n_160),
.B2(n_165),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_175),
.B(n_5),
.Y(n_182)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_166),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_180),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_171),
.A2(n_163),
.B1(n_164),
.B2(n_161),
.Y(n_177)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_177),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_181),
.C(n_182),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_179),
.A2(n_173),
.B1(n_168),
.B2(n_167),
.Y(n_188)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_162),
.C(n_6),
.Y(n_181)
);

OAI21x1_ASAP7_75t_L g189 ( 
.A1(n_183),
.A2(n_170),
.B(n_8),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_R g187 ( 
.A(n_181),
.B(n_174),
.Y(n_187)
);

NAND3xp33_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_189),
.C(n_6),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_190),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_169),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_10),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_186),
.A2(n_185),
.B1(n_184),
.B2(n_172),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_194),
.C(n_195),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_190),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_184),
.A2(n_177),
.B(n_9),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_8),
.C(n_10),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_197),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_11),
.B(n_12),
.Y(n_199)
);

OAI21x1_ASAP7_75t_SL g201 ( 
.A1(n_199),
.A2(n_12),
.B(n_13),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_201),
.A2(n_200),
.B1(n_196),
.B2(n_13),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_12),
.Y(n_203)
);


endmodule