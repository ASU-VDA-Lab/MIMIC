module fake_jpeg_21601_n_103 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_103);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_103;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_13),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_29),
.Y(n_34)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_12),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_23),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_4),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_14),
.B(n_21),
.C(n_22),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_39),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_22),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_17),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_4),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_26),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_43),
.B(n_47),
.Y(n_62)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_50),
.Y(n_70)
);

AO21x1_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_51),
.B(n_55),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_29),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_49),
.Y(n_63)
);

NOR2x1_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_17),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_14),
.B1(n_21),
.B2(n_20),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_57),
.B1(n_61),
.B2(n_5),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_22),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_10),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_53),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_25),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_59),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_33),
.A2(n_25),
.B1(n_24),
.B2(n_18),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_19),
.B1(n_16),
.B2(n_7),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_36),
.B(n_38),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_55),
.B(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_71),
.A2(n_48),
.B1(n_61),
.B2(n_47),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_41),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_72),
.B(n_49),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_60),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_74),
.B(n_76),
.Y(n_87)
);

AOI221xp5_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_66),
.B1(n_65),
.B2(n_64),
.C(n_62),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_52),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_77),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_78),
.A2(n_64),
.B1(n_57),
.B2(n_55),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_81),
.A2(n_44),
.B1(n_69),
.B2(n_68),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_63),
.C(n_72),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_84),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_85),
.Y(n_89)
);

NOR2xp67_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_77),
.Y(n_88)
);

NOR3xp33_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_6),
.C(n_7),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_86),
.A2(n_81),
.B1(n_71),
.B2(n_74),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_85),
.B1(n_51),
.B2(n_79),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_80),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_63),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_91),
.Y(n_98)
);

AOI321xp33_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_62),
.A3(n_82),
.B1(n_65),
.B2(n_67),
.C(n_11),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_95),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_90),
.B(n_89),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_97),
.A2(n_98),
.B(n_16),
.Y(n_100)
);

MAJx2_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_8),
.C(n_9),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_101),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_19),
.B1(n_41),
.B2(n_38),
.Y(n_103)
);


endmodule