module real_jpeg_14198_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx2_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_2),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_4),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_51),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_5),
.A2(n_47),
.B1(n_48),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_5),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_32),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_7),
.A2(n_32),
.B1(n_47),
.B2(n_48),
.Y(n_139)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_9),
.A2(n_47),
.B1(n_48),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_9),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_10),
.B(n_41),
.Y(n_40)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_10),
.A2(n_24),
.B(n_30),
.C(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_10),
.B(n_85),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_75),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_10),
.B(n_48),
.C(n_62),
.Y(n_124)
);

NAND2x1_ASAP7_75t_SL g128 ( 
.A(n_10),
.B(n_23),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_L g148 ( 
.A1(n_10),
.A2(n_52),
.B(n_134),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_75),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_11),
.A2(n_43),
.B1(n_85),
.B2(n_86),
.Y(n_92)
);

NAND2xp33_ASAP7_75t_SL g107 ( 
.A(n_11),
.B(n_31),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_12),
.A2(n_30),
.B1(n_31),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_35),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_12),
.A2(n_35),
.B1(n_47),
.B2(n_48),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_12),
.A2(n_35),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_13),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_67),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_13),
.A2(n_47),
.B1(n_48),
.B2(n_67),
.Y(n_133)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_115),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_113),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_79),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_18),
.B(n_79),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_58),
.C(n_71),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_19),
.A2(n_20),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_38),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_21),
.B(n_39),
.C(n_45),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_29),
.B(n_33),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_22),
.A2(n_29),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2x1_ASAP7_75t_R g36 ( 
.A(n_23),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_23),
.B(n_34),
.Y(n_161)
);

AO22x1_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_23)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_24),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_25),
.A2(n_26),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_L g74 ( 
.A1(n_25),
.A2(n_28),
.B(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_26),
.B(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI32xp33_ASAP7_75t_L g106 ( 
.A1(n_30),
.A2(n_43),
.A3(n_86),
.B1(n_90),
.B2(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_44),
.B2(n_45),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_42),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_42),
.B(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_52),
.B1(n_55),
.B2(n_57),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_57),
.B(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_54),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_48),
.B1(n_62),
.B2(n_63),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_47),
.B(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_52),
.A2(n_55),
.B1(n_57),
.B2(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_52),
.A2(n_133),
.B(n_134),
.Y(n_132)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_53),
.A2(n_54),
.B1(n_138),
.B2(n_140),
.Y(n_137)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_54),
.B(n_78),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_57),
.A2(n_77),
.B(n_139),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_57),
.B(n_75),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_58),
.A2(n_71),
.B1(n_72),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_58),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_65),
.B(n_68),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_SL g121 ( 
.A1(n_59),
.A2(n_68),
.B(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_60),
.B(n_70),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_60),
.A2(n_66),
.B1(n_69),
.B2(n_163),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_64),
.A2(n_98),
.B(n_100),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_64),
.A2(n_100),
.B(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_64),
.B(n_75),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_73),
.B(n_76),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_86),
.B(n_89),
.C(n_91),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_102),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_93),
.B2(n_101),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_88),
.Y(n_82)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_97),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_95),
.A2(n_160),
.B(n_161),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_108),
.B2(n_109),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_167),
.B(n_173),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_154),
.B(n_166),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_135),
.B(n_153),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_125),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_119),
.B(n_125),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_123),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_120),
.A2(n_121),
.B1(n_123),
.B2(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_123),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_132),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_130),
.C(n_132),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_133),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_143),
.B(n_152),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_141),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_137),
.B(n_141),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_147),
.B(n_151),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_145),
.B(n_146),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_155),
.B(n_156),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_162),
.C(n_165),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_162),
.B1(n_164),
.B2(n_165),
.Y(n_158)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_159),
.Y(n_165)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_162),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_168),
.B(n_169),
.Y(n_173)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);


endmodule