module fake_jpeg_3602_n_177 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_177);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_51),
.B(n_0),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_65),
.Y(n_74)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_42),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_47),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

CKINVDCx12_ASAP7_75t_R g78 ( 
.A(n_67),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_66),
.A2(n_60),
.B1(n_53),
.B2(n_44),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_63),
.B(n_49),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_71),
.B(n_52),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_58),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_57),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_65),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_54),
.B1(n_48),
.B2(n_42),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_60),
.B1(n_47),
.B2(n_61),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_54),
.B1(n_48),
.B2(n_46),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_76),
.A2(n_75),
.B(n_66),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_45),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_78),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_88),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_77),
.B1(n_79),
.B2(n_68),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_83),
.B(n_56),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_50),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_84),
.B(n_91),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_73),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_92),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_90),
.A2(n_67),
.B1(n_62),
.B2(n_68),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_46),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_49),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_94),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_0),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_86),
.A2(n_76),
.B1(n_62),
.B2(n_79),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_100),
.B1(n_106),
.B2(n_107),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_98),
.A2(n_110),
.B1(n_1),
.B2(n_2),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_86),
.A2(n_62),
.B1(n_52),
.B2(n_47),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_103),
.B(n_1),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_94),
.Y(n_104)
);

NAND3xp33_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_4),
.C(n_5),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_55),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_3),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_83),
.A2(n_67),
.B1(n_43),
.B2(n_56),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_109),
.B(n_18),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_83),
.A2(n_56),
.B1(n_2),
.B2(n_3),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_113),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_88),
.B(n_82),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_126),
.B(n_100),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_118),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_85),
.C(n_19),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_124),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_121),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_41),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_123),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_21),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_4),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_129),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_5),
.B(n_7),
.Y(n_126)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_25),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_27),
.Y(n_143)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_128),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_38),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_131),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_8),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_133),
.A2(n_141),
.B1(n_146),
.B2(n_14),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_SL g136 ( 
.A1(n_132),
.A2(n_96),
.B(n_112),
.C(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_138),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_121),
.B(n_9),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_145),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_129),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_114),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_123),
.B(n_13),
.Y(n_147)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_122),
.A2(n_30),
.B(n_35),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_28),
.C(n_34),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_148),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

OAI32xp33_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_128),
.A3(n_126),
.B1(n_118),
.B2(n_127),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_152),
.A2(n_139),
.B(n_134),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_140),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_154),
.A2(n_159),
.B1(n_137),
.B2(n_141),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_24),
.C(n_33),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_137),
.C(n_135),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_161),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_162),
.A2(n_163),
.B1(n_150),
.B2(n_156),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_157),
.C(n_155),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_153),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_167),
.C(n_168),
.Y(n_171)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_169),
.A2(n_165),
.B(n_136),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_170),
.A2(n_136),
.B(n_154),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_136),
.B1(n_171),
.B2(n_167),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_173),
.B(n_37),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_14),
.B(n_15),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_16),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_16),
.Y(n_177)
);


endmodule