module fake_jpeg_23395_n_224 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_224);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_2),
.B(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_0),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_0),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_2),
.Y(n_79)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_24),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_22),
.B(n_1),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_46),
.B(n_35),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_44),
.A2(n_31),
.B1(n_25),
.B2(n_24),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_48),
.A2(n_71),
.B1(n_76),
.B2(n_5),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_34),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_23),
.Y(n_81)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_20),
.B1(n_27),
.B2(n_31),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_61),
.Y(n_88)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_17),
.Y(n_59)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_64),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_20),
.B1(n_25),
.B2(n_34),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_72),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_45),
.B(n_19),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_69),
.B(n_2),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_19),
.B1(n_33),
.B2(n_35),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_37),
.A2(n_33),
.B1(n_29),
.B2(n_23),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_38),
.B(n_29),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_74),
.Y(n_105)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_37),
.A2(n_32),
.B1(n_30),
.B2(n_26),
.Y(n_76)
);

BUFx4f_ASAP7_75t_SL g78 ( 
.A(n_36),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_21),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_81),
.B(n_100),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_32),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_89),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_32),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_96),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_49),
.A2(n_30),
.B(n_26),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_93),
.C(n_99),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_78),
.B(n_30),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_26),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_101),
.Y(n_129)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_98),
.B(n_6),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_66),
.A2(n_21),
.B(n_4),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_66),
.B(n_3),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_4),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_108),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_103),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_51),
.B(n_5),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_13),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_109),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_61),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_112),
.Y(n_151)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_114),
.B(n_116),
.Y(n_142)
);

AO22x1_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_76),
.B1(n_77),
.B2(n_54),
.Y(n_115)
);

AO22x1_ASAP7_75t_L g147 ( 
.A1(n_115),
.A2(n_58),
.B1(n_93),
.B2(n_92),
.Y(n_147)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_60),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_118),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_107),
.A2(n_54),
.B1(n_77),
.B2(n_67),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_119),
.A2(n_123),
.B1(n_124),
.B2(n_127),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_122),
.Y(n_156)
);

OAI22x1_ASAP7_75t_SL g123 ( 
.A1(n_87),
.A2(n_58),
.B1(n_62),
.B2(n_75),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_84),
.A2(n_94),
.B1(n_89),
.B2(n_86),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_99),
.A2(n_52),
.B1(n_74),
.B2(n_72),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

INVxp67_ASAP7_75t_SL g144 ( 
.A(n_128),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_95),
.B(n_50),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

HAxp5_ASAP7_75t_SL g143 ( 
.A(n_132),
.B(n_135),
.CON(n_143),
.SN(n_143)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_91),
.A2(n_92),
.B1(n_102),
.B2(n_93),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_95),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_50),
.Y(n_134)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_81),
.B(n_7),
.Y(n_136)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_101),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_146),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_121),
.C(n_133),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_145),
.C(n_159),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_113),
.A2(n_93),
.B(n_98),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_145),
.A2(n_152),
.B(n_116),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_100),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_147),
.A2(n_126),
.B1(n_115),
.B2(n_123),
.Y(n_169)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_150),
.B(n_154),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_SL g152 ( 
.A1(n_115),
.A2(n_100),
.B(n_90),
.C(n_106),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_129),
.Y(n_165)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_82),
.Y(n_155)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_111),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_158),
.B(n_160),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_127),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g164 ( 
.A1(n_146),
.A2(n_161),
.B(n_139),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_164),
.A2(n_178),
.B(n_149),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_175),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_172),
.C(n_174),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_169),
.A2(n_179),
.B1(n_180),
.B2(n_157),
.Y(n_192)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_142),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_173),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_124),
.C(n_135),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_120),
.C(n_129),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_132),
.Y(n_176)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_114),
.C(n_110),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_148),
.C(n_152),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_151),
.A2(n_128),
.B(n_110),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_97),
.B1(n_80),
.B2(n_106),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_80),
.B1(n_97),
.B2(n_137),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_152),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_188),
.Y(n_199)
);

OAI321xp33_ASAP7_75t_L g182 ( 
.A1(n_175),
.A2(n_152),
.A3(n_138),
.B1(n_143),
.B2(n_144),
.C(n_154),
.Y(n_182)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

OAI22x1_ASAP7_75t_SL g185 ( 
.A1(n_177),
.A2(n_152),
.B1(n_148),
.B2(n_162),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_185),
.A2(n_191),
.B1(n_192),
.B2(n_163),
.Y(n_195)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_82),
.C(n_85),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_171),
.A2(n_150),
.B1(n_149),
.B2(n_156),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_157),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_141),
.B(n_112),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_197),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_185),
.A2(n_163),
.B1(n_173),
.B2(n_172),
.Y(n_196)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_174),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_165),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_165),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_202),
.Y(n_204)
);

MAJx2_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_170),
.C(n_179),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_193),
.C(n_186),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_194),
.C(n_184),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_207),
.Y(n_214)
);

AOI31xp67_ASAP7_75t_SL g207 ( 
.A1(n_198),
.A2(n_191),
.A3(n_186),
.B(n_187),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_7),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_210),
.Y(n_212)
);

AOI31xp67_ASAP7_75t_L g211 ( 
.A1(n_206),
.A2(n_199),
.A3(n_202),
.B(n_209),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_204),
.Y(n_215)
);

NAND2xp33_ASAP7_75t_SL g213 ( 
.A(n_208),
.B(n_197),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_8),
.Y(n_216)
);

NAND3xp33_ASAP7_75t_SL g218 ( 
.A(n_215),
.B(n_217),
.C(n_212),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_9),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_9),
.Y(n_217)
);

NOR3xp33_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_219),
.C(n_11),
.Y(n_221)
);

AOI21x1_ASAP7_75t_L g220 ( 
.A1(n_218),
.A2(n_213),
.B(n_12),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_220),
.A2(n_12),
.B(n_13),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_221),
.B(n_12),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_223),
.Y(n_224)
);


endmodule