module fake_jpeg_959_n_56 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_56);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_56;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx4_ASAP7_75t_L g8 ( 
.A(n_7),
.Y(n_8)
);

INVx6_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

OAI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_18),
.A2(n_15),
.B1(n_16),
.B2(n_11),
.Y(n_27)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_2),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_22),
.Y(n_28)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_11),
.B(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_3),
.B(n_4),
.C(n_6),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_12),
.B(n_15),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_21),
.A2(n_14),
.B1(n_16),
.B2(n_9),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_27),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_18),
.B(n_22),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_38),
.C(n_26),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_37),
.B(n_39),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_30),
.A2(n_23),
.B(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_9),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_30),
.C(n_29),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_17),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_45),
.C(n_19),
.Y(n_48)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_47),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_48),
.A2(n_49),
.B1(n_43),
.B2(n_19),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g49 ( 
.A(n_44),
.B(n_12),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_47),
.C(n_40),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_53),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_51),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_55),
.B(n_0),
.Y(n_56)
);


endmodule