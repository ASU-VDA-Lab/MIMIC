module fake_netlist_6_2220_n_124 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_25, n_124);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_25;

output n_124;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_68;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_121;
wire n_47;
wire n_62;
wire n_75;
wire n_109;
wire n_122;
wire n_45;
wire n_34;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_61;
wire n_112;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_55;
wire n_97;
wire n_94;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_60;
wire n_35;
wire n_115;
wire n_69;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVxp67_ASAP7_75t_SL g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp67_ASAP7_75t_L g38 ( 
.A(n_11),
.B(n_25),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

INVxp67_ASAP7_75t_SL g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_9),
.B(n_30),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_28),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_4),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_0),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_2),
.Y(n_59)
);

AND2x4_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_2),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

AND2x6_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_15),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_17),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

AND2x6_ASAP7_75t_L g66 ( 
.A(n_33),
.B(n_22),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_40),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_35),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_68),
.B(n_47),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_59),
.B(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_55),
.B(n_54),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_60),
.B(n_44),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g73 ( 
.A(n_60),
.B(n_52),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_65),
.B(n_37),
.Y(n_74)
);

NAND2xp33_ASAP7_75t_R g75 ( 
.A(n_63),
.B(n_36),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_67),
.B(n_42),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_31),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_57),
.B(n_45),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_61),
.B(n_38),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_61),
.B(n_49),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

OAI21x1_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_64),
.B(n_48),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

AO21x2_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_46),
.B(n_66),
.Y(n_86)
);

OAI21x1_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_66),
.B(n_62),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_69),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_58),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_66),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_74),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

NAND3xp33_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_81),
.C(n_84),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_89),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_96),
.Y(n_103)
);

AO221x2_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_88),
.B1(n_85),
.B2(n_81),
.C(n_84),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_96),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_85),
.B(n_91),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);

AND2x4_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_101),
.Y(n_112)
);

NOR2x1_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_108),
.Y(n_113)
);

AOI211xp5_ASAP7_75t_SL g114 ( 
.A1(n_112),
.A2(n_110),
.B(n_92),
.C(n_93),
.Y(n_114)
);

AOI322xp5_ASAP7_75t_L g115 ( 
.A1(n_112),
.A2(n_107),
.A3(n_93),
.B1(n_66),
.B2(n_58),
.C1(n_56),
.C2(n_86),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_83),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_86),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_116),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_117),
.A2(n_115),
.B1(n_82),
.B2(n_96),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

AOI31xp33_ASAP7_75t_L g121 ( 
.A1(n_119),
.A2(n_23),
.A3(n_26),
.B(n_27),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_86),
.B1(n_62),
.B2(n_87),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g123 ( 
.A1(n_121),
.A2(n_118),
.B(n_87),
.Y(n_123)
);

AOI221xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_56),
.B1(n_62),
.B2(n_122),
.C(n_121),
.Y(n_124)
);


endmodule