module real_aes_4983_n_7 (n_4, n_0, n_3, n_5, n_2, n_6, n_1, n_7);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_6;
input n_1;
output n_7;
wire n_17;
wire n_16;
wire n_13;
wire n_15;
wire n_8;
wire n_9;
wire n_12;
wire n_14;
wire n_10;
wire n_11;
NOR2xp33_ASAP7_75t_L g8 ( .A(n_0), .B(n_9), .Y(n_8) );
AOI221xp5_ASAP7_75t_L g7 ( .A1(n_1), .A2(n_8), .B1(n_11), .B2(n_12), .C(n_15), .Y(n_7) );
OAI22xp5_ASAP7_75t_L g12 ( .A1(n_2), .A2(n_4), .B1(n_13), .B2(n_14), .Y(n_12) );
INVx1_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
AND2x2_ASAP7_75t_L g16 ( .A(n_3), .B(n_17), .Y(n_16) );
INVx2_ASAP7_75t_L g13 ( .A(n_4), .Y(n_13) );
BUFx3_ASAP7_75t_L g10 ( .A(n_5), .Y(n_10) );
INVx1_ASAP7_75t_L g17 ( .A(n_6), .Y(n_17) );
CKINVDCx14_ASAP7_75t_R g11 ( .A(n_8), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g9 ( .A(n_10), .Y(n_9) );
CKINVDCx16_ASAP7_75t_R g15 ( .A(n_16), .Y(n_15) );
endmodule