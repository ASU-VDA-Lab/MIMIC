module real_jpeg_4828_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx1_ASAP7_75t_SL g30 ( 
.A(n_0),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_0),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_0),
.B(n_35),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_0),
.B(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_SL g224 ( 
.A(n_0),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_0),
.B(n_398),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_1),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_2),
.Y(n_91)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_2),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_2),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_2),
.Y(n_287)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_2),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_3),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_3),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_3),
.B(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_SL g221 ( 
.A(n_3),
.B(n_222),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_3),
.B(n_236),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_3),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_3),
.B(n_253),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_3),
.B(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_4),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_4),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_4),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_4),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_4),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_5),
.B(n_49),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_5),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_5),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_5),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_5),
.B(n_174),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_5),
.B(n_259),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_5),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_5),
.B(n_409),
.Y(n_408)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_6),
.Y(n_95)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_6),
.Y(n_110)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_6),
.Y(n_266)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_7),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_8),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_8),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_8),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_8),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_8),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_8),
.B(n_387),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_8),
.B(n_427),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g225 ( 
.A(n_9),
.Y(n_225)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_9),
.Y(n_239)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_9),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_9),
.Y(n_325)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_11),
.Y(n_162)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_11),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_12),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_12),
.B(n_100),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_12),
.B(n_42),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_12),
.B(n_49),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_12),
.B(n_238),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_12),
.B(n_289),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_12),
.B(n_259),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_12),
.B(n_136),
.Y(n_410)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_14),
.B(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_14),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_14),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g112 ( 
.A(n_14),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_14),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_15),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_15),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_15),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_15),
.B(n_299),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_15),
.B(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_15),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_15),
.B(n_219),
.Y(n_380)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_17),
.B(n_32),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_17),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_17),
.B(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_17),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_17),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_17),
.B(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_17),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_18),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_18),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_18),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_18),
.B(n_161),
.Y(n_160)
);

AND2x2_ASAP7_75t_SL g383 ( 
.A(n_18),
.B(n_384),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_19),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_19),
.B(n_211),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_19),
.B(n_233),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_19),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_19),
.B(n_301),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_19),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_19),
.B(n_238),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_19),
.B(n_404),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_478),
.B(n_480),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_180),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_179),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_144),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_25),
.B(n_144),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_104),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_72),
.C(n_86),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_27),
.B(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_47),
.C(n_57),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_28),
.B(n_47),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_33),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_29),
.B(n_39),
.C(n_46),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_30),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_30),
.B(n_256),
.Y(n_255)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_32),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_39),
.B1(n_40),
.B2(n_46),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_36),
.Y(n_234)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_38),
.Y(n_125)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_38),
.Y(n_346)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_44),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_44),
.Y(n_341)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_45),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_45),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_52),
.C(n_54),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_48),
.B(n_54),
.Y(n_164)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_52),
.B(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_57),
.B(n_470),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_63),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_58),
.B(n_64),
.C(n_71),
.Y(n_142)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_61),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_62),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_62),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_66),
.B2(n_71),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_108),
.C(n_111),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_64),
.A2(n_65),
.B1(n_111),
.B2(n_112),
.Y(n_141)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_89),
.C(n_92),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_66),
.A2(n_71),
.B1(n_89),
.B2(n_90),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_70),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_70),
.Y(n_299)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_70),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_72),
.A2(n_86),
.B1(n_87),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_77),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_73),
.B(n_78),
.C(n_81),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_96),
.C(n_101),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_88),
.B(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_89),
.B(n_157),
.C(n_160),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_89),
.A2(n_90),
.B1(n_160),
.B2(n_441),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_92),
.B(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_96),
.A2(n_97),
.B1(n_101),
.B2(n_102),
.Y(n_166)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_101),
.A2(n_102),
.B1(n_177),
.B2(n_178),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_102),
.B(n_168),
.C(n_177),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_139),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_129),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_114),
.B1(n_127),
.B2(n_128),
.Y(n_106)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_141),
.Y(n_140)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_111),
.A2(n_112),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_113),
.Y(n_312)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_119),
.B1(n_120),
.B2(n_126),
.Y(n_114)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_124),
.Y(n_253)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_134),
.B1(n_135),
.B2(n_138),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_132),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_137),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.C(n_143),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_143),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.C(n_150),
.Y(n_144)
);

FAx1_ASAP7_75t_L g474 ( 
.A(n_145),
.B(n_148),
.CI(n_150),
.CON(n_474),
.SN(n_474)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_165),
.C(n_167),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_151),
.A2(n_152),
.B1(n_467),
.B2(n_468),
.Y(n_466)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.C(n_163),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_153),
.A2(n_154),
.B1(n_450),
.B2(n_451),
.Y(n_449)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_156),
.B(n_163),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_157),
.A2(n_158),
.B1(n_439),
.B2(n_440),
.Y(n_438)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_160),
.Y(n_441)
);

BUFx8_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_162),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_162),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_165),
.B(n_167),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_169),
.B(n_458),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.C(n_176),
.Y(n_169)
);

FAx1_ASAP7_75t_SL g435 ( 
.A(n_170),
.B(n_173),
.CI(n_176),
.CON(n_435),
.SN(n_435)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AO21x1_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_473),
.B(n_476),
.Y(n_180)
);

OAI21x1_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_462),
.B(n_472),
.Y(n_181)
);

AOI21x1_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_445),
.B(n_461),
.Y(n_182)
);

OAI21x1_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_414),
.B(n_444),
.Y(n_183)
);

AOI21x1_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_373),
.B(n_413),
.Y(n_184)
);

AO21x1_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_292),
.B(n_372),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_277),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_187),
.B(n_277),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_228),
.B2(n_276),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_188),
.B(n_229),
.C(n_260),
.Y(n_412)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_205),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_190),
.B(n_206),
.C(n_227),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_202),
.C(n_204),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_191),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_196),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_192),
.A2(n_193),
.B1(n_196),
.B2(n_197),
.Y(n_282)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_201),
.Y(n_209)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_201),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_202),
.B(n_204),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_215),
.B1(n_226),
.B2(n_227),
.Y(n_205)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_210),
.B(n_214),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_210),
.Y(n_214)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_214),
.B(n_391),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_214),
.B(n_378),
.C(n_391),
.Y(n_421)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_220),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_216),
.B(n_221),
.C(n_224),
.Y(n_411)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_224),
.Y(n_220)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_228),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_260),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_241),
.C(n_254),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_230),
.B(n_279),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_240),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_235),
.Y(n_231)
);

MAJx2_ASAP7_75t_L g275 ( 
.A(n_232),
.B(n_235),
.C(n_240),
.Y(n_275)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_239),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_241),
.A2(n_242),
.B1(n_254),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

MAJx2_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_246),
.C(n_251),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_243),
.A2(n_244),
.B1(n_251),
.B2(n_252),
.Y(n_365)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_246),
.B(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_249),
.Y(n_400)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_258),
.Y(n_274)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_259),
.Y(n_329)
);

XOR2x1_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_273),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_261),
.B(n_274),
.C(n_275),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

MAJx2_ASAP7_75t_L g391 ( 
.A(n_262),
.B(n_267),
.C(n_271),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_267),
.B1(n_271),
.B2(n_272),
.Y(n_263)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_264),
.Y(n_271)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_266),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_267),
.Y(n_272)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_270),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_281),
.C(n_290),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_278),
.B(n_370),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_281),
.B(n_290),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.C(n_284),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_282),
.B(n_283),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_284),
.B(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_288),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_285),
.B(n_288),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI21x1_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_367),
.B(n_371),
.Y(n_292)
);

OA21x2_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_352),
.B(n_366),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_332),
.B(n_351),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_296),
.A2(n_319),
.B(n_331),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_303),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_303),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_298),
.B(n_300),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_298),
.B(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_313),
.B2(n_314),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_310),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_306),
.B(n_310),
.C(n_313),
.Y(n_350)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

BUFx5_ASAP7_75t_L g428 ( 
.A(n_309),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_318),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_315),
.B(n_318),
.Y(n_336)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_326),
.B(n_330),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_322),
.Y(n_330)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_350),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_333),
.B(n_350),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_337),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_336),
.C(n_354),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_337),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_342),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_338),
.B(n_347),
.C(n_349),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

INVx11_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_347),
.B1(n_348),
.B2(n_349),
.Y(n_342)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_343),
.Y(n_349)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_355),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_353),
.B(n_355),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_356),
.A2(n_357),
.B1(n_359),
.B2(n_360),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_356),
.B(n_362),
.C(n_363),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_362),
.B1(n_363),
.B2(n_364),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_364),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_368),
.B(n_369),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_374),
.B(n_412),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_374),
.B(n_412),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_393),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_376),
.B(n_377),
.C(n_393),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_379),
.B1(n_390),
.B2(n_392),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_380),
.B(n_383),
.C(n_385),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_382),
.A2(n_383),
.B1(n_385),
.B2(n_386),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_390),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_394),
.B(n_395),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_394),
.B(n_396),
.C(n_406),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_406),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_401),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_397),
.B(n_402),
.C(n_403),
.Y(n_437)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_403),
.Y(n_401)
);

INVx6_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_411),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_410),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_408),
.B(n_410),
.C(n_411),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_416),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_415),
.B(n_416),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_417),
.B(n_434),
.C(n_442),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_419),
.A2(n_434),
.B1(n_442),
.B2(n_443),
.Y(n_418)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_419),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_420),
.A2(n_421),
.B1(n_422),
.B2(n_433),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_420),
.B(n_423),
.C(n_424),
.Y(n_447)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_422),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_432),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_429),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_426),
.B(n_429),
.C(n_432),
.Y(n_456)
);

INVx8_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx6_ASAP7_75t_SL g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_434),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_436),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_435),
.B(n_437),
.C(n_438),
.Y(n_454)
);

BUFx24_ASAP7_75t_SL g485 ( 
.A(n_435),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_438),
.Y(n_436)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_446),
.B(n_460),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_446),
.B(n_460),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_447),
.B(n_449),
.C(n_452),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_452),
.Y(n_448)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_450),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_453),
.A2(n_454),
.B1(n_455),
.B2(n_459),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_453),
.B(n_456),
.C(n_457),
.Y(n_464)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_455),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_SL g455 ( 
.A(n_456),
.B(n_457),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_463),
.B(n_471),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_463),
.B(n_471),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_465),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_466),
.C(n_469),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_469),
.Y(n_465)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_475),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_474),
.B(n_475),
.Y(n_477)
);

BUFx24_ASAP7_75t_SL g484 ( 
.A(n_474),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx6_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx13_ASAP7_75t_L g482 ( 
.A(n_479),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_483),
.Y(n_480)
);

BUFx12f_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);


endmodule