module fake_jpeg_11658_n_179 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_179);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_32),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx6f_ASAP7_75t_SL g54 ( 
.A(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_18),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_3),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_34),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_37),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_22),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_5),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_15),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_61),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_81),
.Y(n_99)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_75),
.B(n_0),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_1),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_83),
.B(n_59),
.Y(n_89)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

CKINVDCx6p67_ASAP7_75t_R g94 ( 
.A(n_85),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_84),
.A2(n_77),
.B1(n_63),
.B2(n_73),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_90),
.B1(n_91),
.B2(n_62),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_53),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_63),
.B1(n_74),
.B2(n_56),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_80),
.A2(n_73),
.B1(n_62),
.B2(n_74),
.Y(n_91)
);

BUFx4f_ASAP7_75t_SL g92 ( 
.A(n_86),
.Y(n_92)
);

BUFx8_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_81),
.B(n_60),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_95),
.B(n_58),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_60),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_96),
.B(n_65),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_101),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_102),
.B(n_26),
.Y(n_139)
);

AND2x4_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_76),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_103),
.A2(n_14),
.B(n_16),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_82),
.C(n_71),
.Y(n_104)
);

FAx1_ASAP7_75t_SL g132 ( 
.A(n_104),
.B(n_11),
.CI(n_12),
.CON(n_132),
.SN(n_132)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_105),
.B(n_114),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_100),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_108),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_57),
.B1(n_62),
.B2(n_85),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_116),
.B1(n_4),
.B2(n_5),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_55),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_91),
.A2(n_97),
.B1(n_98),
.B2(n_56),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_110),
.A2(n_40),
.B1(n_44),
.B2(n_46),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_70),
.B1(n_58),
.B2(n_55),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_57),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_115),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_88),
.Y(n_113)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_69),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_70),
.B1(n_67),
.B2(n_66),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_2),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_118),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_2),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_4),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_28),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_138),
.B1(n_139),
.B2(n_127),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_108),
.A2(n_6),
.B(n_7),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_136),
.B(n_140),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_6),
.B(n_7),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_124),
.B(n_125),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_8),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_133),
.B1(n_141),
.B2(n_140),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_111),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_131),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_130),
.B(n_134),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_10),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_139),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_13),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_17),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_137),
.B(n_109),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_113),
.A2(n_20),
.B1(n_21),
.B2(n_24),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_109),
.A2(n_29),
.B1(n_30),
.B2(n_36),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_122),
.B(n_133),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_149),
.Y(n_160)
);

AO21x2_ASAP7_75t_L g145 ( 
.A1(n_136),
.A2(n_109),
.B(n_48),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_145),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_146),
.B(n_152),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_151),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_135),
.B(n_47),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_141),
.A2(n_49),
.B(n_51),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_126),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_153),
.B(n_157),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_132),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_158),
.Y(n_165)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_126),
.C(n_105),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_156),
.B(n_155),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_161),
.B(n_152),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_167),
.B(n_168),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_155),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_SL g169 ( 
.A1(n_163),
.A2(n_148),
.B(n_142),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_170),
.Y(n_171)
);

OA21x2_ASAP7_75t_SL g170 ( 
.A1(n_165),
.A2(n_143),
.B(n_144),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_160),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_160),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_171),
.B(n_162),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_159),
.B(n_166),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_163),
.B(n_164),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_169),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_145),
.Y(n_179)
);


endmodule