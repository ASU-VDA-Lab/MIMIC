module real_jpeg_23069_n_16 (n_5, n_4, n_8, n_0, n_12, n_351, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_351;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_2),
.A2(n_70),
.B1(n_72),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_2),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_2),
.A2(n_75),
.B1(n_88),
.B2(n_92),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_75),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_75),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_4),
.A2(n_92),
.B(n_94),
.Y(n_91)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_4),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_4),
.B(n_83),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g170 ( 
.A1(n_4),
.A2(n_35),
.B1(n_36),
.B2(n_96),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_4),
.B(n_30),
.C(n_31),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_4),
.B(n_73),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_4),
.A2(n_45),
.B1(n_198),
.B2(n_203),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_5),
.A2(n_70),
.B1(n_72),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_5),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_77),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_77),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_5),
.A2(n_77),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

INVx8_ASAP7_75t_SL g84 ( 
.A(n_6),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_7),
.A2(n_87),
.B1(n_88),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_7),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_7),
.A2(n_70),
.B1(n_72),
.B2(n_100),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_100),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_100),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_51),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_8),
.A2(n_51),
.B1(n_70),
.B2(n_72),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_8),
.A2(n_51),
.B1(n_89),
.B2(n_239),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_37),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_9),
.A2(n_37),
.B1(n_70),
.B2(n_72),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_9),
.A2(n_37),
.B1(n_88),
.B2(n_240),
.Y(n_303)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_11),
.A2(n_35),
.B1(n_36),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_43),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_11),
.A2(n_43),
.B1(n_70),
.B2(n_72),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_11),
.A2(n_43),
.B1(n_88),
.B2(n_89),
.Y(n_290)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_12),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_14),
.A2(n_35),
.B1(n_36),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_14),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_14),
.A2(n_62),
.B1(n_70),
.B2(n_72),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_62),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_14),
.A2(n_62),
.B1(n_88),
.B2(n_92),
.Y(n_265)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_15),
.Y(n_184)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_15),
.Y(n_203)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_344),
.C(n_348),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_342),
.B(n_347),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_332),
.B(n_341),
.Y(n_18)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_298),
.A3(n_327),
.B1(n_330),
.B2(n_331),
.C(n_351),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_274),
.B(n_297),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_250),
.B(n_273),
.Y(n_21)
);

O2A1O1Ixp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_134),
.B(n_222),
.C(n_249),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_119),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_24),
.B(n_119),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_103),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_58),
.B1(n_101),
.B2(n_102),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_26),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_26),
.B(n_102),
.C(n_103),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_44),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_27),
.B(n_44),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_34),
.B(n_38),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_28),
.B(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_28),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_28),
.B(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_28),
.B(n_96),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_28),
.A2(n_163),
.B(n_314),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_29),
.B(n_205),
.Y(n_204)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_34),
.Y(n_231)
);

AO22x1_ASAP7_75t_L g73 ( 
.A1(n_35),
.A2(n_36),
.B1(n_68),
.B2(n_69),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_35),
.B(n_68),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

OAI32xp33_ASAP7_75t_L g141 ( 
.A1(n_36),
.A2(n_69),
.A3(n_72),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_36),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_38),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_41),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_61),
.B(n_63),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_39),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_39),
.A2(n_151),
.B(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_39),
.A2(n_150),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_39),
.A2(n_149),
.B1(n_150),
.B2(n_171),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_39),
.A2(n_150),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_39),
.A2(n_63),
.B(n_232),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_39),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_49),
.B(n_52),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_45),
.A2(n_52),
.B(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_45),
.A2(n_181),
.B(n_182),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_45),
.A2(n_189),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_45),
.A2(n_145),
.B(n_199),
.Y(n_258)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_46),
.A2(n_50),
.B1(n_56),
.B2(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_46),
.B(n_53),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_46),
.A2(n_188),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_47),
.Y(n_127)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_48),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_57),
.Y(n_207)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_64),
.C(n_79),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_59),
.A2(n_60),
.B1(n_64),
.B2(n_122),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_61),
.Y(n_163)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_74),
.B1(n_76),
.B2(n_78),
.Y(n_64)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_65),
.A2(n_76),
.B(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_65),
.A2(n_74),
.B1(n_78),
.B2(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_65),
.A2(n_243),
.B(n_244),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_65),
.A2(n_78),
.B1(n_268),
.B2(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_66),
.A2(n_73),
.B1(n_133),
.B2(n_142),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_66),
.B(n_245),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_66),
.A2(n_310),
.B(n_311),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_66),
.A2(n_73),
.B(n_111),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_73),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_70),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_72),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_70),
.A2(n_85),
.B(n_95),
.C(n_114),
.Y(n_113)
);

HAxp5_ASAP7_75t_SL g142 ( 
.A(n_70),
.B(n_96),
.CON(n_142),
.SN(n_142)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_84),
.C(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_73),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_73),
.B(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_78),
.A2(n_268),
.B(n_269),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_79),
.B(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_82),
.B1(n_91),
.B2(n_98),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_83),
.B1(n_99),
.B2(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_81),
.A2(n_83),
.B1(n_107),
.B2(n_238),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_81),
.A2(n_238),
.B(n_264),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_81),
.A2(n_288),
.B(n_289),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_81),
.B(n_305),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_81),
.A2(n_83),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_81),
.A2(n_289),
.B(n_321),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_81),
.A2(n_83),
.B(n_288),
.Y(n_348)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_86),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_82),
.B(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_82),
.B(n_290),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_82),
.A2(n_303),
.B(n_304),
.Y(n_302)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_84),
.A2(n_85),
.B1(n_87),
.B2(n_90),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_89),
.Y(n_90)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_92),
.Y(n_239)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_96),
.B(n_206),
.Y(n_205)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_97),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_112),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_108),
.B2(n_109),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_106),
.B(n_108),
.C(n_112),
.Y(n_247)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_110),
.B(n_269),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_111),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_115),
.B1(n_116),
.B2(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.C(n_125),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_120),
.B(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_123),
.B(n_125),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.C(n_131),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_129),
.B1(n_130),
.B2(n_156),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_126),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_128),
.B(n_182),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_217),
.B(n_221),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_165),
.B(n_216),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_152),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_139),
.B(n_152),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_147),
.C(n_148),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_140),
.B(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_144),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_144),
.Y(n_159)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_183),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_147),
.B(n_148),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_157),
.B2(n_158),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_153),
.B(n_160),
.C(n_164),
.Y(n_218)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_164),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_159),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_162),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_211),
.B(n_215),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_185),
.B(n_210),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_174),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_168),
.B(n_174),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_172),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_180),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_179),
.C(n_180),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

AOI21xp33_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_194),
.B(n_209),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_193),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_193),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_201),
.B(n_208),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_196),
.B(n_197),
.Y(n_208)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_212),
.B(n_213),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_218),
.B(n_219),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_224),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_247),
.B2(n_248),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_234),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_234),
.C(n_248),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_230),
.B2(n_233),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_233),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_230),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_246),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_241),
.B2(n_242),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_237),
.B(n_241),
.C(n_246),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_244),
.Y(n_311)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_247),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_251),
.B(n_252),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_272),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_259),
.B1(n_270),
.B2(n_271),
.Y(n_253)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_254),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_271),
.C(n_272),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_257),
.B2(n_258),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_256),
.B(n_257),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_257),
.A2(n_258),
.B1(n_287),
.B2(n_291),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_257),
.A2(n_291),
.B(n_292),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_260),
.B(n_263),
.C(n_266),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_266),
.B2(n_267),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_264),
.Y(n_345)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_275),
.B(n_276),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_295),
.B2(n_296),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_285),
.B1(n_293),
.B2(n_294),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_279),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_279),
.B(n_294),
.C(n_296),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_282),
.B(n_284),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_282),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_283),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_300),
.C(n_315),
.Y(n_299)
);

FAx1_ASAP7_75t_SL g329 ( 
.A(n_284),
.B(n_300),
.CI(n_315),
.CON(n_329),
.SN(n_329)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_285),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_292),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_287),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_290),
.Y(n_305)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_295),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_316),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_299),
.B(n_316),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_306),
.B2(n_307),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_301),
.A2(n_302),
.B1(n_318),
.B2(n_325),
.Y(n_317)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_302),
.B(n_309),
.C(n_312),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_302),
.B(n_325),
.C(n_326),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_303),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_304),
.B(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_312),
.B2(n_313),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_312),
.A2(n_313),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_313),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_313),
.B(n_319),
.C(n_323),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_326),
.Y(n_316)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_318),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_322),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_328),
.B(n_329),
.Y(n_330)
);

BUFx24_ASAP7_75t_SL g349 ( 
.A(n_329),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_333),
.B(n_334),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_340),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_336),
.A2(n_337),
.B1(n_338),
.B2(n_339),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_336),
.B(n_339),
.C(n_340),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_337),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_339),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_346),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_344),
.B(n_346),
.Y(n_347)
);


endmodule