module real_jpeg_6020_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_2),
.A2(n_89),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_2),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_2),
.A2(n_116),
.B1(n_188),
.B2(n_224),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_2),
.A2(n_188),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_2),
.A2(n_22),
.B1(n_188),
.B2(n_353),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_3),
.A2(n_70),
.B1(n_71),
.B2(n_73),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_3),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_3),
.A2(n_70),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_3),
.A2(n_70),
.B1(n_168),
.B2(n_170),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_3),
.A2(n_70),
.B1(n_107),
.B2(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_4),
.A2(n_37),
.B1(n_41),
.B2(n_42),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_4),
.A2(n_41),
.B1(n_112),
.B2(n_116),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_4),
.A2(n_41),
.B1(n_243),
.B2(n_245),
.Y(n_242)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_5),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_6),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_6),
.Y(n_258)
);

BUFx5_ASAP7_75t_L g368 ( 
.A(n_6),
.Y(n_368)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_7),
.Y(n_86)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_7),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_7),
.Y(n_240)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_8),
.Y(n_97)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_9),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_9),
.Y(n_90)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_9),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_9),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_9),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_10),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_10),
.A2(n_33),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_10),
.A2(n_33),
.B1(n_178),
.B2(n_180),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_10),
.B(n_91),
.Y(n_253)
);

O2A1O1Ixp33_ASAP7_75t_L g313 ( 
.A1(n_10),
.A2(n_120),
.B(n_314),
.C(n_321),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_10),
.B(n_343),
.C(n_344),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_10),
.B(n_118),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_10),
.B(n_258),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_10),
.B(n_58),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g343 ( 
.A(n_11),
.Y(n_343)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_211),
.B1(n_409),
.B2(n_410),
.Y(n_13)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_14),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_209),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_189),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_16),
.B(n_189),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_108),
.C(n_157),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_17),
.A2(n_108),
.B1(n_109),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_17),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_75),
.B2(n_76),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_18),
.A2(n_77),
.B(n_79),
.Y(n_208)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_35),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_20),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_20),
.A2(n_35),
.B1(n_77),
.B2(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_20),
.B(n_313),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_20),
.A2(n_77),
.B1(n_313),
.B2(n_392),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_27),
.B(n_29),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_21),
.B(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_21),
.B(n_29),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_21),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_21),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_23),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_24),
.Y(n_345)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_29),
.Y(n_164)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_32),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_33),
.A2(n_83),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_33),
.B(n_106),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g314 ( 
.A1(n_33),
.A2(n_315),
.B(n_318),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_35),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_47),
.B(n_68),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_36),
.A2(n_153),
.B(n_155),
.Y(n_172)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_39),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_39),
.Y(n_151)
);

INVx6_ASAP7_75t_L g320 ( 
.A(n_39),
.Y(n_320)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_40),
.Y(n_123)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_40),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_40),
.Y(n_341)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_47),
.A2(n_148),
.B(n_153),
.Y(n_203)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_48),
.B(n_69),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_48),
.B(n_149),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_48),
.B(n_328),
.Y(n_327)
);

NOR2x1_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_58),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_52),
.B1(n_54),
.B2(n_57),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AO22x2_ASAP7_75t_L g58 ( 
.A1(n_55),
.A2(n_59),
.B1(n_61),
.B2(n_65),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_58),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_58),
.B(n_328),
.Y(n_347)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_64),
.Y(n_169)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_67),
.Y(n_171)
);

AND2x2_ASAP7_75t_SL g265 ( 
.A(n_68),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_68),
.B(n_327),
.Y(n_356)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_102),
.B(n_103),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_81),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_81),
.B(n_104),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_81),
.B(n_196),
.Y(n_285)
);

NOR2x1_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_91),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_85),
.B1(n_87),
.B2(n_89),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_86),
.Y(n_230)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_90),
.Y(n_198)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_91),
.B(n_104),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_91),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_91),
.B(n_186),
.Y(n_218)
);

AO22x2_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_94),
.B1(n_98),
.B2(n_100),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_97),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_97),
.Y(n_179)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_99),
.Y(n_237)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVxp33_ASAP7_75t_L g234 ( 
.A(n_105),
.Y(n_234)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_146),
.B(n_156),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_110),
.B(n_146),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_118),
.B(n_129),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_111),
.A2(n_176),
.B(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_115),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_115),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_115),
.Y(n_323)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_118),
.B(n_140),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_118),
.B(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_118),
.A2(n_176),
.B(n_177),
.Y(n_283)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_119),
.B(n_274),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_122),
.B1(n_124),
.B2(n_125),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

INVx5_ASAP7_75t_L g329 ( 
.A(n_122),
.Y(n_329)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_129),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_139),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_130),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_134),
.B1(n_136),
.B2(n_138),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_133),
.Y(n_317)
);

AOI32xp33_ASAP7_75t_L g229 ( 
.A1(n_134),
.A2(n_230),
.A3(n_231),
.B1(n_234),
.B2(n_235),
.Y(n_229)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_141),
.Y(n_225)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_154),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_147),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_153),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

INVxp67_ASAP7_75t_SL g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_155),
.B(n_347),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_156),
.A2(n_191),
.B1(n_192),
.B2(n_207),
.Y(n_190)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_156),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_157),
.B(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_173),
.C(n_183),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_158),
.A2(n_159),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_172),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_160),
.B(n_172),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_161),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_163),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_165),
.B(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_166),
.A2(n_242),
.B(n_247),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_167),
.B(n_257),
.Y(n_256)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_169),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_169),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_173),
.B(n_183),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_174),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_175),
.B(n_222),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_176),
.B(n_223),
.Y(n_251)
);

INVxp67_ASAP7_75t_SL g274 ( 
.A(n_177),
.Y(n_274)
);

INVx6_ASAP7_75t_SL g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_185),
.B(n_195),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_208),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_200),
.B2(n_201),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_199),
.Y(n_194)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_199),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_202),
.A2(n_203),
.B1(n_220),
.B2(n_226),
.Y(n_219)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_203),
.B(n_217),
.C(n_220),
.Y(n_261)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_211),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_401),
.Y(n_211)
);

NAND3xp33_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_289),
.C(n_303),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_275),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_259),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_215),
.B(n_259),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_227),
.C(n_249),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_216),
.B(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_218),
.B(n_285),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_220),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_227),
.A2(n_228),
.B1(n_249),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_241),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_229),
.B(n_241),
.Y(n_268)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

NAND2xp33_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_242),
.A2(n_256),
.B(n_264),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx8_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_249),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.C(n_254),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_250),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_272),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_254),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_255),
.B(n_366),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_256),
.B(n_351),
.Y(n_379)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_267),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_262),
.C(n_267),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_265),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_266),
.B(n_347),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_270),
.C(n_271),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_275),
.A2(n_404),
.B(n_405),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_288),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_276),
.B(n_288),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_279),
.C(n_280),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_284),
.C(n_286),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_286),
.B2(n_287),
.Y(n_282)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_283),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_284),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_301),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_290),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_298),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_291),
.B(n_302),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_291),
.B(n_302),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_291),
.B(n_298),
.Y(n_408)
);

FAx1_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_295),
.CI(n_297),
.CON(n_291),
.SN(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_301),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_333),
.B(n_400),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_308),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_305),
.B(n_308),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_312),
.C(n_324),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_309),
.B(n_396),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_312),
.A2(n_324),
.B1(n_325),
.B2(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_312),
.Y(n_397)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_313),
.Y(n_392)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx8_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx3_ASAP7_75t_SL g318 ( 
.A(n_319),
.Y(n_318)
);

INVx8_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

BUFx12f_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_394),
.B(n_399),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_335),
.A2(n_384),
.B(n_393),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_360),
.B(n_383),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_348),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_337),
.B(n_348),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_346),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_338),
.A2(n_339),
.B1(n_346),
.B2(n_363),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_342),
.Y(n_339)
);

INVx5_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_346),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_355),
.Y(n_348)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_349),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_352),
.B(n_367),
.Y(n_366)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_356),
.A2(n_357),
.B1(n_358),
.B2(n_359),
.Y(n_355)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_356),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_357),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_357),
.B(n_358),
.C(n_386),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_361),
.A2(n_369),
.B(n_382),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_362),
.B(n_364),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_362),
.B(n_364),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_370),
.A2(n_378),
.B(n_381),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_377),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_376),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx6_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_379),
.B(n_380),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_387),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_385),
.B(n_387),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_391),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_390),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_389),
.B(n_390),
.C(n_391),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_395),
.B(n_398),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_395),
.B(n_398),
.Y(n_399)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g401 ( 
.A1(n_402),
.A2(n_403),
.B(n_406),
.C(n_407),
.D(n_408),
.Y(n_401)
);


endmodule