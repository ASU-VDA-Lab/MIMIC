module fake_jpeg_31183_n_533 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_533);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_533;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_412;
wire n_249;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_16),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_55),
.Y(n_132)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_56),
.B(n_82),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_59),
.Y(n_126)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_64),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_42),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_66),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_20),
.B(n_7),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_67),
.B(n_71),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_69),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_70),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_20),
.B(n_31),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_72),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

NAND2xp33_ASAP7_75t_SL g74 ( 
.A(n_17),
.B(n_8),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_74),
.B(n_79),
.Y(n_158)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_23),
.B(n_6),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

BUFx4f_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_23),
.B(n_10),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_83),
.Y(n_161)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

HAxp5_ASAP7_75t_SL g85 ( 
.A(n_28),
.B(n_10),
.CON(n_85),
.SN(n_85)
);

AOI21xp33_ASAP7_75t_SL g152 ( 
.A1(n_85),
.A2(n_0),
.B(n_1),
.Y(n_152)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_91),
.Y(n_163)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_95),
.Y(n_109)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_31),
.B(n_40),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_94),
.B(n_49),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_38),
.B(n_5),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_48),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_25),
.Y(n_101)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_35),
.Y(n_102)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_18),
.Y(n_103)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_32),
.Y(n_104)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_104),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_43),
.B1(n_51),
.B2(n_49),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_111),
.A2(n_39),
.B1(n_28),
.B2(n_46),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_117),
.B(n_120),
.Y(n_215)
);

BUFx12f_ASAP7_75t_SL g120 ( 
.A(n_85),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_122),
.B(n_149),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_96),
.A2(n_25),
.B1(n_51),
.B2(n_48),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_153),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_95),
.A2(n_30),
.B1(n_52),
.B2(n_41),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_140),
.A2(n_144),
.B1(n_154),
.B2(n_157),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_95),
.A2(n_30),
.B1(n_52),
.B2(n_41),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_79),
.B(n_43),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_148),
.B(n_150),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_56),
.B(n_40),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_69),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_151),
.B(n_164),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_L g205 ( 
.A1(n_152),
.A2(n_39),
.B(n_27),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_54),
.A2(n_25),
.B1(n_38),
.B2(n_52),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_86),
.A2(n_41),
.B1(n_52),
.B2(n_72),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_58),
.Y(n_156)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_72),
.A2(n_41),
.B1(n_46),
.B2(n_50),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_80),
.A2(n_50),
.B1(n_46),
.B2(n_29),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_165),
.A2(n_27),
.B1(n_29),
.B2(n_50),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_59),
.B1(n_100),
.B2(n_99),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_167),
.A2(n_176),
.B1(n_185),
.B2(n_206),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_109),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_169),
.B(n_171),
.Y(n_228)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_170),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_116),
.A2(n_102),
.B1(n_97),
.B2(n_87),
.Y(n_172)
);

OA22x2_ASAP7_75t_L g223 ( 
.A1(n_172),
.A2(n_204),
.B1(n_208),
.B2(n_214),
.Y(n_223)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_174),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_34),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_175),
.B(n_106),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_112),
.A2(n_107),
.B1(n_110),
.B2(n_134),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_177),
.Y(n_252)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_108),
.Y(n_178)
);

INVx11_ASAP7_75t_L g249 ( 
.A(n_178),
.Y(n_249)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_179),
.Y(n_253)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_115),
.Y(n_180)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_180),
.Y(n_259)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_181),
.Y(n_230)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_182),
.Y(n_260)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_183),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_121),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_184),
.B(n_189),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_123),
.A2(n_130),
.B1(n_116),
.B2(n_159),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_186),
.Y(n_250)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_118),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_188),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_113),
.Y(n_191)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_142),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_193),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_196),
.Y(n_233)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_113),
.Y(n_195)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_195),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_34),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_108),
.Y(n_197)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_197),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_121),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_200),
.Y(n_239)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_155),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_129),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_142),
.Y(n_201)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_201),
.Y(n_247)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_124),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_202),
.Y(n_264)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_135),
.Y(n_203)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_203),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_159),
.A2(n_57),
.B1(n_83),
.B2(n_62),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_215),
.Y(n_229)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_138),
.Y(n_207)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_207),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_119),
.A2(n_63),
.B1(n_73),
.B2(n_70),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_132),
.Y(n_209)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_209),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_158),
.B(n_18),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_211),
.Y(n_243)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_135),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_129),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_212),
.B(n_213),
.Y(n_255)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_138),
.Y(n_213)
);

OA22x2_ASAP7_75t_L g214 ( 
.A1(n_157),
.A2(n_64),
.B1(n_22),
.B2(n_37),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_165),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_216),
.B(n_217),
.Y(n_256)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_119),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_218),
.A2(n_221),
.B1(n_161),
.B2(n_137),
.Y(n_226)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_163),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_219),
.Y(n_225)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_124),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_220),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_131),
.A2(n_80),
.B1(n_65),
.B2(n_37),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_226),
.A2(n_251),
.B1(n_262),
.B2(n_224),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_229),
.A2(n_243),
.B(n_257),
.Y(n_277)
);

AO22x1_ASAP7_75t_L g234 ( 
.A1(n_192),
.A2(n_214),
.B1(n_206),
.B2(n_205),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_234),
.B(n_257),
.Y(n_300)
);

O2A1O1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_214),
.A2(n_149),
.B(n_154),
.C(n_140),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_235),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_261),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_173),
.A2(n_161),
.B1(n_147),
.B2(n_128),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_245),
.A2(n_254),
.B1(n_167),
.B2(n_197),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_192),
.A2(n_127),
.B1(n_136),
.B2(n_139),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_221),
.A2(n_144),
.B1(n_147),
.B2(n_128),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_215),
.B(n_127),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_168),
.B(n_126),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_217),
.A2(n_105),
.B1(n_22),
.B2(n_126),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_234),
.A2(n_219),
.B(n_176),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_265),
.A2(n_270),
.B(n_264),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_231),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_266),
.B(n_284),
.Y(n_307)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_261),
.Y(n_268)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_268),
.Y(n_308)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_239),
.Y(n_269)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_269),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_234),
.A2(n_185),
.B(n_170),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_254),
.A2(n_171),
.B1(n_178),
.B2(n_195),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_271),
.Y(n_333)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_239),
.Y(n_272)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_272),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_273),
.A2(n_279),
.B1(n_286),
.B2(n_287),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_228),
.B(n_190),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_274),
.B(n_278),
.Y(n_305)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_247),
.Y(n_275)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_275),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_228),
.A2(n_218),
.B1(n_208),
.B2(n_204),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_276),
.A2(n_223),
.B1(n_242),
.B2(n_235),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_277),
.B(n_295),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_240),
.B(n_187),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_238),
.A2(n_172),
.B1(n_191),
.B2(n_27),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_231),
.B(n_29),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_280),
.B(n_285),
.Y(n_323)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_247),
.Y(n_281)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_281),
.Y(n_336)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_246),
.Y(n_282)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_282),
.Y(n_329)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_248),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_283),
.Y(n_315)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_248),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_233),
.B(n_207),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_238),
.A2(n_213),
.B1(n_47),
.B2(n_32),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_223),
.A2(n_47),
.B1(n_32),
.B2(n_92),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_243),
.B(n_0),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_288),
.B(n_290),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_289),
.A2(n_297),
.B1(n_257),
.B2(n_224),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_256),
.B(n_1),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_256),
.B(n_1),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_291),
.B(n_293),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_233),
.B(n_255),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_255),
.B(n_229),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_294),
.B(n_301),
.Y(n_314)
);

MAJx2_ASAP7_75t_L g295 ( 
.A(n_229),
.B(n_2),
.C(n_3),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_223),
.A2(n_47),
.B1(n_3),
.B2(n_4),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_296),
.A2(n_223),
.B1(n_225),
.B2(n_241),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_235),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_230),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_299),
.Y(n_313)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_237),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_225),
.B(n_2),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_274),
.B(n_230),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_304),
.B(n_335),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_301),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_306),
.B(n_310),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_309),
.A2(n_311),
.B1(n_312),
.B2(n_326),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_280),
.Y(n_310)
);

OAI22x1_ASAP7_75t_SL g312 ( 
.A1(n_292),
.A2(n_270),
.B1(n_265),
.B2(n_296),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_267),
.B(n_263),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_316),
.B(n_300),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_266),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_317),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_244),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_319),
.B(n_320),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_269),
.B(n_272),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_267),
.B(n_241),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_321),
.B(n_288),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_322),
.A2(n_312),
.B1(n_334),
.B2(n_303),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_292),
.A2(n_223),
.B1(n_242),
.B2(n_250),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_290),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_327),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_328),
.A2(n_300),
.B(n_297),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_286),
.A2(n_259),
.B1(n_253),
.B2(n_237),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_330),
.A2(n_276),
.B1(n_268),
.B2(n_299),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_300),
.A2(n_263),
.B(n_222),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_334),
.A2(n_291),
.B(n_271),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_293),
.B(n_244),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_339),
.B(n_321),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_341),
.B(n_344),
.Y(n_387)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_331),
.Y(n_342)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_342),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_319),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_345),
.A2(n_348),
.B(n_349),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_329),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_346),
.Y(n_388)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_331),
.Y(n_347)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_347),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_328),
.A2(n_300),
.B(n_333),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_309),
.A2(n_289),
.B(n_294),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_320),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_350),
.B(n_351),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_307),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_325),
.B(n_316),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_352),
.B(n_366),
.C(n_323),
.Y(n_370)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_329),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g384 ( 
.A1(n_353),
.A2(n_250),
.B1(n_237),
.B2(n_282),
.Y(n_384)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_336),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_354),
.B(n_356),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_307),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_313),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_357),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_313),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_358),
.B(n_362),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_359),
.A2(n_363),
.B(n_314),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_361),
.A2(n_306),
.B1(n_324),
.B2(n_318),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_317),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_312),
.A2(n_287),
.B(n_277),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_322),
.A2(n_279),
.B1(n_273),
.B2(n_285),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_364),
.A2(n_369),
.B1(n_311),
.B2(n_303),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_335),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_365),
.B(n_367),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_325),
.B(n_278),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_336),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_326),
.A2(n_299),
.B1(n_284),
.B2(n_283),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_368),
.A2(n_308),
.B1(n_318),
.B2(n_324),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_370),
.B(n_373),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_352),
.B(n_316),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_371),
.B(n_385),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_366),
.B(n_314),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_377),
.B(n_399),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_379),
.A2(n_393),
.B(n_395),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_350),
.B(n_305),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_380),
.B(n_337),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_339),
.B(n_305),
.C(n_308),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_381),
.B(n_391),
.C(n_400),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_382),
.A2(n_390),
.B1(n_343),
.B2(n_358),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_384),
.B(n_361),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_338),
.B(n_323),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_386),
.A2(n_396),
.B1(n_368),
.B2(n_379),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_349),
.B(n_310),
.C(n_302),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_363),
.A2(n_359),
.B(n_340),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_355),
.A2(n_304),
.B1(n_327),
.B2(n_302),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_394),
.A2(n_342),
.B1(n_353),
.B2(n_275),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_340),
.A2(n_332),
.B(n_315),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_364),
.A2(n_369),
.B1(n_343),
.B2(n_355),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_338),
.B(n_332),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_397),
.B(n_398),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_360),
.B(n_295),
.Y(n_398)
);

XNOR2x1_ASAP7_75t_L g399 ( 
.A(n_348),
.B(n_295),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_360),
.B(n_330),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_357),
.B(n_315),
.C(n_281),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_401),
.B(n_365),
.C(n_337),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_402),
.A2(n_409),
.B1(n_395),
.B2(n_393),
.Y(n_435)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_403),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_376),
.A2(n_345),
.B(n_362),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_405),
.A2(n_383),
.B(n_386),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_406),
.B(n_417),
.C(n_429),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_378),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_407),
.Y(n_441)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_374),
.Y(n_408)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_408),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_410),
.A2(n_422),
.B1(n_400),
.B2(n_390),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_372),
.B(n_354),
.Y(n_411)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_411),
.Y(n_448)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_374),
.Y(n_412)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_412),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_397),
.B(n_232),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_413),
.Y(n_437)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_389),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_415),
.B(n_421),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_370),
.B(n_367),
.C(n_347),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_385),
.B(n_258),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_418),
.B(n_424),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_388),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_419),
.Y(n_444)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_392),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_388),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_423),
.B(n_426),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_387),
.B(n_258),
.Y(n_424)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_375),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_381),
.B(n_236),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_428),
.B(n_401),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_371),
.B(n_253),
.C(n_259),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_420),
.B(n_391),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_432),
.B(n_436),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_434),
.A2(n_438),
.B1(n_446),
.B2(n_402),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_435),
.B(n_440),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_420),
.B(n_377),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_410),
.A2(n_376),
.B1(n_399),
.B2(n_396),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_443),
.A2(n_445),
.B(n_450),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_414),
.A2(n_373),
.B(n_398),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_415),
.A2(n_346),
.B1(n_250),
.B2(n_227),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_407),
.B(n_236),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_449),
.B(n_411),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_414),
.A2(n_227),
.B(n_346),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_427),
.B(n_249),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_452),
.B(n_429),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_438),
.A2(n_405),
.B(n_412),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_453),
.B(n_451),
.Y(n_481)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_447),
.Y(n_454)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_454),
.Y(n_475)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_442),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_455),
.B(n_458),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_431),
.B(n_417),
.C(n_404),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_457),
.B(n_459),
.C(n_470),
.Y(n_473)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_442),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_431),
.B(n_404),
.C(n_406),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_430),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_460),
.B(n_466),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_461),
.B(n_465),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_463),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_448),
.A2(n_408),
.B1(n_421),
.B2(n_427),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_464),
.A2(n_468),
.B1(n_444),
.B2(n_437),
.Y(n_483)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_451),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_448),
.A2(n_425),
.B1(n_426),
.B2(n_423),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_441),
.B(n_419),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_469),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_432),
.B(n_416),
.C(n_425),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_441),
.B(n_416),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_471),
.B(n_249),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_456),
.B(n_433),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_474),
.B(n_483),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_457),
.B(n_436),
.C(n_434),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_479),
.B(n_480),
.C(n_484),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_459),
.B(n_452),
.C(n_443),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_481),
.B(n_469),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_465),
.B(n_445),
.Y(n_482)
);

XNOR2x1_ASAP7_75t_L g492 ( 
.A(n_482),
.B(n_471),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_470),
.B(n_450),
.C(n_439),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_456),
.A2(n_430),
.B1(n_446),
.B2(n_249),
.Y(n_485)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_485),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_462),
.B(n_246),
.C(n_252),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_487),
.B(n_468),
.C(n_463),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_488),
.B(n_2),
.Y(n_502)
);

CKINVDCx14_ASAP7_75t_R g505 ( 
.A(n_489),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_492),
.B(n_480),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_477),
.A2(n_461),
.B1(n_460),
.B2(n_467),
.Y(n_493)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_493),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_494),
.B(n_502),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_473),
.A2(n_453),
.B(n_467),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_495),
.A2(n_499),
.B(n_478),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_473),
.B(n_464),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_496),
.B(n_497),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_486),
.B(n_462),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_484),
.A2(n_252),
.B(n_260),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_472),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_500),
.A2(n_483),
.B1(n_488),
.B2(n_481),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_476),
.B(n_260),
.C(n_5),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_501),
.B(n_503),
.C(n_475),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_476),
.B(n_5),
.C(n_11),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_506),
.B(n_508),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_509),
.B(n_511),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_491),
.B(n_479),
.C(n_494),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_510),
.B(n_492),
.C(n_493),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_491),
.B(n_487),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_512),
.B(n_11),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_498),
.A2(n_482),
.B1(n_12),
.B2(n_13),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_513),
.B(n_16),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_515),
.A2(n_514),
.B(n_507),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_510),
.B(n_490),
.C(n_501),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_517),
.A2(n_518),
.B(n_520),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_512),
.B(n_503),
.C(n_12),
.Y(n_518)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_519),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_521),
.B(n_505),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_522),
.B(n_508),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_523),
.B(n_515),
.C(n_516),
.Y(n_526)
);

AOI21xp33_ASAP7_75t_L g528 ( 
.A1(n_526),
.A2(n_527),
.B(n_504),
.Y(n_528)
);

AOI31xp67_ASAP7_75t_SL g529 ( 
.A1(n_528),
.A2(n_504),
.A3(n_524),
.B(n_509),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_529),
.B(n_525),
.C(n_12),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_530),
.B(n_11),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_531),
.B(n_13),
.C(n_15),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_16),
.Y(n_533)
);


endmodule