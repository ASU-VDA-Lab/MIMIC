module real_jpeg_7516_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_288;
wire n_78;
wire n_83;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_0),
.B(n_35),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_0),
.B(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_0),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_0),
.B(n_292),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_0),
.B(n_327),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_0),
.B(n_343),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_0),
.B(n_408),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_1),
.Y(n_162)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_1),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g262 ( 
.A(n_1),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_1),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_1),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_1),
.Y(n_327)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_2),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_2),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_2),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_3),
.B(n_169),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_3),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_3),
.B(n_307),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_3),
.B(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_3),
.B(n_352),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_3),
.B(n_386),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_3),
.B(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_4),
.B(n_97),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_4),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_4),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_4),
.B(n_310),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_4),
.B(n_323),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_4),
.B(n_189),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_4),
.B(n_380),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_4),
.B(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_5),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_5),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_5),
.B(n_142),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_5),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_5),
.B(n_97),
.Y(n_217)
);

AND2x2_ASAP7_75t_SL g283 ( 
.A(n_5),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_5),
.B(n_310),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_5),
.B(n_414),
.Y(n_413)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_6),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_6),
.Y(n_237)
);

BUFx5_ASAP7_75t_L g399 ( 
.A(n_6),
.Y(n_399)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_8),
.Y(n_189)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_8),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_8),
.Y(n_334)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_10),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_10),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_10),
.Y(n_203)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_12),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_12),
.B(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_12),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_12),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_12),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_12),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_12),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_12),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_13),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_13),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_13),
.B(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_13),
.B(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_13),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_13),
.B(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_13),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_14),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_14),
.B(n_191),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_14),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_14),
.B(n_74),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_14),
.B(n_288),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_14),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_14),
.B(n_372),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_14),
.B(n_189),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_15),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_15),
.B(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_15),
.B(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_15),
.B(n_288),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_15),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_15),
.B(n_383),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_15),
.B(n_399),
.Y(n_398)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_17),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_18),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_18),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_18),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_18),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_18),
.B(n_134),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_18),
.B(n_272),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_18),
.B(n_284),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_18),
.B(n_417),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_19),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_19),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_19),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_19),
.B(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g183 ( 
.A(n_19),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_19),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_19),
.B(n_224),
.Y(n_223)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_119),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_117),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_100),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_28),
.B(n_100),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_80),
.C(n_81),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_29),
.A2(n_30),
.B1(n_525),
.B2(n_526),
.Y(n_524)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_54),
.C(n_69),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_31),
.A2(n_32),
.B1(n_504),
.B2(n_506),
.Y(n_503)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_42),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_37),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_34),
.B(n_37),
.C(n_42),
.Y(n_80)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_36),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_40),
.Y(n_294)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_40),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_40),
.Y(n_397)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_41),
.Y(n_171)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_41),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_41),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_47),
.C(n_52),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_43),
.B(n_494),
.Y(n_493)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_47),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_494)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_50),
.Y(n_356)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_51),
.Y(n_136)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_51),
.Y(n_149)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_51),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_51),
.Y(n_387)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_51),
.Y(n_405)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_54),
.A2(n_69),
.B1(n_70),
.B2(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_54),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_60),
.C(n_64),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_SL g499 ( 
.A(n_55),
.B(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_57),
.Y(n_269)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_60),
.A2(n_61),
.B1(n_201),
.B2(n_204),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_60),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_500)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_61),
.B(n_197),
.C(n_201),
.Y(n_501)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_63),
.Y(n_285)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_63),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_65),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_77),
.C(n_79),
.Y(n_89)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_68),
.Y(n_225)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_68),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_68),
.Y(n_353)
);

BUFx5_ASAP7_75t_L g409 ( 
.A(n_68),
.Y(n_409)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_75),
.B1(n_76),
.B2(n_79),
.Y(n_70)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_78),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_93),
.C(n_96),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g526 ( 
.A(n_80),
.B(n_81),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_90),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_89),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_89),
.C(n_90),
.Y(n_116)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_88),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_96),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_92),
.A2(n_93),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_116),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_114),
.B2(n_115),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_102),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_107),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_113),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_523),
.B(n_528),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_487),
.B(n_520),
.Y(n_120)
);

OAI21x1_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_295),
.B(n_486),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_247),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_123),
.B(n_247),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_194),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_124),
.B(n_195),
.C(n_228),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_164),
.C(n_175),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_125),
.B(n_250),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_138),
.C(n_150),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_126),
.B(n_472),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_132),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_127),
.B(n_133),
.C(n_137),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_131),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_131),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.Y(n_132)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_138),
.A2(n_139),
.B1(n_150),
.B2(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.C(n_146),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_140),
.B(n_146),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_141),
.B(n_462),
.Y(n_461)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_148),
.B(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_150),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_155),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_151),
.B(n_156),
.C(n_161),
.Y(n_244)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_160),
.B1(n_161),
.B2(n_163),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_156),
.Y(n_163)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx8_ASAP7_75t_L g372 ( 
.A(n_158),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_159),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_160),
.B(n_201),
.C(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_160),
.A2(n_161),
.B1(n_201),
.B2(n_204),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_162),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_164),
.B(n_175),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_174),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.Y(n_165)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_170),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_170),
.B(n_172),
.C(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_170),
.A2(n_173),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

INVx6_ASAP7_75t_L g265 ( 
.A(n_171),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_173),
.B(n_233),
.C(n_240),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_174),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_188),
.C(n_190),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_176),
.B(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.C(n_183),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_177),
.B(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_179),
.B(n_183),
.Y(n_259)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_182),
.Y(n_308)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_188),
.B(n_190),
.Y(n_277)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_228),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_205),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_196),
.B(n_206),
.C(n_227),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_201),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx8_ASAP7_75t_L g272 ( 
.A(n_203),
.Y(n_272)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_203),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_216),
.B1(n_226),
.B2(n_227),
.Y(n_205)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.C(n_212),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_207),
.B(n_212),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_217),
.B(n_219),
.C(n_223),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_223),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_241),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_230),
.B(n_232),
.C(n_241),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_238),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_234),
.B(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

INVx3_ASAP7_75t_SL g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_239),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.C(n_245),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_245),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_251),
.C(n_254),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_249),
.B(n_252),
.Y(n_482)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_254),
.B(n_482),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_275),
.C(n_278),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_256),
.B(n_475),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_260),
.C(n_266),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_257),
.A2(n_258),
.B1(n_453),
.B2(n_454),
.Y(n_452)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_260),
.A2(n_261),
.B(n_263),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_260),
.B(n_266),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_263),
.Y(n_260)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_270),
.C(n_273),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_267),
.A2(n_268),
.B1(n_270),
.B2(n_271),
.Y(n_430)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_273),
.B(n_430),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_274),
.B(n_285),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g475 ( 
.A1(n_275),
.A2(n_276),
.B1(n_278),
.B2(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_278),
.Y(n_476)
);

MAJx2_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_290),
.C(n_291),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_280),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_280),
.B(n_464),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_283),
.C(n_286),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_281),
.B(n_442),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_283),
.A2(n_286),
.B1(n_287),
.B2(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_283),
.Y(n_443)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_290),
.B(n_291),
.Y(n_464)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx5_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

AOI21x1_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_480),
.B(n_485),
.Y(n_295)
);

OAI21x1_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_467),
.B(n_479),
.Y(n_296)
);

AOI21x1_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_449),
.B(n_466),
.Y(n_297)
);

OAI21x1_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_423),
.B(n_448),
.Y(n_298)
);

AOI21x1_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_391),
.B(n_422),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_360),
.B(n_390),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_338),
.B(n_359),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_317),
.B(n_337),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_313),
.B(n_316),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_311),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_311),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_309),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_314),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_309),
.Y(n_318)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_315),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_318),
.B(n_319),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_320),
.A2(n_321),
.B1(n_328),
.B2(n_329),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_320),
.B(n_331),
.C(n_335),
.Y(n_358)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_326),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_322),
.B(n_326),
.Y(n_349)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_330),
.A2(n_331),
.B1(n_335),
.B2(n_336),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_358),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_339),
.B(n_358),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_350),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_349),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_341),
.B(n_349),
.C(n_362),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_346),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_342),
.B(n_346),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_345),
.Y(n_415)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_350),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_354),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_351),
.B(n_376),
.C(n_377),
.Y(n_375)
);

INVx5_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_357),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_355),
.Y(n_376)
);

CKINVDCx14_ASAP7_75t_R g377 ( 
.A(n_357),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_363),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_361),
.B(n_363),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_374),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_364),
.B(n_375),
.C(n_378),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_365),
.B(n_367),
.C(n_368),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_369),
.A2(n_370),
.B1(n_371),
.B2(n_373),
.Y(n_368)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_369),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_370),
.B(n_373),
.Y(n_400)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_378),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_381),
.Y(n_378)
);

MAJx2_ASAP7_75t_L g420 ( 
.A(n_379),
.B(n_385),
.C(n_388),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_382),
.A2(n_385),
.B1(n_388),
.B2(n_389),
.Y(n_381)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_382),
.Y(n_388)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_385),
.Y(n_389)
);

INVx6_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_392),
.B(n_421),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_392),
.B(n_421),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_393),
.B(n_402),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_401),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_394),
.B(n_401),
.C(n_447),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_400),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_398),
.Y(n_395)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_396),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_398),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_400),
.B(n_437),
.C(n_438),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_402),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_410),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_403),
.B(n_412),
.C(n_419),
.Y(n_426)
);

BUFx24_ASAP7_75t_SL g530 ( 
.A(n_403),
.Y(n_530)
);

FAx1_ASAP7_75t_SL g403 ( 
.A(n_404),
.B(n_406),
.CI(n_407),
.CON(n_403),
.SN(n_403)
);

MAJx2_ASAP7_75t_L g434 ( 
.A(n_404),
.B(n_406),
.C(n_407),
.Y(n_434)
);

INVx3_ASAP7_75t_SL g408 ( 
.A(n_409),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_411),
.A2(n_412),
.B1(n_419),
.B2(n_420),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_416),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_413),
.B(n_416),
.Y(n_433)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx3_ASAP7_75t_SL g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_420),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_424),
.B(n_446),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_424),
.B(n_446),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_435),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_427),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_426),
.B(n_427),
.C(n_435),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_428),
.A2(n_429),
.B1(n_431),
.B2(n_432),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_428),
.B(n_458),
.C(n_459),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_434),
.Y(n_432)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_433),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_434),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_436),
.B(n_439),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_436),
.B(n_440),
.C(n_445),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_440),
.A2(n_441),
.B1(n_444),
.B2(n_445),
.Y(n_439)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_440),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_441),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_450),
.B(n_465),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_450),
.B(n_465),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_451),
.B(n_456),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_455),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_452),
.B(n_455),
.C(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_453),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_456),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_457),
.B(n_460),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_457),
.B(n_461),
.C(n_463),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_463),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_468),
.B(n_477),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_468),
.B(n_477),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_470),
.Y(n_468)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_469),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_474),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_471),
.B(n_474),
.C(n_484),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_481),
.B(n_483),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_481),
.B(n_483),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_515),
.Y(n_487)
);

OAI21xp33_ASAP7_75t_L g520 ( 
.A1(n_488),
.A2(n_521),
.B(n_522),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_489),
.B(n_508),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_489),
.B(n_508),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_490),
.A2(n_491),
.B1(n_497),
.B2(n_507),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_490),
.B(n_498),
.C(n_503),
.Y(n_527)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_493),
.C(n_495),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_SL g510 ( 
.A(n_492),
.B(n_511),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_493),
.A2(n_495),
.B1(n_496),
.B2(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_493),
.Y(n_512)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_497),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_503),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_501),
.C(n_502),
.Y(n_498)
);

FAx1_ASAP7_75t_SL g513 ( 
.A(n_499),
.B(n_501),
.CI(n_502),
.CON(n_513),
.SN(n_513)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_504),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_513),
.C(n_514),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_509),
.A2(n_510),
.B1(n_513),
.B2(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_513),
.Y(n_518)
);

BUFx24_ASAP7_75t_SL g531 ( 
.A(n_513),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_514),
.B(n_517),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_516),
.B(n_519),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_516),
.B(n_519),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_524),
.B(n_527),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_524),
.B(n_527),
.Y(n_528)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);


endmodule