module fake_netlist_1_935_n_38 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_38);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_30;
wire n_13;
wire n_26;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx3_ASAP7_75t_L g11 ( .A(n_9), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_10), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_4), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_7), .Y(n_16) );
AND2x4_ASAP7_75t_L g17 ( .A(n_5), .B(n_6), .Y(n_17) );
AOI22xp33_ASAP7_75t_SL g18 ( .A1(n_17), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_14), .B(n_0), .Y(n_19) );
AND2x4_ASAP7_75t_L g20 ( .A(n_11), .B(n_2), .Y(n_20) );
BUFx3_ASAP7_75t_L g21 ( .A(n_11), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_11), .B(n_3), .Y(n_22) );
AOI22xp33_ASAP7_75t_SL g23 ( .A1(n_20), .A2(n_12), .B1(n_17), .B2(n_16), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_21), .Y(n_24) );
INVx6_ASAP7_75t_L g25 ( .A(n_20), .Y(n_25) );
OA332x1_ASAP7_75t_L g26 ( .A1(n_23), .A2(n_18), .A3(n_19), .B1(n_14), .B2(n_15), .B3(n_16), .C1(n_13), .C2(n_17), .Y(n_26) );
AND2x2_ASAP7_75t_L g27 ( .A(n_25), .B(n_20), .Y(n_27) );
OAI22xp5_ASAP7_75t_L g28 ( .A1(n_25), .A2(n_19), .B1(n_21), .B2(n_22), .Y(n_28) );
INVx1_ASAP7_75t_SL g29 ( .A(n_27), .Y(n_29) );
NOR2xp67_ASAP7_75t_L g30 ( .A(n_28), .B(n_24), .Y(n_30) );
HB1xp67_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
OR2x2_ASAP7_75t_L g32 ( .A(n_30), .B(n_26), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_32), .Y(n_33) );
NAND2xp5_ASAP7_75t_L g34 ( .A(n_31), .B(n_26), .Y(n_34) );
OAI221xp5_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_30), .B1(n_15), .B2(n_13), .C(n_17), .Y(n_35) );
OAI22xp5_ASAP7_75t_L g36 ( .A1(n_33), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_36) );
INVx2_ASAP7_75t_L g37 ( .A(n_36), .Y(n_37) );
AOI22xp5_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_35), .B1(n_6), .B2(n_7), .Y(n_38) );
endmodule