module fake_jpeg_30159_n_441 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_441);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_441;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_332;
wire n_92;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_13),
.B(n_2),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_45),
.B(n_72),
.Y(n_96)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_48),
.Y(n_117)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_8),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_52),
.B(n_60),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_53),
.Y(n_130)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_55),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_8),
.Y(n_60)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_8),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_62),
.B(n_74),
.Y(n_100)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_23),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_19),
.B(n_9),
.Y(n_74)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_87),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_81),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_124)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_82),
.B(n_86),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_30),
.B(n_7),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_30),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_52),
.A2(n_19),
.B1(n_22),
.B2(n_39),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_99),
.A2(n_36),
.B1(n_41),
.B2(n_38),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_102),
.B(n_115),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_74),
.B(n_22),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_110),
.B(n_111),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_62),
.B(n_39),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_75),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_116),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_86),
.B(n_0),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_42),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_41),
.C(n_36),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_121),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_72),
.B(n_42),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_61),
.A2(n_30),
.B(n_25),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_126),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_53),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_132),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_46),
.B(n_38),
.Y(n_132)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_24),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_137),
.B(n_166),
.Y(n_182)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_138),
.Y(n_197)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_139),
.Y(n_192)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_140),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_149),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_144),
.Y(n_177)
);

BUFx12_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_146),
.Y(n_190)
);

BUFx8_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_147),
.Y(n_194)
);

BUFx8_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_152),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_100),
.B(n_41),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_85),
.B1(n_84),
.B2(n_83),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_153),
.A2(n_124),
.B1(n_131),
.B2(n_81),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_105),
.Y(n_154)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_94),
.Y(n_155)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_109),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_160),
.Y(n_179)
);

BUFx10_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_157),
.Y(n_187)
);

AND2x2_ASAP7_75t_SL g158 ( 
.A(n_115),
.B(n_80),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_135),
.C(n_114),
.Y(n_196)
);

INVx5_ASAP7_75t_SL g160 ( 
.A(n_109),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_104),
.B(n_30),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_163),
.Y(n_186)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_162),
.Y(n_200)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_119),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_91),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_165),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_96),
.B(n_30),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_91),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_168),
.Y(n_185)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_93),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_169),
.A2(n_172),
.B1(n_135),
.B2(n_114),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_98),
.B(n_27),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_27),
.Y(n_198)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_90),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_180),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_148),
.A2(n_115),
.B1(n_126),
.B2(n_123),
.Y(n_180)
);

INVx11_ASAP7_75t_L g224 ( 
.A(n_183),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_137),
.A2(n_124),
.B1(n_78),
.B2(n_134),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_188),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_145),
.A2(n_59),
.B1(n_58),
.B2(n_47),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_158),
.A2(n_97),
.B1(n_125),
.B2(n_65),
.Y(n_191)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_158),
.A2(n_97),
.B1(n_93),
.B2(n_103),
.Y(n_193)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_196),
.B(n_201),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_159),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_103),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_179),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_203),
.Y(n_238)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_204),
.Y(n_227)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_205),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_208),
.B(n_174),
.Y(n_234)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_178),
.Y(n_209)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_209),
.Y(n_239)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

CKINVDCx12_ASAP7_75t_R g211 ( 
.A(n_190),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_211),
.Y(n_245)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_190),
.Y(n_214)
);

INVxp33_ASAP7_75t_L g248 ( 
.A(n_214),
.Y(n_248)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_216),
.Y(n_249)
);

INVx4_ASAP7_75t_SL g217 ( 
.A(n_192),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_219),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_180),
.A2(n_171),
.B(n_150),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_218),
.A2(n_186),
.B(n_199),
.Y(n_231)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

INVx13_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_222),
.Y(n_233)
);

INVx13_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

AND2x6_ASAP7_75t_L g223 ( 
.A(n_182),
.B(n_171),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_223),
.A2(n_201),
.B(n_196),
.Y(n_229)
);

INVx13_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_187),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_206),
.A2(n_179),
.B(n_182),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_226),
.A2(n_156),
.B(n_200),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_229),
.B(n_234),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_231),
.B(n_247),
.Y(n_274)
);

O2A1O1Ixp33_ASAP7_75t_L g232 ( 
.A1(n_221),
.A2(n_187),
.B(n_183),
.C(n_176),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_206),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_184),
.C(n_186),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_237),
.C(n_181),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_207),
.A2(n_191),
.B1(n_173),
.B2(n_175),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_236),
.A2(n_243),
.B1(n_224),
.B2(n_177),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_188),
.C(n_199),
.Y(n_237)
);

AOI32xp33_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_173),
.A3(n_174),
.B1(n_193),
.B2(n_142),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_206),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_221),
.A2(n_198),
.B1(n_177),
.B2(n_168),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_244),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_181),
.Y(n_247)
);

AO22x1_ASAP7_75t_SL g250 ( 
.A1(n_240),
.A2(n_202),
.B1(n_210),
.B2(n_216),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_255),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_253),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g252 ( 
.A(n_229),
.B(n_202),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_252),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_233),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_233),
.Y(n_254)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_254),
.Y(n_284)
);

INVx6_ASAP7_75t_SL g255 ( 
.A(n_248),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_256),
.Y(n_298)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_238),
.Y(n_257)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_257),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_228),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_259),
.B(n_260),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_228),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_240),
.Y(n_261)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_261),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_217),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_266),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_263),
.A2(n_265),
.B1(n_267),
.B2(n_277),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_269),
.C(n_276),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_249),
.A2(n_224),
.B1(n_197),
.B2(n_138),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_219),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_226),
.A2(n_197),
.B1(n_205),
.B2(n_189),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_244),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_239),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_235),
.B(n_200),
.C(n_214),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_234),
.B(n_222),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_270),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_272),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_236),
.A2(n_176),
.B1(n_220),
.B2(n_192),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_242),
.B(n_31),
.Y(n_275)
);

NOR2x1_ASAP7_75t_L g305 ( 
.A(n_275),
.B(n_160),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_235),
.B(n_225),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_231),
.A2(n_237),
.B1(n_232),
.B2(n_243),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_263),
.A2(n_237),
.B1(n_232),
.B2(n_245),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_279),
.A2(n_280),
.B1(n_303),
.B2(n_272),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_255),
.A2(n_227),
.B1(n_230),
.B2(n_241),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_247),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_285),
.B(n_293),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_256),
.A2(n_247),
.B(n_230),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_286),
.A2(n_302),
.B(n_262),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_250),
.B(n_227),
.Y(n_290)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_290),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_246),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_291),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_264),
.B(n_241),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_246),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_267),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_295),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_257),
.B(n_215),
.Y(n_297)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_297),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_275),
.A2(n_239),
.B1(n_189),
.B2(n_169),
.Y(n_301)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_301),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_273),
.A2(n_209),
.B(n_204),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_277),
.A2(n_167),
.B1(n_143),
.B2(n_164),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_250),
.B(n_212),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_304),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_268),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_274),
.B(n_136),
.C(n_140),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_274),
.C(n_252),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_308),
.B(n_321),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_283),
.B(n_281),
.Y(n_310)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_310),
.Y(n_335)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_311),
.Y(n_342)
);

INVxp33_ASAP7_75t_L g312 ( 
.A(n_292),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_312),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_282),
.Y(n_313)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_313),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_314),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_278),
.B(n_252),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_316),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_317),
.A2(n_318),
.B1(n_319),
.B2(n_322),
.Y(n_348)
);

OA22x2_ASAP7_75t_L g318 ( 
.A1(n_287),
.A2(n_254),
.B1(n_259),
.B2(n_260),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_291),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_327),
.C(n_289),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_288),
.A2(n_261),
.B(n_266),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_325),
.B(n_326),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_282),
.B(n_258),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_289),
.B(n_258),
.C(n_265),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_298),
.A2(n_172),
.B1(n_162),
.B2(n_125),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_329),
.A2(n_331),
.B1(n_303),
.B2(n_279),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_284),
.B(n_31),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_330),
.B(n_34),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_288),
.A2(n_286),
.B1(n_291),
.B2(n_287),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_328),
.A2(n_305),
.B1(n_288),
.B2(n_299),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_332),
.A2(n_336),
.B1(n_347),
.B2(n_341),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_333),
.B(n_331),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_334),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_317),
.A2(n_299),
.B1(n_300),
.B2(n_296),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_327),
.B(n_293),
.C(n_294),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_337),
.B(n_338),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_315),
.B(n_285),
.C(n_306),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_315),
.B(n_300),
.C(n_302),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_340),
.A2(n_341),
.B(n_89),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_321),
.B(n_304),
.C(n_290),
.Y(n_341)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_344),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_311),
.A2(n_278),
.B1(n_139),
.B2(n_34),
.Y(n_345)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_345),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_312),
.B(n_7),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_346),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_348),
.A2(n_319),
.B1(n_322),
.B2(n_307),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_320),
.B(n_146),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_349),
.Y(n_369)
);

BUFx24_ASAP7_75t_SL g350 ( 
.A(n_323),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_350),
.B(n_354),
.Y(n_367)
);

BUFx24_ASAP7_75t_SL g354 ( 
.A(n_324),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_308),
.B(n_146),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_355),
.B(n_340),
.Y(n_361)
);

INVx13_ASAP7_75t_L g356 ( 
.A(n_352),
.Y(n_356)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_356),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_357),
.B(n_359),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_358),
.B(n_362),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_348),
.A2(n_309),
.B1(n_342),
.B2(n_307),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_339),
.A2(n_326),
.B1(n_318),
.B2(n_329),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_360),
.B(n_366),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_361),
.B(n_368),
.Y(n_391)
);

A2O1A1O1Ixp25_ASAP7_75t_L g362 ( 
.A1(n_353),
.A2(n_318),
.B(n_325),
.C(n_314),
.D(n_37),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_338),
.B(n_318),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_363),
.B(n_374),
.Y(n_383)
);

INVx13_ASAP7_75t_L g366 ( 
.A(n_351),
.Y(n_366)
);

NAND2x1_ASAP7_75t_L g368 ( 
.A(n_355),
.B(n_157),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_343),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_373),
.B(n_375),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_357),
.A2(n_335),
.B(n_343),
.Y(n_377)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_377),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_372),
.B(n_333),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_378),
.B(n_380),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_363),
.B(n_337),
.C(n_353),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_359),
.A2(n_166),
.B(n_89),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_381),
.A2(n_371),
.B(n_368),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_361),
.B(n_113),
.C(n_122),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_385),
.B(n_386),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_369),
.B(n_154),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_370),
.B(n_113),
.C(n_106),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_387),
.B(n_389),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_358),
.B(n_106),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_360),
.B(n_24),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_390),
.B(n_365),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_382),
.A2(n_370),
.B(n_362),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_393),
.B(n_396),
.Y(n_409)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_394),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_376),
.A2(n_356),
.B1(n_366),
.B2(n_364),
.Y(n_398)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_398),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_379),
.B(n_367),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_399),
.B(n_400),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_388),
.B(n_18),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_376),
.Y(n_401)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_401),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_383),
.B(n_37),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_402),
.B(n_37),
.C(n_107),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_384),
.B(n_18),
.Y(n_404)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_404),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_397),
.A2(n_380),
.B1(n_383),
.B2(n_398),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_405),
.A2(n_406),
.B1(n_95),
.B2(n_92),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_393),
.A2(n_391),
.B1(n_385),
.B2(n_387),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_395),
.B(n_391),
.C(n_107),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_408),
.B(n_411),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_402),
.B(n_90),
.C(n_105),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_414),
.B(n_149),
.Y(n_424)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_392),
.Y(n_415)
);

AOI322xp5_ASAP7_75t_L g418 ( 
.A1(n_415),
.A2(n_101),
.A3(n_95),
.B1(n_157),
.B2(n_147),
.C1(n_149),
.C2(n_105),
.Y(n_418)
);

NAND3xp33_ASAP7_75t_L g417 ( 
.A(n_409),
.B(n_403),
.C(n_17),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_417),
.Y(n_427)
);

AOI21xp33_ASAP7_75t_L g426 ( 
.A1(n_418),
.A2(n_420),
.B(n_425),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_407),
.B(n_25),
.C(n_7),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_419),
.A2(n_424),
.B(n_6),
.Y(n_428)
);

AOI322xp5_ASAP7_75t_L g420 ( 
.A1(n_412),
.A2(n_410),
.A3(n_415),
.B1(n_416),
.B2(n_413),
.C1(n_414),
.C2(n_411),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_422),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_405),
.A2(n_15),
.B(n_18),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_423),
.A2(n_6),
.B(n_16),
.Y(n_431)
);

AOI322xp5_ASAP7_75t_L g425 ( 
.A1(n_407),
.A2(n_92),
.A3(n_147),
.B1(n_13),
.B2(n_16),
.C1(n_17),
.C2(n_14),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_428),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_421),
.A2(n_6),
.B(n_16),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_430),
.A2(n_427),
.B(n_429),
.Y(n_432)
);

AOI322xp5_ASAP7_75t_L g435 ( 
.A1(n_431),
.A2(n_14),
.A3(n_11),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_432),
.B(n_434),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_426),
.B(n_417),
.Y(n_434)
);

OAI311xp33_ASAP7_75t_L g436 ( 
.A1(n_435),
.A2(n_0),
.A3(n_1),
.B1(n_4),
.C1(n_5),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_436),
.B(n_433),
.C(n_4),
.Y(n_438)
);

OAI321xp33_ASAP7_75t_L g439 ( 
.A1(n_438),
.A2(n_437),
.A3(n_4),
.B1(n_1),
.B2(n_130),
.C(n_25),
.Y(n_439)
);

AOI21x1_ASAP7_75t_L g440 ( 
.A1(n_439),
.A2(n_1),
.B(n_25),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_440),
.B(n_25),
.Y(n_441)
);


endmodule