module fake_ibex_692_n_793 (n_151, n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_120, n_93, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_126, n_1, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_132, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_793);

input n_151;
input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_120;
input n_93;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_126;
input n_1;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_132;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_793;

wire n_599;
wire n_778;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_191;
wire n_593;
wire n_153;
wire n_545;
wire n_583;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_738;
wire n_475;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_375;
wire n_280;
wire n_317;
wire n_340;
wire n_708;
wire n_187;
wire n_667;
wire n_154;
wire n_682;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_723;
wire n_170;
wire n_270;
wire n_383;
wire n_346;
wire n_561;
wire n_417;
wire n_471;
wire n_739;
wire n_755;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_674;
wire n_481;
wire n_243;
wire n_287;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_598;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_732;
wire n_673;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_168;
wire n_526;
wire n_785;
wire n_155;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_789;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_355;
wire n_767;
wire n_474;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_689;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_643;
wire n_679;
wire n_772;
wire n_768;
wire n_338;
wire n_173;
wire n_696;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_257;
wire n_718;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_713;
wire n_307;
wire n_192;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_567;
wire n_548;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_546;
wire n_199;
wire n_788;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_308;
wire n_675;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_397;
wire n_366;
wire n_283;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_332;
wire n_517;
wire n_211;
wire n_744;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_415;
wire n_597;
wire n_288;
wire n_320;
wire n_285;
wire n_379;
wire n_247;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_385;
wire n_342;
wire n_414;
wire n_233;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_217;
wire n_324;
wire n_391;
wire n_537;
wire n_728;
wire n_670;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_752;
wire n_668;
wire n_779;
wire n_266;
wire n_294;
wire n_485;
wire n_284;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_693;
wire n_311;
wire n_661;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_687;
wire n_159;
wire n_202;
wire n_298;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_559;
wire n_425;

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_43),
.Y(n_154)
);

INVxp67_ASAP7_75t_SL g155 ( 
.A(n_50),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_99),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_147),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_38),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_62),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_76),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_128),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_113),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_138),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_142),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_98),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_88),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_101),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_134),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_40),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_4),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_49),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_64),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_105),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_120),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_26),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_103),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_0),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_130),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_75),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_96),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_85),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_145),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_65),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_44),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_77),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_135),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_109),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_28),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_74),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_57),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_116),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_11),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_55),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_37),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_118),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_72),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_108),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_71),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_54),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_87),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_24),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_21),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_117),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_68),
.Y(n_208)
);

INVxp67_ASAP7_75t_SL g209 ( 
.A(n_100),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_111),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_137),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_81),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_131),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_73),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_53),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_119),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_79),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_122),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_34),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_78),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_34),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_95),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_115),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_33),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_102),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_56),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_80),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_51),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_106),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_10),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_136),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_149),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_123),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_70),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_69),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_82),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_84),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_89),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_114),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_3),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_35),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_19),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_146),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_129),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_112),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_104),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_133),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_23),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_151),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_3),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_132),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_5),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_42),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_18),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_83),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_25),
.Y(n_256)
);

BUFx12f_ASAP7_75t_L g257 ( 
.A(n_165),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_152),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_205),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_205),
.Y(n_260)
);

AND2x4_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_0),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_196),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_152),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_177),
.B(n_1),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_2),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_153),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_152),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_225),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_154),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_152),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_225),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_160),
.Y(n_272)
);

OAI22x1_ASAP7_75t_R g273 ( 
.A1(n_173),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_179),
.Y(n_274)
);

BUFx8_ASAP7_75t_L g275 ( 
.A(n_157),
.Y(n_275)
);

OAI21x1_ASAP7_75t_L g276 ( 
.A1(n_158),
.A2(n_63),
.B(n_148),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_174),
.B(n_39),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_178),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_220),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_159),
.B(n_7),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_162),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_179),
.Y(n_282)
);

INVx5_ASAP7_75t_L g283 ( 
.A(n_179),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_202),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_227),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_169),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_179),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_180),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_175),
.Y(n_289)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_181),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_176),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_230),
.B(n_11),
.Y(n_292)
);

OA21x2_ASAP7_75t_L g293 ( 
.A1(n_182),
.A2(n_66),
.B(n_144),
.Y(n_293)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_181),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_240),
.Y(n_295)
);

AND2x2_ASAP7_75t_SL g296 ( 
.A(n_189),
.B(n_150),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_192),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_241),
.B(n_12),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_242),
.B(n_13),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_190),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_177),
.B(n_13),
.Y(n_301)
);

BUFx12f_ASAP7_75t_L g302 ( 
.A(n_164),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_191),
.Y(n_303)
);

OA21x2_ASAP7_75t_L g304 ( 
.A1(n_193),
.A2(n_67),
.B(n_139),
.Y(n_304)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_161),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_248),
.Y(n_306)
);

INVx6_ASAP7_75t_L g307 ( 
.A(n_181),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_173),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_199),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_181),
.Y(n_310)
);

BUFx12f_ASAP7_75t_L g311 ( 
.A(n_164),
.Y(n_311)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_223),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_223),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_203),
.Y(n_314)
);

AND2x6_ASAP7_75t_L g315 ( 
.A(n_207),
.B(n_41),
.Y(n_315)
);

INVx6_ASAP7_75t_L g316 ( 
.A(n_223),
.Y(n_316)
);

OAI22x1_ASAP7_75t_R g317 ( 
.A1(n_156),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_211),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_213),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_214),
.Y(n_320)
);

INVx6_ASAP7_75t_L g321 ( 
.A(n_243),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_216),
.Y(n_322)
);

AND2x6_ASAP7_75t_L g323 ( 
.A(n_218),
.B(n_45),
.Y(n_323)
);

AND2x4_ASAP7_75t_L g324 ( 
.A(n_222),
.B(n_17),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_324),
.B(n_234),
.Y(n_325)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_288),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_321),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_324),
.B(n_296),
.Y(n_328)
);

AO21x2_ASAP7_75t_L g329 ( 
.A1(n_276),
.A2(n_244),
.B(n_238),
.Y(n_329)
);

CKINVDCx6p67_ASAP7_75t_R g330 ( 
.A(n_302),
.Y(n_330)
);

BUFx10_ASAP7_75t_L g331 ( 
.A(n_321),
.Y(n_331)
);

NAND2xp33_ASAP7_75t_SL g332 ( 
.A(n_264),
.B(n_301),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_324),
.Y(n_333)
);

INVx6_ASAP7_75t_L g334 ( 
.A(n_305),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_324),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_302),
.B(n_156),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_311),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_313),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_296),
.B(n_249),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_275),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_296),
.B(n_163),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_321),
.B(n_155),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_315),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_258),
.Y(n_344)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_315),
.Y(n_345)
);

OR2x6_ASAP7_75t_L g346 ( 
.A(n_311),
.B(n_171),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_297),
.B(n_206),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_258),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_303),
.B(n_219),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_263),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_266),
.B(n_166),
.Y(n_351)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_323),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_278),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_278),
.Y(n_354)
);

INVx5_ASAP7_75t_L g355 ( 
.A(n_315),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_264),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_263),
.Y(n_357)
);

AND2x4_ASAP7_75t_L g358 ( 
.A(n_261),
.B(n_209),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_257),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_269),
.B(n_167),
.Y(n_360)
);

NOR2x1p5_ASAP7_75t_L g361 ( 
.A(n_257),
.B(n_221),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_269),
.B(n_168),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_319),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_301),
.B(n_256),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_281),
.B(n_224),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_281),
.B(n_170),
.Y(n_366)
);

NAND2xp33_ASAP7_75t_SL g367 ( 
.A(n_261),
.B(n_171),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_261),
.A2(n_215),
.B1(n_253),
.B2(n_184),
.Y(n_368)
);

INVx2_ASAP7_75t_SL g369 ( 
.A(n_261),
.Y(n_369)
);

AND2x6_ASAP7_75t_L g370 ( 
.A(n_320),
.B(n_194),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_295),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_300),
.B(n_250),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_318),
.B(n_252),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_318),
.B(n_254),
.Y(n_374)
);

INVxp33_ASAP7_75t_L g375 ( 
.A(n_265),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_267),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_319),
.Y(n_377)
);

BUFx10_ASAP7_75t_L g378 ( 
.A(n_315),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_275),
.Y(n_379)
);

OAI22xp33_ASAP7_75t_L g380 ( 
.A1(n_308),
.A2(n_253),
.B1(n_172),
.B2(n_185),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_275),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_322),
.B(n_183),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_320),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_306),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_268),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_270),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_270),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_270),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_274),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_274),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_274),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_268),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_286),
.B(n_186),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_271),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_271),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_272),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_375),
.B(n_286),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_375),
.B(n_289),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_383),
.B(n_291),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_328),
.A2(n_277),
.B1(n_212),
.B2(n_185),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g401 ( 
.A(n_326),
.B(n_308),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_358),
.B(n_291),
.Y(n_402)
);

O2A1O1Ixp33_ASAP7_75t_L g403 ( 
.A1(n_339),
.A2(n_284),
.B(n_292),
.C(n_299),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_363),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_353),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_354),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g407 ( 
.A(n_347),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_328),
.A2(n_304),
.B(n_293),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_351),
.B(n_309),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_358),
.B(n_309),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_351),
.B(n_360),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_358),
.B(n_314),
.Y(n_412)
);

O2A1O1Ixp33_ASAP7_75t_L g413 ( 
.A1(n_339),
.A2(n_298),
.B(n_262),
.C(n_259),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_326),
.B(n_259),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_362),
.B(n_280),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_379),
.B(n_212),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_341),
.A2(n_245),
.B1(n_215),
.B2(n_232),
.Y(n_417)
);

INVx2_ASAP7_75t_SL g418 ( 
.A(n_364),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_377),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_365),
.B(n_315),
.Y(n_420)
);

OR2x6_ASAP7_75t_L g421 ( 
.A(n_346),
.B(n_273),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_371),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_352),
.B(n_187),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_372),
.B(n_323),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_332),
.A2(n_232),
.B1(n_245),
.B2(n_323),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_373),
.B(n_323),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_366),
.B(n_260),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_374),
.B(n_323),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_349),
.B(n_323),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_346),
.B(n_260),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_377),
.Y(n_431)
);

NOR2xp67_ASAP7_75t_L g432 ( 
.A(n_359),
.B(n_279),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_385),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_356),
.B(n_285),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_366),
.B(n_382),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_392),
.Y(n_436)
);

BUFx8_ASAP7_75t_L g437 ( 
.A(n_330),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_352),
.B(n_317),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_355),
.B(n_188),
.Y(n_439)
);

O2A1O1Ixp5_ASAP7_75t_L g440 ( 
.A1(n_325),
.A2(n_293),
.B(n_304),
.C(n_312),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_333),
.Y(n_441)
);

NOR2xp67_ASAP7_75t_L g442 ( 
.A(n_337),
.B(n_18),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_394),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_368),
.B(n_20),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_395),
.Y(n_445)
);

OR2x6_ASAP7_75t_L g446 ( 
.A(n_361),
.B(n_317),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_384),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_381),
.B(n_231),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_340),
.A2(n_293),
.B1(n_304),
.B2(n_195),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_396),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_369),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_335),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_355),
.B(n_197),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_382),
.B(n_198),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_L g455 ( 
.A1(n_335),
.A2(n_293),
.B1(n_304),
.B2(n_316),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_367),
.A2(n_239),
.B1(n_201),
.B2(n_204),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_370),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_327),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_393),
.B(n_200),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_334),
.B(n_208),
.Y(n_460)
);

BUFx8_ASAP7_75t_L g461 ( 
.A(n_370),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_370),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_355),
.B(n_210),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_370),
.A2(n_316),
.B1(n_294),
.B2(n_307),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_334),
.B(n_217),
.Y(n_465)
);

NOR3xp33_ASAP7_75t_L g466 ( 
.A(n_380),
.B(n_226),
.C(n_228),
.Y(n_466)
);

NAND2x1_ASAP7_75t_L g467 ( 
.A(n_370),
.B(n_294),
.Y(n_467)
);

OAI321xp33_ASAP7_75t_L g468 ( 
.A1(n_449),
.A2(n_274),
.A3(n_282),
.B1(n_287),
.B2(n_310),
.C(n_342),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_407),
.B(n_367),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_397),
.B(n_398),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_414),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_420),
.A2(n_343),
.B(n_329),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_437),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_397),
.B(n_336),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_437),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_425),
.A2(n_340),
.B1(n_229),
.B2(n_247),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_424),
.A2(n_428),
.B(n_426),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_400),
.A2(n_233),
.B1(n_235),
.B2(n_236),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_467),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_429),
.A2(n_378),
.B(n_338),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_416),
.B(n_370),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_418),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_452),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_438),
.A2(n_378),
.B1(n_331),
.B2(n_246),
.Y(n_484)
);

CKINVDCx10_ASAP7_75t_R g485 ( 
.A(n_421),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_421),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_451),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_411),
.B(n_251),
.Y(n_488)
);

BUFx4f_ASAP7_75t_L g489 ( 
.A(n_421),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_430),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_433),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_441),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_436),
.Y(n_493)
);

AOI21x1_ASAP7_75t_L g494 ( 
.A1(n_408),
.A2(n_357),
.B(n_390),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_441),
.Y(n_495)
);

AND2x6_ASAP7_75t_L g496 ( 
.A(n_457),
.B(n_282),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_401),
.B(n_417),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_443),
.Y(n_498)
);

NOR2x1p5_ASAP7_75t_L g499 ( 
.A(n_444),
.B(n_22),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_448),
.B(n_22),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_435),
.B(n_23),
.Y(n_501)
);

INVx11_ASAP7_75t_L g502 ( 
.A(n_461),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_445),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_440),
.A2(n_357),
.B(n_389),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_450),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_402),
.B(n_25),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_399),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_410),
.B(n_26),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_458),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_412),
.B(n_27),
.Y(n_510)
);

A2O1A1Ixp33_ASAP7_75t_L g511 ( 
.A1(n_409),
.A2(n_310),
.B(n_290),
.C(n_283),
.Y(n_511)
);

AOI221xp5_ASAP7_75t_SL g512 ( 
.A1(n_403),
.A2(n_376),
.B1(n_388),
.B2(n_387),
.C(n_386),
.Y(n_512)
);

CKINVDCx11_ASAP7_75t_R g513 ( 
.A(n_446),
.Y(n_513)
);

AO32x2_ASAP7_75t_L g514 ( 
.A1(n_462),
.A2(n_283),
.A3(n_290),
.B1(n_312),
.B2(n_31),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_446),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_SL g516 ( 
.A1(n_446),
.A2(n_290),
.B1(n_312),
.B2(n_31),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_427),
.B(n_29),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_456),
.B(n_30),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_432),
.B(n_30),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_405),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_415),
.B(n_32),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_406),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_434),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_403),
.B(n_33),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_422),
.B(n_35),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_447),
.Y(n_526)
);

NOR3xp33_ASAP7_75t_L g527 ( 
.A(n_454),
.B(n_350),
.C(n_348),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_455),
.A2(n_348),
.B1(n_391),
.B2(n_344),
.Y(n_528)
);

AOI21x1_ASAP7_75t_L g529 ( 
.A1(n_439),
.A2(n_391),
.B(n_344),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_459),
.B(n_36),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_460),
.B(n_465),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_455),
.A2(n_391),
.B1(n_344),
.B2(n_36),
.Y(n_532)
);

O2A1O1Ixp33_ASAP7_75t_L g533 ( 
.A1(n_423),
.A2(n_46),
.B(n_47),
.C(n_48),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_477),
.A2(n_453),
.B(n_463),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_507),
.B(n_442),
.Y(n_535)
);

NAND2x1p5_ASAP7_75t_L g536 ( 
.A(n_473),
.B(n_404),
.Y(n_536)
);

AO22x2_ASAP7_75t_L g537 ( 
.A1(n_486),
.A2(n_464),
.B1(n_431),
.B2(n_419),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_507),
.B(n_471),
.Y(n_538)
);

NAND3xp33_ASAP7_75t_L g539 ( 
.A(n_512),
.B(n_391),
.C(n_344),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_471),
.B(n_470),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_475),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_523),
.B(n_52),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_497),
.B(n_58),
.Y(n_543)
);

A2O1A1Ixp33_ASAP7_75t_L g544 ( 
.A1(n_531),
.A2(n_59),
.B(n_60),
.C(n_61),
.Y(n_544)
);

CKINVDCx6p67_ASAP7_75t_R g545 ( 
.A(n_485),
.Y(n_545)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_502),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_490),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_469),
.B(n_90),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_474),
.B(n_91),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_480),
.A2(n_92),
.B(n_93),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_520),
.Y(n_551)
);

NAND2x1p5_ASAP7_75t_L g552 ( 
.A(n_489),
.B(n_94),
.Y(n_552)
);

BUFx4_ASAP7_75t_SL g553 ( 
.A(n_515),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_L g554 ( 
.A1(n_532),
.A2(n_107),
.B(n_110),
.Y(n_554)
);

CKINVDCx11_ASAP7_75t_R g555 ( 
.A(n_513),
.Y(n_555)
);

AO22x2_ASAP7_75t_L g556 ( 
.A1(n_486),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_487),
.B(n_140),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_522),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_479),
.Y(n_559)
);

BUFx4f_ASAP7_75t_L g560 ( 
.A(n_481),
.Y(n_560)
);

A2O1A1Ixp33_ASAP7_75t_SL g561 ( 
.A1(n_468),
.A2(n_518),
.B(n_533),
.C(n_527),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_526),
.B(n_500),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_503),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_492),
.B(n_495),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_499),
.B(n_482),
.Y(n_565)
);

CKINVDCx6p67_ASAP7_75t_R g566 ( 
.A(n_509),
.Y(n_566)
);

INVx6_ASAP7_75t_SL g567 ( 
.A(n_489),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_476),
.B(n_516),
.Y(n_568)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_519),
.Y(n_569)
);

HAxp5_ASAP7_75t_L g570 ( 
.A(n_478),
.B(n_525),
.CON(n_570),
.SN(n_570)
);

OAI21xp5_ASAP7_75t_L g571 ( 
.A1(n_517),
.A2(n_506),
.B(n_508),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_510),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_L g573 ( 
.A1(n_511),
.A2(n_483),
.B(n_530),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_491),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_484),
.B(n_493),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_498),
.Y(n_576)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_505),
.B(n_488),
.Y(n_577)
);

OAI22x1_ASAP7_75t_L g578 ( 
.A1(n_514),
.A2(n_499),
.B1(n_368),
.B2(n_417),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_514),
.A2(n_507),
.B1(n_425),
.B2(n_328),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_496),
.B(n_507),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_473),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_507),
.B(n_471),
.Y(n_582)
);

A2O1A1Ixp33_ASAP7_75t_L g583 ( 
.A1(n_531),
.A2(n_524),
.B(n_501),
.C(n_521),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_520),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_507),
.A2(n_425),
.B1(n_328),
.B2(n_470),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_SL g586 ( 
.A(n_507),
.B(n_345),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_507),
.B(n_471),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_473),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_507),
.B(n_471),
.Y(n_589)
);

OAI21x1_ASAP7_75t_L g590 ( 
.A1(n_494),
.A2(n_504),
.B(n_529),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_SL g591 ( 
.A1(n_486),
.A2(n_421),
.B1(n_446),
.B2(n_173),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_507),
.A2(n_425),
.B1(n_328),
.B2(n_470),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_497),
.A2(n_507),
.B1(n_328),
.B2(n_332),
.Y(n_593)
);

OAI21x1_ASAP7_75t_L g594 ( 
.A1(n_494),
.A2(n_504),
.B(n_529),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_507),
.B(n_471),
.Y(n_595)
);

NOR2xp67_ASAP7_75t_SL g596 ( 
.A(n_473),
.B(n_475),
.Y(n_596)
);

NAND2x1p5_ASAP7_75t_L g597 ( 
.A(n_473),
.B(n_475),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_L g598 ( 
.A1(n_477),
.A2(n_408),
.B(n_472),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_L g599 ( 
.A1(n_477),
.A2(n_408),
.B(n_472),
.Y(n_599)
);

OR2x2_ASAP7_75t_L g600 ( 
.A(n_490),
.B(n_401),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_507),
.B(n_416),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_507),
.B(n_471),
.Y(n_602)
);

INVxp67_ASAP7_75t_SL g603 ( 
.A(n_507),
.Y(n_603)
);

OAI22xp33_ASAP7_75t_L g604 ( 
.A1(n_593),
.A2(n_603),
.B1(n_602),
.B2(n_582),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_545),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_551),
.Y(n_606)
);

AOI221xp5_ASAP7_75t_L g607 ( 
.A1(n_578),
.A2(n_591),
.B1(n_540),
.B2(n_558),
.C(n_584),
.Y(n_607)
);

OA21x2_ASAP7_75t_L g608 ( 
.A1(n_539),
.A2(n_594),
.B(n_590),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_538),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_587),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_589),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_595),
.Y(n_612)
);

OR2x2_ASAP7_75t_L g613 ( 
.A(n_600),
.B(n_547),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_566),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_568),
.A2(n_591),
.B1(n_572),
.B2(n_585),
.Y(n_615)
);

OR3x4_ASAP7_75t_SL g616 ( 
.A(n_555),
.B(n_567),
.C(n_553),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_559),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_593),
.B(n_592),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_SL g619 ( 
.A1(n_556),
.A2(n_557),
.B1(n_579),
.B2(n_554),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_567),
.Y(n_620)
);

OR2x6_ASAP7_75t_L g621 ( 
.A(n_597),
.B(n_588),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_583),
.B(n_569),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_581),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_601),
.A2(n_565),
.B1(n_562),
.B2(n_541),
.Y(n_624)
);

OAI221xp5_ASAP7_75t_L g625 ( 
.A1(n_571),
.A2(n_564),
.B1(n_577),
.B2(n_535),
.C(n_561),
.Y(n_625)
);

OAI21x1_ASAP7_75t_L g626 ( 
.A1(n_573),
.A2(n_550),
.B(n_534),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_563),
.A2(n_575),
.B1(n_571),
.B2(n_543),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_536),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_542),
.B(n_576),
.Y(n_629)
);

BUFx6f_ASAP7_75t_SL g630 ( 
.A(n_596),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_580),
.Y(n_631)
);

CKINVDCx6p67_ASAP7_75t_R g632 ( 
.A(n_574),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_552),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_549),
.A2(n_560),
.B1(n_537),
.B2(n_548),
.Y(n_634)
);

OA21x2_ASAP7_75t_L g635 ( 
.A1(n_544),
.A2(n_570),
.B(n_586),
.Y(n_635)
);

CKINVDCx8_ASAP7_75t_R g636 ( 
.A(n_581),
.Y(n_636)
);

NAND2x1p5_ASAP7_75t_L g637 ( 
.A(n_546),
.B(n_507),
.Y(n_637)
);

AO32x2_ASAP7_75t_L g638 ( 
.A1(n_579),
.A2(n_449),
.A3(n_532),
.B1(n_528),
.B2(n_585),
.Y(n_638)
);

A2O1A1Ixp33_ASAP7_75t_L g639 ( 
.A1(n_583),
.A2(n_571),
.B(n_593),
.C(n_554),
.Y(n_639)
);

AND2x4_ASAP7_75t_SL g640 ( 
.A(n_566),
.B(n_546),
.Y(n_640)
);

INVxp67_ASAP7_75t_SL g641 ( 
.A(n_603),
.Y(n_641)
);

AO21x2_ASAP7_75t_L g642 ( 
.A1(n_539),
.A2(n_599),
.B(n_598),
.Y(n_642)
);

AOI221xp5_ASAP7_75t_L g643 ( 
.A1(n_578),
.A2(n_380),
.B1(n_413),
.B2(n_403),
.C(n_466),
.Y(n_643)
);

BUFx8_ASAP7_75t_SL g644 ( 
.A(n_581),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_566),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_545),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_545),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_603),
.A2(n_367),
.B1(n_466),
.B2(n_336),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_551),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_606),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_641),
.Y(n_651)
);

BUFx12f_ASAP7_75t_L g652 ( 
.A(n_646),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_637),
.Y(n_653)
);

BUFx12f_ASAP7_75t_L g654 ( 
.A(n_646),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_642),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_613),
.B(n_610),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_649),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_615),
.A2(n_607),
.B1(n_643),
.B2(n_619),
.Y(n_658)
);

AND2x6_ASAP7_75t_L g659 ( 
.A(n_618),
.B(n_617),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_633),
.B(n_629),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_611),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_616),
.Y(n_662)
);

BUFx12f_ASAP7_75t_L g663 ( 
.A(n_621),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_629),
.B(n_609),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_612),
.Y(n_665)
);

AO22x1_ASAP7_75t_L g666 ( 
.A1(n_616),
.A2(n_645),
.B1(n_614),
.B2(n_641),
.Y(n_666)
);

OAI21xp5_ASAP7_75t_L g667 ( 
.A1(n_627),
.A2(n_625),
.B(n_639),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_607),
.B(n_648),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_624),
.B(n_625),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_637),
.Y(n_670)
);

HB1xp67_ASAP7_75t_L g671 ( 
.A(n_631),
.Y(n_671)
);

INVx5_ASAP7_75t_L g672 ( 
.A(n_621),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_640),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_SL g674 ( 
.A1(n_630),
.A2(n_622),
.B1(n_618),
.B2(n_623),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_623),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_630),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_628),
.Y(n_677)
);

BUFx10_ASAP7_75t_L g678 ( 
.A(n_640),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_628),
.B(n_632),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_621),
.Y(n_680)
);

INVx8_ASAP7_75t_L g681 ( 
.A(n_644),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_636),
.B(n_604),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_620),
.B(n_604),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_631),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_627),
.B(n_619),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_645),
.B(n_614),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_634),
.B(n_644),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_605),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_672),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_655),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_655),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_651),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_671),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_667),
.B(n_638),
.Y(n_694)
);

INVx4_ASAP7_75t_L g695 ( 
.A(n_659),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_659),
.Y(n_696)
);

BUFx2_ASAP7_75t_L g697 ( 
.A(n_659),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_685),
.B(n_638),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_684),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_650),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_661),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_658),
.B(n_635),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_657),
.B(n_608),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_665),
.B(n_626),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_703),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_689),
.B(n_672),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_698),
.B(n_669),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_690),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_699),
.B(n_656),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_692),
.Y(n_710)
);

OR2x2_ASAP7_75t_L g711 ( 
.A(n_693),
.B(n_683),
.Y(n_711)
);

OR2x2_ASAP7_75t_L g712 ( 
.A(n_693),
.B(n_687),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_694),
.A2(n_669),
.B1(n_682),
.B2(n_668),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_700),
.B(n_688),
.Y(n_714)
);

OR2x6_ASAP7_75t_L g715 ( 
.A(n_695),
.B(n_666),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_704),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_704),
.Y(n_717)
);

INVx5_ASAP7_75t_L g718 ( 
.A(n_695),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_691),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_710),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_719),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_709),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_707),
.B(n_701),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_712),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_716),
.B(n_717),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_718),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_712),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_711),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_711),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_708),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_714),
.B(n_676),
.Y(n_731)
);

AOI211xp5_ASAP7_75t_SL g732 ( 
.A1(n_726),
.A2(n_682),
.B(n_702),
.C(n_694),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_720),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_728),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_729),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_725),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_SL g737 ( 
.A(n_726),
.B(n_662),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_725),
.Y(n_738)
);

AND3x2_ASAP7_75t_L g739 ( 
.A(n_731),
.B(n_697),
.C(n_696),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_724),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_727),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_730),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_723),
.B(n_705),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_721),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_742),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_743),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_743),
.A2(n_726),
.B1(n_715),
.B2(n_662),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_737),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_733),
.B(n_722),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_736),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_738),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_742),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_744),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_L g754 ( 
.A1(n_734),
.A2(n_715),
.B1(n_713),
.B2(n_718),
.Y(n_754)
);

INVxp33_ASAP7_75t_L g755 ( 
.A(n_749),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_746),
.B(n_735),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_752),
.B(n_732),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_752),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_754),
.A2(n_694),
.B1(n_707),
.B2(n_698),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_745),
.B(n_740),
.Y(n_760)
);

NAND3xp33_ASAP7_75t_L g761 ( 
.A(n_757),
.B(n_749),
.C(n_747),
.Y(n_761)
);

NOR3xp33_ASAP7_75t_L g762 ( 
.A(n_757),
.B(n_688),
.C(n_686),
.Y(n_762)
);

NAND3xp33_ASAP7_75t_L g763 ( 
.A(n_758),
.B(n_674),
.C(n_751),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_761),
.B(n_755),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_762),
.B(n_758),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_765),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_764),
.B(n_763),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_766),
.B(n_760),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_767),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_768),
.B(n_756),
.Y(n_770)
);

NOR2x1p5_ASAP7_75t_L g771 ( 
.A(n_769),
.B(n_652),
.Y(n_771)
);

OAI21xp33_ASAP7_75t_L g772 ( 
.A1(n_770),
.A2(n_605),
.B(n_647),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_771),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_771),
.Y(n_774)
);

OR4x1_ASAP7_75t_L g775 ( 
.A(n_774),
.B(n_647),
.C(n_673),
.D(n_654),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_772),
.A2(n_654),
.B1(n_652),
.B2(n_681),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_773),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_772),
.Y(n_778)
);

NOR2x1_ASAP7_75t_L g779 ( 
.A(n_773),
.B(n_679),
.Y(n_779)
);

AO22x2_ASAP7_75t_L g780 ( 
.A1(n_778),
.A2(n_677),
.B1(n_681),
.B2(n_748),
.Y(n_780)
);

OAI22x1_ASAP7_75t_L g781 ( 
.A1(n_777),
.A2(n_681),
.B1(n_672),
.B2(n_680),
.Y(n_781)
);

A2O1A1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_779),
.A2(n_760),
.B(n_750),
.C(n_745),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_776),
.A2(n_775),
.B1(n_759),
.B2(n_715),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_778),
.A2(n_741),
.B1(n_753),
.B2(n_663),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_775),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_785),
.A2(n_678),
.B(n_715),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_780),
.A2(n_663),
.B1(n_678),
.B2(n_715),
.Y(n_787)
);

OAI21xp5_ASAP7_75t_SL g788 ( 
.A1(n_784),
.A2(n_739),
.B(n_674),
.Y(n_788)
);

NAND3xp33_ASAP7_75t_L g789 ( 
.A(n_783),
.B(n_675),
.C(n_670),
.Y(n_789)
);

OAI222xp33_ASAP7_75t_L g790 ( 
.A1(n_786),
.A2(n_781),
.B1(n_782),
.B2(n_653),
.C1(n_660),
.C2(n_706),
.Y(n_790)
);

AOI21xp33_ASAP7_75t_SL g791 ( 
.A1(n_790),
.A2(n_789),
.B(n_788),
.Y(n_791)
);

OR2x2_ASAP7_75t_L g792 ( 
.A(n_791),
.B(n_787),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_792),
.A2(n_660),
.B1(n_653),
.B2(n_664),
.Y(n_793)
);


endmodule