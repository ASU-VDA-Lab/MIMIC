module fake_jpeg_7415_n_80 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_80);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_80;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_8),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx8_ASAP7_75t_SL g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx4_ASAP7_75t_SL g20 ( 
.A(n_18),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_23),
.Y(n_26)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_9),
.B(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_23),
.A2(n_17),
.B1(n_10),
.B2(n_13),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_17),
.B1(n_10),
.B2(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_28),
.B(n_2),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_14),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_31),
.B(n_12),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_30),
.B(n_29),
.C(n_26),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_29),
.Y(n_35)
);

NOR2x1_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_38),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_13),
.B1(n_22),
.B2(n_12),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_19),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_40),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_26),
.A2(n_11),
.B1(n_16),
.B2(n_20),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_43),
.Y(n_52)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_2),
.Y(n_45)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_2),
.Y(n_46)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_58),
.Y(n_65)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_40),
.C(n_36),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_60),
.C(n_55),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_45),
.C(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_56),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_53),
.Y(n_64)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_33),
.B1(n_53),
.B2(n_52),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_59),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_63),
.B(n_64),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_49),
.C(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_67),
.B(n_48),
.Y(n_70)
);

OAI321xp33_ASAP7_75t_L g68 ( 
.A1(n_64),
.A2(n_48),
.A3(n_55),
.B1(n_49),
.B2(n_46),
.C(n_42),
.Y(n_68)
);

OAI321xp33_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_16),
.A3(n_41),
.B1(n_54),
.B2(n_25),
.C(n_51),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_66),
.B1(n_65),
.B2(n_44),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_71),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_73),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_69),
.C(n_54),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_76),
.B(n_51),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_77),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_78),
.B(n_75),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_4),
.Y(n_80)
);


endmodule