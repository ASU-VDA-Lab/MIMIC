module fake_jpeg_1863_n_198 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_198);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_198;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_33),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_34),
.Y(n_65)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

CKINVDCx9p33_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_24),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_17),
.B(n_14),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_9),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_21),
.Y(n_48)
);

NAND2xp33_ASAP7_75t_SL g82 ( 
.A(n_48),
.B(n_61),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_24),
.B1(n_23),
.B2(n_31),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_52),
.A2(n_23),
.B1(n_24),
.B2(n_29),
.Y(n_83)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_56),
.B(n_20),
.Y(n_78)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_21),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_18),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_31),
.Y(n_86)
);

NAND2xp33_ASAP7_75t_SL g64 ( 
.A(n_40),
.B(n_32),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_61),
.B(n_48),
.Y(n_72)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_37),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_67),
.B(n_69),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_36),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_83),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_25),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_74),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_25),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_20),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_78),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_61),
.B(n_17),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_38),
.B1(n_40),
.B2(n_43),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_80),
.A2(n_57),
.B1(n_47),
.B2(n_35),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_21),
.Y(n_81)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_88),
.Y(n_106)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx6_ASAP7_75t_SL g88 ( 
.A(n_60),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_34),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_89),
.A2(n_72),
.B1(n_83),
.B2(n_82),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_95),
.B1(n_109),
.B2(n_112),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_89),
.A2(n_47),
.B1(n_59),
.B2(n_58),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_46),
.B1(n_64),
.B2(n_42),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_99),
.B1(n_100),
.B2(n_66),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_46),
.B1(n_42),
.B2(n_49),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_29),
.B1(n_18),
.B2(n_32),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_35),
.B1(n_71),
.B2(n_27),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_70),
.A2(n_29),
.B1(n_19),
.B2(n_30),
.Y(n_109)
);

INVxp33_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_70),
.A2(n_75),
.B1(n_91),
.B2(n_68),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_116),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_76),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_107),
.C(n_39),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_113),
.A2(n_68),
.B1(n_76),
.B2(n_22),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_122),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_88),
.B(n_87),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_118),
.A2(n_131),
.B(n_127),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_104),
.B(n_85),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_119),
.B(n_121),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_22),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_110),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_130),
.Y(n_136)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_93),
.A2(n_113),
.B1(n_98),
.B2(n_99),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_90),
.Y(n_127)
);

A2O1A1O1Ixp25_ASAP7_75t_L g134 ( 
.A1(n_127),
.A2(n_102),
.B(n_100),
.C(n_103),
.D(n_26),
.Y(n_134)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_113),
.A2(n_30),
.B1(n_19),
.B2(n_27),
.Y(n_132)
);

AOI221xp5_ASAP7_75t_L g138 ( 
.A1(n_132),
.A2(n_133),
.B1(n_92),
.B2(n_109),
.C(n_71),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_103),
.A2(n_30),
.B1(n_19),
.B2(n_26),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_137),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_92),
.B(n_107),
.Y(n_137)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_147),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_149),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_SL g143 ( 
.A(n_132),
.B(n_8),
.C(n_14),
.Y(n_143)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_39),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_144),
.B(n_120),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_126),
.A2(n_90),
.B(n_1),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_118),
.C(n_122),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_137),
.C(n_146),
.Y(n_167)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

MAJx2_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_145),
.C(n_150),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_158),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_149),
.A2(n_148),
.B1(n_145),
.B2(n_135),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_159),
.A2(n_145),
.B1(n_136),
.B2(n_124),
.Y(n_170)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_161),
.B(n_162),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_129),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_120),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_163),
.B(n_133),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_141),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_167),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_173),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_170),
.A2(n_172),
.B1(n_159),
.B2(n_163),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_13),
.C(n_10),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_174),
.B(n_176),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_167),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_171),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_164),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_152),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_152),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_168),
.A2(n_162),
.B(n_158),
.C(n_153),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_180),
.B(n_166),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_176),
.A2(n_161),
.B(n_151),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_182),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_173),
.C(n_169),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_185),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_186),
.A2(n_178),
.B1(n_170),
.B2(n_155),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_188),
.A2(n_190),
.B1(n_9),
.B2(n_2),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_184),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_187),
.A2(n_184),
.B(n_13),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_191),
.A2(n_192),
.B(n_193),
.Y(n_194)
);

NAND3xp33_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_0),
.C(n_4),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_L g195 ( 
.A1(n_192),
.A2(n_190),
.B1(n_5),
.B2(n_6),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_195),
.Y(n_196)
);

OAI31xp33_ASAP7_75t_L g197 ( 
.A1(n_196),
.A2(n_194),
.A3(n_0),
.B(n_6),
.Y(n_197)
);

BUFx24_ASAP7_75t_SL g198 ( 
.A(n_197),
.Y(n_198)
);


endmodule