module fake_jpeg_27122_n_224 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_224);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_SL g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_35),
.B(n_38),
.Y(n_51)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_17),
.B(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_16),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_46),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_24),
.B1(n_26),
.B2(n_29),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_58),
.B1(n_63),
.B2(n_18),
.Y(n_68)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_29),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_30),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_53),
.B(n_39),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_23),
.B(n_19),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_52),
.B1(n_46),
.B2(n_23),
.Y(n_67)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_55),
.B(n_61),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_41),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_24),
.B1(n_22),
.B2(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_36),
.A2(n_22),
.B1(n_30),
.B2(n_27),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_65),
.B(n_75),
.Y(n_98)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_66),
.B(n_74),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_47),
.B1(n_62),
.B2(n_64),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_68),
.A2(n_78),
.B1(n_60),
.B2(n_47),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_81),
.Y(n_94)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_40),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_50),
.A2(n_18),
.B1(n_20),
.B2(n_31),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_79),
.Y(n_109)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_20),
.B1(n_31),
.B2(n_19),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_82),
.A2(n_19),
.B(n_43),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_14),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_86),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_53),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

AND2x6_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_15),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_87),
.B(n_100),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_95),
.B1(n_99),
.B2(n_79),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_90),
.A2(n_101),
.B1(n_81),
.B2(n_82),
.Y(n_123)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_93),
.Y(n_112)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_60),
.B1(n_43),
.B2(n_61),
.Y(n_95)
);

BUFx12_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_66),
.A2(n_64),
.B1(n_60),
.B2(n_40),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_70),
.A2(n_43),
.B1(n_40),
.B2(n_42),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_76),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_69),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_108),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_111),
.A2(n_113),
.B1(n_128),
.B2(n_125),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_98),
.B1(n_108),
.B2(n_99),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_120),
.Y(n_144)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_107),
.B(n_70),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_116),
.B(n_122),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_65),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_121),
.Y(n_134)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_75),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_103),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_123),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_74),
.Y(n_124)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_127),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_98),
.B(n_75),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_126),
.A2(n_95),
.B(n_87),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_69),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_90),
.A2(n_80),
.B1(n_73),
.B2(n_86),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_41),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_88),
.C(n_96),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_96),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_130),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_132),
.Y(n_156)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_138),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_127),
.C(n_129),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_95),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_141),
.A2(n_120),
.B(n_123),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_88),
.C(n_105),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_143),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_102),
.B(n_105),
.C(n_91),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_110),
.A2(n_113),
.B(n_114),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_13),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_147),
.A2(n_149),
.B1(n_133),
.B2(n_139),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_91),
.C(n_96),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_151),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_72),
.C(n_109),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_158),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_155),
.A2(n_157),
.B1(n_160),
.B2(n_163),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_140),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_151),
.A2(n_128),
.B1(n_119),
.B2(n_109),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_143),
.A2(n_92),
.B1(n_32),
.B2(n_49),
.Y(n_163)
);

AO21x1_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_168),
.B(n_11),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_28),
.B1(n_42),
.B2(n_34),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_165),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_134),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_166),
.Y(n_169)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_167),
.Y(n_177)
);

FAx1_ASAP7_75t_SL g168 ( 
.A(n_138),
.B(n_42),
.CI(n_34),
.CON(n_168),
.SN(n_168)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_137),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_176),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_134),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_172),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_135),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_132),
.C(n_145),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_180),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_131),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_178),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_49),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_154),
.B(n_13),
.Y(n_178)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_156),
.Y(n_180)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_182),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_11),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_183),
.B(n_2),
.Y(n_185)
);

NOR3xp33_ASAP7_75t_SL g184 ( 
.A(n_179),
.B(n_155),
.C(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_184),
.B(n_185),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_181),
.A2(n_175),
.B1(n_161),
.B2(n_160),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_187),
.A2(n_193),
.B1(n_157),
.B2(n_162),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_194),
.A2(n_168),
.B1(n_177),
.B2(n_169),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_193),
.B(n_172),
.C(n_174),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_196),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_201),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_192),
.A2(n_161),
.B(n_168),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_199),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_171),
.C(n_163),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_4),
.C(n_5),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_184),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_5),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_191),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_208),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_190),
.Y(n_208)
);

NOR2xp67_ASAP7_75t_SL g209 ( 
.A(n_199),
.B(n_188),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_209),
.B(n_210),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_195),
.C(n_202),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_212),
.B(n_214),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_210),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_215),
.A2(n_6),
.B(n_7),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_213),
.A2(n_200),
.B(n_7),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_216),
.A2(n_218),
.B(n_217),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_220),
.C(n_6),
.Y(n_221)
);

AOI322xp5_ASAP7_75t_L g220 ( 
.A1(n_217),
.A2(n_214),
.A3(n_211),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_7),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_10),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_8),
.Y(n_223)
);

HAxp5_ASAP7_75t_SL g224 ( 
.A(n_223),
.B(n_8),
.CON(n_224),
.SN(n_224)
);


endmodule