module real_aes_8872_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_548;
wire n_678;
wire n_427;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_234;
wire n_284;
wire n_656;
wire n_316;
wire n_532;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_504;
wire n_455;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_691;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_681;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_224;
wire n_639;
wire n_587;
wire n_546;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI22xp33_ASAP7_75t_SL g299 ( .A1(n_0), .A2(n_204), .B1(n_300), .B2(n_305), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g347 ( .A1(n_1), .A2(n_212), .B1(n_348), .B2(n_349), .Y(n_347) );
AOI22xp33_ASAP7_75t_SL g574 ( .A1(n_2), .A2(n_194), .B1(n_450), .B2(n_575), .Y(n_574) );
AOI22xp33_ASAP7_75t_SL g576 ( .A1(n_3), .A2(n_85), .B1(n_315), .B2(n_521), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_4), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_5), .B(n_540), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g612 ( .A(n_6), .Y(n_612) );
AOI222xp33_ASAP7_75t_L g702 ( .A1(n_7), .A2(n_64), .B1(n_203), .B2(n_262), .C1(n_269), .C2(n_703), .Y(n_702) );
AOI22xp5_ASAP7_75t_SL g601 ( .A1(n_8), .A2(n_47), .B1(n_329), .B2(n_438), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_9), .B(n_700), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_10), .A2(n_137), .B1(n_322), .B2(n_388), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_11), .B(n_540), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_12), .A2(n_58), .B1(n_429), .B2(n_614), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_13), .A2(n_101), .B1(n_281), .B2(n_457), .Y(n_456) );
AOI22xp33_ASAP7_75t_SL g578 ( .A1(n_14), .A2(n_181), .B1(n_355), .B2(n_579), .Y(n_578) );
AOI22xp33_ASAP7_75t_SL g259 ( .A1(n_15), .A2(n_116), .B1(n_260), .B2(n_268), .Y(n_259) );
AOI22xp33_ASAP7_75t_SL g369 ( .A1(n_16), .A2(n_111), .B1(n_370), .B2(n_371), .Y(n_369) );
AOI222xp33_ASAP7_75t_L g357 ( .A1(n_17), .A2(n_89), .B1(n_105), .B2(n_244), .C1(n_358), .C2(n_361), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_18), .A2(n_28), .B1(n_294), .B2(n_360), .Y(n_669) );
INVx1_ASAP7_75t_L g543 ( .A(n_19), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_20), .A2(n_213), .B1(n_269), .B2(n_294), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_21), .A2(n_606), .B1(n_638), .B2(n_639), .Y(n_605) );
INVx1_ASAP7_75t_L g639 ( .A(n_21), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_22), .A2(n_147), .B1(n_450), .B2(n_451), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g628 ( .A(n_23), .Y(n_628) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_24), .Y(n_480) );
AO22x2_ASAP7_75t_L g247 ( .A1(n_25), .A2(n_65), .B1(n_248), .B2(n_249), .Y(n_247) );
INVx1_ASAP7_75t_L g654 ( .A(n_25), .Y(n_654) );
AOI22xp5_ASAP7_75t_SL g600 ( .A1(n_26), .A2(n_217), .B1(n_305), .B2(n_492), .Y(n_600) );
AOI22xp33_ASAP7_75t_SL g318 ( .A1(n_27), .A2(n_49), .B1(n_319), .B2(n_322), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_29), .B(n_591), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_30), .A2(n_129), .B1(n_320), .B2(n_355), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_31), .A2(n_61), .B1(n_310), .B2(n_435), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_32), .A2(n_195), .B1(n_302), .B2(n_579), .Y(n_691) );
AOI22xp5_ASAP7_75t_SL g595 ( .A1(n_33), .A2(n_115), .B1(n_486), .B2(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_34), .A2(n_215), .B1(n_289), .B2(n_384), .Y(n_383) );
AO22x2_ASAP7_75t_L g251 ( .A1(n_35), .A2(n_68), .B1(n_248), .B2(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g655 ( .A(n_35), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_36), .A2(n_158), .B1(n_438), .B2(n_439), .Y(n_437) );
AOI22xp33_ASAP7_75t_SL g432 ( .A1(n_37), .A2(n_80), .B1(n_433), .B2(n_435), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_38), .A2(n_51), .B1(n_294), .B2(n_460), .Y(n_459) );
AOI222xp33_ASAP7_75t_L g461 ( .A1(n_39), .A2(n_131), .B1(n_175), .B2(n_462), .C1(n_463), .C2(n_464), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_40), .A2(n_134), .B1(n_340), .B2(n_341), .Y(n_339) );
CKINVDCx20_ASAP7_75t_R g634 ( .A(n_41), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_42), .A2(n_221), .B1(n_340), .B2(n_374), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g558 ( .A(n_43), .Y(n_558) );
AOI22xp33_ASAP7_75t_SL g286 ( .A1(n_44), .A2(n_63), .B1(n_287), .B2(n_292), .Y(n_286) );
XOR2xp5_ASAP7_75t_L g334 ( .A(n_45), .B(n_335), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_46), .A2(n_239), .B1(n_240), .B2(n_332), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_46), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_48), .Y(n_513) );
AOI22xp33_ASAP7_75t_SL g483 ( .A1(n_50), .A2(n_103), .B1(n_484), .B2(n_486), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_52), .A2(n_157), .B1(n_320), .B2(n_512), .Y(n_511) );
AOI22xp33_ASAP7_75t_SL g487 ( .A1(n_53), .A2(n_93), .B1(n_488), .B2(n_489), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_54), .B(n_281), .Y(n_506) );
AOI22xp33_ASAP7_75t_SL g664 ( .A1(n_55), .A2(n_120), .B1(n_348), .B2(n_665), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_56), .A2(n_183), .B1(n_388), .B2(n_690), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_57), .Y(n_524) );
AOI22xp33_ASAP7_75t_SL g593 ( .A1(n_59), .A2(n_206), .B1(n_349), .B2(n_542), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_60), .A2(n_66), .B1(n_345), .B2(n_346), .Y(n_344) );
INVxp67_ASAP7_75t_L g685 ( .A(n_62), .Y(n_685) );
XNOR2x2_ASAP7_75t_L g686 ( .A(n_62), .B(n_687), .Y(n_686) );
CKINVDCx20_ASAP7_75t_R g390 ( .A(n_67), .Y(n_390) );
AOI22xp33_ASAP7_75t_SL g428 ( .A1(n_69), .A2(n_150), .B1(n_429), .B2(n_431), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_70), .B(n_280), .Y(n_592) );
CKINVDCx20_ASAP7_75t_R g668 ( .A(n_71), .Y(n_668) );
INVx1_ASAP7_75t_L g230 ( .A(n_72), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_73), .A2(n_97), .B1(n_320), .B2(n_322), .Y(n_693) );
AOI22xp33_ASAP7_75t_SL g672 ( .A1(n_74), .A2(n_127), .B1(n_454), .B2(n_492), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_75), .A2(n_91), .B1(n_352), .B2(n_353), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_76), .A2(n_113), .B1(n_262), .B2(n_360), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g410 ( .A(n_77), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_78), .A2(n_156), .B1(n_302), .B2(n_371), .Y(n_500) );
INVx1_ASAP7_75t_L g226 ( .A(n_79), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_81), .A2(n_146), .B1(n_435), .B2(n_676), .Y(n_694) );
AOI22xp33_ASAP7_75t_SL g677 ( .A1(n_82), .A2(n_92), .B1(n_489), .B2(n_519), .Y(n_677) );
CKINVDCx20_ASAP7_75t_R g414 ( .A(n_83), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_84), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_86), .A2(n_117), .B1(n_338), .B2(n_435), .Y(n_447) );
OA22x2_ASAP7_75t_L g467 ( .A1(n_87), .A2(n_468), .B1(n_469), .B2(n_470), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_87), .Y(n_468) );
AOI22xp33_ASAP7_75t_SL g309 ( .A1(n_88), .A2(n_90), .B1(n_310), .B2(n_315), .Y(n_309) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_94), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_95), .A2(n_100), .B1(n_353), .B2(n_446), .Y(n_445) );
AOI22xp33_ASAP7_75t_SL g588 ( .A1(n_96), .A2(n_143), .B1(n_260), .B2(n_360), .Y(n_588) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_98), .Y(n_534) );
AOI22xp33_ASAP7_75t_SL g499 ( .A1(n_99), .A2(n_178), .B1(n_331), .B2(n_434), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_102), .Y(n_527) );
XOR2x2_ASAP7_75t_L g394 ( .A(n_104), .B(n_395), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_106), .A2(n_180), .B1(n_439), .B2(n_451), .Y(n_580) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_107), .Y(n_570) );
XNOR2x2_ASAP7_75t_L g442 ( .A(n_108), .B(n_443), .Y(n_442) );
AOI22xp33_ASAP7_75t_SL g675 ( .A1(n_109), .A2(n_128), .B1(n_329), .B2(n_676), .Y(n_675) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_110), .Y(n_528) );
AND2x2_ASAP7_75t_L g229 ( .A(n_112), .B(n_230), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g587 ( .A(n_114), .Y(n_587) );
CKINVDCx20_ASAP7_75t_R g629 ( .A(n_118), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_119), .A2(n_177), .B1(n_431), .B2(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_121), .B(n_462), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_122), .B(n_275), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_123), .B(n_345), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_124), .A2(n_167), .B1(n_287), .B2(n_542), .Y(n_701) );
AND2x6_ASAP7_75t_L g225 ( .A(n_125), .B(n_226), .Y(n_225) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_125), .Y(n_648) );
AO22x2_ASAP7_75t_L g255 ( .A1(n_126), .A2(n_188), .B1(n_248), .B2(n_252), .Y(n_255) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_130), .Y(n_403) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_132), .A2(n_223), .B(n_231), .C(n_656), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_133), .A2(n_208), .B1(n_269), .B2(n_294), .Y(n_379) );
AOI22xp5_ASAP7_75t_SL g597 ( .A1(n_135), .A2(n_187), .B1(n_489), .B2(n_598), .Y(n_597) );
AOI22xp33_ASAP7_75t_SL g491 ( .A1(n_136), .A2(n_196), .B1(n_374), .B2(n_492), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_138), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_139), .A2(n_205), .B1(n_460), .B2(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_140), .B(n_538), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_141), .A2(n_174), .B1(n_263), .B2(n_289), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_142), .B(n_280), .Y(n_279) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_144), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_145), .A2(n_202), .B1(n_342), .B2(n_521), .Y(n_520) );
AOI22xp33_ASAP7_75t_SL g493 ( .A1(n_148), .A2(n_153), .B1(n_326), .B2(n_337), .Y(n_493) );
AO22x2_ASAP7_75t_L g257 ( .A1(n_149), .A2(n_198), .B1(n_248), .B2(n_249), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_151), .A2(n_219), .B1(n_320), .B2(n_338), .Y(n_389) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_152), .Y(n_473) );
AOI22xp33_ASAP7_75t_SL g535 ( .A1(n_154), .A2(n_171), .B1(n_262), .B2(n_464), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_155), .B(n_274), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_159), .A2(n_176), .B1(n_305), .B2(n_596), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_160), .A2(n_179), .B1(n_329), .B2(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g602 ( .A(n_161), .Y(n_602) );
CKINVDCx20_ASAP7_75t_R g632 ( .A(n_162), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_163), .Y(n_565) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_164), .Y(n_420) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_165), .A2(n_658), .B1(n_659), .B2(n_678), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g678 ( .A(n_165), .Y(n_678) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_166), .Y(n_636) );
AOI22xp33_ASAP7_75t_SL g325 ( .A1(n_168), .A2(n_169), .B1(n_326), .B2(n_329), .Y(n_325) );
AOI22xp33_ASAP7_75t_SL g386 ( .A1(n_170), .A2(n_218), .B1(n_387), .B2(n_388), .Y(n_386) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_172), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_173), .B(n_275), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g610 ( .A(n_182), .Y(n_610) );
CKINVDCx20_ASAP7_75t_R g617 ( .A(n_184), .Y(n_617) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_185), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g623 ( .A(n_186), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_188), .B(n_653), .Y(n_652) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_189), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g398 ( .A(n_190), .Y(n_398) );
CKINVDCx20_ASAP7_75t_R g377 ( .A(n_191), .Y(n_377) );
AOI22xp33_ASAP7_75t_SL g510 ( .A1(n_192), .A2(n_220), .B1(n_323), .B2(n_328), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_193), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_197), .Y(n_503) );
INVx1_ASAP7_75t_L g651 ( .A(n_198), .Y(n_651) );
CKINVDCx20_ASAP7_75t_R g417 ( .A(n_199), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_200), .B(n_262), .Y(n_415) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_201), .Y(n_258) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_207), .Y(n_557) );
INVx1_ASAP7_75t_L g248 ( .A(n_209), .Y(n_248) );
INVx1_ASAP7_75t_L g250 ( .A(n_209), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g567 ( .A(n_210), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_211), .A2(n_214), .B1(n_337), .B2(n_338), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_216), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_227), .Y(n_224) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_226), .Y(n_647) );
OAI21xp5_ASAP7_75t_L g683 ( .A1(n_227), .A2(n_646), .B(n_684), .Y(n_683) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_228), .Y(n_227) );
INVxp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AOI221xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_548), .B1(n_641), .B2(n_642), .C(n_643), .Y(n_231) );
INVxp67_ASAP7_75t_L g641 ( .A(n_232), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B1(n_363), .B2(n_547), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
OAI22xp5_ASAP7_75t_SL g234 ( .A1(n_235), .A2(n_236), .B1(n_333), .B2(n_362), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
BUFx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g332 ( .A(n_240), .Y(n_332) );
NAND3x1_ASAP7_75t_L g240 ( .A(n_241), .B(n_298), .C(n_317), .Y(n_240) );
NOR2x1_ASAP7_75t_L g241 ( .A(n_242), .B(n_272), .Y(n_241) );
OAI21xp5_ASAP7_75t_SL g242 ( .A1(n_243), .A2(n_258), .B(n_259), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx4_ASAP7_75t_L g378 ( .A(n_245), .Y(n_378) );
INVx2_ASAP7_75t_L g409 ( .A(n_245), .Y(n_409) );
BUFx3_ASAP7_75t_L g462 ( .A(n_245), .Y(n_462) );
INVx2_ASAP7_75t_SL g564 ( .A(n_245), .Y(n_564) );
AND2x6_ASAP7_75t_L g245 ( .A(n_246), .B(n_253), .Y(n_245) );
AND2x4_ASAP7_75t_L g295 ( .A(n_246), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g424 ( .A(n_246), .Y(n_424) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_251), .Y(n_246) );
AND2x2_ASAP7_75t_L g267 ( .A(n_247), .B(n_255), .Y(n_267) );
INVx2_ASAP7_75t_L g277 ( .A(n_247), .Y(n_277) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g252 ( .A(n_250), .Y(n_252) );
INVx2_ASAP7_75t_L g266 ( .A(n_251), .Y(n_266) );
AND2x2_ASAP7_75t_L g276 ( .A(n_251), .B(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g285 ( .A(n_251), .B(n_277), .Y(n_285) );
INVx1_ASAP7_75t_L g291 ( .A(n_251), .Y(n_291) );
AND2x2_ASAP7_75t_L g321 ( .A(n_253), .B(n_304), .Y(n_321) );
AND2x6_ASAP7_75t_L g328 ( .A(n_253), .B(n_284), .Y(n_328) );
AND2x4_ASAP7_75t_L g331 ( .A(n_253), .B(n_276), .Y(n_331) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_256), .Y(n_253) );
AND2x2_ASAP7_75t_L g278 ( .A(n_254), .B(n_257), .Y(n_278) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_255), .B(n_257), .Y(n_308) );
AND2x2_ASAP7_75t_L g314 ( .A(n_255), .B(n_297), .Y(n_314) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g265 ( .A(n_257), .Y(n_265) );
INVx1_ASAP7_75t_L g297 ( .A(n_257), .Y(n_297) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx4_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_263), .Y(n_348) );
BUFx4f_ASAP7_75t_SL g384 ( .A(n_263), .Y(n_384) );
BUFx2_ASAP7_75t_L g463 ( .A(n_263), .Y(n_463) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_263), .Y(n_562) );
AND2x4_ASAP7_75t_L g263 ( .A(n_264), .B(n_267), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx1_ASAP7_75t_L g271 ( .A(n_265), .Y(n_271) );
AND2x2_ASAP7_75t_L g304 ( .A(n_266), .B(n_277), .Y(n_304) );
INVx1_ASAP7_75t_L g372 ( .A(n_266), .Y(n_372) );
AND2x4_ASAP7_75t_L g270 ( .A(n_267), .B(n_271), .Y(n_270) );
AND2x4_ASAP7_75t_L g289 ( .A(n_267), .B(n_290), .Y(n_289) );
NAND2x1p5_ASAP7_75t_L g419 ( .A(n_267), .B(n_372), .Y(n_419) );
INVx1_ASAP7_75t_L g566 ( .A(n_268), .Y(n_566) );
BUFx4f_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
BUFx12f_ASAP7_75t_L g360 ( .A(n_270), .Y(n_360) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_270), .Y(n_413) );
NAND3xp33_ASAP7_75t_L g272 ( .A(n_273), .B(n_279), .C(n_286), .Y(n_272) );
BUFx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
BUFx4f_ASAP7_75t_L g346 ( .A(n_275), .Y(n_346) );
INVx1_ASAP7_75t_SL g458 ( .A(n_275), .Y(n_458) );
BUFx2_ASAP7_75t_L g538 ( .A(n_275), .Y(n_538) );
AND2x6_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
AND2x2_ASAP7_75t_L g313 ( .A(n_276), .B(n_314), .Y(n_313) );
NAND2x1p5_ASAP7_75t_L g407 ( .A(n_276), .B(n_278), .Y(n_407) );
AND2x4_ASAP7_75t_L g283 ( .A(n_278), .B(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g303 ( .A(n_278), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g402 ( .A(n_278), .Y(n_402) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx5_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g345 ( .A(n_282), .Y(n_345) );
INVx2_ASAP7_75t_L g540 ( .A(n_282), .Y(n_540) );
INVx2_ASAP7_75t_L g700 ( .A(n_282), .Y(n_700) );
INVx4_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g401 ( .A(n_285), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g460 ( .A(n_288), .Y(n_460) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx3_ASAP7_75t_L g349 ( .A(n_289), .Y(n_349) );
BUFx2_ASAP7_75t_L g665 ( .A(n_289), .Y(n_665) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x6_ASAP7_75t_L g316 ( .A(n_291), .B(n_308), .Y(n_316) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
BUFx6f_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
BUFx3_ASAP7_75t_L g361 ( .A(n_295), .Y(n_361) );
BUFx2_ASAP7_75t_SL g542 ( .A(n_295), .Y(n_542) );
INVx1_ASAP7_75t_L g425 ( .A(n_296), .Y(n_425) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_309), .Y(n_298) );
INVx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx4_ASAP7_75t_L g446 ( .A(n_301), .Y(n_446) );
INVx4_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
BUFx3_ASAP7_75t_L g340 ( .A(n_303), .Y(n_340) );
BUFx3_ASAP7_75t_L g486 ( .A(n_303), .Y(n_486) );
BUFx3_ASAP7_75t_L g519 ( .A(n_303), .Y(n_519) );
INVx2_ASAP7_75t_L g616 ( .A(n_303), .Y(n_616) );
AND2x4_ASAP7_75t_L g306 ( .A(n_304), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g324 ( .A(n_304), .B(n_314), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_304), .B(n_314), .Y(n_531) );
BUFx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx3_ASAP7_75t_L g353 ( .A(n_306), .Y(n_353) );
BUFx3_ASAP7_75t_L g374 ( .A(n_306), .Y(n_374) );
BUFx2_ASAP7_75t_SL g431 ( .A(n_306), .Y(n_431) );
BUFx3_ASAP7_75t_L g512 ( .A(n_306), .Y(n_512) );
BUFx2_ASAP7_75t_SL g579 ( .A(n_306), .Y(n_579) );
INVx1_ASAP7_75t_L g618 ( .A(n_306), .Y(n_618) );
AND2x2_ASAP7_75t_L g371 ( .A(n_307), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx3_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
BUFx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx3_ASAP7_75t_L g338 ( .A(n_312), .Y(n_338) );
INVx4_ASAP7_75t_L g434 ( .A(n_312), .Y(n_434) );
INVx5_ASAP7_75t_L g488 ( .A(n_312), .Y(n_488) );
INVx1_ASAP7_75t_L g676 ( .A(n_312), .Y(n_676) );
INVx8_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
INVx6_ASAP7_75t_SL g342 ( .A(n_316), .Y(n_342) );
INVx1_ASAP7_75t_L g435 ( .A(n_316), .Y(n_435) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_325), .Y(n_317) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx3_ASAP7_75t_L g430 ( .A(n_320), .Y(n_430) );
BUFx3_ASAP7_75t_L g450 ( .A(n_320), .Y(n_450) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g485 ( .A(n_321), .Y(n_485) );
BUFx2_ASAP7_75t_SL g596 ( .A(n_321), .Y(n_596) );
BUFx4f_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g452 ( .A(n_323), .Y(n_452) );
BUFx3_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
BUFx3_ASAP7_75t_L g352 ( .A(n_324), .Y(n_352) );
BUFx3_ASAP7_75t_L g370 ( .A(n_324), .Y(n_370) );
BUFx3_ASAP7_75t_L g492 ( .A(n_324), .Y(n_492) );
INVx4_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_SL g438 ( .A(n_327), .Y(n_438) );
INVx11_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx11_ASAP7_75t_L g356 ( .A(n_328), .Y(n_356) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_330), .A2(n_356), .B1(n_524), .B2(n_525), .Y(n_523) );
INVx6_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx3_ASAP7_75t_L g337 ( .A(n_331), .Y(n_337) );
BUFx3_ASAP7_75t_L g388 ( .A(n_331), .Y(n_388) );
BUFx3_ASAP7_75t_L g575 ( .A(n_331), .Y(n_575) );
CKINVDCx16_ASAP7_75t_R g362 ( .A(n_333), .Y(n_362) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND5xp2_ASAP7_75t_SL g335 ( .A(n_336), .B(n_339), .C(n_343), .D(n_350), .E(n_357), .Y(n_335) );
BUFx2_ASAP7_75t_L g439 ( .A(n_340), .Y(n_439) );
BUFx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx2_ASAP7_75t_L g489 ( .A(n_342), .Y(n_489) );
AND2x2_ASAP7_75t_SL g343 ( .A(n_344), .B(n_347), .Y(n_343) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_354), .Y(n_350) );
BUFx3_ASAP7_75t_L g614 ( .A(n_352), .Y(n_614) );
INVx5_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_SL g387 ( .A(n_356), .Y(n_387) );
INVx4_ASAP7_75t_L g454 ( .A(n_356), .Y(n_454) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_356), .Y(n_609) );
INVx1_ASAP7_75t_L g690 ( .A(n_356), .Y(n_690) );
INVx3_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx4f_ASAP7_75t_SL g464 ( .A(n_360), .Y(n_464) );
INVx1_ASAP7_75t_L g547 ( .A(n_363), .Y(n_547) );
XOR2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_465), .Y(n_363) );
XOR2xp5_ASAP7_75t_L g364 ( .A(n_365), .B(n_391), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
XOR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_390), .Y(n_366) );
NAND3x1_ASAP7_75t_L g367 ( .A(n_368), .B(n_375), .C(n_385), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_373), .Y(n_368) );
NOR2x1_ASAP7_75t_L g375 ( .A(n_376), .B(n_380), .Y(n_375) );
OAI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_378), .B(n_379), .Y(n_376) );
OAI21xp5_ASAP7_75t_L g502 ( .A1(n_378), .A2(n_503), .B(n_504), .Y(n_502) );
OAI21xp5_ASAP7_75t_SL g533 ( .A1(n_378), .A2(n_534), .B(n_535), .Y(n_533) );
OAI21xp5_ASAP7_75t_SL g586 ( .A1(n_378), .A2(n_587), .B(n_588), .Y(n_586) );
BUFx2_ASAP7_75t_L g667 ( .A(n_378), .Y(n_667) );
INVx4_ASAP7_75t_L g703 ( .A(n_378), .Y(n_703) );
NAND3xp33_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .C(n_383), .Y(n_380) );
INVx1_ASAP7_75t_L g627 ( .A(n_384), .Y(n_627) );
AND2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_389), .Y(n_385) );
INVx3_ASAP7_75t_L g611 ( .A(n_388), .Y(n_611) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OAI22xp5_ASAP7_75t_SL g392 ( .A1(n_393), .A2(n_394), .B1(n_441), .B2(n_442), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_426), .Y(n_395) );
NOR3xp33_ASAP7_75t_L g396 ( .A(n_397), .B(n_408), .C(n_416), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B1(n_403), .B2(n_404), .Y(n_397) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g624 ( .A(n_400), .Y(n_624) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx3_ASAP7_75t_L g474 ( .A(n_401), .Y(n_474) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_401), .Y(n_556) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_406), .A2(n_473), .B1(n_474), .B2(n_475), .Y(n_472) );
OAI22xp5_ASAP7_75t_SL g555 ( .A1(n_406), .A2(n_556), .B1(n_557), .B2(n_558), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_406), .A2(n_623), .B1(n_624), .B2(n_625), .Y(n_622) );
BUFx3_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g698 ( .A(n_407), .Y(n_698) );
OAI221xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B1(n_411), .B2(n_414), .C(n_415), .Y(n_408) );
OAI222xp33_ASAP7_75t_L g626 ( .A1(n_409), .A2(n_627), .B1(n_628), .B2(n_629), .C1(n_630), .C2(n_632), .Y(n_626) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx3_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B1(n_420), .B2(n_421), .Y(n_416) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_419), .A2(n_423), .B1(n_480), .B2(n_481), .Y(n_479) );
BUFx3_ASAP7_75t_L g569 ( .A(n_419), .Y(n_569) );
INVx4_ASAP7_75t_L g631 ( .A(n_419), .Y(n_631) );
OAI22xp5_ASAP7_75t_SL g568 ( .A1(n_421), .A2(n_569), .B1(n_570), .B2(n_571), .Y(n_568) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
CKINVDCx16_ASAP7_75t_R g422 ( .A(n_423), .Y(n_422) );
BUFx2_ASAP7_75t_L g637 ( .A(n_423), .Y(n_637) );
OR2x6_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_436), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_432), .Y(n_427) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_430), .A2(n_527), .B1(n_528), .B2(n_529), .Y(n_526) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g522 ( .A(n_434), .Y(n_522) );
BUFx2_ASAP7_75t_L g598 ( .A(n_434), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_440), .Y(n_436) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NAND4xp75_ASAP7_75t_L g443 ( .A(n_444), .B(n_448), .C(n_455), .D(n_461), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_447), .Y(n_444) );
AND2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_453), .Y(n_448) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_SL g455 ( .A(n_456), .B(n_459), .Y(n_455) );
INVx1_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_SL g591 ( .A(n_458), .Y(n_591) );
INVx1_ASAP7_75t_L g635 ( .A(n_464), .Y(n_635) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_494), .B1(n_545), .B2(n_546), .Y(n_466) );
INVx2_ASAP7_75t_SL g545 ( .A(n_467), .Y(n_545) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND3x1_ASAP7_75t_L g470 ( .A(n_471), .B(n_482), .C(n_490), .Y(n_470) );
NOR3xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_476), .C(n_479), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_487), .Y(n_482) );
INVx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_493), .Y(n_490) );
INVx1_ASAP7_75t_L g546 ( .A(n_494), .Y(n_546) );
OA22x2_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B1(n_514), .B2(n_544), .Y(n_494) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
XOR2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_513), .Y(n_496) );
NAND3x1_ASAP7_75t_SL g497 ( .A(n_498), .B(n_501), .C(n_509), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
NOR2x1_ASAP7_75t_L g501 ( .A(n_502), .B(n_505), .Y(n_501) );
NAND3xp33_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .C(n_508), .Y(n_505) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
INVx1_ASAP7_75t_L g544 ( .A(n_514), .Y(n_544) );
XOR2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_543), .Y(n_514) );
AND2x2_ASAP7_75t_SL g515 ( .A(n_516), .B(n_532), .Y(n_515) );
NOR3xp33_ASAP7_75t_L g516 ( .A(n_517), .B(n_523), .C(n_526), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_520), .Y(n_517) );
INVx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_533), .B(n_536), .Y(n_532) );
NAND3xp33_ASAP7_75t_L g536 ( .A(n_537), .B(n_539), .C(n_541), .Y(n_536) );
INVx1_ASAP7_75t_L g642 ( .A(n_548), .Y(n_642) );
AOI22xp5_ASAP7_75t_SL g548 ( .A1(n_549), .A2(n_550), .B1(n_604), .B2(n_640), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
OAI22xp5_ASAP7_75t_SL g550 ( .A1(n_551), .A2(n_581), .B1(n_582), .B2(n_603), .Y(n_550) );
INVx2_ASAP7_75t_L g603 ( .A(n_551), .Y(n_603) );
XNOR2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_572), .Y(n_553) );
NOR3xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_559), .C(n_568), .Y(n_554) );
OAI222xp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_563), .B1(n_564), .B2(n_565), .C1(n_566), .C2(n_567), .Y(n_559) );
INVx2_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_577), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .Y(n_577) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
XOR2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_602), .Y(n_583) );
NAND3x1_ASAP7_75t_L g584 ( .A(n_585), .B(n_594), .C(n_599), .Y(n_584) );
NOR2x1_ASAP7_75t_L g585 ( .A(n_586), .B(n_589), .Y(n_585) );
NAND3xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .C(n_593), .Y(n_589) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .Y(n_594) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g640 ( .A(n_604), .Y(n_640) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g638 ( .A(n_606), .Y(n_638) );
AND2x2_ASAP7_75t_SL g606 ( .A(n_607), .B(n_621), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_615), .Y(n_607) );
OAI221xp5_ASAP7_75t_SL g608 ( .A1(n_609), .A2(n_610), .B1(n_611), .B2(n_612), .C(n_613), .Y(n_608) );
OAI221xp5_ASAP7_75t_SL g615 ( .A1(n_616), .A2(n_617), .B1(n_618), .B2(n_619), .C(n_620), .Y(n_615) );
NOR3xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_626), .C(n_633), .Y(n_621) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_635), .B1(n_636), .B2(n_637), .Y(n_633) );
INVx1_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
NOR2x1_ASAP7_75t_L g644 ( .A(n_645), .B(n_649), .Y(n_644) );
OR2x2_ASAP7_75t_SL g706 ( .A(n_645), .B(n_650), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_648), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_647), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_647), .B(n_681), .Y(n_684) );
CKINVDCx16_ASAP7_75t_R g681 ( .A(n_648), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
OAI322xp33_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_679), .A3(n_680), .B1(n_682), .B2(n_685), .C1(n_686), .C2(n_704), .Y(n_656) );
INVx2_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
NAND2x1p5_ASAP7_75t_L g659 ( .A(n_660), .B(n_670), .Y(n_659) );
NOR2xp67_ASAP7_75t_SL g660 ( .A(n_661), .B(n_666), .Y(n_660) );
NAND3xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .C(n_664), .Y(n_661) );
OAI21xp5_ASAP7_75t_SL g666 ( .A1(n_667), .A2(n_668), .B(n_669), .Y(n_666) );
NOR2x1_ASAP7_75t_L g670 ( .A(n_671), .B(n_674), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_677), .Y(n_674) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
CKINVDCx16_ASAP7_75t_R g682 ( .A(n_683), .Y(n_682) );
NAND4xp75_ASAP7_75t_L g687 ( .A(n_688), .B(n_692), .C(n_695), .D(n_702), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_691), .Y(n_688) );
AND2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
OA211x2_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B(n_699), .C(n_701), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_705), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_706), .Y(n_705) );
endmodule