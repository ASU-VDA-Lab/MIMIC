module real_jpeg_5863_n_32 (n_17, n_8, n_0, n_21, n_2, n_188, n_185, n_29, n_180, n_10, n_31, n_9, n_186, n_12, n_24, n_189, n_187, n_6, n_28, n_183, n_23, n_11, n_14, n_25, n_7, n_22, n_18, n_3, n_5, n_4, n_181, n_1, n_26, n_27, n_20, n_19, n_182, n_184, n_30, n_16, n_15, n_13, n_32);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_188;
input n_185;
input n_29;
input n_180;
input n_10;
input n_31;
input n_9;
input n_186;
input n_12;
input n_24;
input n_189;
input n_187;
input n_6;
input n_28;
input n_183;
input n_23;
input n_11;
input n_14;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_181;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_182;
input n_184;
input n_30;
input n_16;
input n_15;
input n_13;

output n_32;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_174;
wire n_87;
wire n_173;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_164;
wire n_48;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_150;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

INVx5_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_0),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_1),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_2),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_2),
.B(n_61),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_3),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_4),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_5),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_5),
.B(n_122),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_6),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_6),
.B(n_108),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_7),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_8),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_8),
.B(n_76),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_9),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_9),
.B(n_137),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_10),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_11),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_12),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_13),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_13),
.B(n_161),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_14),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_14),
.B(n_85),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_15),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_16),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_16),
.B(n_67),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_17),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_18),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_19),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_21),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_21),
.B(n_164),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_22),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_22),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_22),
.B(n_53),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_22),
.A2(n_50),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_23),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_23),
.B(n_147),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_24),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_24),
.B(n_88),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_25),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_25),
.B(n_73),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_26),
.B(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_28),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_29),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_30),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_31),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_175),
.Y(n_32)
);

AO21x1_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_42),
.B(n_173),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_36),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

AO21x1_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_51),
.B(n_172),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_50),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_44),
.B(n_50),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_49),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_50),
.B(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_56),
.B(n_171),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_159),
.B(n_168),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_139),
.B(n_153),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_80),
.B(n_127),
.C(n_136),
.Y(n_58)
);

NOR4xp25_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_66),
.C(n_72),
.D(n_75),
.Y(n_59)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_64),
.Y(n_125)
);

BUFx8_ASAP7_75t_L g144 ( 
.A(n_64),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_72),
.A2(n_131),
.B(n_132),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_78),
.B(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_121),
.B(n_126),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_115),
.B(n_120),
.Y(n_81)
);

AO221x1_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_91),
.B1(n_112),
.B2(n_113),
.C(n_114),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_90),
.B(n_109),
.Y(n_108)
);

AO21x1_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_96),
.B(n_111),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_95),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_107),
.B(n_110),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_101),
.B(n_106),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_105),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_119),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_119),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_151),
.Y(n_150)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

A2O1A1O1Ixp25_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B(n_133),
.C(n_134),
.D(n_135),
.Y(n_128)
);

NAND3xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_145),
.C(n_149),
.Y(n_139)
);

A2O1A1O1Ixp25_ASAP7_75t_L g153 ( 
.A1(n_140),
.A2(n_149),
.B(n_154),
.C(n_157),
.D(n_158),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_142),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_146),
.A2(n_155),
.B(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_152),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_180),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_181),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_182),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_183),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_184),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_185),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_186),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_187),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_188),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_189),
.Y(n_123)
);


endmodule