module fake_jpeg_2664_n_545 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_545);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_545;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_14),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_48),
.B(n_64),
.Y(n_103)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_52),
.Y(n_141)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_53),
.Y(n_137)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_55),
.Y(n_130)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_18),
.B(n_11),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_59),
.B(n_87),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_62),
.Y(n_149)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_31),
.B(n_11),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_68),
.Y(n_104)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_66),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_69),
.Y(n_161)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_70),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_72),
.B(n_86),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_73),
.Y(n_145)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_76),
.Y(n_140)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_15),
.Y(n_79)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_82),
.Y(n_157)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx11_ASAP7_75t_SL g85 ( 
.A(n_37),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_85),
.Y(n_138)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_17),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_18),
.B(n_11),
.Y(n_87)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_15),
.Y(n_88)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_25),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_95),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_92),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_27),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_22),
.B(n_10),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_96),
.B(n_16),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_48),
.B(n_39),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_112),
.B(n_143),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_85),
.A2(n_19),
.B1(n_40),
.B2(n_34),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_113),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_118),
.Y(n_187)
);

BUFx2_ASAP7_75t_R g122 ( 
.A(n_74),
.Y(n_122)
);

INVx6_ASAP7_75t_SL g193 ( 
.A(n_122),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_65),
.A2(n_20),
.B1(n_34),
.B2(n_42),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_123),
.A2(n_43),
.B1(n_20),
.B2(n_34),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_126),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_57),
.B(n_43),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_15),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g183 ( 
.A1(n_131),
.A2(n_33),
.B(n_32),
.Y(n_183)
);

INVx6_ASAP7_75t_SL g133 ( 
.A(n_83),
.Y(n_133)
);

CKINVDCx9p33_ASAP7_75t_R g186 ( 
.A(n_133),
.Y(n_186)
);

INVx6_ASAP7_75t_SL g139 ( 
.A(n_89),
.Y(n_139)
);

CKINVDCx12_ASAP7_75t_R g170 ( 
.A(n_139),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_79),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_158),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_94),
.Y(n_143)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_146),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_46),
.B(n_39),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_154),
.B(n_155),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_55),
.B(n_22),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_58),
.B(n_17),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_70),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_166),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_167),
.Y(n_222)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_168),
.Y(n_239)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_171),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_128),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_183),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_136),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_173),
.B(n_175),
.Y(n_220)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_121),
.Y(n_174)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_174),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_132),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_176),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_126),
.A2(n_43),
.B(n_32),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_177),
.A2(n_182),
.B(n_208),
.Y(n_229)
);

CKINVDCx12_ASAP7_75t_R g178 ( 
.A(n_121),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_178),
.Y(n_213)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_137),
.Y(n_179)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

INVx11_ASAP7_75t_L g181 ( 
.A(n_129),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_181),
.A2(n_206),
.B1(n_207),
.B2(n_129),
.Y(n_238)
);

OR2x2_ASAP7_75t_SL g182 ( 
.A(n_103),
.B(n_63),
.Y(n_182)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_129),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_184),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_104),
.B(n_34),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_195),
.Y(n_223)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_117),
.Y(n_188)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_188),
.Y(n_230)
);

AND2x6_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_10),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_194),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_190),
.A2(n_20),
.B1(n_140),
.B2(n_107),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_101),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_191),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_105),
.A2(n_16),
.B1(n_92),
.B2(n_90),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_192),
.A2(n_199),
.B1(n_38),
.B2(n_33),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_109),
.B(n_34),
.Y(n_195)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_106),
.Y(n_196)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_196),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_132),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_202),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_141),
.A2(n_97),
.B1(n_84),
.B2(n_82),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_150),
.Y(n_200)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_200),
.Y(n_218)
);

INVx3_ASAP7_75t_SL g201 ( 
.A(n_119),
.Y(n_201)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_201),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_140),
.B(n_56),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_117),
.Y(n_204)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_106),
.Y(n_205)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_205),
.Y(n_212)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_119),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_120),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_131),
.A2(n_19),
.B1(n_29),
.B2(n_23),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_108),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_125),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_116),
.Y(n_210)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_210),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_180),
.A2(n_113),
.B1(n_73),
.B2(n_71),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_190),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_234),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_232),
.A2(n_236),
.B1(n_243),
.B2(n_246),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_180),
.A2(n_151),
.B1(n_145),
.B2(n_147),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_164),
.A2(n_98),
.B1(n_110),
.B2(n_102),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_240),
.A2(n_242),
.B(n_245),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_177),
.A2(n_98),
.B(n_110),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_185),
.A2(n_151),
.B1(n_145),
.B2(n_147),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_193),
.A2(n_175),
.B1(n_186),
.B2(n_200),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_193),
.A2(n_130),
.B1(n_99),
.B2(n_40),
.Y(n_246)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_218),
.Y(n_248)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_248),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_249),
.A2(n_120),
.B1(n_81),
.B2(n_75),
.Y(n_306)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_214),
.Y(n_250)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_250),
.Y(n_294)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_214),
.Y(n_251)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_251),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_223),
.B(n_169),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_252),
.B(n_266),
.Y(n_280)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_253),
.Y(n_281)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_254),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_186),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_255),
.A2(n_222),
.B(n_142),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_220),
.B(n_162),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_256),
.B(n_262),
.Y(n_286)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_218),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_257),
.B(n_259),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_173),
.Y(n_258)
);

INVxp33_ASAP7_75t_L g291 ( 
.A(n_258),
.Y(n_291)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_225),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_223),
.A2(n_165),
.B1(n_195),
.B2(n_208),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_261),
.A2(n_268),
.B1(n_263),
.B2(n_266),
.Y(n_289)
);

AND2x6_ASAP7_75t_L g262 ( 
.A(n_216),
.B(n_189),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_211),
.B(n_179),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_264),
.B(n_277),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_167),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_265),
.A2(n_271),
.B(n_203),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_224),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_229),
.B(n_182),
.C(n_170),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_204),
.C(n_188),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_229),
.B(n_176),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_270),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_225),
.B(n_168),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_269),
.B(n_273),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_221),
.B(n_239),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_232),
.B(n_236),
.Y(n_271)
);

AND2x6_ASAP7_75t_L g273 ( 
.A(n_219),
.B(n_181),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_221),
.B(n_171),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_275),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_239),
.B(n_207),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_239),
.B(n_228),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_276),
.B(n_241),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_213),
.B(n_167),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_263),
.A2(n_234),
.B1(n_196),
.B2(n_212),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_278),
.A2(n_247),
.B1(n_257),
.B2(n_254),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_213),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_279),
.B(n_285),
.C(n_292),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_272),
.A2(n_222),
.B(n_228),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_282),
.A2(n_265),
.B(n_271),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_255),
.A2(n_187),
.B(n_231),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_283),
.A2(n_290),
.B(n_295),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_227),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_289),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_255),
.A2(n_187),
.B(n_231),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_293),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_263),
.A2(n_235),
.B1(n_226),
.B2(n_166),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_249),
.A2(n_244),
.B1(n_217),
.B2(n_163),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_296),
.A2(n_306),
.B1(n_271),
.B2(n_217),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_298),
.A2(n_299),
.B(n_303),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_272),
.A2(n_222),
.B(n_235),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_267),
.B(n_227),
.C(n_230),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_300),
.B(n_302),
.C(n_275),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_250),
.B(n_230),
.C(n_226),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_251),
.A2(n_184),
.B(n_241),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_270),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_274),
.Y(n_309)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_309),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_310),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_307),
.Y(n_311)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_311),
.Y(n_353)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_307),
.Y(n_312)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_312),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_276),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_313),
.B(n_322),
.C(n_330),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_305),
.Y(n_314)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_314),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_315),
.B(n_327),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_248),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_316),
.B(n_318),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_317),
.A2(n_284),
.B(n_281),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_280),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_287),
.A2(n_247),
.B1(n_265),
.B2(n_273),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_319),
.A2(n_331),
.B1(n_287),
.B2(n_317),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_308),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_320),
.B(n_338),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_285),
.B(n_259),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_321),
.B(n_293),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_300),
.B(n_262),
.Y(n_322)
);

AND2x6_ASAP7_75t_L g323 ( 
.A(n_286),
.B(n_260),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_323),
.B(n_326),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_281),
.Y(n_325)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_325),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_303),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_294),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_328),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_280),
.B(n_253),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_332),
.B(n_336),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_298),
.B(n_260),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_333),
.B(n_337),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_308),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_335),
.B(n_302),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_288),
.B(n_167),
.Y(n_336)
);

OR2x2_ASAP7_75t_L g337 ( 
.A(n_288),
.B(n_198),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_279),
.B(n_35),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_292),
.B(n_206),
.C(n_130),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_339),
.B(n_340),
.C(n_304),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_285),
.B(n_174),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_342),
.B(n_349),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_346),
.A2(n_350),
.B1(n_366),
.B2(n_340),
.Y(n_389)
);

INVx5_ASAP7_75t_L g347 ( 
.A(n_325),
.Y(n_347)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_347),
.Y(n_383)
);

AO22x1_ASAP7_75t_SL g348 ( 
.A1(n_327),
.A2(n_315),
.B1(n_278),
.B2(n_312),
.Y(n_348)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_348),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_322),
.B(n_286),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_319),
.A2(n_299),
.B1(n_290),
.B2(n_283),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_329),
.B(n_282),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_351),
.B(n_321),
.Y(n_396)
);

CKINVDCx14_ASAP7_75t_R g378 ( 
.A(n_355),
.Y(n_378)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_325),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_359),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_360),
.B(n_367),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_318),
.B(n_330),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_363),
.B(n_364),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_338),
.B(n_301),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_326),
.A2(n_295),
.B1(n_296),
.B2(n_306),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_329),
.B(n_282),
.C(n_301),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_333),
.B(n_311),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_368),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_309),
.B(n_294),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_369),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_332),
.B(n_304),
.Y(n_370)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_370),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_336),
.B(n_284),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_371),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_374),
.A2(n_324),
.B(n_341),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_375),
.A2(n_397),
.B(n_403),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_344),
.A2(n_337),
.B1(n_314),
.B2(n_323),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_376),
.A2(n_386),
.B1(n_399),
.B2(n_400),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_352),
.A2(n_337),
.B1(n_313),
.B2(n_316),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_380),
.A2(n_381),
.B1(n_389),
.B2(n_392),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_344),
.A2(n_310),
.B1(n_323),
.B2(n_328),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_373),
.Y(n_382)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_382),
.Y(n_415)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_373),
.Y(n_385)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_385),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_344),
.A2(n_333),
.B1(n_334),
.B2(n_324),
.Y(n_386)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_372),
.Y(n_388)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_388),
.Y(n_424)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_372),
.Y(n_390)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_390),
.Y(n_425)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_358),
.Y(n_391)
);

BUFx4f_ASAP7_75t_SL g422 ( 
.A(n_391),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_346),
.A2(n_350),
.B1(n_365),
.B2(n_354),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_357),
.A2(n_362),
.B1(n_365),
.B2(n_354),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_393),
.A2(n_394),
.B1(n_348),
.B2(n_366),
.Y(n_419)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_361),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_396),
.B(n_356),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_345),
.A2(n_341),
.B(n_339),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_361),
.A2(n_260),
.B1(n_281),
.B2(n_212),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_345),
.A2(n_260),
.B1(n_215),
.B2(n_212),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_345),
.A2(n_215),
.B1(n_217),
.B2(n_244),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_401),
.A2(n_343),
.B1(n_205),
.B2(n_191),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_368),
.A2(n_198),
.B(n_215),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_407),
.B(n_414),
.Y(n_457)
);

FAx1_ASAP7_75t_SL g408 ( 
.A(n_376),
.B(n_367),
.CI(n_349),
.CON(n_408),
.SN(n_408)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_408),
.B(n_409),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_378),
.B(n_356),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_379),
.B(n_360),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_410),
.B(n_420),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_405),
.B(n_353),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_411),
.B(n_416),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_386),
.A2(n_377),
.B1(n_387),
.B2(n_368),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_413),
.A2(n_426),
.B1(n_433),
.B2(n_403),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_402),
.B(n_351),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_396),
.B(n_342),
.C(n_374),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_392),
.A2(n_347),
.B(n_359),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_417),
.B(n_427),
.Y(n_436)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_419),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_348),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_377),
.A2(n_343),
.B1(n_244),
.B2(n_210),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_423),
.A2(n_401),
.B1(n_383),
.B2(n_400),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_397),
.B(n_201),
.C(n_99),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_387),
.B(n_146),
.C(n_115),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_428),
.B(n_429),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_404),
.B(n_115),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_382),
.B(n_161),
.C(n_149),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_430),
.B(n_431),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_385),
.B(n_161),
.C(n_149),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_384),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_432),
.B(n_124),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_389),
.A2(n_134),
.B1(n_116),
.B2(n_157),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_421),
.A2(n_413),
.B1(n_424),
.B2(n_425),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_435),
.B(n_441),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_437),
.Y(n_463)
);

AOI322xp5_ASAP7_75t_L g438 ( 
.A1(n_415),
.A2(n_398),
.A3(n_394),
.B1(n_395),
.B2(n_388),
.C1(n_390),
.C2(n_391),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_438),
.B(n_431),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_422),
.Y(n_441)
);

AOI21x1_ASAP7_75t_L g442 ( 
.A1(n_412),
.A2(n_375),
.B(n_383),
.Y(n_442)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_442),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_443),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_406),
.A2(n_399),
.B1(n_134),
.B2(n_153),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_444),
.A2(n_426),
.B1(n_433),
.B2(n_422),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_410),
.B(n_69),
.C(n_62),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_445),
.B(n_452),
.C(n_455),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_420),
.B(n_60),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_447),
.B(n_449),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_412),
.B(n_416),
.Y(n_449)
);

NOR2xp67_ASAP7_75t_SL g450 ( 
.A(n_407),
.B(n_127),
.Y(n_450)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_450),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_414),
.B(n_51),
.C(n_50),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_418),
.B(n_47),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_453),
.B(n_458),
.Y(n_461)
);

INVx13_ASAP7_75t_L g454 ( 
.A(n_422),
.Y(n_454)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_454),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_427),
.B(n_35),
.C(n_33),
.Y(n_455)
);

CKINVDCx14_ASAP7_75t_R g471 ( 
.A(n_456),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_421),
.B(n_157),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_439),
.B(n_408),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_460),
.B(n_478),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_464),
.A2(n_468),
.B1(n_470),
.B2(n_111),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_435),
.A2(n_434),
.B(n_440),
.Y(n_467)
);

NAND3xp33_ASAP7_75t_SL g482 ( 
.A(n_467),
.B(n_455),
.C(n_23),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_443),
.A2(n_408),
.B1(n_423),
.B2(n_430),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_453),
.B(n_428),
.Y(n_469)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_469),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_444),
.A2(n_436),
.B1(n_451),
.B2(n_458),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_446),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_472),
.B(n_473),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_439),
.B(n_124),
.Y(n_475)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_475),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_449),
.B(n_457),
.C(n_447),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_477),
.B(n_470),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_445),
.B(n_160),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_465),
.A2(n_457),
.B(n_448),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_480),
.A2(n_476),
.B(n_474),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_463),
.B(n_452),
.C(n_454),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_481),
.B(n_484),
.Y(n_510)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_482),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_479),
.B(n_93),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_467),
.A2(n_93),
.B1(n_29),
.B2(n_23),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_485),
.B(n_486),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_477),
.B(n_135),
.C(n_100),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_466),
.B(n_135),
.C(n_100),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_487),
.B(n_495),
.C(n_464),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_459),
.B(n_29),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_488),
.B(n_494),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_490),
.B(n_496),
.C(n_474),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_459),
.B(n_114),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_491),
.B(n_492),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_462),
.B(n_15),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_468),
.B(n_38),
.C(n_41),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_460),
.B(n_40),
.Y(n_496)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_500),
.Y(n_516)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_502),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_503),
.B(n_507),
.Y(n_515)
);

FAx1_ASAP7_75t_L g504 ( 
.A(n_493),
.B(n_461),
.CI(n_471),
.CON(n_504),
.SN(n_504)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_504),
.A2(n_505),
.B(n_506),
.Y(n_514)
);

A2O1A1Ixp33_ASAP7_75t_L g505 ( 
.A1(n_483),
.A2(n_469),
.B(n_461),
.C(n_478),
.Y(n_505)
);

A2O1A1Ixp33_ASAP7_75t_L g506 ( 
.A1(n_493),
.A2(n_10),
.B(n_9),
.C(n_38),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_489),
.A2(n_10),
.B(n_9),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_481),
.B(n_41),
.C(n_9),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_509),
.B(n_0),
.Y(n_517)
);

AOI31xp67_ASAP7_75t_L g511 ( 
.A1(n_495),
.A2(n_0),
.A3(n_1),
.B(n_2),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_511),
.A2(n_512),
.B1(n_1),
.B2(n_2),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_L g512 ( 
.A1(n_497),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_504),
.A2(n_496),
.B1(n_491),
.B2(n_488),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_513),
.B(n_518),
.Y(n_525)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_517),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g518 ( 
.A(n_504),
.Y(n_518)
);

AOI322xp5_ASAP7_75t_L g519 ( 
.A1(n_510),
.A2(n_487),
.A3(n_486),
.B1(n_3),
.B2(n_4),
.C1(n_1),
.C2(n_6),
.Y(n_519)
);

AO21x1_ASAP7_75t_L g531 ( 
.A1(n_519),
.A2(n_3),
.B(n_4),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_520),
.B(n_524),
.Y(n_529)
);

NOR2xp67_ASAP7_75t_L g521 ( 
.A(n_501),
.B(n_2),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_521),
.A2(n_522),
.B(n_506),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_505),
.A2(n_3),
.B(n_4),
.Y(n_522)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_499),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_516),
.B(n_508),
.C(n_503),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_526),
.B(n_527),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_523),
.B(n_508),
.C(n_498),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_528),
.A2(n_531),
.B(n_522),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_515),
.B(n_512),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_530),
.A2(n_514),
.B(n_5),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_533),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_525),
.A2(n_514),
.B1(n_513),
.B2(n_6),
.Y(n_534)
);

OAI21xp33_ASAP7_75t_L g540 ( 
.A1(n_534),
.A2(n_535),
.B(n_5),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_529),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_537)
);

OAI31xp33_ASAP7_75t_L g539 ( 
.A1(n_537),
.A2(n_532),
.A3(n_529),
.B(n_8),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_539),
.A2(n_540),
.B(n_536),
.Y(n_541)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_541),
.Y(n_543)
);

MAJx2_ASAP7_75t_L g542 ( 
.A(n_538),
.B(n_5),
.C(n_8),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_543),
.B(n_542),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_544),
.B(n_5),
.Y(n_545)
);


endmodule