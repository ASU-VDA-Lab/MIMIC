module real_jpeg_26526_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_327, n_1, n_328, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_327;
input n_1;
input n_328;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_0),
.A2(n_55),
.B1(n_57),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_0),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_0),
.A2(n_38),
.B1(n_39),
.B2(n_87),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_0),
.A2(n_31),
.B1(n_32),
.B2(n_87),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_0),
.A2(n_64),
.B1(n_70),
.B2(n_87),
.Y(n_295)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_1),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_2),
.A2(n_55),
.B1(n_57),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_2),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_2),
.A2(n_38),
.B1(n_39),
.B2(n_83),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_83),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_2),
.A2(n_64),
.B1(n_70),
.B2(n_83),
.Y(n_280)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_4),
.A2(n_55),
.B1(n_57),
.B2(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_4),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_4),
.A2(n_38),
.B1(n_39),
.B2(n_129),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_129),
.Y(n_298)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_5),
.A2(n_38),
.B1(n_39),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_5),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_5),
.A2(n_55),
.B1(n_57),
.B2(n_60),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_60),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_5),
.A2(n_60),
.B1(n_64),
.B2(n_70),
.Y(n_258)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_7),
.A2(n_64),
.B1(n_70),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_7),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_74),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_7),
.A2(n_38),
.B1(n_39),
.B2(n_74),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_7),
.A2(n_55),
.B1(n_57),
.B2(n_74),
.Y(n_175)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_9),
.A2(n_38),
.B1(n_39),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_49),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_9),
.A2(n_49),
.B1(n_55),
.B2(n_57),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_9),
.A2(n_49),
.B1(n_64),
.B2(n_70),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_10),
.A2(n_44),
.B1(n_64),
.B2(n_70),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_10),
.A2(n_44),
.B1(n_55),
.B2(n_57),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_10),
.A2(n_38),
.B1(n_39),
.B2(n_44),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_42),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_11),
.A2(n_42),
.B1(n_64),
.B2(n_70),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_11),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_11),
.A2(n_42),
.B1(n_55),
.B2(n_57),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_12),
.A2(n_55),
.B1(n_57),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_12),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_12),
.A2(n_38),
.B1(n_39),
.B2(n_108),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_108),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_12),
.A2(n_64),
.B1(n_70),
.B2(n_108),
.Y(n_319)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_14),
.A2(n_64),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_14),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_SL g77 ( 
.A1(n_14),
.A2(n_32),
.B(n_65),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_14),
.B(n_67),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_14),
.A2(n_38),
.B(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_14),
.B(n_38),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_14),
.B(n_94),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_14),
.A2(n_81),
.B1(n_105),
.B2(n_175),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_14),
.A2(n_31),
.B(n_190),
.Y(n_189)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_16),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

INVx11_ASAP7_75t_SL g56 ( 
.A(n_17),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_307),
.Y(n_18)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_275),
.A3(n_302),
.B1(n_305),
.B2(n_306),
.C(n_327),
.Y(n_19)
);

AOI321xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_226),
.A3(n_264),
.B1(n_269),
.B2(n_274),
.C(n_328),
.Y(n_20)
);

NOR3xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_121),
.C(n_140),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_98),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_23),
.B(n_98),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_75),
.C(n_88),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_24),
.B(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_62),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_45),
.B2(n_46),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_26),
.B(n_46),
.C(n_62),
.Y(n_109)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_37),
.B1(n_40),
.B2(n_43),
.Y(n_27)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_28),
.A2(n_37),
.B1(n_43),
.B2(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_28),
.A2(n_37),
.B1(n_92),
.B2(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_28),
.A2(n_37),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_28),
.A2(n_37),
.B(n_315),
.Y(n_314)
);

A2O1A1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_31),
.B(n_34),
.C(n_37),
.Y(n_28)
);

OAI32xp33_ASAP7_75t_L g198 ( 
.A1(n_29),
.A2(n_31),
.A3(n_39),
.B1(n_191),
.B2(n_199),
.Y(n_198)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_29),
.Y(n_200)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_35),
.Y(n_34)
);

AO22x1_ASAP7_75t_L g67 ( 
.A1(n_31),
.A2(n_32),
.B1(n_65),
.B2(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_32),
.B(n_71),
.Y(n_191)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_39),
.B1(n_53),
.B2(n_54),
.Y(n_58)
);

OAI32xp33_ASAP7_75t_L g152 ( 
.A1(n_38),
.A2(n_53),
.A3(n_57),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_38),
.B(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_41),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_90)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B1(n_59),
.B2(n_61),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_48),
.A2(n_51),
.B1(n_52),
.B2(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_50),
.A2(n_61),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_50),
.A2(n_61),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_51),
.A2(n_52),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_51),
.A2(n_52),
.B1(n_103),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_51),
.A2(n_52),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_51),
.A2(n_52),
.B1(n_150),
.B2(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_51),
.A2(n_52),
.B1(n_239),
.B2(n_251),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_51),
.A2(n_52),
.B(n_251),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_58),
.Y(n_51)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_52),
.B(n_71),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_54),
.B(n_55),
.Y(n_154)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_55),
.B(n_180),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_59),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_67),
.B1(n_69),
.B2(n_72),
.Y(n_62)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_63),
.A2(n_67),
.B1(n_116),
.B2(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_63),
.A2(n_67),
.B1(n_136),
.B2(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_63),
.A2(n_67),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

O2A1O1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B(n_66),
.C(n_67),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_SL g66 ( 
.A(n_64),
.B(n_65),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_64),
.Y(n_70)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_67),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_70),
.B(n_71),
.C(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_71),
.B(n_85),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_73),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_75),
.A2(n_88),
.B1(n_89),
.B2(n_224),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_75),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_76),
.B(n_78),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B1(n_84),
.B2(n_86),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_80),
.B1(n_82),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_79),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_79),
.A2(n_80),
.B1(n_168),
.B2(n_170),
.Y(n_167)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_85),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_85),
.A2(n_105),
.B1(n_107),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_85),
.A2(n_105),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_85),
.A2(n_105),
.B1(n_169),
.B2(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_85),
.A2(n_105),
.B1(n_164),
.B2(n_202),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_85),
.A2(n_105),
.B(n_128),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_86),
.Y(n_106)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_95),
.C(n_97),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_90),
.B(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_93),
.A2(n_94),
.B1(n_119),
.B2(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_93),
.A2(n_94),
.B1(n_138),
.B2(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_93),
.A2(n_94),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_93),
.A2(n_94),
.B1(n_284),
.B2(n_298),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_95),
.B(n_97),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_96),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_110),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_109),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_109),
.C(n_110),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_104),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_120),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_117),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_117),
.C(n_120),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_113),
.A2(n_114),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_113),
.A2(n_114),
.B1(n_258),
.B2(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_113),
.A2(n_114),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_L g270 ( 
.A1(n_122),
.A2(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_123),
.B(n_124),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_139),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_132),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_126),
.B(n_132),
.C(n_139),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_127),
.B(n_130),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_131),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_133),
.B(n_135),
.C(n_137),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_220),
.B(n_225),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_206),
.B(n_219),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_184),
.B(n_205),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_165),
.B(n_183),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_155),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_145),
.B(n_155),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_151),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_146),
.A2(n_147),
.B1(n_151),
.B2(n_152),
.Y(n_171)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_149),
.Y(n_153)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_162),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_160),
.C(n_162),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_161),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_163),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_172),
.B(n_182),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_171),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_167),
.B(n_171),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_177),
.B(n_181),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_174),
.B(n_176),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_185),
.B(n_186),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_197),
.B1(n_203),
.B2(n_204),
.Y(n_186)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_192),
.B1(n_195),
.B2(n_196),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_188),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_192),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_196),
.C(n_204),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_194),
.Y(n_216)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_197),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_201),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_207),
.B(n_208),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_212),
.B2(n_213),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_215),
.C(n_217),
.Y(n_221)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_217),
.B2(n_218),
.Y(n_213)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_214),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_221),
.B(n_222),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_243),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_227),
.B(n_243),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_234),
.C(n_242),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_228),
.B(n_234),
.Y(n_268)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_228),
.Y(n_324)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_231),
.CI(n_233),
.CON(n_228),
.SN(n_228)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_231),
.C(n_233),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_230),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_232),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_240),
.B2(n_241),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_235),
.B(n_241),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_240),
.A2(n_241),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_240),
.A2(n_256),
.B(n_259),
.Y(n_289)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_268),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_262),
.B2(n_263),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_253),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_246),
.B(n_253),
.C(n_263),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_250),
.B(n_252),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_250),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_249),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_277),
.C(n_289),
.Y(n_276)
);

FAx1_ASAP7_75t_SL g304 ( 
.A(n_252),
.B(n_277),
.CI(n_289),
.CON(n_304),
.SN(n_304)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_259),
.B1(n_260),
.B2(n_261),
.Y(n_253)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_254),
.Y(n_261)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_262),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_265),
.A2(n_270),
.B(n_273),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_266),
.B(n_267),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_290),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_276),
.B(n_290),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_281),
.B2(n_288),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_278),
.A2(n_279),
.B1(n_292),
.B2(n_300),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_282),
.C(n_287),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_279),
.B(n_300),
.C(n_301),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_280),
.Y(n_294)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_281),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_281)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_282),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_285),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_285),
.A2(n_287),
.B1(n_297),
.B2(n_299),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_285),
.B(n_293),
.C(n_297),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_301),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_292),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_296),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_295),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_297),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_298),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_303),
.B(n_304),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_304),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_322),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_310),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_312),
.B1(n_320),
.B2(n_321),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_316),
.B2(n_317),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_314),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_317),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_321),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);


endmodule