module fake_jpeg_13740_n_110 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_3),
.B(n_4),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_5),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_29),
.B(n_30),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_7),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_32),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_0),
.C(n_1),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_L g35 ( 
.A1(n_20),
.A2(n_1),
.B(n_3),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_35),
.B(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_37),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_7),
.Y(n_37)
);

NAND2xp33_ASAP7_75t_SL g38 ( 
.A(n_23),
.B(n_8),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_41),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_11),
.C(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_15),
.B(n_19),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_13),
.B(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_44),
.Y(n_53)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_46),
.B(n_24),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_22),
.A2(n_20),
.B1(n_24),
.B2(n_23),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_22),
.B1(n_27),
.B2(n_12),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_16),
.B(n_21),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_30),
.B(n_43),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_60),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_62),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_36),
.B1(n_34),
.B2(n_33),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_32),
.B(n_18),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_64),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_44),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_38),
.B(n_28),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_65),
.B(n_67),
.Y(n_90)
);

FAx1_ASAP7_75t_SL g70 ( 
.A(n_56),
.B(n_53),
.CI(n_60),
.CON(n_70),
.SN(n_70)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_50),
.C(n_54),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_77),
.B1(n_80),
.B2(n_81),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_57),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_74),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_40),
.B1(n_45),
.B2(n_52),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_65),
.B1(n_67),
.B2(n_51),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_52),
.A2(n_54),
.B1(n_55),
.B2(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_58),
.Y(n_78)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_82),
.B(n_84),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_70),
.C(n_77),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_70),
.B1(n_74),
.B2(n_69),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_89),
.B1(n_73),
.B2(n_80),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_90),
.B(n_71),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_71),
.B1(n_76),
.B2(n_72),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_92),
.A2(n_94),
.B(n_90),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_86),
.B(n_72),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_96),
.C(n_92),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_100),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_82),
.C(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_83),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_85),
.B1(n_96),
.B2(n_88),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_103),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_101),
.A2(n_87),
.B1(n_83),
.B2(n_81),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_102),
.C(n_51),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_106),
.Y(n_108)
);

FAx1_ASAP7_75t_SL g107 ( 
.A(n_104),
.B(n_66),
.CI(n_105),
.CON(n_107),
.SN(n_107)
);

AOI322xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_66),
.A3(n_106),
.B1(n_107),
.B2(n_93),
.C1(n_101),
.C2(n_98),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_106),
.Y(n_110)
);


endmodule