module fake_jpeg_30373_n_178 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_178);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_7),
.B(n_35),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_30),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_72),
.Y(n_86)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_75),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_49),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_68),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_0),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_55),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_81),
.Y(n_96)
);

BUFx8_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_93),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_46),
.B1(n_59),
.B2(n_61),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_59),
.B1(n_61),
.B2(n_65),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_55),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_88),
.B(n_92),
.Y(n_111)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_71),
.A2(n_52),
.B1(n_65),
.B2(n_50),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_90),
.A2(n_52),
.B1(n_53),
.B2(n_64),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_74),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_56),
.B(n_62),
.C(n_63),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_95),
.B(n_100),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_97),
.A2(n_106),
.B1(n_96),
.B2(n_109),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_87),
.B(n_66),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_47),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_86),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_58),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_105),
.A2(n_1),
.B(n_2),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_81),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_106),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_90),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_110),
.Y(n_123)
);

BUFx4f_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_67),
.C(n_57),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_121),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_19),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_115),
.A2(n_124),
.B1(n_134),
.B2(n_16),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_99),
.B(n_22),
.Y(n_116)
);

NOR3xp33_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_6),
.C(n_9),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_1),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_98),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

BUFx24_ASAP7_75t_SL g130 ( 
.A(n_111),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_130),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_96),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_11),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_3),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_133),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_4),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_108),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_138),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_119),
.B(n_10),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_141),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_13),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_142),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_120),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_146),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_116),
.B(n_127),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_149),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_128),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_148),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_17),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_152),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_SL g151 ( 
.A1(n_125),
.A2(n_118),
.B(n_122),
.C(n_23),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_151),
.A2(n_153),
.B1(n_125),
.B2(n_21),
.Y(n_159)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_140),
.C(n_135),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_157),
.B(n_161),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_159),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_20),
.C(n_25),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_163),
.B(n_33),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_156),
.A2(n_151),
.B1(n_149),
.B2(n_143),
.Y(n_164)
);

OA21x2_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_166),
.B(n_154),
.Y(n_169)
);

XNOR2x1_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_147),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_168),
.A2(n_159),
.B(n_160),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_169),
.B(n_170),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_171),
.B(n_139),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_165),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_167),
.B(n_155),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_167),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_162),
.C(n_151),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_161),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_37),
.Y(n_178)
);


endmodule