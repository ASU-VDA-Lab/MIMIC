module fake_ariane_2186_n_2106 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_598, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_587, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_588, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_579, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_601, n_565, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_575, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_606, n_213, n_110, n_304, n_67, n_509, n_583, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_573, n_127, n_531, n_2106);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_587;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_588;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_601;
input n_565;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_575;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_583;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;

output n_2106;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_1383;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_1713;
wire n_1436;
wire n_690;
wire n_1109;
wire n_1430;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_1682;
wire n_1836;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_813;
wire n_1985;
wire n_995;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_770;
wire n_1514;
wire n_1528;
wire n_901;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_1703;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_661;
wire n_2098;
wire n_1751;
wire n_1917;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_1432;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_652;
wire n_1819;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_696;
wire n_1442;
wire n_798;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_2087;
wire n_931;
wire n_669;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_632;
wire n_650;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_1578;
wire n_1455;
wire n_836;
wire n_1279;
wire n_1029;
wire n_1247;
wire n_760;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_706;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_670;
wire n_1826;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_2059;
wire n_1439;
wire n_814;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_1899;
wire n_1467;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_677;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_727;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_1156;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_1402;
wire n_957;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_1005;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_1708;
wire n_1222;
wire n_1844;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_890;
wire n_842;
wire n_1898;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_1783;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_1406;
wire n_1405;
wire n_1757;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_1281;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_1154;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_802;
wire n_1151;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_2020;
wire n_748;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_1165;
wire n_1641;
wire n_1517;
wire n_2036;
wire n_843;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_1362;
wire n_1559;
wire n_683;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_1038;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_1695;
wire n_1164;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_1789;
wire n_763;
wire n_1986;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_1579;
wire n_2014;
wire n_975;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_1775;
wire n_908;
wire n_788;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_1537;
wire n_2065;
wire n_1077;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_917;
wire n_1271;
wire n_2096;
wire n_1530;
wire n_631;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_1813;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_1344;
wire n_1390;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_1150;
wire n_977;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_1136;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_1967;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_768;
wire n_1091;
wire n_2052;
wire n_1063;
wire n_991;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_937;
wire n_1474;
wire n_2081;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_849;
wire n_2095;
wire n_1820;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_796;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_292),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_127),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_159),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_564),
.Y(n_615)
);

CKINVDCx16_ASAP7_75t_R g616 ( 
.A(n_607),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_211),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_595),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_246),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_308),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_358),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_462),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_387),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_31),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_216),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_588),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_535),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_516),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g629 ( 
.A(n_296),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_585),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_374),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_72),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_517),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_489),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_169),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_380),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_65),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_439),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_547),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_321),
.Y(n_640)
);

CKINVDCx16_ASAP7_75t_R g641 ( 
.A(n_415),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_286),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_537),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_417),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_179),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_575),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_217),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_567),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_82),
.Y(n_649)
);

INVx1_ASAP7_75t_SL g650 ( 
.A(n_130),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_252),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_221),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_172),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_475),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_555),
.Y(n_655)
);

INVxp67_ASAP7_75t_SL g656 ( 
.A(n_501),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_105),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_337),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_457),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_260),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_531),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_509),
.Y(n_662)
);

BUFx10_ASAP7_75t_L g663 ( 
.A(n_566),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_583),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_505),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_278),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_129),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_83),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_574),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_0),
.Y(n_670)
);

BUFx6f_ASAP7_75t_L g671 ( 
.A(n_277),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_422),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_361),
.Y(n_673)
);

CKINVDCx16_ASAP7_75t_R g674 ( 
.A(n_478),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_573),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_399),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_210),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_571),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_552),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_437),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_391),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_606),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_587),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_601),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_550),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_108),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_579),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_539),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_440),
.Y(n_689)
);

CKINVDCx14_ASAP7_75t_R g690 ( 
.A(n_251),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_504),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_568),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_580),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_448),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_519),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_597),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_312),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_102),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_594),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_590),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_70),
.Y(n_701)
);

CKINVDCx20_ASAP7_75t_R g702 ( 
.A(n_178),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_610),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_490),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_514),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_543),
.Y(n_706)
);

INVx1_ASAP7_75t_SL g707 ( 
.A(n_364),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_542),
.Y(n_708)
);

CKINVDCx20_ASAP7_75t_R g709 ( 
.A(n_548),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_185),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_313),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_429),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_551),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_194),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_416),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_70),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_463),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_545),
.Y(n_718)
);

BUFx2_ASAP7_75t_L g719 ( 
.A(n_599),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_190),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_577),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_294),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_522),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_32),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_268),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_556),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_538),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_559),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_395),
.Y(n_729)
);

CKINVDCx20_ASAP7_75t_R g730 ( 
.A(n_226),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_565),
.Y(n_731)
);

BUFx10_ASAP7_75t_L g732 ( 
.A(n_234),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_372),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_609),
.Y(n_734)
);

INVx1_ASAP7_75t_SL g735 ( 
.A(n_561),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_282),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_512),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_549),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_46),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_335),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_602),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_405),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_608),
.Y(n_743)
);

INVx1_ASAP7_75t_SL g744 ( 
.A(n_524),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_491),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_347),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_289),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_503),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_584),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_371),
.Y(n_750)
);

BUFx5_ASAP7_75t_L g751 ( 
.A(n_467),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_215),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_344),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_600),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_122),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_397),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_160),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_231),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_438),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_582),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_339),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_558),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_246),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_560),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_240),
.Y(n_765)
);

INVx1_ASAP7_75t_SL g766 ( 
.A(n_61),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_557),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_404),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_591),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_593),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_136),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_510),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_569),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_541),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_605),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_56),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_544),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_142),
.Y(n_778)
);

BUFx10_ASAP7_75t_L g779 ( 
.A(n_481),
.Y(n_779)
);

CKINVDCx16_ASAP7_75t_R g780 ( 
.A(n_527),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_520),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_145),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_518),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_123),
.Y(n_784)
);

CKINVDCx20_ASAP7_75t_R g785 ( 
.A(n_497),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_495),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_423),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_532),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_411),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_332),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_611),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_554),
.Y(n_792)
);

BUFx2_ASAP7_75t_L g793 ( 
.A(n_435),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_521),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_170),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_506),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_563),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_471),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_148),
.Y(n_799)
);

CKINVDCx16_ASAP7_75t_R g800 ( 
.A(n_359),
.Y(n_800)
);

INVxp67_ASAP7_75t_L g801 ( 
.A(n_586),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_298),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_403),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_47),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_576),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_578),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_250),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_333),
.Y(n_808)
);

CKINVDCx16_ASAP7_75t_R g809 ( 
.A(n_534),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_581),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_249),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_528),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_49),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_128),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_1),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_418),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_493),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_562),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_572),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_492),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_459),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_445),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_446),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_540),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_553),
.Y(n_825)
);

CKINVDCx16_ASAP7_75t_R g826 ( 
.A(n_125),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_432),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_8),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_598),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_264),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_135),
.Y(n_831)
);

BUFx5_ASAP7_75t_L g832 ( 
.A(n_187),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_447),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_181),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_409),
.Y(n_835)
);

CKINVDCx20_ASAP7_75t_R g836 ( 
.A(n_208),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_536),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_44),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_368),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_570),
.Y(n_840)
);

BUFx10_ASAP7_75t_L g841 ( 
.A(n_592),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_596),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_201),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_376),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_589),
.Y(n_845)
);

CKINVDCx16_ASAP7_75t_R g846 ( 
.A(n_276),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_603),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_460),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_108),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_309),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_287),
.Y(n_851)
);

CKINVDCx20_ASAP7_75t_R g852 ( 
.A(n_266),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_45),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_456),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_30),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_267),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_103),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_507),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_523),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_455),
.Y(n_860)
);

BUFx10_ASAP7_75t_L g861 ( 
.A(n_172),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_494),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_533),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_236),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_499),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_444),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_525),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_234),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_280),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_198),
.Y(n_870)
);

INVx1_ASAP7_75t_SL g871 ( 
.A(n_604),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_267),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_205),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_546),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_684),
.Y(n_875)
);

INVxp67_ASAP7_75t_SL g876 ( 
.A(n_671),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_832),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_832),
.Y(n_878)
);

CKINVDCx16_ASAP7_75t_R g879 ( 
.A(n_690),
.Y(n_879)
);

CKINVDCx20_ASAP7_75t_R g880 ( 
.A(n_695),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_826),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_832),
.Y(n_882)
);

CKINVDCx20_ASAP7_75t_R g883 ( 
.A(n_706),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_677),
.Y(n_884)
);

CKINVDCx20_ASAP7_75t_R g885 ( 
.A(n_709),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_785),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_846),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_832),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_613),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_614),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_617),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_832),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_625),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_619),
.Y(n_894)
);

INVxp33_ASAP7_75t_L g895 ( 
.A(n_624),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_765),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_635),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_632),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_637),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_652),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_876),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_895),
.B(n_616),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_877),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_879),
.B(n_641),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_878),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_882),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_888),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_892),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_894),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_897),
.Y(n_910)
);

AND2x6_ASAP7_75t_L g911 ( 
.A(n_899),
.B(n_712),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_896),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_875),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_889),
.B(n_674),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_875),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_890),
.B(n_891),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_893),
.Y(n_917)
);

OR2x2_ASAP7_75t_L g918 ( 
.A(n_884),
.B(n_645),
.Y(n_918)
);

NAND2x1_ASAP7_75t_L g919 ( 
.A(n_898),
.B(n_712),
.Y(n_919)
);

BUFx8_ASAP7_75t_L g920 ( 
.A(n_900),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_881),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_887),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_880),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_883),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_885),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_886),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_L g927 ( 
.A1(n_903),
.A2(n_703),
.B1(n_793),
.B2(n_719),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_917),
.B(n_780),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_901),
.B(n_800),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_905),
.B(n_809),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_908),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_L g932 ( 
.A1(n_914),
.A2(n_647),
.B1(n_815),
.B2(n_799),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_906),
.B(n_773),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_902),
.B(n_702),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_907),
.B(n_850),
.Y(n_935)
);

OR2x2_ASAP7_75t_L g936 ( 
.A(n_918),
.B(n_650),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_908),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_911),
.B(n_629),
.Y(n_938)
);

OR2x6_ASAP7_75t_L g939 ( 
.A(n_923),
.B(n_667),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_911),
.B(n_707),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_921),
.B(n_801),
.Y(n_941)
);

OR2x6_ASAP7_75t_L g942 ( 
.A(n_924),
.B(n_925),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_916),
.B(n_642),
.Y(n_943)
);

AOI22xp33_ASAP7_75t_L g944 ( 
.A1(n_911),
.A2(n_758),
.B1(n_778),
.B2(n_736),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_922),
.B(n_732),
.Y(n_945)
);

OR2x6_ASAP7_75t_L g946 ( 
.A(n_926),
.B(n_843),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_915),
.B(n_730),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_910),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_915),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_909),
.B(n_913),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_912),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_919),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_904),
.B(n_735),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_920),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_908),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_916),
.B(n_649),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_902),
.B(n_732),
.Y(n_957)
);

AND2x6_ASAP7_75t_L g958 ( 
.A(n_916),
.B(n_630),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_915),
.Y(n_959)
);

INVx2_ASAP7_75t_SL g960 ( 
.A(n_902),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_915),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_902),
.B(n_836),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_910),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_910),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_902),
.B(n_852),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_910),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_929),
.B(n_928),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_948),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_963),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_964),
.Y(n_970)
);

AO22x2_ASAP7_75t_L g971 ( 
.A1(n_934),
.A2(n_776),
.B1(n_766),
.B2(n_651),
.Y(n_971)
);

INVx4_ASAP7_75t_L g972 ( 
.A(n_949),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_966),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_945),
.B(n_861),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_958),
.A2(n_656),
.B1(n_774),
.B2(n_633),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_959),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_950),
.Y(n_977)
);

NAND2x1p5_ASAP7_75t_L g978 ( 
.A(n_961),
.B(n_744),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_937),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_954),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_941),
.B(n_871),
.Y(n_981)
);

AO22x2_ASAP7_75t_L g982 ( 
.A1(n_962),
.A2(n_653),
.B1(n_670),
.B2(n_657),
.Y(n_982)
);

INVxp67_ASAP7_75t_L g983 ( 
.A(n_936),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_931),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_931),
.Y(n_985)
);

INVxp67_ASAP7_75t_L g986 ( 
.A(n_957),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_955),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_933),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_960),
.B(n_864),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_935),
.Y(n_990)
);

AO22x2_ASAP7_75t_L g991 ( 
.A1(n_965),
.A2(n_716),
.B1(n_757),
.B2(n_710),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_952),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_930),
.B(n_671),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_951),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_958),
.B(n_724),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_938),
.Y(n_996)
);

AND2x6_ASAP7_75t_L g997 ( 
.A(n_940),
.B(n_631),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_947),
.B(n_784),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_953),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_958),
.B(n_724),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_939),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_944),
.B(n_724),
.Y(n_1002)
);

AO22x2_ASAP7_75t_L g1003 ( 
.A1(n_932),
.A2(n_943),
.B1(n_956),
.B2(n_927),
.Y(n_1003)
);

AO22x2_ASAP7_75t_L g1004 ( 
.A1(n_939),
.A2(n_814),
.B1(n_828),
.B2(n_813),
.Y(n_1004)
);

CKINVDCx20_ASAP7_75t_R g1005 ( 
.A(n_942),
.Y(n_1005)
);

AO22x2_ASAP7_75t_L g1006 ( 
.A1(n_946),
.A2(n_849),
.B1(n_853),
.B2(n_831),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_946),
.Y(n_1007)
);

NAND2x1p5_ASAP7_75t_L g1008 ( 
.A(n_949),
.B(n_855),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_948),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_948),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_958),
.A2(n_779),
.B1(n_841),
.B2(n_663),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_948),
.Y(n_1012)
);

BUFx12f_ASAP7_75t_SL g1013 ( 
.A(n_945),
.Y(n_1013)
);

AO22x2_ASAP7_75t_L g1014 ( 
.A1(n_934),
.A2(n_872),
.B1(n_873),
.B2(n_868),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_948),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_945),
.B(n_660),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_947),
.Y(n_1017)
);

AO22x2_ASAP7_75t_L g1018 ( 
.A1(n_934),
.A2(n_644),
.B1(n_783),
.B2(n_689),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_948),
.Y(n_1019)
);

OAI221xp5_ASAP7_75t_L g1020 ( 
.A1(n_927),
.A2(n_686),
.B1(n_698),
.B2(n_668),
.C(n_666),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_948),
.Y(n_1021)
);

OAI22xp33_ASAP7_75t_SL g1022 ( 
.A1(n_936),
.A2(n_714),
.B1(n_720),
.B2(n_701),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_948),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_949),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_948),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_948),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_948),
.Y(n_1027)
);

OAI221xp5_ASAP7_75t_L g1028 ( 
.A1(n_927),
.A2(n_752),
.B1(n_755),
.B2(n_739),
.C(n_725),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_948),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_948),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_929),
.B(n_763),
.Y(n_1031)
);

AO22x2_ASAP7_75t_L g1032 ( 
.A1(n_934),
.A2(n_646),
.B1(n_713),
.B2(n_662),
.Y(n_1032)
);

INVxp67_ASAP7_75t_L g1033 ( 
.A(n_945),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_958),
.A2(n_663),
.B1(n_841),
.B2(n_779),
.Y(n_1034)
);

AO22x2_ASAP7_75t_L g1035 ( 
.A1(n_934),
.A2(n_688),
.B1(n_733),
.B2(n_680),
.Y(n_1035)
);

AO22x2_ASAP7_75t_L g1036 ( 
.A1(n_934),
.A2(n_723),
.B1(n_738),
.B2(n_692),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_948),
.Y(n_1037)
);

NAND2x1p5_ASAP7_75t_L g1038 ( 
.A(n_949),
.B(n_678),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_949),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_945),
.B(n_771),
.Y(n_1040)
);

AO22x2_ASAP7_75t_L g1041 ( 
.A1(n_934),
.A2(n_835),
.B1(n_859),
.B2(n_741),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_948),
.Y(n_1042)
);

BUFx8_ASAP7_75t_L g1043 ( 
.A(n_954),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_929),
.B(n_782),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_948),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_958),
.A2(n_679),
.B1(n_682),
.B2(n_638),
.Y(n_1046)
);

NAND2x1p5_ASAP7_75t_L g1047 ( 
.A(n_949),
.B(n_743),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_948),
.Y(n_1048)
);

INVxp67_ASAP7_75t_L g1049 ( 
.A(n_945),
.Y(n_1049)
);

NAND2x1p5_ASAP7_75t_L g1050 ( 
.A(n_949),
.B(n_798),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_949),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_948),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_948),
.Y(n_1053)
);

AO22x2_ASAP7_75t_L g1054 ( 
.A1(n_934),
.A2(n_756),
.B1(n_746),
.B2(n_745),
.Y(n_1054)
);

INVxp67_ASAP7_75t_L g1055 ( 
.A(n_945),
.Y(n_1055)
);

NAND2xp33_ASAP7_75t_SL g1056 ( 
.A(n_1016),
.B(n_795),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_994),
.B(n_804),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_999),
.B(n_807),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_1024),
.B(n_697),
.Y(n_1059)
);

NAND2xp33_ASAP7_75t_SL g1060 ( 
.A(n_1040),
.B(n_811),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_1033),
.B(n_830),
.Y(n_1061)
);

NAND2xp33_ASAP7_75t_SL g1062 ( 
.A(n_1031),
.B(n_834),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_1049),
.B(n_838),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_974),
.B(n_748),
.Y(n_1064)
);

NAND2xp33_ASAP7_75t_SL g1065 ( 
.A(n_1044),
.B(n_851),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_1055),
.B(n_856),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_988),
.B(n_857),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_990),
.B(n_869),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_986),
.B(n_870),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_1046),
.B(n_612),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_975),
.B(n_618),
.Y(n_1071)
);

NAND2xp33_ASAP7_75t_SL g1072 ( 
.A(n_981),
.B(n_847),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_977),
.B(n_620),
.Y(n_1073)
);

NAND2xp33_ASAP7_75t_SL g1074 ( 
.A(n_976),
.B(n_854),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_1051),
.B(n_621),
.Y(n_1075)
);

NAND2xp33_ASAP7_75t_SL g1076 ( 
.A(n_1051),
.B(n_860),
.Y(n_1076)
);

NAND2xp33_ASAP7_75t_SL g1077 ( 
.A(n_1011),
.B(n_623),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_1039),
.B(n_626),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_996),
.B(n_867),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_995),
.B(n_628),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_998),
.B(n_0),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_972),
.B(n_760),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_1000),
.B(n_634),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_997),
.B(n_768),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_1022),
.B(n_636),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_989),
.B(n_639),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_993),
.B(n_640),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_1034),
.B(n_643),
.Y(n_1088)
);

NAND2xp33_ASAP7_75t_SL g1089 ( 
.A(n_992),
.B(n_842),
.Y(n_1089)
);

NAND2xp33_ASAP7_75t_SL g1090 ( 
.A(n_980),
.B(n_844),
.Y(n_1090)
);

NAND2xp33_ASAP7_75t_SL g1091 ( 
.A(n_1005),
.B(n_984),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_997),
.B(n_848),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_997),
.B(n_863),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_968),
.B(n_648),
.Y(n_1094)
);

NAND2xp33_ASAP7_75t_SL g1095 ( 
.A(n_985),
.B(n_969),
.Y(n_1095)
);

NAND2xp33_ASAP7_75t_SL g1096 ( 
.A(n_970),
.B(n_973),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1009),
.B(n_781),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_1012),
.B(n_654),
.Y(n_1098)
);

NAND2xp33_ASAP7_75t_SL g1099 ( 
.A(n_1015),
.B(n_866),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1019),
.B(n_791),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_1023),
.B(n_655),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1025),
.B(n_1026),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_1029),
.B(n_659),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_1007),
.B(n_792),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_1030),
.B(n_661),
.Y(n_1105)
);

NAND2xp33_ASAP7_75t_SL g1106 ( 
.A(n_1042),
.B(n_833),
.Y(n_1106)
);

NAND2xp33_ASAP7_75t_SL g1107 ( 
.A(n_1052),
.B(n_837),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_1053),
.B(n_664),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_978),
.B(n_1010),
.Y(n_1109)
);

NAND2xp33_ASAP7_75t_SL g1110 ( 
.A(n_1013),
.B(n_840),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_1021),
.B(n_665),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1027),
.B(n_803),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_1037),
.B(n_669),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1045),
.B(n_812),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_1048),
.B(n_672),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_1008),
.B(n_673),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1003),
.B(n_820),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_1001),
.B(n_676),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_979),
.B(n_681),
.Y(n_1119)
);

NAND2xp33_ASAP7_75t_SL g1120 ( 
.A(n_987),
.B(n_845),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_1017),
.B(n_683),
.Y(n_1121)
);

NAND2xp33_ASAP7_75t_SL g1122 ( 
.A(n_1002),
.B(n_824),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_1038),
.B(n_1047),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_1050),
.B(n_685),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_1043),
.B(n_687),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_1018),
.B(n_691),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_1032),
.B(n_693),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_1035),
.B(n_694),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1036),
.B(n_825),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_1041),
.B(n_696),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_1054),
.B(n_699),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_1006),
.B(n_700),
.Y(n_1132)
);

NAND2xp33_ASAP7_75t_SL g1133 ( 
.A(n_1020),
.B(n_874),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_1004),
.B(n_704),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_982),
.B(n_705),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_1028),
.B(n_708),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_991),
.B(n_711),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_1014),
.B(n_715),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_971),
.B(n_718),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_994),
.B(n_808),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_967),
.B(n_721),
.Y(n_1141)
);

NAND2xp33_ASAP7_75t_SL g1142 ( 
.A(n_967),
.B(n_829),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_967),
.B(n_722),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_967),
.B(n_726),
.Y(n_1144)
);

NAND2xp33_ASAP7_75t_SL g1145 ( 
.A(n_967),
.B(n_858),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_967),
.B(n_727),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_967),
.B(n_728),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_967),
.B(n_731),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_967),
.B(n_734),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_967),
.B(n_737),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_967),
.B(n_740),
.Y(n_1151)
);

AND2x6_ASAP7_75t_L g1152 ( 
.A(n_974),
.B(n_675),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_967),
.B(n_747),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_983),
.B(n_1),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_967),
.B(n_749),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_967),
.B(n_750),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_967),
.B(n_753),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_967),
.B(n_754),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_967),
.B(n_761),
.Y(n_1159)
);

NAND2xp33_ASAP7_75t_SL g1160 ( 
.A(n_967),
.B(n_762),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_967),
.B(n_764),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_967),
.B(n_767),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_967),
.B(n_769),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_967),
.B(n_770),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_983),
.B(n_2),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_967),
.B(n_772),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_967),
.B(n_775),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_967),
.B(n_777),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_967),
.B(n_786),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_967),
.B(n_787),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_967),
.B(n_788),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_967),
.B(n_789),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_967),
.B(n_790),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_967),
.B(n_794),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_967),
.B(n_796),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_967),
.B(n_797),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_967),
.B(n_802),
.Y(n_1177)
);

NAND2xp33_ASAP7_75t_SL g1178 ( 
.A(n_967),
.B(n_805),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_967),
.B(n_810),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_983),
.B(n_2),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_967),
.B(n_816),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_967),
.B(n_817),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_967),
.B(n_818),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_967),
.B(n_819),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_967),
.B(n_821),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_983),
.B(n_3),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_967),
.B(n_823),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1102),
.A2(n_862),
.B(n_622),
.Y(n_1188)
);

NAND2x1_ASAP7_75t_L g1189 ( 
.A(n_1152),
.B(n_675),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1112),
.A2(n_627),
.B(n_615),
.Y(n_1190)
);

AO32x2_ASAP7_75t_L g1191 ( 
.A1(n_1117),
.A2(n_5),
.A3(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1081),
.B(n_4),
.Y(n_1192)
);

NAND3xp33_ASAP7_75t_SL g1193 ( 
.A(n_1136),
.B(n_839),
.C(n_827),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1114),
.Y(n_1194)
);

NAND2x1p5_ASAP7_75t_L g1195 ( 
.A(n_1123),
.B(n_675),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1097),
.A2(n_717),
.B(n_658),
.Y(n_1196)
);

OAI22x1_ASAP7_75t_L g1197 ( 
.A1(n_1126),
.A2(n_742),
.B1(n_759),
.B2(n_729),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1143),
.B(n_6),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1100),
.A2(n_822),
.B(n_806),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_1091),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_1090),
.B(n_865),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1079),
.Y(n_1202)
);

NAND2x1_ASAP7_75t_L g1203 ( 
.A(n_1152),
.B(n_290),
.Y(n_1203)
);

AO21x2_ASAP7_75t_L g1204 ( 
.A1(n_1087),
.A2(n_1083),
.B(n_1080),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1084),
.Y(n_1205)
);

AOI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1141),
.A2(n_1146),
.B(n_1144),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1109),
.A2(n_751),
.B(n_293),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1119),
.A2(n_751),
.B(n_295),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1096),
.A2(n_297),
.B(n_291),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_1059),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1059),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1151),
.A2(n_1172),
.B(n_1168),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1092),
.A2(n_751),
.B(n_300),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1181),
.B(n_7),
.Y(n_1214)
);

CKINVDCx6p67_ASAP7_75t_R g1215 ( 
.A(n_1125),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1104),
.Y(n_1216)
);

CKINVDCx12_ASAP7_75t_R g1217 ( 
.A(n_1154),
.Y(n_1217)
);

OR2x2_ASAP7_75t_L g1218 ( 
.A(n_1064),
.B(n_7),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1093),
.Y(n_1219)
);

INVx4_ASAP7_75t_SL g1220 ( 
.A(n_1152),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1062),
.A2(n_11),
.B(n_9),
.C(n_10),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1064),
.B(n_9),
.Y(n_1222)
);

AOI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1147),
.A2(n_1149),
.B(n_1148),
.Y(n_1223)
);

BUFx10_ASAP7_75t_L g1224 ( 
.A(n_1082),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1150),
.A2(n_301),
.B(n_299),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1104),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1058),
.Y(n_1227)
);

INVxp67_ASAP7_75t_SL g1228 ( 
.A(n_1165),
.Y(n_1228)
);

AO31x2_ASAP7_75t_L g1229 ( 
.A1(n_1129),
.A2(n_1067),
.A3(n_1122),
.B(n_1095),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_SL g1230 ( 
.A(n_1152),
.B(n_10),
.Y(n_1230)
);

CKINVDCx8_ASAP7_75t_R g1231 ( 
.A(n_1152),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1180),
.B(n_11),
.Y(n_1232)
);

AOI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1153),
.A2(n_303),
.B(n_302),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1086),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_1234)
);

OA21x2_ASAP7_75t_L g1235 ( 
.A1(n_1155),
.A2(n_305),
.B(n_304),
.Y(n_1235)
);

AO31x2_ASAP7_75t_L g1236 ( 
.A1(n_1134),
.A2(n_307),
.A3(n_310),
.B(n_306),
.Y(n_1236)
);

OAI21xp33_ASAP7_75t_SL g1237 ( 
.A1(n_1156),
.A2(n_20),
.B(n_12),
.Y(n_1237)
);

NOR2x1_ASAP7_75t_SL g1238 ( 
.A(n_1124),
.B(n_311),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1186),
.B(n_13),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1068),
.B(n_14),
.Y(n_1240)
);

AOI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1157),
.A2(n_315),
.B(n_314),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1082),
.B(n_15),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1065),
.A2(n_17),
.B(n_15),
.C(n_16),
.Y(n_1243)
);

NAND2xp33_ASAP7_75t_R g1244 ( 
.A(n_1140),
.B(n_316),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1158),
.A2(n_318),
.B(n_317),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1140),
.B(n_16),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1088),
.B(n_17),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1111),
.A2(n_1115),
.B(n_1113),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1094),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1159),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1071),
.B(n_19),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1161),
.A2(n_1187),
.B(n_1170),
.Y(n_1252)
);

A2O1A1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1133),
.A2(n_23),
.B(n_21),
.C(n_22),
.Y(n_1253)
);

BUFx12f_ASAP7_75t_L g1254 ( 
.A(n_1110),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1098),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1101),
.A2(n_320),
.B(n_319),
.Y(n_1256)
);

CKINVDCx20_ASAP7_75t_R g1257 ( 
.A(n_1074),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_1116),
.B(n_21),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1103),
.A2(n_323),
.B(n_322),
.Y(n_1259)
);

INVx1_ASAP7_75t_SL g1260 ( 
.A(n_1076),
.Y(n_1260)
);

INVxp67_ASAP7_75t_L g1261 ( 
.A(n_1069),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1162),
.A2(n_325),
.B(n_324),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1105),
.A2(n_327),
.B(n_326),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1163),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1164),
.A2(n_329),
.B(n_328),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1108),
.A2(n_331),
.B(n_330),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1056),
.Y(n_1267)
);

AO31x2_ASAP7_75t_L g1268 ( 
.A1(n_1085),
.A2(n_1132),
.A3(n_1127),
.B(n_1130),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1121),
.B(n_24),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1073),
.B(n_25),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1057),
.Y(n_1271)
);

O2A1O1Ixp5_ASAP7_75t_SL g1272 ( 
.A1(n_1128),
.A2(n_1131),
.B(n_1137),
.C(n_1135),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1078),
.A2(n_336),
.B(n_334),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_1075),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1166),
.A2(n_340),
.B(n_338),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_SL g1276 ( 
.A(n_1060),
.B(n_25),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1167),
.B(n_26),
.Y(n_1277)
);

INVx4_ASAP7_75t_L g1278 ( 
.A(n_1099),
.Y(n_1278)
);

NAND2xp33_ASAP7_75t_L g1279 ( 
.A(n_1142),
.B(n_1145),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1169),
.B(n_26),
.Y(n_1280)
);

AOI21xp33_ASAP7_75t_L g1281 ( 
.A1(n_1070),
.A2(n_27),
.B(n_28),
.Y(n_1281)
);

BUFx10_ASAP7_75t_L g1282 ( 
.A(n_1118),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1138),
.B(n_29),
.Y(n_1283)
);

AO31x2_ASAP7_75t_L g1284 ( 
.A1(n_1089),
.A2(n_342),
.A3(n_343),
.B(n_341),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1061),
.Y(n_1285)
);

AO21x2_ASAP7_75t_L g1286 ( 
.A1(n_1171),
.A2(n_346),
.B(n_345),
.Y(n_1286)
);

OR2x6_ASAP7_75t_L g1287 ( 
.A(n_1139),
.B(n_30),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1063),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1173),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1174),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_1290)
);

INVx1_ASAP7_75t_SL g1291 ( 
.A(n_1211),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1216),
.Y(n_1292)
);

AOI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1276),
.A2(n_1077),
.B1(n_1107),
.B2(n_1106),
.Y(n_1293)
);

INVx6_ASAP7_75t_SL g1294 ( 
.A(n_1224),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1216),
.A2(n_1066),
.B1(n_1120),
.B2(n_1072),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1228),
.A2(n_1176),
.B1(n_1177),
.B2(n_1175),
.Y(n_1296)
);

NOR2xp67_ASAP7_75t_L g1297 ( 
.A(n_1278),
.B(n_1179),
.Y(n_1297)
);

BUFx3_ASAP7_75t_L g1298 ( 
.A(n_1254),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1205),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1219),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1190),
.A2(n_1183),
.B(n_1182),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1210),
.B(n_1184),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_1226),
.Y(n_1303)
);

NAND3xp33_ASAP7_75t_L g1304 ( 
.A(n_1253),
.B(n_1243),
.C(n_1221),
.Y(n_1304)
);

INVx2_ASAP7_75t_SL g1305 ( 
.A(n_1226),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1217),
.Y(n_1306)
);

AOI21xp33_ASAP7_75t_L g1307 ( 
.A1(n_1198),
.A2(n_1185),
.B(n_1160),
.Y(n_1307)
);

NOR2xp67_ASAP7_75t_L g1308 ( 
.A(n_1227),
.B(n_348),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1194),
.Y(n_1309)
);

OAI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1218),
.A2(n_1178),
.B1(n_42),
.B2(n_50),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1202),
.Y(n_1311)
);

OAI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1214),
.A2(n_36),
.B(n_37),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1242),
.B(n_37),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1196),
.A2(n_350),
.B(n_349),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1251),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1249),
.Y(n_1316)
);

NAND2x1p5_ASAP7_75t_L g1317 ( 
.A(n_1260),
.B(n_351),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1193),
.A2(n_38),
.B(n_39),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1255),
.Y(n_1319)
);

O2A1O1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1240),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_1320)
);

NOR2x1_ASAP7_75t_SL g1321 ( 
.A(n_1204),
.B(n_40),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1229),
.Y(n_1322)
);

AOI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1199),
.A2(n_353),
.B(n_352),
.Y(n_1323)
);

AOI332xp33_ASAP7_75t_L g1324 ( 
.A1(n_1239),
.A2(n_46),
.A3(n_45),
.B1(n_43),
.B2(n_47),
.B3(n_48),
.C1(n_42),
.C2(n_44),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1200),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1285),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1288),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1209),
.A2(n_355),
.B(n_354),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1287),
.A2(n_48),
.B1(n_41),
.B2(n_43),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1247),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1267),
.B(n_41),
.Y(n_1331)
);

OA21x2_ASAP7_75t_L g1332 ( 
.A1(n_1213),
.A2(n_357),
.B(n_356),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1229),
.Y(n_1333)
);

INVx2_ASAP7_75t_SL g1334 ( 
.A(n_1282),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1271),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1222),
.B(n_49),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1192),
.B(n_50),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1191),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1207),
.A2(n_362),
.B(n_360),
.Y(n_1339)
);

AO21x2_ASAP7_75t_L g1340 ( 
.A1(n_1188),
.A2(n_365),
.B(n_363),
.Y(n_1340)
);

OR2x6_ASAP7_75t_L g1341 ( 
.A(n_1274),
.B(n_51),
.Y(n_1341)
);

OAI211xp5_ASAP7_75t_L g1342 ( 
.A1(n_1237),
.A2(n_54),
.B(n_52),
.C(n_53),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1270),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1246),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_1230),
.B(n_54),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1261),
.B(n_55),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1274),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1208),
.A2(n_367),
.B(n_366),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1277),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_1215),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1280),
.Y(n_1351)
);

A2O1A1Ixp33_ASAP7_75t_L g1352 ( 
.A1(n_1252),
.A2(n_57),
.B(n_58),
.C(n_56),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1257),
.B(n_55),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1232),
.B(n_57),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1269),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1283),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1248),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1258),
.B(n_59),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1220),
.B(n_369),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1256),
.A2(n_373),
.B(n_370),
.Y(n_1360)
);

OR2x6_ASAP7_75t_L g1361 ( 
.A(n_1195),
.B(n_60),
.Y(n_1361)
);

INVx2_ASAP7_75t_SL g1362 ( 
.A(n_1268),
.Y(n_1362)
);

INVx3_ASAP7_75t_L g1363 ( 
.A(n_1231),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1268),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1250),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1264),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1272),
.A2(n_61),
.B(n_62),
.Y(n_1367)
);

INVx3_ASAP7_75t_L g1368 ( 
.A(n_1206),
.Y(n_1368)
);

AOI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1223),
.A2(n_1241),
.B(n_1233),
.Y(n_1369)
);

OA21x2_ASAP7_75t_L g1370 ( 
.A1(n_1259),
.A2(n_377),
.B(n_375),
.Y(n_1370)
);

OAI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1234),
.A2(n_63),
.B(n_64),
.Y(n_1371)
);

BUFx8_ASAP7_75t_L g1372 ( 
.A(n_1244),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1289),
.Y(n_1373)
);

INVxp67_ASAP7_75t_L g1374 ( 
.A(n_1197),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1235),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_SL g1376 ( 
.A1(n_1238),
.A2(n_65),
.B(n_64),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1290),
.Y(n_1377)
);

AO31x2_ASAP7_75t_L g1378 ( 
.A1(n_1225),
.A2(n_379),
.A3(n_381),
.B(n_378),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1263),
.A2(n_383),
.B(n_382),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1281),
.B(n_63),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1266),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1201),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1273),
.A2(n_385),
.B(n_384),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1279),
.B(n_66),
.Y(n_1384)
);

OR2x6_ASAP7_75t_L g1385 ( 
.A(n_1203),
.B(n_67),
.Y(n_1385)
);

INVx3_ASAP7_75t_L g1386 ( 
.A(n_1236),
.Y(n_1386)
);

OA21x2_ASAP7_75t_L g1387 ( 
.A1(n_1245),
.A2(n_388),
.B(n_386),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_SL g1388 ( 
.A1(n_1189),
.A2(n_1220),
.B1(n_1284),
.B2(n_71),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1262),
.B(n_68),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1286),
.A2(n_72),
.B1(n_69),
.B2(n_71),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1265),
.A2(n_390),
.B(n_389),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_1275),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1284),
.Y(n_1393)
);

OAI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1212),
.A2(n_69),
.B(n_73),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1190),
.A2(n_393),
.B(n_392),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1205),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1202),
.B(n_74),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1190),
.A2(n_396),
.B(n_394),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1190),
.A2(n_400),
.B(n_398),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1369),
.A2(n_402),
.B(n_401),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_1292),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1325),
.B(n_74),
.Y(n_1402)
);

NAND2x1p5_ASAP7_75t_L g1403 ( 
.A(n_1363),
.B(n_406),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1300),
.Y(n_1404)
);

AND2x4_ASAP7_75t_L g1405 ( 
.A(n_1298),
.B(n_75),
.Y(n_1405)
);

OA21x2_ASAP7_75t_L g1406 ( 
.A1(n_1393),
.A2(n_408),
.B(n_407),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1309),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1311),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1299),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1347),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1396),
.Y(n_1411)
);

AOI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1323),
.A2(n_412),
.B(n_410),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1357),
.Y(n_1413)
);

INVx3_ASAP7_75t_L g1414 ( 
.A(n_1292),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1291),
.B(n_75),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1316),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1327),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1314),
.A2(n_414),
.B(n_413),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1313),
.B(n_76),
.Y(n_1419)
);

OA21x2_ASAP7_75t_L g1420 ( 
.A1(n_1322),
.A2(n_420),
.B(n_419),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1395),
.A2(n_424),
.B(n_421),
.Y(n_1421)
);

BUFx3_ASAP7_75t_L g1422 ( 
.A(n_1347),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1326),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1319),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1335),
.Y(n_1425)
);

AOI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1333),
.A2(n_426),
.B(n_425),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1330),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1344),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1315),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1349),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1343),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1351),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1364),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1397),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1368),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1356),
.B(n_76),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1362),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1302),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1372),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_1439)
);

AND2x4_ASAP7_75t_SL g1440 ( 
.A(n_1303),
.B(n_427),
.Y(n_1440)
);

BUFx2_ASAP7_75t_L g1441 ( 
.A(n_1386),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1303),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1328),
.A2(n_1392),
.B(n_1394),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1305),
.B(n_77),
.Y(n_1444)
);

OA21x2_ASAP7_75t_L g1445 ( 
.A1(n_1375),
.A2(n_430),
.B(n_428),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1321),
.Y(n_1446)
);

INVx2_ASAP7_75t_SL g1447 ( 
.A(n_1350),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1381),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_1294),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1384),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1371),
.A2(n_1304),
.B1(n_1318),
.B2(n_1374),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1338),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1331),
.B(n_78),
.Y(n_1453)
);

AOI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1398),
.A2(n_1399),
.B(n_1366),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1334),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1365),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1336),
.B(n_1354),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1373),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1306),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1377),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1367),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1312),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1378),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1297),
.B(n_79),
.Y(n_1464)
);

INVx3_ASAP7_75t_L g1465 ( 
.A(n_1359),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1348),
.A2(n_433),
.B(n_431),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1308),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1455),
.Y(n_1468)
);

NAND2xp33_ASAP7_75t_R g1469 ( 
.A(n_1464),
.B(n_1341),
.Y(n_1469)
);

XNOR2xp5_ASAP7_75t_L g1470 ( 
.A(n_1419),
.B(n_1341),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_R g1471 ( 
.A(n_1465),
.B(n_1353),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_R g1472 ( 
.A(n_1449),
.B(n_1346),
.Y(n_1472)
);

AND2x4_ASAP7_75t_L g1473 ( 
.A(n_1438),
.B(n_1385),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1428),
.B(n_1358),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1410),
.B(n_1385),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1422),
.B(n_1361),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1417),
.B(n_1361),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1453),
.B(n_1337),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1404),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1459),
.B(n_1345),
.Y(n_1480)
);

NAND2xp33_ASAP7_75t_R g1481 ( 
.A(n_1444),
.B(n_1436),
.Y(n_1481)
);

NAND2xp33_ASAP7_75t_R g1482 ( 
.A(n_1444),
.B(n_1380),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1442),
.B(n_1293),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_R g1484 ( 
.A(n_1447),
.B(n_1295),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1429),
.B(n_1329),
.Y(n_1485)
);

INVxp67_ASAP7_75t_L g1486 ( 
.A(n_1401),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_1401),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1416),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_R g1489 ( 
.A(n_1414),
.B(n_1389),
.Y(n_1489)
);

NAND2xp33_ASAP7_75t_R g1490 ( 
.A(n_1402),
.B(n_1332),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1405),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1427),
.B(n_1352),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1431),
.B(n_1301),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1424),
.B(n_1355),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1425),
.B(n_1340),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_R g1496 ( 
.A(n_1457),
.B(n_1390),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_R g1497 ( 
.A(n_1434),
.B(n_80),
.Y(n_1497)
);

INVxp67_ASAP7_75t_L g1498 ( 
.A(n_1430),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1432),
.B(n_1320),
.Y(n_1499)
);

INVxp67_ASAP7_75t_L g1500 ( 
.A(n_1450),
.Y(n_1500)
);

NAND2xp33_ASAP7_75t_R g1501 ( 
.A(n_1415),
.B(n_1370),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1408),
.Y(n_1502)
);

NAND2xp33_ASAP7_75t_R g1503 ( 
.A(n_1420),
.B(n_1387),
.Y(n_1503)
);

NAND2xp33_ASAP7_75t_R g1504 ( 
.A(n_1420),
.B(n_1324),
.Y(n_1504)
);

NAND2xp33_ASAP7_75t_R g1505 ( 
.A(n_1406),
.B(n_81),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_1440),
.Y(n_1506)
);

INVxp67_ASAP7_75t_L g1507 ( 
.A(n_1409),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1456),
.B(n_1317),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1498),
.Y(n_1509)
);

INVxp67_ASAP7_75t_SL g1510 ( 
.A(n_1500),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1507),
.B(n_1433),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1479),
.B(n_1452),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1488),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1474),
.B(n_1452),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1502),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_1468),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1493),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1471),
.Y(n_1518)
);

BUFx2_ASAP7_75t_L g1519 ( 
.A(n_1489),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1477),
.B(n_1435),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1478),
.A2(n_1451),
.B1(n_1439),
.B2(n_1462),
.Y(n_1521)
);

INVxp67_ASAP7_75t_SL g1522 ( 
.A(n_1503),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1499),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1492),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1508),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1495),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1486),
.B(n_1458),
.Y(n_1527)
);

BUFx3_ASAP7_75t_L g1528 ( 
.A(n_1487),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1485),
.B(n_1460),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1480),
.B(n_1423),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1496),
.A2(n_1467),
.B1(n_1461),
.B2(n_1307),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1470),
.A2(n_1310),
.B1(n_1342),
.B2(n_1382),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1473),
.B(n_1413),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1483),
.B(n_1413),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1494),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_1475),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1497),
.B(n_1448),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1491),
.B(n_1448),
.Y(n_1538)
);

NOR2x1_ASAP7_75t_SL g1539 ( 
.A(n_1501),
.B(n_1446),
.Y(n_1539)
);

INVx2_ASAP7_75t_SL g1540 ( 
.A(n_1476),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1506),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1484),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1470),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1472),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1482),
.Y(n_1545)
);

AND2x4_ASAP7_75t_SL g1546 ( 
.A(n_1469),
.B(n_1407),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1505),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1481),
.B(n_1441),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1490),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1504),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1498),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1479),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1514),
.B(n_1441),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1515),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1509),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1548),
.B(n_1437),
.Y(n_1556)
);

OAI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1550),
.A2(n_1443),
.B1(n_1403),
.B2(n_1296),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1551),
.B(n_1437),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1552),
.Y(n_1559)
);

NOR2xp67_ASAP7_75t_SL g1560 ( 
.A(n_1519),
.B(n_1406),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1512),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1513),
.Y(n_1562)
);

AOI222xp33_ASAP7_75t_L g1563 ( 
.A1(n_1521),
.A2(n_1388),
.B1(n_1376),
.B2(n_1463),
.C1(n_1411),
.C2(n_1391),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1510),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1538),
.B(n_1454),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1533),
.B(n_1454),
.Y(n_1566)
);

BUFx3_ASAP7_75t_L g1567 ( 
.A(n_1516),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1523),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1511),
.B(n_80),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1511),
.B(n_81),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1536),
.B(n_1400),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1525),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1535),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1528),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1520),
.B(n_1466),
.Y(n_1575)
);

OAI33xp33_ASAP7_75t_L g1576 ( 
.A1(n_1532),
.A2(n_85),
.A3(n_87),
.B1(n_83),
.B2(n_84),
.B3(n_86),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1547),
.A2(n_1549),
.B1(n_1545),
.B2(n_1522),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1533),
.B(n_1426),
.Y(n_1578)
);

OR2x6_ASAP7_75t_L g1579 ( 
.A(n_1537),
.B(n_1426),
.Y(n_1579)
);

INVxp67_ASAP7_75t_SL g1580 ( 
.A(n_1539),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1534),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1529),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1544),
.B(n_1418),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1541),
.B(n_1540),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1527),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1539),
.B(n_1421),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1542),
.B(n_1412),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1524),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1518),
.B(n_1412),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1530),
.Y(n_1590)
);

OAI221xp5_ASAP7_75t_L g1591 ( 
.A1(n_1531),
.A2(n_1445),
.B1(n_86),
.B2(n_84),
.C(n_85),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1526),
.Y(n_1592)
);

NOR2xp67_ASAP7_75t_L g1593 ( 
.A(n_1517),
.B(n_87),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1546),
.Y(n_1594)
);

OAI31xp33_ASAP7_75t_SL g1595 ( 
.A1(n_1543),
.A2(n_1383),
.A3(n_1379),
.B(n_1360),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1514),
.B(n_88),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1514),
.B(n_88),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1515),
.Y(n_1598)
);

INVx1_ASAP7_75t_SL g1599 ( 
.A(n_1519),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1515),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1514),
.B(n_1445),
.Y(n_1601)
);

INVx1_ASAP7_75t_SL g1602 ( 
.A(n_1519),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1509),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1514),
.B(n_1339),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1514),
.B(n_89),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_SL g1606 ( 
.A1(n_1550),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_1606)
);

INVx2_ASAP7_75t_SL g1607 ( 
.A(n_1528),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1523),
.B(n_90),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1515),
.Y(n_1609)
);

OAI31xp33_ASAP7_75t_L g1610 ( 
.A1(n_1550),
.A2(n_93),
.A3(n_91),
.B(n_92),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1514),
.B(n_92),
.Y(n_1611)
);

INVx1_ASAP7_75t_SL g1612 ( 
.A(n_1599),
.Y(n_1612)
);

AND2x4_ASAP7_75t_L g1613 ( 
.A(n_1556),
.B(n_94),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1554),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1603),
.B(n_95),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1558),
.B(n_96),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1602),
.B(n_1574),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1568),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1561),
.B(n_96),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1564),
.B(n_97),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1590),
.B(n_1588),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1556),
.B(n_1581),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1584),
.B(n_97),
.Y(n_1623)
);

INVx1_ASAP7_75t_SL g1624 ( 
.A(n_1567),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1582),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1565),
.B(n_1607),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1582),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1587),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1559),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1566),
.B(n_98),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1572),
.B(n_98),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1562),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1566),
.B(n_99),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1601),
.B(n_99),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1585),
.B(n_100),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1594),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1598),
.B(n_1600),
.Y(n_1637)
);

BUFx2_ASAP7_75t_L g1638 ( 
.A(n_1580),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1571),
.B(n_100),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1609),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1604),
.B(n_101),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1589),
.B(n_102),
.Y(n_1642)
);

INVxp67_ASAP7_75t_L g1643 ( 
.A(n_1608),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1575),
.B(n_103),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1573),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1583),
.B(n_104),
.Y(n_1646)
);

NAND2x1p5_ASAP7_75t_L g1647 ( 
.A(n_1593),
.B(n_104),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1596),
.B(n_105),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1597),
.B(n_106),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1605),
.B(n_1611),
.Y(n_1650)
);

NOR2x1_ASAP7_75t_L g1651 ( 
.A(n_1569),
.B(n_106),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1577),
.B(n_107),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1579),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1586),
.B(n_109),
.Y(n_1654)
);

INVx3_ASAP7_75t_L g1655 ( 
.A(n_1578),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1592),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1570),
.B(n_109),
.Y(n_1657)
);

OR2x6_ASAP7_75t_L g1658 ( 
.A(n_1557),
.B(n_110),
.Y(n_1658)
);

INVxp67_ASAP7_75t_L g1659 ( 
.A(n_1576),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1560),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1591),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1560),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1563),
.B(n_111),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1610),
.B(n_111),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1595),
.B(n_112),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1606),
.B(n_113),
.Y(n_1666)
);

INVxp67_ASAP7_75t_SL g1667 ( 
.A(n_1555),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1553),
.B(n_113),
.Y(n_1668)
);

AND2x4_ASAP7_75t_L g1669 ( 
.A(n_1556),
.B(n_114),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1555),
.B(n_114),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1561),
.B(n_115),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1599),
.B(n_115),
.Y(n_1672)
);

AND2x4_ASAP7_75t_SL g1673 ( 
.A(n_1607),
.B(n_116),
.Y(n_1673)
);

NAND4xp25_ASAP7_75t_L g1674 ( 
.A(n_1610),
.B(n_118),
.C(n_116),
.D(n_117),
.Y(n_1674)
);

INVx3_ASAP7_75t_L g1675 ( 
.A(n_1574),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1555),
.B(n_117),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1554),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1554),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1554),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1553),
.B(n_119),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1553),
.B(n_120),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1561),
.B(n_120),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1588),
.Y(n_1683)
);

AO221x2_ASAP7_75t_L g1684 ( 
.A1(n_1665),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.C(n_124),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1621),
.B(n_121),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1643),
.B(n_124),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1667),
.B(n_125),
.Y(n_1687)
);

AOI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1661),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_1688)
);

AO221x2_ASAP7_75t_L g1689 ( 
.A1(n_1670),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.C(n_134),
.Y(n_1689)
);

NAND2xp33_ASAP7_75t_SL g1690 ( 
.A(n_1638),
.B(n_131),
.Y(n_1690)
);

AO221x2_ASAP7_75t_L g1691 ( 
.A1(n_1676),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.C(n_135),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1642),
.B(n_137),
.Y(n_1692)
);

AOI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1658),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1634),
.B(n_138),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1654),
.B(n_139),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1625),
.B(n_140),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1627),
.B(n_141),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1653),
.B(n_143),
.Y(n_1698)
);

INVxp67_ASAP7_75t_L g1699 ( 
.A(n_1651),
.Y(n_1699)
);

NAND2xp33_ASAP7_75t_SL g1700 ( 
.A(n_1638),
.B(n_144),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1618),
.B(n_144),
.Y(n_1701)
);

OAI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1658),
.A2(n_148),
.B1(n_149),
.B2(n_147),
.Y(n_1702)
);

INVxp67_ASAP7_75t_L g1703 ( 
.A(n_1617),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_1624),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1637),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1612),
.B(n_146),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_1673),
.Y(n_1707)
);

AO221x2_ASAP7_75t_L g1708 ( 
.A1(n_1666),
.A2(n_1662),
.B1(n_1660),
.B2(n_1649),
.C(n_1648),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1641),
.B(n_1644),
.Y(n_1709)
);

NOR2x1_ASAP7_75t_L g1710 ( 
.A(n_1639),
.B(n_1613),
.Y(n_1710)
);

OAI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1674),
.A2(n_152),
.B1(n_153),
.B2(n_151),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1614),
.Y(n_1712)
);

NAND2xp33_ASAP7_75t_SL g1713 ( 
.A(n_1615),
.B(n_150),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_R g1714 ( 
.A(n_1672),
.B(n_151),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1646),
.B(n_152),
.Y(n_1715)
);

OAI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1663),
.A2(n_155),
.B1(n_156),
.B2(n_154),
.Y(n_1716)
);

OAI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1652),
.A2(n_156),
.B1(n_157),
.B2(n_155),
.Y(n_1717)
);

INVxp67_ASAP7_75t_L g1718 ( 
.A(n_1630),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1677),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1678),
.Y(n_1720)
);

AOI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1664),
.A2(n_162),
.B1(n_158),
.B2(n_161),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1679),
.B(n_163),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1632),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1629),
.B(n_163),
.Y(n_1724)
);

NOR2xp67_ASAP7_75t_L g1725 ( 
.A(n_1655),
.B(n_164),
.Y(n_1725)
);

NAND2xp33_ASAP7_75t_SL g1726 ( 
.A(n_1668),
.B(n_164),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1640),
.B(n_165),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1620),
.B(n_165),
.Y(n_1728)
);

AOI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1647),
.A2(n_168),
.B1(n_166),
.B2(n_167),
.Y(n_1729)
);

NOR2x1_ASAP7_75t_R g1730 ( 
.A(n_1669),
.B(n_166),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1633),
.B(n_167),
.Y(n_1731)
);

OAI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1635),
.A2(n_171),
.B1(n_173),
.B2(n_170),
.Y(n_1732)
);

INVx2_ASAP7_75t_SL g1733 ( 
.A(n_1636),
.Y(n_1733)
);

OAI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1631),
.A2(n_174),
.B1(n_175),
.B2(n_173),
.Y(n_1734)
);

NOR2x1_ASAP7_75t_L g1735 ( 
.A(n_1657),
.B(n_168),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_1623),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1626),
.B(n_174),
.Y(n_1737)
);

OAI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1671),
.A2(n_177),
.B1(n_178),
.B2(n_176),
.Y(n_1738)
);

OAI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1682),
.A2(n_177),
.B1(n_179),
.B2(n_176),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1650),
.B(n_175),
.Y(n_1740)
);

AOI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1683),
.A2(n_1619),
.B1(n_1645),
.B2(n_1616),
.Y(n_1741)
);

NAND2xp33_ASAP7_75t_SL g1742 ( 
.A(n_1680),
.B(n_180),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1681),
.B(n_180),
.Y(n_1743)
);

NOR2xp33_ASAP7_75t_L g1744 ( 
.A(n_1622),
.B(n_182),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1628),
.B(n_183),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1656),
.B(n_184),
.Y(n_1746)
);

NAND2xp33_ASAP7_75t_SL g1747 ( 
.A(n_1638),
.B(n_185),
.Y(n_1747)
);

NOR2x1_ASAP7_75t_L g1748 ( 
.A(n_1675),
.B(n_186),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1643),
.B(n_188),
.Y(n_1749)
);

AO221x2_ASAP7_75t_L g1750 ( 
.A1(n_1665),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.C(n_191),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1643),
.B(n_189),
.Y(n_1751)
);

NAND2xp33_ASAP7_75t_R g1752 ( 
.A(n_1639),
.B(n_191),
.Y(n_1752)
);

INVx3_ASAP7_75t_L g1753 ( 
.A(n_1675),
.Y(n_1753)
);

BUFx2_ASAP7_75t_L g1754 ( 
.A(n_1667),
.Y(n_1754)
);

NAND2xp33_ASAP7_75t_SL g1755 ( 
.A(n_1638),
.B(n_192),
.Y(n_1755)
);

CKINVDCx14_ASAP7_75t_R g1756 ( 
.A(n_1650),
.Y(n_1756)
);

OAI221xp5_ASAP7_75t_L g1757 ( 
.A1(n_1659),
.A2(n_194),
.B1(n_192),
.B2(n_193),
.C(n_195),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1614),
.Y(n_1758)
);

NAND2xp33_ASAP7_75t_SL g1759 ( 
.A(n_1638),
.B(n_193),
.Y(n_1759)
);

OAI221xp5_ASAP7_75t_L g1760 ( 
.A1(n_1659),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.C(n_199),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1667),
.B(n_200),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1643),
.B(n_202),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1667),
.B(n_203),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1667),
.B(n_204),
.Y(n_1764)
);

INVx2_ASAP7_75t_SL g1765 ( 
.A(n_1675),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1626),
.B(n_206),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_R g1767 ( 
.A(n_1704),
.B(n_206),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1756),
.B(n_207),
.Y(n_1768)
);

INVx1_ASAP7_75t_SL g1769 ( 
.A(n_1707),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1723),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1708),
.B(n_208),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1712),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1708),
.B(n_209),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1753),
.B(n_209),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1754),
.B(n_210),
.Y(n_1775)
);

INVx1_ASAP7_75t_SL g1776 ( 
.A(n_1736),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1705),
.B(n_211),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1719),
.Y(n_1778)
);

AOI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1684),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1699),
.B(n_213),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1720),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_SL g1782 ( 
.A(n_1730),
.B(n_214),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1685),
.B(n_215),
.Y(n_1783)
);

INVx1_ASAP7_75t_SL g1784 ( 
.A(n_1714),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1758),
.B(n_216),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1733),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1746),
.Y(n_1787)
);

AOI22x1_ASAP7_75t_L g1788 ( 
.A1(n_1765),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1718),
.B(n_218),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1703),
.A2(n_222),
.B1(n_219),
.B2(n_220),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1737),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1766),
.Y(n_1792)
);

AND2x4_ASAP7_75t_L g1793 ( 
.A(n_1741),
.B(n_1709),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1740),
.B(n_220),
.Y(n_1794)
);

AND2x4_ASAP7_75t_SL g1795 ( 
.A(n_1743),
.B(n_222),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1745),
.B(n_223),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1722),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1696),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1697),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1701),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1735),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1687),
.B(n_223),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1724),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1727),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1698),
.B(n_224),
.Y(n_1805)
);

INVx5_ASAP7_75t_L g1806 ( 
.A(n_1689),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1748),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1761),
.B(n_224),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1763),
.B(n_225),
.Y(n_1809)
);

AO21x2_ASAP7_75t_L g1810 ( 
.A1(n_1764),
.A2(n_227),
.B(n_228),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1728),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1750),
.B(n_229),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_SL g1813 ( 
.A(n_1725),
.B(n_230),
.Y(n_1813)
);

NOR2xp33_ASAP7_75t_L g1814 ( 
.A(n_1686),
.B(n_1749),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1744),
.B(n_230),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1706),
.B(n_231),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1750),
.A2(n_235),
.B1(n_232),
.B2(n_233),
.Y(n_1817)
);

INVx1_ASAP7_75t_SL g1818 ( 
.A(n_1726),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1751),
.B(n_232),
.Y(n_1819)
);

INVx2_ASAP7_75t_SL g1820 ( 
.A(n_1689),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1692),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1695),
.B(n_233),
.Y(n_1822)
);

INVxp67_ASAP7_75t_SL g1823 ( 
.A(n_1762),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_L g1824 ( 
.A(n_1715),
.B(n_235),
.Y(n_1824)
);

OAI22xp5_ASAP7_75t_L g1825 ( 
.A1(n_1693),
.A2(n_238),
.B1(n_236),
.B2(n_237),
.Y(n_1825)
);

AND2x4_ASAP7_75t_L g1826 ( 
.A(n_1694),
.B(n_237),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1731),
.Y(n_1827)
);

INVx2_ASAP7_75t_SL g1828 ( 
.A(n_1691),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1690),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1700),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1747),
.Y(n_1831)
);

AOI222xp33_ASAP7_75t_L g1832 ( 
.A1(n_1757),
.A2(n_241),
.B1(n_243),
.B2(n_239),
.C1(n_240),
.C2(n_242),
.Y(n_1832)
);

INVx4_ASAP7_75t_L g1833 ( 
.A(n_1742),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1721),
.Y(n_1834)
);

INVx1_ASAP7_75t_SL g1835 ( 
.A(n_1713),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1729),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1755),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1716),
.B(n_1759),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1734),
.B(n_239),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1717),
.B(n_241),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1732),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1738),
.B(n_1739),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1688),
.Y(n_1843)
);

OAI21xp5_ASAP7_75t_L g1844 ( 
.A1(n_1760),
.A2(n_242),
.B(n_243),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1702),
.B(n_244),
.Y(n_1845)
);

BUFx2_ASAP7_75t_L g1846 ( 
.A(n_1711),
.Y(n_1846)
);

NOR2x1p5_ASAP7_75t_L g1847 ( 
.A(n_1753),
.B(n_245),
.Y(n_1847)
);

INVx1_ASAP7_75t_SL g1848 ( 
.A(n_1704),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1712),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1708),
.B(n_247),
.Y(n_1850)
);

CKINVDCx14_ASAP7_75t_R g1851 ( 
.A(n_1714),
.Y(n_1851)
);

INVx3_ASAP7_75t_L g1852 ( 
.A(n_1753),
.Y(n_1852)
);

BUFx3_ASAP7_75t_L g1853 ( 
.A(n_1704),
.Y(n_1853)
);

AO21x2_ASAP7_75t_L g1854 ( 
.A1(n_1687),
.A2(n_248),
.B(n_250),
.Y(n_1854)
);

CKINVDCx16_ASAP7_75t_R g1855 ( 
.A(n_1752),
.Y(n_1855)
);

INVx1_ASAP7_75t_SL g1856 ( 
.A(n_1704),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1705),
.B(n_251),
.Y(n_1857)
);

AO21x2_ASAP7_75t_L g1858 ( 
.A1(n_1687),
.A2(n_252),
.B(n_253),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1712),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1756),
.B(n_253),
.Y(n_1860)
);

BUFx3_ASAP7_75t_L g1861 ( 
.A(n_1704),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1712),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1705),
.B(n_254),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1756),
.B(n_255),
.Y(n_1864)
);

INVx1_ASAP7_75t_SL g1865 ( 
.A(n_1704),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1712),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1712),
.Y(n_1867)
);

AND2x4_ASAP7_75t_L g1868 ( 
.A(n_1710),
.B(n_256),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1756),
.B(n_257),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1756),
.B(n_258),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1708),
.B(n_259),
.Y(n_1871)
);

AOI222xp33_ASAP7_75t_L g1872 ( 
.A1(n_1757),
.A2(n_261),
.B1(n_263),
.B2(n_259),
.C1(n_260),
.C2(n_262),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1756),
.B(n_261),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1756),
.B(n_264),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1708),
.B(n_265),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1712),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1712),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1712),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1708),
.B(n_265),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1712),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1712),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1705),
.B(n_266),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1712),
.Y(n_1883)
);

OR2x2_ASAP7_75t_L g1884 ( 
.A(n_1705),
.B(n_269),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1712),
.Y(n_1885)
);

CKINVDCx16_ASAP7_75t_R g1886 ( 
.A(n_1855),
.Y(n_1886)
);

INVx1_ASAP7_75t_SL g1887 ( 
.A(n_1848),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1852),
.B(n_270),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1791),
.Y(n_1889)
);

AOI22xp33_ASAP7_75t_L g1890 ( 
.A1(n_1806),
.A2(n_273),
.B1(n_271),
.B2(n_272),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1786),
.B(n_273),
.Y(n_1891)
);

OAI322xp33_ASAP7_75t_L g1892 ( 
.A1(n_1850),
.A2(n_279),
.A3(n_278),
.B1(n_276),
.B2(n_274),
.C1(n_275),
.C2(n_277),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1803),
.B(n_274),
.Y(n_1893)
);

INVx1_ASAP7_75t_SL g1894 ( 
.A(n_1856),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1823),
.B(n_280),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1772),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1778),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1792),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1781),
.Y(n_1899)
);

INVx1_ASAP7_75t_SL g1900 ( 
.A(n_1865),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1771),
.B(n_1773),
.Y(n_1901)
);

AOI221xp5_ASAP7_75t_L g1902 ( 
.A1(n_1871),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.C(n_284),
.Y(n_1902)
);

O2A1O1Ixp33_ASAP7_75t_L g1903 ( 
.A1(n_1875),
.A2(n_284),
.B(n_281),
.C(n_283),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1806),
.B(n_285),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1849),
.Y(n_1905)
);

OAI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1806),
.A2(n_287),
.B1(n_288),
.B2(n_434),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_SL g1907 ( 
.A(n_1833),
.B(n_288),
.Y(n_1907)
);

NOR2x1_ASAP7_75t_L g1908 ( 
.A(n_1879),
.B(n_436),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1859),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1820),
.B(n_441),
.Y(n_1910)
);

NOR2xp33_ASAP7_75t_SL g1911 ( 
.A(n_1769),
.B(n_442),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1828),
.B(n_443),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1862),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1866),
.Y(n_1914)
);

HB1xp67_ASAP7_75t_L g1915 ( 
.A(n_1811),
.Y(n_1915)
);

INVx1_ASAP7_75t_SL g1916 ( 
.A(n_1767),
.Y(n_1916)
);

O2A1O1Ixp33_ASAP7_75t_L g1917 ( 
.A1(n_1846),
.A2(n_451),
.B(n_449),
.C(n_450),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1867),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1876),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1807),
.Y(n_1920)
);

AOI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1779),
.A2(n_454),
.B1(n_452),
.B2(n_453),
.Y(n_1921)
);

INVx1_ASAP7_75t_SL g1922 ( 
.A(n_1853),
.Y(n_1922)
);

INVxp67_ASAP7_75t_SL g1923 ( 
.A(n_1838),
.Y(n_1923)
);

AND2x4_ASAP7_75t_L g1924 ( 
.A(n_1793),
.B(n_458),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1821),
.B(n_461),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1877),
.Y(n_1926)
);

NAND2x1_ASAP7_75t_L g1927 ( 
.A(n_1868),
.B(n_464),
.Y(n_1927)
);

AOI21xp33_ASAP7_75t_L g1928 ( 
.A1(n_1832),
.A2(n_465),
.B(n_466),
.Y(n_1928)
);

OAI22xp33_ASAP7_75t_SL g1929 ( 
.A1(n_1812),
.A2(n_470),
.B1(n_468),
.B2(n_469),
.Y(n_1929)
);

OAI22xp5_ASAP7_75t_L g1930 ( 
.A1(n_1817),
.A2(n_1829),
.B1(n_1831),
.B2(n_1830),
.Y(n_1930)
);

AOI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1844),
.A2(n_474),
.B1(n_472),
.B2(n_473),
.Y(n_1931)
);

INVxp67_ASAP7_75t_SL g1932 ( 
.A(n_1861),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1800),
.B(n_476),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_SL g1934 ( 
.A(n_1837),
.B(n_477),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1878),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1880),
.Y(n_1936)
);

AOI22xp5_ASAP7_75t_L g1937 ( 
.A1(n_1834),
.A2(n_1814),
.B1(n_1843),
.B2(n_1836),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1804),
.B(n_1797),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1798),
.B(n_479),
.Y(n_1939)
);

AOI22xp33_ASAP7_75t_SL g1940 ( 
.A1(n_1782),
.A2(n_483),
.B1(n_480),
.B2(n_482),
.Y(n_1940)
);

AOI21xp5_ASAP7_75t_L g1941 ( 
.A1(n_1842),
.A2(n_484),
.B(n_485),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1881),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1801),
.Y(n_1943)
);

NOR4xp25_ASAP7_75t_L g1944 ( 
.A(n_1780),
.B(n_488),
.C(n_486),
.D(n_487),
.Y(n_1944)
);

AOI22xp5_ASAP7_75t_L g1945 ( 
.A1(n_1835),
.A2(n_500),
.B1(n_496),
.B2(n_498),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1799),
.B(n_502),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1787),
.B(n_1827),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1857),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1863),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1883),
.Y(n_1950)
);

INVxp67_ASAP7_75t_L g1951 ( 
.A(n_1768),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1885),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1882),
.Y(n_1953)
);

INVx1_ASAP7_75t_SL g1954 ( 
.A(n_1860),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1864),
.B(n_508),
.Y(n_1955)
);

AOI21xp5_ASAP7_75t_L g1956 ( 
.A1(n_1818),
.A2(n_511),
.B(n_513),
.Y(n_1956)
);

NOR2xp33_ASAP7_75t_L g1957 ( 
.A(n_1776),
.B(n_515),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1884),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1785),
.Y(n_1959)
);

INVxp67_ASAP7_75t_L g1960 ( 
.A(n_1869),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1841),
.Y(n_1961)
);

OAI21xp5_ASAP7_75t_SL g1962 ( 
.A1(n_1872),
.A2(n_526),
.B(n_529),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1789),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1810),
.B(n_530),
.Y(n_1964)
);

INVxp67_ASAP7_75t_L g1965 ( 
.A(n_1870),
.Y(n_1965)
);

INVx3_ASAP7_75t_L g1966 ( 
.A(n_1886),
.Y(n_1966)
);

INVx1_ASAP7_75t_SL g1967 ( 
.A(n_1916),
.Y(n_1967)
);

INVx1_ASAP7_75t_SL g1968 ( 
.A(n_1954),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1923),
.B(n_1854),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1915),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1963),
.B(n_1858),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1932),
.B(n_1873),
.Y(n_1972)
);

INVxp67_ASAP7_75t_L g1973 ( 
.A(n_1904),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1959),
.B(n_1775),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1938),
.Y(n_1975)
);

HB1xp67_ASAP7_75t_L g1976 ( 
.A(n_1887),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1924),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1893),
.B(n_1895),
.Y(n_1978)
);

NAND3xp33_ASAP7_75t_L g1979 ( 
.A(n_1902),
.B(n_1788),
.C(n_1825),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1947),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1961),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1901),
.B(n_1874),
.Y(n_1982)
);

OR2x2_ASAP7_75t_L g1983 ( 
.A(n_1889),
.B(n_1783),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1894),
.B(n_1774),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1951),
.B(n_1794),
.Y(n_1985)
);

INVxp67_ASAP7_75t_L g1986 ( 
.A(n_1907),
.Y(n_1986)
);

INVxp67_ASAP7_75t_L g1987 ( 
.A(n_1908),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1960),
.B(n_1965),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1900),
.B(n_1808),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1903),
.B(n_1824),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1898),
.B(n_1796),
.Y(n_1991)
);

NAND3xp33_ASAP7_75t_L g1992 ( 
.A(n_1962),
.B(n_1840),
.C(n_1790),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1922),
.B(n_1822),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1896),
.Y(n_1994)
);

CKINVDCx16_ASAP7_75t_R g1995 ( 
.A(n_1911),
.Y(n_1995)
);

AND2x4_ASAP7_75t_L g1996 ( 
.A(n_1891),
.B(n_1847),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1888),
.B(n_1816),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1897),
.Y(n_1998)
);

OAI22xp5_ASAP7_75t_L g1999 ( 
.A1(n_1930),
.A2(n_1851),
.B1(n_1839),
.B2(n_1819),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_SL g2000 ( 
.A(n_1924),
.B(n_1815),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1899),
.B(n_1805),
.Y(n_2001)
);

INVx1_ASAP7_75t_SL g2002 ( 
.A(n_1955),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1905),
.B(n_1826),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1953),
.B(n_1777),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1909),
.Y(n_2005)
);

INVx2_ASAP7_75t_SL g2006 ( 
.A(n_1927),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1913),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1914),
.B(n_1795),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1918),
.Y(n_2009)
);

INVxp67_ASAP7_75t_SL g2010 ( 
.A(n_1941),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1919),
.Y(n_2011)
);

INVxp67_ASAP7_75t_SL g2012 ( 
.A(n_1934),
.Y(n_2012)
);

AND2x4_ASAP7_75t_L g2013 ( 
.A(n_1920),
.B(n_1784),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1926),
.B(n_1802),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1935),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1936),
.B(n_1809),
.Y(n_2016)
);

AND2x4_ASAP7_75t_L g2017 ( 
.A(n_1942),
.B(n_1845),
.Y(n_2017)
);

NAND2xp33_ASAP7_75t_SL g2018 ( 
.A(n_1950),
.B(n_1813),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1952),
.B(n_1948),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1943),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1949),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1958),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1964),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_SL g2024 ( 
.A(n_1929),
.B(n_1770),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1976),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1966),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1988),
.Y(n_2027)
);

AND2x4_ASAP7_75t_SL g2028 ( 
.A(n_1972),
.B(n_1957),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1997),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1993),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_2019),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1981),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1982),
.B(n_1984),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1996),
.Y(n_2034)
);

CKINVDCx20_ASAP7_75t_R g2035 ( 
.A(n_1967),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2021),
.Y(n_2036)
);

BUFx2_ASAP7_75t_L g2037 ( 
.A(n_1989),
.Y(n_2037)
);

INVx1_ASAP7_75t_SL g2038 ( 
.A(n_1978),
.Y(n_2038)
);

INVx1_ASAP7_75t_SL g2039 ( 
.A(n_1968),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_2022),
.Y(n_2040)
);

HB1xp67_ASAP7_75t_L g2041 ( 
.A(n_1985),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_2001),
.B(n_1937),
.Y(n_2042)
);

BUFx2_ASAP7_75t_L g2043 ( 
.A(n_2018),
.Y(n_2043)
);

HB1xp67_ASAP7_75t_L g2044 ( 
.A(n_1986),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1994),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1998),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2005),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2007),
.Y(n_2048)
);

CKINVDCx5p33_ASAP7_75t_R g2049 ( 
.A(n_1995),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_2009),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2011),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2015),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1983),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1970),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2004),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1974),
.Y(n_2056)
);

NOR2x1_ASAP7_75t_L g2057 ( 
.A(n_2035),
.B(n_1992),
.Y(n_2057)
);

NOR2x1_ASAP7_75t_L g2058 ( 
.A(n_2025),
.B(n_1979),
.Y(n_2058)
);

NAND3xp33_ASAP7_75t_L g2059 ( 
.A(n_2043),
.B(n_2049),
.C(n_2025),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_2039),
.B(n_2003),
.Y(n_2060)
);

OAI22xp5_ASAP7_75t_L g2061 ( 
.A1(n_2044),
.A2(n_2010),
.B1(n_2012),
.B2(n_1990),
.Y(n_2061)
);

AOI21xp5_ASAP7_75t_L g2062 ( 
.A1(n_2042),
.A2(n_2024),
.B(n_1987),
.Y(n_2062)
);

NOR3xp33_ASAP7_75t_L g2063 ( 
.A(n_2037),
.B(n_1969),
.C(n_1973),
.Y(n_2063)
);

NAND3xp33_ASAP7_75t_L g2064 ( 
.A(n_2026),
.B(n_1999),
.C(n_1890),
.Y(n_2064)
);

NAND3xp33_ASAP7_75t_L g2065 ( 
.A(n_2030),
.B(n_1917),
.C(n_2023),
.Y(n_2065)
);

AND2x4_ASAP7_75t_L g2066 ( 
.A(n_2033),
.B(n_2013),
.Y(n_2066)
);

NAND4xp25_ASAP7_75t_L g2067 ( 
.A(n_2038),
.B(n_1980),
.C(n_1975),
.D(n_1971),
.Y(n_2067)
);

OAI22xp5_ASAP7_75t_L g2068 ( 
.A1(n_2029),
.A2(n_2006),
.B1(n_2002),
.B2(n_2017),
.Y(n_2068)
);

OAI21xp33_ASAP7_75t_L g2069 ( 
.A1(n_2034),
.A2(n_2016),
.B(n_2014),
.Y(n_2069)
);

NOR2x1_ASAP7_75t_L g2070 ( 
.A(n_2027),
.B(n_2008),
.Y(n_2070)
);

AOI211xp5_ASAP7_75t_L g2071 ( 
.A1(n_2031),
.A2(n_1906),
.B(n_1892),
.C(n_1944),
.Y(n_2071)
);

AOI222xp33_ASAP7_75t_L g2072 ( 
.A1(n_2036),
.A2(n_2020),
.B1(n_2040),
.B2(n_2053),
.C1(n_2054),
.C2(n_2056),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2041),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_SL g2074 ( 
.A(n_2028),
.B(n_2017),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_2066),
.Y(n_2075)
);

NOR4xp25_ASAP7_75t_L g2076 ( 
.A(n_2059),
.B(n_2032),
.C(n_2046),
.D(n_2045),
.Y(n_2076)
);

AOI21xp33_ASAP7_75t_SL g2077 ( 
.A1(n_2060),
.A2(n_2055),
.B(n_2048),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_2066),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_SL g2079 ( 
.A(n_2057),
.B(n_1991),
.Y(n_2079)
);

HB1xp67_ASAP7_75t_L g2080 ( 
.A(n_2058),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2073),
.Y(n_2081)
);

NOR3x1_ASAP7_75t_L g2082 ( 
.A(n_2064),
.B(n_2052),
.C(n_2050),
.Y(n_2082)
);

OAI31xp33_ASAP7_75t_L g2083 ( 
.A1(n_2062),
.A2(n_1928),
.A3(n_2051),
.B(n_2047),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2080),
.B(n_2069),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2075),
.Y(n_2085)
);

NOR4xp25_ASAP7_75t_L g2086 ( 
.A(n_2079),
.B(n_2061),
.C(n_2067),
.D(n_2074),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2078),
.B(n_2070),
.Y(n_2087)
);

INVx3_ASAP7_75t_L g2088 ( 
.A(n_2081),
.Y(n_2088)
);

AND3x1_ASAP7_75t_L g2089 ( 
.A(n_2076),
.B(n_2063),
.C(n_2071),
.Y(n_2089)
);

NOR2x1_ASAP7_75t_L g2090 ( 
.A(n_2082),
.B(n_2068),
.Y(n_2090)
);

HB1xp67_ASAP7_75t_L g2091 ( 
.A(n_2077),
.Y(n_2091)
);

NAND3xp33_ASAP7_75t_L g2092 ( 
.A(n_2089),
.B(n_2083),
.C(n_2072),
.Y(n_2092)
);

NOR2xp33_ASAP7_75t_R g2093 ( 
.A(n_2087),
.B(n_1910),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_SL g2094 ( 
.A(n_2086),
.B(n_2065),
.Y(n_2094)
);

NOR2xp33_ASAP7_75t_R g2095 ( 
.A(n_2088),
.B(n_1912),
.Y(n_2095)
);

XNOR2x1_ASAP7_75t_L g2096 ( 
.A(n_2090),
.B(n_1977),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2096),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_2094),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_2098),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2099),
.B(n_2091),
.Y(n_2100)
);

AOI31xp33_ASAP7_75t_L g2101 ( 
.A1(n_2100),
.A2(n_2084),
.A3(n_2097),
.B(n_2092),
.Y(n_2101)
);

OAI22xp5_ASAP7_75t_SL g2102 ( 
.A1(n_2101),
.A2(n_2085),
.B1(n_2093),
.B2(n_2095),
.Y(n_2102)
);

OAI211xp5_ASAP7_75t_L g2103 ( 
.A1(n_2102),
.A2(n_2000),
.B(n_1939),
.C(n_1946),
.Y(n_2103)
);

INVxp67_ASAP7_75t_L g2104 ( 
.A(n_2103),
.Y(n_2104)
);

OAI221xp5_ASAP7_75t_R g2105 ( 
.A1(n_2104),
.A2(n_1945),
.B1(n_1940),
.B2(n_1921),
.C(n_1931),
.Y(n_2105)
);

AOI211xp5_ASAP7_75t_L g2106 ( 
.A1(n_2105),
.A2(n_1956),
.B(n_1933),
.C(n_1925),
.Y(n_2106)
);


endmodule