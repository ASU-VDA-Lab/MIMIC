module fake_jpeg_2724_n_437 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_437);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_437;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_6),
.B(n_5),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_1),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_19),
.A2(n_9),
.B1(n_14),
.B2(n_2),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_48),
.A2(n_25),
.B1(n_32),
.B2(n_38),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_19),
.B(n_8),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_54),
.B(n_57),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_31),
.B(n_8),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_59),
.Y(n_146)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_21),
.B(n_8),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_62),
.B(n_72),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_63),
.Y(n_129)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_64),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_67),
.Y(n_124)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_68),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_46),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_90),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_70),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_71),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_37),
.B(n_6),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_37),
.B(n_31),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_75),
.B(n_80),
.Y(n_135)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_33),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_34),
.B(n_43),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_24),
.B(n_6),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_83),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_10),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_82),
.B(n_93),
.Y(n_106)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_24),
.B(n_10),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_86),
.Y(n_111)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_16),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_89),
.B(n_25),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_39),
.B(n_10),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_23),
.Y(n_91)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_16),
.Y(n_92)
);

AOI21xp33_ASAP7_75t_SL g110 ( 
.A1(n_92),
.A2(n_44),
.B(n_40),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_39),
.B(n_15),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_73),
.A2(n_44),
.B1(n_45),
.B2(n_42),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_107),
.A2(n_63),
.B1(n_71),
.B2(n_70),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_110),
.A2(n_126),
.B(n_116),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_87),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_113),
.B(n_114),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_91),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_69),
.A2(n_45),
.B1(n_44),
.B2(n_26),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_116),
.A2(n_130),
.B1(n_132),
.B2(n_77),
.Y(n_153)
);

NAND2xp67_ASAP7_75t_SL g125 ( 
.A(n_48),
.B(n_45),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_SL g192 ( 
.A(n_125),
.B(n_142),
.C(n_122),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_52),
.B(n_38),
.C(n_26),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_50),
.A2(n_38),
.B1(n_60),
.B2(n_61),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_51),
.A2(n_38),
.B1(n_42),
.B2(n_28),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g136 ( 
.A(n_67),
.B(n_38),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_136),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_78),
.A2(n_32),
.B1(n_28),
.B2(n_36),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_138),
.A2(n_79),
.B1(n_68),
.B2(n_49),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_59),
.B(n_36),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_139),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_84),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_140),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_141),
.A2(n_0),
.B1(n_1),
.B2(n_15),
.Y(n_163)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_51),
.Y(n_142)
);

INVx11_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_77),
.B(n_12),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_145),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_149),
.A2(n_159),
.B1(n_129),
.B2(n_112),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_92),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_150),
.B(n_156),
.Y(n_207)
);

OA22x2_ASAP7_75t_L g223 ( 
.A1(n_153),
.A2(n_134),
.B1(n_149),
.B2(n_191),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_123),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_155),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_88),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_157),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_158),
.A2(n_174),
.B1(n_161),
.B2(n_165),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_100),
.A2(n_56),
.B1(n_66),
.B2(n_55),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_141),
.A2(n_47),
.B1(n_58),
.B2(n_40),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_160),
.A2(n_166),
.B1(n_193),
.B2(n_121),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_125),
.A2(n_53),
.B1(n_74),
.B2(n_35),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_161),
.A2(n_163),
.B1(n_165),
.B2(n_168),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_103),
.A2(n_35),
.B(n_29),
.C(n_2),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_162),
.A2(n_184),
.B(n_147),
.C(n_131),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_107),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_108),
.A2(n_11),
.B1(n_13),
.B2(n_3),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_94),
.Y(n_167)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_167),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_L g168 ( 
.A1(n_132),
.A2(n_3),
.B1(n_4),
.B2(n_11),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_96),
.Y(n_169)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_169),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_118),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_104),
.Y(n_204)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_94),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_171),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_95),
.A2(n_3),
.B1(n_4),
.B2(n_12),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_173),
.A2(n_181),
.B1(n_183),
.B2(n_191),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_130),
.A2(n_12),
.B1(n_15),
.B2(n_0),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_95),
.B(n_1),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_179),
.Y(n_210)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_178),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_111),
.B(n_1),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_115),
.Y(n_180)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_126),
.A2(n_106),
.B1(n_127),
.B2(n_102),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_119),
.Y(n_182)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_99),
.A2(n_120),
.B1(n_97),
.B2(n_133),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_135),
.A2(n_109),
.B(n_118),
.C(n_124),
.Y(n_184)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_105),
.Y(n_185)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

AO22x1_ASAP7_75t_L g186 ( 
.A1(n_108),
.A2(n_122),
.B1(n_98),
.B2(n_137),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_186),
.A2(n_105),
.B(n_146),
.Y(n_197)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_97),
.B(n_143),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_188),
.B(n_194),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_189),
.Y(n_213)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_98),
.Y(n_190)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_96),
.A2(n_128),
.B1(n_134),
.B2(n_131),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_192),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_137),
.A2(n_146),
.B1(n_104),
.B2(n_121),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_101),
.B(n_102),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_101),
.Y(n_195)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_197),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_198),
.A2(n_175),
.B1(n_155),
.B2(n_185),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_164),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_208),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_202),
.B(n_223),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_204),
.Y(n_262)
);

AOI32xp33_ASAP7_75t_L g208 ( 
.A1(n_150),
.A2(n_104),
.A3(n_112),
.B1(n_117),
.B2(n_128),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_152),
.B(n_117),
.C(n_129),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_194),
.C(n_195),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_148),
.B(n_147),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_219),
.B(n_225),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_220),
.B(n_235),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_148),
.B(n_154),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_154),
.B(n_172),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_228),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_227),
.A2(n_232),
.B1(n_162),
.B2(n_163),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_172),
.B(n_179),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_188),
.Y(n_230)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_230),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_177),
.B(n_181),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_175),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_189),
.A2(n_151),
.B1(n_152),
.B2(n_156),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_164),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_234),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_151),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_184),
.B(n_173),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_236),
.B(n_255),
.C(n_260),
.Y(n_273)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_240),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_200),
.B(n_170),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_241),
.B(n_244),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_243),
.A2(n_266),
.B1(n_270),
.B2(n_210),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_190),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_219),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_246),
.B(n_263),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_167),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_247),
.B(n_254),
.Y(n_287)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_249),
.Y(n_290)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_221),
.Y(n_250)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_250),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_213),
.A2(n_186),
.B1(n_180),
.B2(n_178),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_251),
.A2(n_252),
.B(n_259),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_213),
.A2(n_186),
.B(n_178),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_171),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_187),
.C(n_176),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_207),
.B(n_183),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_256),
.B(n_203),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_215),
.A2(n_182),
.B1(n_169),
.B2(n_157),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_257),
.A2(n_214),
.B1(n_201),
.B2(n_203),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_207),
.B(n_155),
.C(n_169),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_261),
.B(n_256),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_204),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_212),
.Y(n_264)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_230),
.B(n_209),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_268),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_209),
.A2(n_227),
.B1(n_199),
.B2(n_222),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_197),
.B(n_218),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_267),
.B(n_269),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_210),
.B(n_220),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_235),
.B(n_222),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_199),
.A2(n_223),
.B1(n_208),
.B2(n_215),
.Y(n_270)
);

OA22x2_ASAP7_75t_L g271 ( 
.A1(n_251),
.A2(n_223),
.B1(n_214),
.B2(n_221),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_271),
.B(n_281),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_236),
.B(n_265),
.C(n_267),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_293),
.C(n_263),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_237),
.A2(n_223),
.B1(n_228),
.B2(n_226),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_275),
.A2(n_211),
.B1(n_217),
.B2(n_196),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_278),
.A2(n_296),
.B1(n_257),
.B2(n_248),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_252),
.A2(n_223),
.B(n_216),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_279),
.A2(n_243),
.B(n_264),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_238),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_245),
.B(n_211),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_283),
.B(n_286),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_285),
.A2(n_262),
.B1(n_258),
.B2(n_264),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_238),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_289),
.B(n_300),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_247),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_297),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_253),
.C(n_255),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_294),
.B(n_289),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_248),
.A2(n_212),
.B1(n_201),
.B2(n_216),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_295),
.A2(n_249),
.B1(n_250),
.B2(n_248),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_270),
.A2(n_212),
.B1(n_217),
.B2(n_196),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_244),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_240),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_298),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_246),
.B(n_239),
.Y(n_299)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_299),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_241),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_239),
.B(n_245),
.Y(n_301)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_301),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_302),
.A2(n_306),
.B1(n_325),
.B2(n_297),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_303),
.B(n_309),
.C(n_311),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_304),
.B(n_287),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_278),
.A2(n_237),
.B1(n_268),
.B2(n_242),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_279),
.A2(n_242),
.B(n_269),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_307),
.B(n_277),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_SL g308 ( 
.A(n_275),
.B(n_248),
.C(n_266),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_308),
.B(n_272),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_273),
.B(n_267),
.C(n_253),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_310),
.A2(n_317),
.B1(n_326),
.B2(n_329),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_273),
.B(n_269),
.C(n_260),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_274),
.B(n_254),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_312),
.B(n_313),
.C(n_321),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_261),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_258),
.C(n_262),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_294),
.B(n_256),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_322),
.B(n_327),
.C(n_291),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_299),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_281),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_282),
.Y(n_324)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_324),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_272),
.B(n_205),
.C(n_206),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_296),
.A2(n_205),
.B1(n_229),
.B2(n_206),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_328),
.A2(n_285),
.B1(n_291),
.B2(n_290),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_300),
.A2(n_229),
.B1(n_282),
.B2(n_286),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_330),
.A2(n_335),
.B(n_322),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_331),
.A2(n_345),
.B1(n_348),
.B2(n_353),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_332),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_312),
.B(n_311),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_333),
.B(n_337),
.C(n_352),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_301),
.Y(n_334)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_334),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_309),
.B(n_288),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_315),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_338),
.B(n_327),
.Y(n_371)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_314),
.Y(n_341)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_341),
.Y(n_374)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_314),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_342),
.B(n_346),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_306),
.B(n_288),
.Y(n_344)
);

NAND3xp33_ASAP7_75t_L g366 ( 
.A(n_344),
.B(n_351),
.C(n_284),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_302),
.A2(n_292),
.B1(n_277),
.B2(n_295),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_318),
.B(n_283),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_318),
.B(n_287),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_347),
.B(n_320),
.Y(n_361)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_329),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_320),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_349),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_350),
.B(n_313),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_324),
.B(n_229),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_348),
.A2(n_316),
.B1(n_325),
.B2(n_310),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_354),
.A2(n_355),
.B1(n_358),
.B2(n_368),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_339),
.A2(n_316),
.B1(n_319),
.B2(n_326),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_341),
.A2(n_308),
.B1(n_319),
.B2(n_307),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_360),
.B(n_350),
.Y(n_388)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_361),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_345),
.A2(n_305),
.B1(n_271),
.B2(n_276),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_362),
.B(n_369),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_333),
.B(n_303),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_365),
.B(n_373),
.Y(n_376)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_366),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_336),
.B(n_321),
.C(n_304),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_367),
.B(n_343),
.C(n_336),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_331),
.A2(n_342),
.B1(n_332),
.B2(n_334),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_330),
.A2(n_271),
.B1(n_276),
.B2(n_290),
.Y(n_369)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_371),
.Y(n_385)
);

NOR2x1_ASAP7_75t_L g389 ( 
.A(n_372),
.B(n_358),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_347),
.A2(n_271),
.B1(n_284),
.B2(n_298),
.Y(n_373)
);

NAND4xp25_ASAP7_75t_L g377 ( 
.A(n_368),
.B(n_340),
.C(n_353),
.D(n_280),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_377),
.B(n_386),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_364),
.B(n_352),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_378),
.B(n_388),
.C(n_390),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_379),
.B(n_384),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_357),
.A2(n_340),
.B(n_346),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_381),
.A2(n_374),
.B(n_370),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_365),
.B(n_343),
.C(n_337),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_364),
.B(n_372),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_359),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_387),
.A2(n_370),
.B1(n_374),
.B2(n_359),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_389),
.B(n_362),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_360),
.B(n_271),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_391),
.A2(n_397),
.B(n_363),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_381),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_SL g411 ( 
.A1(n_392),
.A2(n_393),
.B1(n_403),
.B2(n_363),
.Y(n_411)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_382),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_378),
.B(n_367),
.C(n_356),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_395),
.B(n_398),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_380),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_399),
.A2(n_376),
.B(n_328),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_389),
.A2(n_354),
.B(n_355),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_400),
.A2(n_384),
.B(n_379),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_385),
.B(n_349),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_401),
.Y(n_409)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_380),
.Y(n_403)
);

INVx11_ASAP7_75t_L g404 ( 
.A(n_396),
.Y(n_404)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_404),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_403),
.A2(n_375),
.B1(n_373),
.B2(n_369),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_406),
.B(n_407),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_393),
.B(n_383),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_392),
.A2(n_375),
.B1(n_376),
.B2(n_390),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_408),
.B(n_400),
.Y(n_416)
);

AO21x1_ASAP7_75t_L g419 ( 
.A1(n_410),
.A2(n_411),
.B(n_413),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_402),
.B(n_386),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_412),
.B(n_394),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_414),
.A2(n_280),
.B(n_388),
.Y(n_423)
);

BUFx24_ASAP7_75t_SL g415 ( 
.A(n_405),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_415),
.B(n_420),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_416),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_414),
.B(n_395),
.C(n_401),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g424 ( 
.A(n_417),
.B(n_418),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_410),
.B(n_394),
.C(n_399),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_423),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_419),
.A2(n_409),
.B(n_408),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_425),
.A2(n_421),
.B(n_406),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_422),
.B(n_419),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_427),
.B(n_404),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_424),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_430),
.Y(n_433)
);

AOI21x1_ASAP7_75t_L g434 ( 
.A1(n_431),
.A2(n_432),
.B(n_429),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_434),
.B(n_428),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_435),
.A2(n_433),
.B(n_426),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_436),
.B(n_426),
.Y(n_437)
);


endmodule