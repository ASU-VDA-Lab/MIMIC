module fake_netlist_6_2381_n_1925 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1925);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1925;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx10_ASAP7_75t_L g185 ( 
.A(n_9),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_7),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_73),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_77),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_166),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_163),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_80),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_2),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_180),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_5),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_139),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_111),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_138),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_29),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_39),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_24),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_8),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_64),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_171),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_120),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_130),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_45),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_88),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_36),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_47),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_134),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_61),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_172),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_108),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_169),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_14),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_43),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_95),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_10),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_48),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_36),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_37),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_156),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_183),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_29),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_81),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_178),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_132),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_104),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_174),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_84),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_117),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_116),
.Y(n_233)
);

BUFx8_ASAP7_75t_SL g234 ( 
.A(n_168),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_47),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_157),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_94),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_114),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_127),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_87),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_136),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_72),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_20),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_31),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_17),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_18),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_63),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_158),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_23),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_106),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_122),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_121),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_44),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_3),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_154),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_41),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_57),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_79),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_75),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_8),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_50),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_149),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_142),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_23),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_110),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_68),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_2),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_59),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_18),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_48),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_102),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_15),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_0),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_56),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_173),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_10),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_129),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_12),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_19),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_70),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_153),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_119),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_89),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_165),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_37),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_105),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_7),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_60),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_49),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_33),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_3),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_83),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_21),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_9),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_66),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_144),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_133),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_34),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_97),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_148),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_51),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_176),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_164),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_6),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g305 ( 
.A(n_41),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_46),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_54),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_35),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_43),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_5),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_82),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_175),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_35),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_22),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_91),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_15),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_92),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_99),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_150),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_135),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_159),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_30),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_93),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_112),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_160),
.Y(n_325)
);

BUFx10_ASAP7_75t_L g326 ( 
.A(n_40),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_4),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_0),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_20),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_151),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_123),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_22),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_55),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_107),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_52),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_128),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_62),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_69),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_113),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_67),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_51),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_19),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_118),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_181),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_147),
.Y(n_345)
);

INVx2_ASAP7_75t_SL g346 ( 
.A(n_14),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_25),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_34),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_115),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_71),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_103),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_54),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_137),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_12),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_55),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_17),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_1),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_30),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_126),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_182),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_125),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_33),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_141),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_86),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_46),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_109),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_11),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_162),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_228),
.Y(n_369)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_301),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_301),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_301),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_301),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_301),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_234),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_227),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_357),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_357),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_357),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_357),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_261),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_228),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_357),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_195),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_240),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_247),
.Y(n_386)
);

INVxp33_ASAP7_75t_SL g387 ( 
.A(n_332),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_313),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_313),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_229),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_233),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_324),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_231),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_192),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_328),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_236),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_206),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_208),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_217),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_221),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_238),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_241),
.Y(n_402)
);

INVxp67_ASAP7_75t_SL g403 ( 
.A(n_233),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_242),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_225),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_243),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_244),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_245),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_350),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_253),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_267),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_278),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_350),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_279),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_210),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_254),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_289),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_255),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_186),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_257),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_293),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_298),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_306),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_259),
.Y(n_424)
);

INVxp33_ASAP7_75t_L g425 ( 
.A(n_307),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_308),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_262),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_333),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_246),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_335),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_353),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_347),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_265),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_271),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_355),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_275),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_281),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_194),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_194),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_239),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_216),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_282),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_284),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_286),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_216),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_292),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_346),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_185),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_296),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_239),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_186),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_299),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_302),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_198),
.Y(n_454)
);

INVxp33_ASAP7_75t_SL g455 ( 
.A(n_198),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_303),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_256),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_311),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_346),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_348),
.Y(n_460)
);

NAND2xp33_ASAP7_75t_L g461 ( 
.A(n_376),
.B(n_199),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_371),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_382),
.B(n_348),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_371),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_383),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_370),
.B(n_353),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_383),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_370),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_370),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_416),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_372),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_451),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_390),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_372),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_375),
.B(n_263),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_415),
.A2(n_354),
.B1(n_358),
.B2(n_273),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_373),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_373),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_391),
.B(n_431),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_374),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_393),
.B(n_204),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_429),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_374),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_391),
.B(n_204),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_391),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_457),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_396),
.B(n_300),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_377),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_377),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_378),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_378),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_379),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_379),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_403),
.B(n_263),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_431),
.B(n_300),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_380),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_440),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_431),
.B(n_187),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_401),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_387),
.A2(n_362),
.B1(n_367),
.B2(n_199),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_380),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_422),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_440),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_422),
.Y(n_504)
);

BUFx2_ASAP7_75t_L g505 ( 
.A(n_395),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_409),
.B(n_263),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_402),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_450),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_455),
.B(n_187),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_450),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_394),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_394),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_397),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_397),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_398),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_381),
.A2(n_362),
.B1(n_367),
.B2(n_200),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_413),
.B(n_232),
.Y(n_517)
);

BUFx8_ASAP7_75t_L g518 ( 
.A(n_419),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_369),
.B(n_336),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_369),
.B(n_188),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_404),
.B(n_351),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_398),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_399),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_424),
.B(n_336),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_427),
.Y(n_525)
);

OA21x2_ASAP7_75t_L g526 ( 
.A1(n_399),
.A2(n_211),
.B(n_209),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_388),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_400),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_388),
.B(n_188),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_400),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_384),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_407),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_433),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_407),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_389),
.B(n_223),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_434),
.B(n_437),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_389),
.B(n_226),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_408),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_385),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_465),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_489),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_463),
.B(n_419),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_523),
.Y(n_543)
);

NOR2x1p5_ASAP7_75t_L g544 ( 
.A(n_473),
.B(n_200),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_489),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_489),
.Y(n_546)
);

AND3x2_ASAP7_75t_L g547 ( 
.A(n_470),
.B(n_448),
.C(n_414),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_523),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_523),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_517),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_523),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_485),
.B(n_442),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_521),
.B(n_444),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_485),
.B(n_449),
.Y(n_554)
);

NAND2xp33_ASAP7_75t_L g555 ( 
.A(n_487),
.B(n_230),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_482),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_527),
.Y(n_557)
);

INVxp33_ASAP7_75t_L g558 ( 
.A(n_486),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_527),
.Y(n_559)
);

BUFx6f_ASAP7_75t_SL g560 ( 
.A(n_519),
.Y(n_560)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_498),
.B(n_520),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_485),
.B(n_452),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_498),
.B(n_454),
.Y(n_563)
);

NAND2xp33_ASAP7_75t_L g564 ( 
.A(n_524),
.B(n_237),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_491),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_485),
.B(n_456),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_523),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_491),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_468),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_531),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_491),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_496),
.Y(n_572)
);

AOI21x1_ASAP7_75t_L g573 ( 
.A1(n_462),
.A2(n_250),
.B(n_248),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_496),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_465),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_523),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_517),
.B(n_458),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_496),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_463),
.A2(n_405),
.B1(n_406),
.B2(n_425),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_481),
.B(n_312),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_528),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_528),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_465),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_468),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_528),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_479),
.B(n_315),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_468),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_R g588 ( 
.A(n_499),
.B(n_418),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_503),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_507),
.B(n_420),
.Y(n_590)
);

OR2x6_ASAP7_75t_L g591 ( 
.A(n_536),
.B(n_438),
.Y(n_591)
);

BUFx6f_ASAP7_75t_SL g592 ( 
.A(n_519),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_479),
.B(n_318),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_527),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_525),
.B(n_436),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_503),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_503),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_497),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_497),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_468),
.Y(n_600)
);

INVx8_ASAP7_75t_L g601 ( 
.A(n_484),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_497),
.Y(n_602)
);

INVx4_ASAP7_75t_L g603 ( 
.A(n_468),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_533),
.B(n_443),
.Y(n_604)
);

INVx8_ASAP7_75t_L g605 ( 
.A(n_484),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_497),
.Y(n_606)
);

CKINVDCx6p67_ASAP7_75t_R g607 ( 
.A(n_539),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_494),
.B(n_446),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_494),
.B(n_453),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_497),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_518),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_518),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_497),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_469),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_506),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_465),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_509),
.B(n_392),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_506),
.Y(n_618)
);

AO22x2_ASAP7_75t_L g619 ( 
.A1(n_472),
.A2(n_264),
.B1(n_291),
.B2(n_320),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_528),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_479),
.B(n_319),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g622 ( 
.A(n_520),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_466),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_512),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_465),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_465),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_469),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_469),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_512),
.Y(n_629)
);

BUFx6f_ASAP7_75t_SL g630 ( 
.A(n_519),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_467),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_468),
.Y(n_632)
);

BUFx10_ASAP7_75t_L g633 ( 
.A(n_519),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_466),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_479),
.B(n_321),
.Y(n_635)
);

AND3x2_ASAP7_75t_L g636 ( 
.A(n_505),
.B(n_252),
.C(n_251),
.Y(n_636)
);

AND2x6_ASAP7_75t_L g637 ( 
.A(n_484),
.B(n_258),
.Y(n_637)
);

NOR3xp33_ASAP7_75t_SL g638 ( 
.A(n_500),
.B(n_219),
.C(n_201),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_462),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_466),
.B(n_408),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_467),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_466),
.B(n_484),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_461),
.A2(n_386),
.B1(n_207),
.B2(n_193),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_464),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_467),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_528),
.Y(n_646)
);

INVxp33_ASAP7_75t_L g647 ( 
.A(n_500),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_535),
.B(n_438),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_495),
.B(n_535),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_495),
.B(n_323),
.Y(n_650)
);

NAND2xp33_ASAP7_75t_L g651 ( 
.A(n_529),
.B(n_266),
.Y(n_651)
);

AND3x2_ASAP7_75t_L g652 ( 
.A(n_505),
.B(n_274),
.C(n_268),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_464),
.Y(n_653)
);

AND3x1_ASAP7_75t_L g654 ( 
.A(n_516),
.B(n_441),
.C(n_439),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_471),
.Y(n_655)
);

AND3x1_ASAP7_75t_L g656 ( 
.A(n_516),
.B(n_441),
.C(n_439),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_529),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_471),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_528),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_467),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_475),
.B(n_445),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_477),
.Y(n_662)
);

INVxp33_ASAP7_75t_L g663 ( 
.A(n_476),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_477),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_478),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_467),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_495),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_467),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_534),
.B(n_445),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_495),
.Y(n_670)
);

BUFx6f_ASAP7_75t_L g671 ( 
.A(n_474),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_518),
.Y(n_672)
);

XNOR2x2_ASAP7_75t_R g673 ( 
.A(n_476),
.B(n_1),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_478),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_483),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_513),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_483),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_535),
.B(n_447),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_488),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_535),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_488),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_534),
.B(n_447),
.Y(n_682)
);

NAND2xp33_ASAP7_75t_L g683 ( 
.A(n_534),
.B(n_280),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_518),
.B(n_189),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_537),
.B(n_189),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_490),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_490),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_537),
.B(n_190),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_534),
.B(n_459),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_474),
.Y(n_690)
);

OR2x2_ASAP7_75t_L g691 ( 
.A(n_537),
.B(n_460),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_537),
.B(n_492),
.Y(n_692)
);

INVxp67_ASAP7_75t_SL g693 ( 
.A(n_671),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_561),
.A2(n_526),
.B1(n_345),
.B2(n_283),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_622),
.B(n_526),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_614),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_550),
.B(n_288),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_623),
.Y(n_698)
);

AO22x2_ASAP7_75t_L g699 ( 
.A1(n_673),
.A2(n_295),
.B1(n_297),
.B2(n_317),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_561),
.B(n_190),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_657),
.B(n_191),
.Y(n_701)
);

INVxp33_ASAP7_75t_L g702 ( 
.A(n_558),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_556),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_550),
.B(n_191),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_615),
.B(n_193),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_615),
.B(n_325),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_618),
.B(n_331),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_640),
.B(n_513),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_542),
.B(n_514),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_553),
.B(n_618),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_563),
.B(n_196),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_542),
.B(n_556),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_680),
.B(n_334),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_614),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_680),
.B(n_339),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_667),
.B(n_526),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_667),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_627),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_678),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_670),
.B(n_526),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_627),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_670),
.B(n_492),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_563),
.B(n_196),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_579),
.B(n_514),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_557),
.B(n_493),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_628),
.Y(n_726)
);

OAI21xp5_ASAP7_75t_L g727 ( 
.A1(n_642),
.A2(n_493),
.B(n_340),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_678),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_559),
.B(n_474),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_577),
.B(n_522),
.Y(n_730)
);

HB1xp67_ASAP7_75t_L g731 ( 
.A(n_591),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_648),
.B(n_522),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_648),
.B(n_608),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_691),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_591),
.B(n_197),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_623),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_594),
.B(n_474),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_628),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_SL g739 ( 
.A1(n_647),
.A2(n_663),
.B1(n_673),
.B2(n_570),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_634),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_634),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_624),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_629),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_691),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_676),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_552),
.B(n_480),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_640),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_640),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_591),
.B(n_197),
.Y(n_749)
);

INVx5_ASAP7_75t_L g750 ( 
.A(n_637),
.Y(n_750)
);

NOR3xp33_ASAP7_75t_L g751 ( 
.A(n_609),
.B(n_530),
.C(n_459),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_554),
.B(n_480),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_562),
.B(n_480),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_566),
.B(n_480),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_633),
.B(n_330),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_649),
.Y(n_756)
);

OAI22xp33_ASAP7_75t_L g757 ( 
.A1(n_591),
.A2(n_201),
.B1(n_219),
.B2(n_365),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_580),
.B(n_202),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_589),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_674),
.B(n_501),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_589),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_643),
.B(n_202),
.Y(n_762)
);

OAI22xp33_ASAP7_75t_L g763 ( 
.A1(n_586),
.A2(n_220),
.B1(n_365),
.B2(n_356),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_674),
.B(n_501),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_675),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_633),
.B(n_337),
.Y(n_766)
);

AOI221xp5_ASAP7_75t_L g767 ( 
.A1(n_619),
.A2(n_222),
.B1(n_220),
.B2(n_352),
.C(n_356),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_617),
.B(n_530),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_675),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_681),
.Y(n_770)
);

O2A1O1Ixp33_ASAP7_75t_L g771 ( 
.A1(n_651),
.A2(n_538),
.B(n_532),
.C(n_515),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_661),
.B(n_203),
.Y(n_772)
);

INVxp33_ASAP7_75t_L g773 ( 
.A(n_588),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_L g774 ( 
.A1(n_601),
.A2(n_224),
.B1(n_205),
.B2(n_366),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_681),
.B(n_410),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_619),
.A2(n_222),
.B1(n_352),
.B2(n_305),
.Y(n_776)
);

BUFx6f_ASAP7_75t_SL g777 ( 
.A(n_607),
.Y(n_777)
);

AND2x4_ASAP7_75t_SL g778 ( 
.A(n_607),
.B(n_185),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_686),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_633),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_596),
.Y(n_781)
);

NOR3xp33_ASAP7_75t_L g782 ( 
.A(n_590),
.B(n_460),
.C(n_411),
.Y(n_782)
);

NAND2xp33_ASAP7_75t_L g783 ( 
.A(n_601),
.B(n_338),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_601),
.A2(n_218),
.B1(n_205),
.B2(n_366),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_671),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_555),
.A2(n_368),
.B1(n_218),
.B2(n_364),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_596),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_601),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_636),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_692),
.B(n_203),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_686),
.B(n_501),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_605),
.B(n_501),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_597),
.Y(n_793)
);

OR2x6_ASAP7_75t_L g794 ( 
.A(n_595),
.B(n_410),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_555),
.A2(n_215),
.B1(n_364),
.B2(n_363),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_671),
.B(n_207),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_685),
.B(n_411),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_671),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_593),
.B(n_212),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_619),
.A2(n_651),
.B1(n_683),
.B2(n_637),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_671),
.B(n_212),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_690),
.B(n_213),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_621),
.B(n_412),
.Y(n_803)
);

NOR2xp67_ASAP7_75t_L g804 ( 
.A(n_611),
.B(n_511),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_605),
.B(n_669),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_605),
.B(n_682),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_597),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_635),
.B(n_213),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_605),
.B(n_510),
.Y(n_809)
);

OR2x2_ASAP7_75t_L g810 ( 
.A(n_688),
.B(n_412),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_650),
.B(n_214),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_689),
.B(n_510),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_639),
.B(n_508),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_564),
.B(n_560),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_544),
.B(n_185),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_604),
.B(n_305),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_639),
.B(n_508),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_652),
.Y(n_818)
);

CKINVDCx20_ASAP7_75t_R g819 ( 
.A(n_570),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_644),
.B(n_508),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_644),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_653),
.B(n_508),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_541),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_653),
.Y(n_824)
);

AO221x1_ASAP7_75t_L g825 ( 
.A1(n_619),
.A2(n_430),
.B1(n_417),
.B2(n_421),
.C(n_423),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_655),
.B(n_538),
.Y(n_826)
);

INVx8_ASAP7_75t_L g827 ( 
.A(n_560),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_655),
.A2(n_538),
.B(n_532),
.C(n_515),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_611),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_658),
.B(n_511),
.Y(n_830)
);

OAI22xp33_ASAP7_75t_L g831 ( 
.A1(n_612),
.A2(n_316),
.B1(n_249),
.B2(n_260),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_683),
.A2(n_637),
.B1(n_564),
.B2(n_679),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_690),
.B(n_214),
.Y(n_833)
);

OAI221xp5_ASAP7_75t_L g834 ( 
.A1(n_654),
.A2(n_532),
.B1(n_515),
.B2(n_511),
.C(n_432),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_560),
.B(n_215),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_690),
.B(n_224),
.Y(n_836)
);

INVxp67_ASAP7_75t_L g837 ( 
.A(n_656),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_690),
.B(n_277),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_658),
.B(n_502),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_662),
.B(n_502),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_662),
.B(n_504),
.Y(n_841)
);

AND2x6_ASAP7_75t_SL g842 ( 
.A(n_638),
.B(n_435),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_664),
.B(n_277),
.Y(n_843)
);

NOR2xp67_ASAP7_75t_L g844 ( 
.A(n_612),
.B(n_343),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_690),
.B(n_343),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_665),
.B(n_344),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_665),
.B(n_677),
.Y(n_847)
);

NAND2xp33_ASAP7_75t_L g848 ( 
.A(n_637),
.B(n_344),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_684),
.B(n_305),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_679),
.B(n_349),
.Y(n_850)
);

NAND2xp33_ASAP7_75t_L g851 ( 
.A(n_637),
.B(n_349),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_687),
.B(n_359),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_569),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_687),
.B(n_359),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_541),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_543),
.B(n_360),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_545),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_592),
.B(n_360),
.Y(n_858)
);

NAND2x1p5_ASAP7_75t_L g859 ( 
.A(n_584),
.B(n_417),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_545),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_546),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_719),
.B(n_547),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_703),
.Y(n_863)
);

NAND3xp33_ASAP7_75t_SL g864 ( 
.A(n_762),
.B(n_672),
.C(n_363),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_821),
.Y(n_865)
);

INVx5_ASAP7_75t_L g866 ( 
.A(n_788),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_R g867 ( 
.A(n_819),
.B(n_672),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_710),
.B(n_592),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_756),
.B(n_758),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_694),
.A2(n_637),
.B1(n_592),
.B2(n_630),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_758),
.B(n_548),
.Y(n_871)
);

NOR3xp33_ASAP7_75t_SL g872 ( 
.A(n_757),
.B(n_309),
.C(n_235),
.Y(n_872)
);

NAND2x1p5_ASAP7_75t_L g873 ( 
.A(n_788),
.B(n_584),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_712),
.B(n_630),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_824),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_765),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_768),
.B(n_630),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_728),
.B(n_421),
.Y(n_878)
);

INVx8_ASAP7_75t_L g879 ( 
.A(n_827),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_769),
.Y(n_880)
);

INVx4_ASAP7_75t_L g881 ( 
.A(n_788),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_770),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_759),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_709),
.B(n_361),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_788),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_700),
.B(n_548),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_700),
.B(n_549),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_794),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_794),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_734),
.Y(n_890)
);

AND3x1_ASAP7_75t_L g891 ( 
.A(n_767),
.B(n_423),
.C(n_426),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_694),
.A2(n_326),
.B1(n_546),
.B2(n_565),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_761),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_803),
.B(n_549),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_853),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_837),
.B(n_551),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_779),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_825),
.A2(n_326),
.B1(n_565),
.B2(n_568),
.Y(n_898)
);

BUFx8_ASAP7_75t_L g899 ( 
.A(n_777),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_781),
.Y(n_900)
);

BUFx4f_ASAP7_75t_L g901 ( 
.A(n_827),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_847),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_698),
.Y(n_903)
);

NAND2xp33_ASAP7_75t_SL g904 ( 
.A(n_773),
.B(n_731),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_750),
.B(n_551),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_717),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_742),
.Y(n_907)
);

INVx5_ASAP7_75t_L g908 ( 
.A(n_853),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_733),
.A2(n_585),
.B1(n_567),
.B2(n_576),
.Y(n_909)
);

AND2x6_ASAP7_75t_SL g910 ( 
.A(n_762),
.B(n_426),
.Y(n_910)
);

NOR2xp67_ASAP7_75t_L g911 ( 
.A(n_829),
.B(n_567),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_711),
.B(n_326),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_743),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_745),
.Y(n_914)
);

INVx3_ASAP7_75t_SL g915 ( 
.A(n_827),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_787),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_839),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_840),
.Y(n_918)
);

INVx5_ASAP7_75t_L g919 ( 
.A(n_853),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_731),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_794),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_698),
.Y(n_922)
);

INVxp67_ASAP7_75t_L g923 ( 
.A(n_730),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_708),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_695),
.A2(n_571),
.B1(n_568),
.B2(n_572),
.Y(n_925)
);

INVxp67_ASAP7_75t_L g926 ( 
.A(n_704),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_793),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_841),
.Y(n_928)
);

INVx6_ASAP7_75t_L g929 ( 
.A(n_708),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_803),
.B(n_576),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_744),
.B(n_747),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_808),
.B(n_569),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_777),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_716),
.A2(n_620),
.B(n_581),
.Y(n_934)
);

INVx5_ASAP7_75t_L g935 ( 
.A(n_853),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_732),
.B(n_581),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_780),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_711),
.B(n_582),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_807),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_808),
.A2(n_620),
.B1(n_582),
.B2(n_585),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_811),
.B(n_646),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_804),
.B(n_569),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_748),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_780),
.B(n_569),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_811),
.B(n_646),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_696),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_704),
.B(n_659),
.Y(n_947)
);

O2A1O1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_834),
.A2(n_571),
.B(n_572),
.C(n_574),
.Y(n_948)
);

OAI22xp33_ASAP7_75t_L g949 ( 
.A1(n_797),
.A2(n_269),
.B1(n_270),
.B2(n_272),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_736),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_714),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_718),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_785),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_723),
.B(n_659),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_721),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_726),
.Y(n_956)
);

NAND2xp33_ASAP7_75t_SL g957 ( 
.A(n_849),
.B(n_276),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_738),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_823),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_785),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_855),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_L g962 ( 
.A1(n_800),
.A2(n_578),
.B1(n_574),
.B2(n_290),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_857),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_775),
.B(n_740),
.Y(n_964)
);

BUFx8_ASAP7_75t_L g965 ( 
.A(n_789),
.Y(n_965)
);

INVx5_ASAP7_75t_L g966 ( 
.A(n_750),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_842),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_778),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_741),
.Y(n_969)
);

NOR2x2_ASAP7_75t_L g970 ( 
.A(n_699),
.B(n_598),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_818),
.Y(n_971)
);

INVx5_ASAP7_75t_L g972 ( 
.A(n_750),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_860),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_723),
.B(n_540),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_706),
.A2(n_578),
.B(n_428),
.C(n_598),
.Y(n_975)
);

OR2x6_ASAP7_75t_L g976 ( 
.A(n_739),
.B(n_584),
.Y(n_976)
);

HB1xp67_ASAP7_75t_L g977 ( 
.A(n_702),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_705),
.B(n_540),
.Y(n_978)
);

AOI22xp33_ASAP7_75t_L g979 ( 
.A1(n_800),
.A2(n_285),
.B1(n_287),
.B2(n_294),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_701),
.A2(n_599),
.B(n_602),
.C(n_606),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_705),
.B(n_540),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_701),
.B(n_603),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_724),
.B(n_304),
.Y(n_983)
);

NOR3xp33_ASAP7_75t_SL g984 ( 
.A(n_757),
.B(n_310),
.C(n_314),
.Y(n_984)
);

NOR3xp33_ASAP7_75t_SL g985 ( 
.A(n_831),
.B(n_322),
.C(n_327),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_776),
.A2(n_329),
.B1(n_341),
.B2(n_342),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_775),
.B(n_575),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_722),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_812),
.B(n_575),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_727),
.B(n_575),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_861),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_805),
.B(n_583),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_755),
.A2(n_613),
.B1(n_599),
.B2(n_602),
.Y(n_993)
);

AND2x6_ASAP7_75t_L g994 ( 
.A(n_814),
.B(n_606),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_SL g995 ( 
.A1(n_771),
.A2(n_610),
.B(n_613),
.C(n_616),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_798),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_815),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_725),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_798),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_826),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_735),
.B(n_569),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_806),
.B(n_668),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_832),
.A2(n_610),
.B1(n_666),
.B2(n_616),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_830),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_832),
.A2(n_668),
.B1(n_666),
.B2(n_583),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_735),
.B(n_587),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_810),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_697),
.B(n_668),
.Y(n_1008)
);

OR2x2_ASAP7_75t_L g1009 ( 
.A(n_697),
.B(n_4),
.Y(n_1009)
);

INVxp67_ASAP7_75t_L g1010 ( 
.A(n_706),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_707),
.B(n_666),
.Y(n_1011)
);

NOR2x1p5_ASAP7_75t_L g1012 ( 
.A(n_816),
.B(n_843),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_760),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_750),
.Y(n_1014)
);

AND2x6_ASAP7_75t_SL g1015 ( 
.A(n_749),
.B(n_6),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_835),
.Y(n_1016)
);

AOI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_776),
.A2(n_625),
.B1(n_645),
.B2(n_641),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_713),
.Y(n_1018)
);

OR2x2_ASAP7_75t_L g1019 ( 
.A(n_707),
.B(n_772),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_749),
.B(n_573),
.Y(n_1020)
);

AO22x1_ASAP7_75t_L g1021 ( 
.A1(n_835),
.A2(n_583),
.B1(n_616),
.B2(n_625),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_729),
.Y(n_1022)
);

NAND3xp33_ASAP7_75t_SL g1023 ( 
.A(n_782),
.B(n_603),
.C(n_632),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_790),
.B(n_626),
.Y(n_1024)
);

BUFx3_ASAP7_75t_L g1025 ( 
.A(n_858),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_790),
.B(n_632),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_764),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_791),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_713),
.B(n_626),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_751),
.B(n_573),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_715),
.B(n_626),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_831),
.B(n_587),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_844),
.B(n_632),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_737),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_699),
.A2(n_625),
.B1(n_645),
.B2(n_641),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_715),
.B(n_645),
.Y(n_1036)
);

NAND2x1p5_ASAP7_75t_L g1037 ( 
.A(n_755),
.B(n_603),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_846),
.B(n_641),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_858),
.B(n_631),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_813),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_SL g1041 ( 
.A1(n_699),
.A2(n_11),
.B1(n_13),
.B2(n_16),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_814),
.B(n_600),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_R g1043 ( 
.A(n_783),
.B(n_78),
.Y(n_1043)
);

INVx3_ASAP7_75t_SL g1044 ( 
.A(n_799),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_850),
.B(n_631),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_763),
.B(n_600),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_856),
.B(n_631),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_852),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_859),
.Y(n_1049)
);

AND2x6_ASAP7_75t_SL g1050 ( 
.A(n_854),
.B(n_13),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_763),
.B(n_600),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_856),
.B(n_600),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_859),
.B(n_600),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_766),
.B(n_587),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_876),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_983),
.B(n_795),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_926),
.A2(n_766),
.B(n_802),
.C(n_796),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_926),
.B(n_774),
.Y(n_1058)
);

BUFx8_ASAP7_75t_SL g1059 ( 
.A(n_933),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_977),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_966),
.A2(n_720),
.B(n_792),
.Y(n_1061)
);

NAND2x1_ASAP7_75t_L g1062 ( 
.A(n_881),
.B(n_885),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_966),
.A2(n_809),
.B(n_693),
.Y(n_1063)
);

O2A1O1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_864),
.A2(n_833),
.B(n_801),
.C(n_845),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_961),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_998),
.B(n_802),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_966),
.A2(n_746),
.B(n_752),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_963),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_966),
.A2(n_754),
.B(n_753),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_988),
.B(n_796),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_877),
.B(n_784),
.Y(n_1071)
);

OAI22x1_ASAP7_75t_L g1072 ( 
.A1(n_1012),
.A2(n_786),
.B1(n_801),
.B2(n_833),
.Y(n_1072)
);

CKINVDCx6p67_ASAP7_75t_R g1073 ( 
.A(n_915),
.Y(n_1073)
);

OAI22x1_ASAP7_75t_L g1074 ( 
.A1(n_888),
.A2(n_836),
.B1(n_838),
.B2(n_845),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_880),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_SL g1076 ( 
.A(n_901),
.B(n_828),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_863),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_923),
.B(n_838),
.Y(n_1078)
);

NAND2x1p5_ASAP7_75t_L g1079 ( 
.A(n_866),
.B(n_836),
.Y(n_1079)
);

HB1xp67_ASAP7_75t_L g1080 ( 
.A(n_977),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_917),
.B(n_822),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_918),
.B(n_820),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_1007),
.B(n_817),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_979),
.A2(n_587),
.B1(n_660),
.B2(n_848),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_979),
.A2(n_864),
.B1(n_1018),
.B2(n_912),
.Y(n_1085)
);

CKINVDCx11_ASAP7_75t_R g1086 ( 
.A(n_915),
.Y(n_1086)
);

AOI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_877),
.A2(n_851),
.B1(n_587),
.B2(n_660),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_962),
.A2(n_660),
.B1(n_21),
.B2(n_24),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_928),
.B(n_660),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_962),
.A2(n_660),
.B1(n_25),
.B2(n_26),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_920),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_1018),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_1092)
);

INVx4_ASAP7_75t_L g1093 ( 
.A(n_866),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_923),
.B(n_27),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_971),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1007),
.B(n_28),
.Y(n_1096)
);

OAI22x1_ASAP7_75t_L g1097 ( 
.A1(n_889),
.A2(n_31),
.B1(n_32),
.B2(n_38),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_885),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_973),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_972),
.A2(n_96),
.B(n_177),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_885),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_1016),
.B(n_32),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_R g1103 ( 
.A(n_968),
.B(n_90),
.Y(n_1103)
);

NAND2x1p5_ASAP7_75t_L g1104 ( 
.A(n_866),
.B(n_98),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_885),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_924),
.B(n_868),
.Y(n_1106)
);

AOI21xp33_ASAP7_75t_L g1107 ( 
.A1(n_1019),
.A2(n_38),
.B(n_39),
.Y(n_1107)
);

BUFx12f_ASAP7_75t_L g1108 ( 
.A(n_899),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_R g1109 ( 
.A(n_904),
.B(n_100),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_1025),
.B(n_40),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_972),
.A2(n_919),
.B(n_908),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_882),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_991),
.Y(n_1113)
);

INVx2_ASAP7_75t_SL g1114 ( 
.A(n_890),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_972),
.A2(n_101),
.B(n_170),
.Y(n_1115)
);

INVx1_ASAP7_75t_SL g1116 ( 
.A(n_890),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_875),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_972),
.A2(n_85),
.B(n_167),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_897),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_907),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_902),
.B(n_42),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_883),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_924),
.B(n_76),
.Y(n_1123)
);

NOR2x1_ASAP7_75t_L g1124 ( 
.A(n_881),
.B(n_124),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_964),
.B(n_74),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_913),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_893),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_914),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_895),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_868),
.B(n_131),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_934),
.A2(n_1003),
.B(n_1005),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_1048),
.B(n_65),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_938),
.B(n_42),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_870),
.A2(n_44),
.B1(n_45),
.B2(n_49),
.Y(n_1134)
);

AOI21x1_ASAP7_75t_L g1135 ( 
.A1(n_1021),
.A2(n_145),
.B(n_161),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_938),
.B(n_50),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_908),
.A2(n_143),
.B(n_155),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_1010),
.A2(n_52),
.B(n_53),
.C(n_58),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_874),
.B(n_140),
.Y(n_1139)
);

AOI21x1_ASAP7_75t_L g1140 ( 
.A1(n_932),
.A2(n_146),
.B(n_152),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_908),
.A2(n_179),
.B(n_53),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_931),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_870),
.A2(n_1010),
.B1(n_1035),
.B2(n_892),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_874),
.B(n_964),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_903),
.B(n_922),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_982),
.B(n_1004),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_SL g1147 ( 
.A1(n_1041),
.A2(n_967),
.B1(n_986),
.B2(n_976),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_903),
.B(n_922),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1035),
.A2(n_892),
.B1(n_1009),
.B2(n_886),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_878),
.B(n_997),
.Y(n_1150)
);

OA22x2_ASAP7_75t_L g1151 ( 
.A1(n_921),
.A2(n_862),
.B1(n_976),
.B2(n_1044),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_937),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_908),
.A2(n_919),
.B(n_935),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_957),
.A2(n_929),
.B1(n_931),
.B2(n_896),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_982),
.B(n_896),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_887),
.A2(n_986),
.B1(n_872),
.B2(n_984),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_872),
.A2(n_984),
.B1(n_936),
.B2(n_976),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_934),
.A2(n_873),
.B(n_948),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_1046),
.A2(n_1051),
.B(n_884),
.C(n_949),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_900),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_919),
.A2(n_935),
.B(n_992),
.Y(n_1161)
);

AO32x1_ASAP7_75t_L g1162 ( 
.A1(n_1020),
.A2(n_1030),
.A3(n_1039),
.B1(n_1047),
.B2(n_865),
.Y(n_1162)
);

INVx3_ASAP7_75t_L g1163 ( 
.A(n_937),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_943),
.Y(n_1164)
);

BUFx3_ASAP7_75t_L g1165 ( 
.A(n_879),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_919),
.A2(n_935),
.B(n_1002),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_911),
.B(n_937),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1044),
.B(n_891),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_954),
.A2(n_871),
.B1(n_898),
.B2(n_930),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_895),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_898),
.A2(n_894),
.B1(n_947),
.B2(n_985),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1000),
.B(n_1013),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_985),
.A2(n_941),
.B1(n_945),
.B2(n_1028),
.Y(n_1173)
);

NOR3xp33_ASAP7_75t_SL g1174 ( 
.A(n_949),
.B(n_950),
.C(n_969),
.Y(n_1174)
);

AOI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1042),
.A2(n_981),
.B(n_978),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_916),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_927),
.Y(n_1177)
);

O2A1O1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1032),
.A2(n_1006),
.B(n_1001),
.C(n_906),
.Y(n_1178)
);

AOI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_929),
.A2(n_1026),
.B1(n_994),
.B2(n_1054),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_939),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_946),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_873),
.A2(n_948),
.B(n_925),
.Y(n_1182)
);

AOI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_929),
.A2(n_1026),
.B1(n_994),
.B2(n_987),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_937),
.B(n_935),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_925),
.A2(n_993),
.B(n_1024),
.Y(n_1185)
);

INVx5_ASAP7_75t_L g1186 ( 
.A(n_1014),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_951),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_990),
.A2(n_1053),
.B(n_989),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1027),
.B(n_1034),
.Y(n_1189)
);

BUFx5_ASAP7_75t_L g1190 ( 
.A(n_994),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_909),
.A2(n_1017),
.B1(n_1049),
.B2(n_1022),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_952),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1017),
.A2(n_1049),
.B1(n_974),
.B2(n_940),
.Y(n_1193)
);

AOI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_994),
.A2(n_1052),
.B1(n_1033),
.B2(n_862),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_955),
.Y(n_1195)
);

BUFx4f_ASAP7_75t_L g1196 ( 
.A(n_879),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1040),
.B(n_994),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1049),
.A2(n_1052),
.B1(n_1037),
.B2(n_895),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1049),
.B(n_901),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_956),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1037),
.A2(n_895),
.B1(n_980),
.B2(n_1008),
.Y(n_1201)
);

AO32x2_ASAP7_75t_L g1202 ( 
.A1(n_970),
.A2(n_995),
.A3(n_910),
.B1(n_975),
.B2(n_1043),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1011),
.A2(n_996),
.B1(n_960),
.B2(n_953),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1033),
.B(n_867),
.Y(n_1204)
);

AOI21xp33_ASAP7_75t_SL g1205 ( 
.A1(n_879),
.A2(n_1015),
.B(n_1050),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_867),
.B(n_1043),
.Y(n_1206)
);

O2A1O1Ixp5_ASAP7_75t_SL g1207 ( 
.A1(n_944),
.A2(n_942),
.B(n_960),
.C(n_996),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_958),
.B(n_959),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_SL g1209 ( 
.A(n_1014),
.B(n_953),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_999),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_899),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1029),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1038),
.A2(n_1045),
.B1(n_1036),
.B2(n_1031),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_1014),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_975),
.Y(n_1215)
);

O2A1O1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_995),
.A2(n_1023),
.B(n_905),
.C(n_965),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1014),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1188),
.A2(n_905),
.B(n_1023),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1146),
.A2(n_965),
.B(n_1067),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1155),
.B(n_1172),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1131),
.A2(n_1159),
.B(n_1173),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1158),
.A2(n_1182),
.B(n_1061),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1064),
.A2(n_1057),
.B(n_1174),
.C(n_1078),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1120),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1091),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1069),
.A2(n_1193),
.B(n_1084),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_1077),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1126),
.Y(n_1228)
);

NOR2x1_ASAP7_75t_L g1229 ( 
.A(n_1206),
.B(n_1093),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1128),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1058),
.B(n_1060),
.Y(n_1231)
);

AO21x2_ASAP7_75t_L g1232 ( 
.A1(n_1201),
.A2(n_1175),
.B(n_1198),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1185),
.A2(n_1201),
.B(n_1203),
.Y(n_1233)
);

AO31x2_ASAP7_75t_L g1234 ( 
.A1(n_1193),
.A2(n_1074),
.A3(n_1169),
.B(n_1173),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_1098),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1189),
.B(n_1083),
.Y(n_1236)
);

OAI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1154),
.A2(n_1151),
.B1(n_1156),
.B2(n_1090),
.Y(n_1237)
);

INVxp67_ASAP7_75t_SL g1238 ( 
.A(n_1080),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1056),
.B(n_1066),
.Y(n_1239)
);

AOI221x1_ASAP7_75t_L g1240 ( 
.A1(n_1156),
.A2(n_1090),
.B1(n_1088),
.B2(n_1171),
.C(n_1072),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1169),
.A2(n_1171),
.A3(n_1213),
.B(n_1198),
.Y(n_1241)
);

NAND3xp33_ASAP7_75t_SL g1242 ( 
.A(n_1085),
.B(n_1071),
.C(n_1102),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1063),
.A2(n_1178),
.B(n_1191),
.Y(n_1243)
);

NAND2x1_ASAP7_75t_L g1244 ( 
.A(n_1093),
.B(n_1214),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1055),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1203),
.A2(n_1207),
.B(n_1161),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1070),
.B(n_1081),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1075),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1082),
.B(n_1149),
.Y(n_1249)
);

OA22x2_ASAP7_75t_L g1250 ( 
.A1(n_1147),
.A2(n_1097),
.B1(n_1134),
.B2(n_1088),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1150),
.B(n_1096),
.Y(n_1251)
);

AO31x2_ASAP7_75t_L g1252 ( 
.A1(n_1191),
.A2(n_1215),
.A3(n_1149),
.B(n_1143),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1112),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1157),
.A2(n_1134),
.B1(n_1143),
.B2(n_1168),
.Y(n_1254)
);

AO21x2_ASAP7_75t_L g1255 ( 
.A1(n_1179),
.A2(n_1135),
.B(n_1183),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1197),
.A2(n_1166),
.B(n_1106),
.Y(n_1256)
);

BUFx10_ASAP7_75t_L g1257 ( 
.A(n_1110),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1153),
.A2(n_1089),
.B(n_1111),
.Y(n_1258)
);

A2O1A1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1216),
.A2(n_1157),
.B(n_1194),
.C(n_1094),
.Y(n_1259)
);

A2O1A1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1121),
.A2(n_1107),
.B(n_1130),
.C(n_1138),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1212),
.A2(n_1087),
.B(n_1139),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1140),
.A2(n_1076),
.B(n_1141),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1186),
.A2(n_1144),
.B(n_1167),
.Y(n_1263)
);

OA21x2_ASAP7_75t_L g1264 ( 
.A1(n_1123),
.A2(n_1132),
.B(n_1137),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_R g1265 ( 
.A(n_1086),
.B(n_1196),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1119),
.B(n_1164),
.Y(n_1266)
);

INVxp67_ASAP7_75t_L g1267 ( 
.A(n_1116),
.Y(n_1267)
);

AO31x2_ASAP7_75t_L g1268 ( 
.A1(n_1162),
.A2(n_1210),
.A3(n_1099),
.B(n_1065),
.Y(n_1268)
);

OR2x6_ASAP7_75t_L g1269 ( 
.A(n_1204),
.B(n_1125),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_1098),
.Y(n_1270)
);

INVx1_ASAP7_75t_SL g1271 ( 
.A(n_1116),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1142),
.B(n_1117),
.Y(n_1272)
);

NAND2x1p5_ASAP7_75t_L g1273 ( 
.A(n_1196),
.B(n_1186),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1186),
.A2(n_1076),
.B(n_1162),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_1114),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1068),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1151),
.B(n_1095),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1113),
.B(n_1208),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1176),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1079),
.A2(n_1209),
.B(n_1104),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1079),
.A2(n_1104),
.B(n_1062),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1125),
.B(n_1208),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1098),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1165),
.B(n_1199),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1187),
.B(n_1200),
.Y(n_1285)
);

BUFx12f_ASAP7_75t_L g1286 ( 
.A(n_1108),
.Y(n_1286)
);

BUFx12f_ASAP7_75t_L g1287 ( 
.A(n_1211),
.Y(n_1287)
);

NOR2x1_ASAP7_75t_SL g1288 ( 
.A(n_1186),
.B(n_1101),
.Y(n_1288)
);

NAND3xp33_ASAP7_75t_L g1289 ( 
.A(n_1092),
.B(n_1177),
.C(n_1122),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1162),
.A2(n_1184),
.B(n_1148),
.Y(n_1290)
);

AO22x1_ASAP7_75t_L g1291 ( 
.A1(n_1124),
.A2(n_1180),
.B1(n_1195),
.B2(n_1192),
.Y(n_1291)
);

AO31x2_ASAP7_75t_L g1292 ( 
.A1(n_1100),
.A2(n_1118),
.A3(n_1115),
.B(n_1127),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1160),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1145),
.A2(n_1152),
.B(n_1163),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1152),
.A2(n_1163),
.B(n_1181),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1190),
.B(n_1217),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1214),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1103),
.B(n_1205),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1073),
.B(n_1059),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_SL g1300 ( 
.A(n_1109),
.B(n_1190),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1129),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1170),
.A2(n_1105),
.B(n_1190),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_1105),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1202),
.A2(n_1156),
.B1(n_762),
.B2(n_864),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1155),
.B(n_926),
.Y(n_1305)
);

BUFx2_ASAP7_75t_L g1306 ( 
.A(n_1091),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1155),
.A2(n_979),
.B1(n_962),
.B2(n_1146),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1158),
.A2(n_1182),
.B(n_934),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1120),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1155),
.B(n_926),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1158),
.A2(n_1182),
.B(n_934),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1188),
.A2(n_972),
.B(n_966),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_SL g1313 ( 
.A(n_1088),
.B(n_1090),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_1165),
.B(n_1125),
.Y(n_1314)
);

CKINVDCx12_ASAP7_75t_R g1315 ( 
.A(n_1150),
.Y(n_1315)
);

AO21x2_ASAP7_75t_L g1316 ( 
.A1(n_1131),
.A2(n_1201),
.B(n_1188),
.Y(n_1316)
);

NOR2x1_ASAP7_75t_SL g1317 ( 
.A(n_1093),
.B(n_866),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1120),
.Y(n_1318)
);

AO31x2_ASAP7_75t_L g1319 ( 
.A1(n_1201),
.A2(n_1193),
.A3(n_1074),
.B(n_1169),
.Y(n_1319)
);

AOI21xp33_ASAP7_75t_L g1320 ( 
.A1(n_1159),
.A2(n_1155),
.B(n_1156),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1186),
.Y(n_1321)
);

A2O1A1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1159),
.A2(n_1064),
.B(n_1057),
.C(n_1174),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1158),
.A2(n_1182),
.B(n_934),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1120),
.Y(n_1324)
);

AO22x2_ASAP7_75t_L g1325 ( 
.A1(n_1088),
.A2(n_1090),
.B1(n_1134),
.B2(n_1156),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1056),
.B(n_712),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1155),
.B(n_1146),
.Y(n_1327)
);

O2A1O1Ixp33_ASAP7_75t_L g1328 ( 
.A1(n_1156),
.A2(n_926),
.B(n_1071),
.C(n_553),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1059),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1155),
.B(n_1146),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1158),
.A2(n_1182),
.B(n_934),
.Y(n_1331)
);

NAND3x1_ASAP7_75t_L g1332 ( 
.A(n_1168),
.B(n_673),
.C(n_762),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1155),
.B(n_1146),
.Y(n_1333)
);

INVx2_ASAP7_75t_SL g1334 ( 
.A(n_1077),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1116),
.B(n_869),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1155),
.B(n_1146),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1120),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_1098),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1165),
.B(n_1125),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1158),
.A2(n_1182),
.B(n_934),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1158),
.A2(n_1182),
.B(n_934),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1155),
.B(n_926),
.Y(n_1342)
);

AND2x4_ASAP7_75t_L g1343 ( 
.A(n_1165),
.B(n_1125),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1120),
.Y(n_1344)
);

OAI22x1_ASAP7_75t_L g1345 ( 
.A1(n_1154),
.A2(n_1058),
.B1(n_1168),
.B2(n_1194),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1120),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1056),
.B(n_712),
.Y(n_1347)
);

AO31x2_ASAP7_75t_L g1348 ( 
.A1(n_1201),
.A2(n_1193),
.A3(n_1074),
.B(n_1169),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_SL g1349 ( 
.A1(n_1193),
.A2(n_788),
.B(n_1084),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_1059),
.Y(n_1350)
);

AO21x2_ASAP7_75t_L g1351 ( 
.A1(n_1131),
.A2(n_1201),
.B(n_1188),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1091),
.Y(n_1352)
);

INVx4_ASAP7_75t_L g1353 ( 
.A(n_1186),
.Y(n_1353)
);

INVxp67_ASAP7_75t_SL g1354 ( 
.A(n_1080),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1060),
.Y(n_1355)
);

INVxp67_ASAP7_75t_L g1356 ( 
.A(n_1080),
.Y(n_1356)
);

INVx1_ASAP7_75t_SL g1357 ( 
.A(n_1116),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1155),
.B(n_926),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_SL g1359 ( 
.A(n_1116),
.B(n_869),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1155),
.A2(n_979),
.B1(n_962),
.B2(n_1146),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1155),
.B(n_926),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1188),
.A2(n_972),
.B(n_966),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1155),
.B(n_926),
.Y(n_1363)
);

AO32x2_ASAP7_75t_L g1364 ( 
.A1(n_1088),
.A2(n_1090),
.A3(n_1156),
.B1(n_1171),
.B2(n_1173),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_SL g1365 ( 
.A1(n_1193),
.A2(n_788),
.B(n_1084),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1188),
.A2(n_972),
.B(n_966),
.Y(n_1366)
);

O2A1O1Ixp33_ASAP7_75t_SL g1367 ( 
.A1(n_1155),
.A2(n_1133),
.B(n_1136),
.C(n_1146),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1155),
.B(n_926),
.Y(n_1368)
);

BUFx12f_ASAP7_75t_L g1369 ( 
.A(n_1086),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_1116),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1165),
.B(n_1125),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_SL g1372 ( 
.A1(n_1193),
.A2(n_788),
.B(n_1084),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1120),
.Y(n_1373)
);

NAND3xp33_ASAP7_75t_SL g1374 ( 
.A(n_1085),
.B(n_588),
.C(n_553),
.Y(n_1374)
);

OAI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1131),
.A2(n_1188),
.B(n_1155),
.Y(n_1375)
);

NAND2xp33_ASAP7_75t_R g1376 ( 
.A(n_1269),
.B(n_1264),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1266),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1344),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1269),
.B(n_1282),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1308),
.A2(n_1323),
.B(n_1311),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_1329),
.Y(n_1381)
);

BUFx6f_ASAP7_75t_L g1382 ( 
.A(n_1235),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1346),
.Y(n_1383)
);

AND2x2_ASAP7_75t_SL g1384 ( 
.A(n_1313),
.B(n_1304),
.Y(n_1384)
);

INVxp67_ASAP7_75t_SL g1385 ( 
.A(n_1249),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_SL g1386 ( 
.A1(n_1219),
.A2(n_1261),
.B(n_1328),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1224),
.Y(n_1387)
);

AOI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1291),
.A2(n_1274),
.B(n_1258),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1228),
.Y(n_1389)
);

NOR2x1_ASAP7_75t_SL g1390 ( 
.A(n_1300),
.B(n_1269),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1239),
.B(n_1236),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1331),
.A2(n_1341),
.B(n_1340),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1319),
.Y(n_1393)
);

INVxp67_ASAP7_75t_SL g1394 ( 
.A(n_1327),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1230),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1245),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1242),
.B(n_1326),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1220),
.B(n_1305),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1222),
.A2(n_1256),
.B(n_1312),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1327),
.A2(n_1333),
.B1(n_1336),
.B2(n_1330),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1310),
.B(n_1342),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1314),
.B(n_1339),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1347),
.B(n_1251),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1225),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1248),
.Y(n_1405)
);

OA21x2_ASAP7_75t_L g1406 ( 
.A1(n_1221),
.A2(n_1240),
.B(n_1226),
.Y(n_1406)
);

NAND3xp33_ASAP7_75t_L g1407 ( 
.A(n_1223),
.B(n_1322),
.C(n_1260),
.Y(n_1407)
);

CKINVDCx9p33_ASAP7_75t_R g1408 ( 
.A(n_1299),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1313),
.A2(n_1250),
.B1(n_1325),
.B2(n_1374),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1253),
.Y(n_1410)
);

OA21x2_ASAP7_75t_L g1411 ( 
.A1(n_1221),
.A2(n_1243),
.B(n_1375),
.Y(n_1411)
);

INVx6_ASAP7_75t_L g1412 ( 
.A(n_1353),
.Y(n_1412)
);

CKINVDCx6p67_ASAP7_75t_R g1413 ( 
.A(n_1286),
.Y(n_1413)
);

AND2x4_ASAP7_75t_L g1414 ( 
.A(n_1314),
.B(n_1339),
.Y(n_1414)
);

NAND2x1p5_ASAP7_75t_L g1415 ( 
.A(n_1353),
.B(n_1321),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1343),
.B(n_1371),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1231),
.B(n_1358),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1309),
.Y(n_1418)
);

BUFx8_ASAP7_75t_L g1419 ( 
.A(n_1369),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_SL g1420 ( 
.A1(n_1315),
.A2(n_1332),
.B1(n_1254),
.B2(n_1277),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1318),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1325),
.A2(n_1307),
.B1(n_1360),
.B2(n_1237),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1324),
.Y(n_1423)
);

AOI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1218),
.A2(n_1366),
.B(n_1362),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1319),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1271),
.B(n_1357),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1321),
.Y(n_1427)
);

AO31x2_ASAP7_75t_L g1428 ( 
.A1(n_1290),
.A2(n_1259),
.A3(n_1307),
.B(n_1360),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1233),
.A2(n_1246),
.B(n_1262),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1337),
.Y(n_1430)
);

CKINVDCx8_ASAP7_75t_R g1431 ( 
.A(n_1350),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1262),
.A2(n_1281),
.B(n_1280),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_SL g1433 ( 
.A1(n_1261),
.A2(n_1263),
.B(n_1333),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1373),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_1227),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_SL g1436 ( 
.A(n_1287),
.B(n_1298),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1330),
.A2(n_1336),
.B1(n_1368),
.B2(n_1363),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1320),
.A2(n_1345),
.B1(n_1361),
.B2(n_1247),
.Y(n_1438)
);

OA21x2_ASAP7_75t_L g1439 ( 
.A1(n_1289),
.A2(n_1295),
.B(n_1296),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1302),
.A2(n_1294),
.B(n_1264),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1235),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1271),
.B(n_1370),
.Y(n_1442)
);

AO21x2_ASAP7_75t_L g1443 ( 
.A1(n_1316),
.A2(n_1351),
.B(n_1255),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1285),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1257),
.A2(n_1359),
.B1(n_1335),
.B2(n_1289),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1357),
.B(n_1370),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1279),
.Y(n_1447)
);

OAI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1367),
.A2(n_1278),
.B(n_1272),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1244),
.A2(n_1273),
.B(n_1297),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_SL g1450 ( 
.A1(n_1267),
.A2(n_1371),
.B1(n_1343),
.B2(n_1284),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_SL g1451 ( 
.A1(n_1317),
.A2(n_1288),
.B(n_1301),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1270),
.Y(n_1452)
);

AND2x6_ASAP7_75t_L g1453 ( 
.A(n_1284),
.B(n_1338),
.Y(n_1453)
);

OAI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1276),
.A2(n_1293),
.B(n_1356),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1355),
.B(n_1354),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1238),
.A2(n_1306),
.B1(n_1352),
.B2(n_1334),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1292),
.A2(n_1351),
.B(n_1316),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1275),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1268),
.Y(n_1459)
);

AO21x2_ASAP7_75t_L g1460 ( 
.A1(n_1255),
.A2(n_1232),
.B(n_1364),
.Y(n_1460)
);

CKINVDCx11_ASAP7_75t_R g1461 ( 
.A(n_1257),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1268),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1303),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_SL g1464 ( 
.A1(n_1364),
.A2(n_1234),
.B(n_1348),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_1265),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1292),
.A2(n_1232),
.B(n_1348),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1292),
.A2(n_1348),
.B(n_1319),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1234),
.A2(n_1252),
.B(n_1241),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1252),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1270),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1252),
.B(n_1234),
.Y(n_1471)
);

OR2x6_ASAP7_75t_L g1472 ( 
.A(n_1270),
.B(n_1283),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1241),
.B(n_1283),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1241),
.B(n_1283),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1338),
.B(n_1364),
.Y(n_1475)
);

BUFx2_ASAP7_75t_SL g1476 ( 
.A(n_1225),
.Y(n_1476)
);

NAND3xp33_ASAP7_75t_L g1477 ( 
.A(n_1328),
.B(n_553),
.C(n_985),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1308),
.A2(n_1323),
.B(n_1311),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1319),
.Y(n_1479)
);

INVx6_ASAP7_75t_L g1480 ( 
.A(n_1353),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_SL g1481 ( 
.A1(n_1219),
.A2(n_1216),
.B(n_1159),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1327),
.A2(n_1330),
.B1(n_1336),
.B2(n_1333),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1239),
.B(n_1236),
.Y(n_1483)
);

O2A1O1Ixp33_ASAP7_75t_L g1484 ( 
.A1(n_1223),
.A2(n_1242),
.B(n_1374),
.C(n_1322),
.Y(n_1484)
);

OAI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1308),
.A2(n_1323),
.B(n_1311),
.Y(n_1485)
);

AND2x4_ASAP7_75t_L g1486 ( 
.A(n_1269),
.B(n_1282),
.Y(n_1486)
);

OA21x2_ASAP7_75t_L g1487 ( 
.A1(n_1221),
.A2(n_1240),
.B(n_1226),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1308),
.A2(n_1323),
.B(n_1311),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1266),
.Y(n_1489)
);

NOR2x1_ASAP7_75t_L g1490 ( 
.A(n_1229),
.B(n_1206),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1269),
.B(n_1282),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1239),
.B(n_1326),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1308),
.A2(n_1323),
.B(n_1311),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1308),
.A2(n_1323),
.B(n_1311),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1266),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1260),
.A2(n_553),
.B(n_1223),
.Y(n_1496)
);

INVxp67_ASAP7_75t_L g1497 ( 
.A(n_1355),
.Y(n_1497)
);

BUFx2_ASAP7_75t_SL g1498 ( 
.A(n_1225),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1308),
.A2(n_1323),
.B(n_1311),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1239),
.B(n_1236),
.Y(n_1500)
);

NAND2x1p5_ASAP7_75t_L g1501 ( 
.A(n_1353),
.B(n_866),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1269),
.B(n_1282),
.Y(n_1502)
);

OR2x6_ASAP7_75t_L g1503 ( 
.A(n_1349),
.B(n_1365),
.Y(n_1503)
);

OAI211xp5_ASAP7_75t_L g1504 ( 
.A1(n_1304),
.A2(n_776),
.B(n_767),
.C(n_986),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1313),
.A2(n_1242),
.B1(n_1250),
.B2(n_1325),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_1329),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1225),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1349),
.A2(n_1372),
.B(n_1365),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1266),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1374),
.A2(n_385),
.B1(n_386),
.B2(n_384),
.Y(n_1510)
);

OAI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1308),
.A2(n_1323),
.B(n_1311),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1319),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1266),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1326),
.B(n_1347),
.Y(n_1514)
);

CKINVDCx6p67_ASAP7_75t_R g1515 ( 
.A(n_1286),
.Y(n_1515)
);

AOI221xp5_ASAP7_75t_L g1516 ( 
.A1(n_1242),
.A2(n_663),
.B1(n_1320),
.B2(n_767),
.C(n_476),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_SL g1517 ( 
.A1(n_1313),
.A2(n_1041),
.B1(n_1250),
.B2(n_1090),
.Y(n_1517)
);

OA21x2_ASAP7_75t_L g1518 ( 
.A1(n_1221),
.A2(n_1240),
.B(n_1226),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1313),
.A2(n_1242),
.B1(n_1250),
.B2(n_1325),
.Y(n_1519)
);

OAI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1260),
.A2(n_553),
.B(n_1223),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1225),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1308),
.A2(n_1323),
.B(n_1311),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1313),
.A2(n_1242),
.B1(n_1250),
.B2(n_1325),
.Y(n_1523)
);

OAI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1308),
.A2(n_1323),
.B(n_1311),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1404),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1395),
.Y(n_1526)
);

CKINVDCx20_ASAP7_75t_R g1527 ( 
.A(n_1381),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1517),
.A2(n_1407),
.B1(n_1519),
.B2(n_1505),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1514),
.B(n_1403),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1391),
.B(n_1483),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1517),
.A2(n_1519),
.B1(n_1523),
.B2(n_1505),
.Y(n_1531)
);

INVx1_ASAP7_75t_SL g1532 ( 
.A(n_1426),
.Y(n_1532)
);

O2A1O1Ixp5_ASAP7_75t_L g1533 ( 
.A1(n_1496),
.A2(n_1520),
.B(n_1508),
.C(n_1504),
.Y(n_1533)
);

INVxp67_ASAP7_75t_L g1534 ( 
.A(n_1442),
.Y(n_1534)
);

INVxp33_ASAP7_75t_L g1535 ( 
.A(n_1442),
.Y(n_1535)
);

O2A1O1Ixp33_ASAP7_75t_L g1536 ( 
.A1(n_1484),
.A2(n_1477),
.B(n_1516),
.C(n_1437),
.Y(n_1536)
);

CKINVDCx6p67_ASAP7_75t_R g1537 ( 
.A(n_1381),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1523),
.A2(n_1417),
.B1(n_1384),
.B2(n_1409),
.Y(n_1538)
);

AOI221xp5_ASAP7_75t_L g1539 ( 
.A1(n_1422),
.A2(n_1409),
.B1(n_1438),
.B2(n_1397),
.C(n_1482),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1500),
.B(n_1417),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1384),
.A2(n_1510),
.B1(n_1445),
.B2(n_1420),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1422),
.B(n_1428),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1445),
.A2(n_1398),
.B1(n_1401),
.B2(n_1503),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1404),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1492),
.B(n_1397),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1400),
.B(n_1394),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1394),
.B(n_1377),
.Y(n_1547)
);

O2A1O1Ixp5_ASAP7_75t_L g1548 ( 
.A1(n_1385),
.A2(n_1388),
.B(n_1448),
.C(n_1471),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1503),
.A2(n_1438),
.B1(n_1450),
.B2(n_1489),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1495),
.A2(n_1509),
.B1(n_1513),
.B2(n_1497),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1497),
.A2(n_1458),
.B1(n_1444),
.B2(n_1490),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1379),
.B(n_1486),
.Y(n_1552)
);

A2O1A1Ixp33_ASAP7_75t_L g1553 ( 
.A1(n_1454),
.A2(n_1468),
.B(n_1434),
.C(n_1421),
.Y(n_1553)
);

AOI21x1_ASAP7_75t_SL g1554 ( 
.A1(n_1474),
.A2(n_1475),
.B(n_1393),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1446),
.B(n_1455),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1378),
.B(n_1383),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1428),
.B(n_1393),
.Y(n_1557)
);

BUFx3_ASAP7_75t_L g1558 ( 
.A(n_1507),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_R g1559 ( 
.A(n_1465),
.B(n_1461),
.Y(n_1559)
);

OA21x2_ASAP7_75t_L g1560 ( 
.A1(n_1457),
.A2(n_1429),
.B(n_1466),
.Y(n_1560)
);

BUFx10_ASAP7_75t_L g1561 ( 
.A(n_1506),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1423),
.B(n_1430),
.Y(n_1562)
);

AOI21x1_ASAP7_75t_SL g1563 ( 
.A1(n_1425),
.A2(n_1479),
.B(n_1512),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_SL g1564 ( 
.A1(n_1465),
.A2(n_1402),
.B1(n_1414),
.B2(n_1416),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_1521),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_1507),
.Y(n_1566)
);

BUFx3_ASAP7_75t_L g1567 ( 
.A(n_1458),
.Y(n_1567)
);

NOR2xp67_ASAP7_75t_L g1568 ( 
.A(n_1435),
.B(n_1506),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_1431),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1491),
.B(n_1502),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1491),
.A2(n_1502),
.B1(n_1456),
.B2(n_1476),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1498),
.A2(n_1447),
.B1(n_1418),
.B2(n_1410),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1402),
.B(n_1414),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1416),
.B(n_1430),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1473),
.B(n_1428),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1387),
.A2(n_1405),
.B1(n_1396),
.B2(n_1389),
.Y(n_1576)
);

O2A1O1Ixp33_ASAP7_75t_L g1577 ( 
.A1(n_1386),
.A2(n_1481),
.B(n_1433),
.C(n_1436),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1390),
.B(n_1427),
.Y(n_1578)
);

OAI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1416),
.A2(n_1463),
.B1(n_1480),
.B2(n_1412),
.Y(n_1579)
);

OAI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1412),
.A2(n_1480),
.B1(n_1518),
.B2(n_1487),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1412),
.A2(n_1480),
.B1(n_1518),
.B2(n_1487),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1428),
.B(n_1425),
.Y(n_1582)
);

O2A1O1Ixp5_ASAP7_75t_L g1583 ( 
.A1(n_1469),
.A2(n_1424),
.B(n_1427),
.C(n_1459),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1406),
.A2(n_1415),
.B1(n_1512),
.B2(n_1470),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1469),
.B(n_1406),
.Y(n_1585)
);

CKINVDCx20_ASAP7_75t_R g1586 ( 
.A(n_1419),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1472),
.B(n_1452),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1415),
.A2(n_1501),
.B1(n_1515),
.B2(n_1413),
.Y(n_1588)
);

O2A1O1Ixp5_ASAP7_75t_L g1589 ( 
.A1(n_1462),
.A2(n_1376),
.B(n_1411),
.C(n_1464),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1460),
.B(n_1467),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1460),
.B(n_1439),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1432),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1439),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1440),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1382),
.A2(n_1441),
.B1(n_1408),
.B2(n_1453),
.Y(n_1595)
);

O2A1O1Ixp33_ASAP7_75t_L g1596 ( 
.A1(n_1451),
.A2(n_1443),
.B(n_1453),
.C(n_1419),
.Y(n_1596)
);

AOI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1419),
.A2(n_1449),
.B1(n_1443),
.B2(n_1399),
.Y(n_1597)
);

BUFx6f_ASAP7_75t_L g1598 ( 
.A(n_1380),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1392),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1478),
.B(n_1485),
.Y(n_1600)
);

O2A1O1Ixp5_ASAP7_75t_L g1601 ( 
.A1(n_1493),
.A2(n_1494),
.B(n_1499),
.C(n_1511),
.Y(n_1601)
);

OA21x2_ASAP7_75t_L g1602 ( 
.A1(n_1524),
.A2(n_1488),
.B(n_1522),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1514),
.B(n_1403),
.Y(n_1603)
);

OA21x2_ASAP7_75t_L g1604 ( 
.A1(n_1457),
.A2(n_1429),
.B(n_1466),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1384),
.B(n_1422),
.Y(n_1605)
);

O2A1O1Ixp33_ASAP7_75t_L g1606 ( 
.A1(n_1496),
.A2(n_1520),
.B(n_1374),
.C(n_1242),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1391),
.B(n_1483),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1492),
.B(n_1446),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1514),
.B(n_1403),
.Y(n_1609)
);

NOR2xp67_ASAP7_75t_R g1610 ( 
.A(n_1412),
.B(n_1369),
.Y(n_1610)
);

INVx1_ASAP7_75t_SL g1611 ( 
.A(n_1403),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1391),
.B(n_1483),
.Y(n_1612)
);

AND2x4_ASAP7_75t_L g1613 ( 
.A(n_1379),
.B(n_1486),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1514),
.B(n_1403),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_1506),
.Y(n_1615)
);

BUFx3_ASAP7_75t_L g1616 ( 
.A(n_1404),
.Y(n_1616)
);

OAI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1517),
.A2(n_1332),
.B1(n_1407),
.B2(n_1505),
.Y(n_1617)
);

OA21x2_ASAP7_75t_L g1618 ( 
.A1(n_1457),
.A2(n_1429),
.B(n_1466),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1514),
.B(n_1403),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1395),
.Y(n_1620)
);

INVx1_ASAP7_75t_SL g1621 ( 
.A(n_1403),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1492),
.B(n_1446),
.Y(n_1622)
);

BUFx6f_ASAP7_75t_L g1623 ( 
.A(n_1598),
.Y(n_1623)
);

AND2x4_ASAP7_75t_SL g1624 ( 
.A(n_1578),
.B(n_1552),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1542),
.B(n_1557),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1575),
.B(n_1557),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1546),
.B(n_1547),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1542),
.B(n_1582),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1592),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1582),
.B(n_1545),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1593),
.Y(n_1631)
);

AOI21xp33_ASAP7_75t_L g1632 ( 
.A1(n_1606),
.A2(n_1536),
.B(n_1533),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1526),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1540),
.B(n_1555),
.Y(n_1634)
);

AO31x2_ASAP7_75t_L g1635 ( 
.A1(n_1553),
.A2(n_1581),
.A3(n_1580),
.B(n_1584),
.Y(n_1635)
);

OAI21x1_ASAP7_75t_L g1636 ( 
.A1(n_1601),
.A2(n_1583),
.B(n_1560),
.Y(n_1636)
);

OA21x2_ASAP7_75t_L g1637 ( 
.A1(n_1589),
.A2(n_1548),
.B(n_1553),
.Y(n_1637)
);

OR2x6_ASAP7_75t_L g1638 ( 
.A(n_1577),
.B(n_1596),
.Y(n_1638)
);

OAI21x1_ASAP7_75t_L g1639 ( 
.A1(n_1560),
.A2(n_1604),
.B(n_1618),
.Y(n_1639)
);

OAI222xp33_ASAP7_75t_L g1640 ( 
.A1(n_1531),
.A2(n_1528),
.B1(n_1538),
.B2(n_1617),
.C1(n_1541),
.C2(n_1605),
.Y(n_1640)
);

BUFx4f_ASAP7_75t_SL g1641 ( 
.A(n_1527),
.Y(n_1641)
);

OA21x2_ASAP7_75t_L g1642 ( 
.A1(n_1591),
.A2(n_1590),
.B(n_1594),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1585),
.B(n_1532),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_1569),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1620),
.B(n_1574),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1530),
.B(n_1607),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1539),
.A2(n_1543),
.B1(n_1605),
.B2(n_1549),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1599),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1562),
.Y(n_1649)
);

OAI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1551),
.A2(n_1612),
.B(n_1597),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1576),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1550),
.B(n_1534),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1572),
.Y(n_1653)
);

INVx4_ASAP7_75t_L g1654 ( 
.A(n_1578),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1556),
.Y(n_1655)
);

OAI21x1_ASAP7_75t_L g1656 ( 
.A1(n_1560),
.A2(n_1618),
.B(n_1604),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1535),
.B(n_1552),
.Y(n_1657)
);

OR2x6_ASAP7_75t_L g1658 ( 
.A(n_1600),
.B(n_1571),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1535),
.B(n_1622),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1600),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1618),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1602),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1608),
.B(n_1613),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1633),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1625),
.B(n_1570),
.Y(n_1665)
);

INVxp67_ASAP7_75t_SL g1666 ( 
.A(n_1631),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1626),
.B(n_1621),
.Y(n_1667)
);

AO21x2_ASAP7_75t_L g1668 ( 
.A1(n_1639),
.A2(n_1656),
.B(n_1636),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1631),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1628),
.B(n_1619),
.Y(n_1670)
);

INVx2_ASAP7_75t_SL g1671 ( 
.A(n_1660),
.Y(n_1671)
);

INVxp67_ASAP7_75t_L g1672 ( 
.A(n_1648),
.Y(n_1672)
);

INVx1_ASAP7_75t_SL g1673 ( 
.A(n_1643),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1642),
.B(n_1609),
.Y(n_1674)
);

OAI21x1_ASAP7_75t_L g1675 ( 
.A1(n_1639),
.A2(n_1563),
.B(n_1554),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1632),
.A2(n_1611),
.B1(n_1603),
.B2(n_1529),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1627),
.B(n_1614),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1627),
.B(n_1565),
.Y(n_1678)
);

OR2x6_ASAP7_75t_L g1679 ( 
.A(n_1658),
.B(n_1564),
.Y(n_1679)
);

INVx1_ASAP7_75t_SL g1680 ( 
.A(n_1643),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1655),
.B(n_1567),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1630),
.B(n_1635),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1632),
.A2(n_1537),
.B1(n_1586),
.B2(n_1525),
.Y(n_1683)
);

BUFx6f_ASAP7_75t_L g1684 ( 
.A(n_1623),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1635),
.B(n_1587),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1655),
.B(n_1544),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1635),
.B(n_1573),
.Y(n_1687)
);

BUFx8_ASAP7_75t_L g1688 ( 
.A(n_1667),
.Y(n_1688)
);

AOI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1682),
.A2(n_1640),
.B1(n_1650),
.B2(n_1647),
.C(n_1646),
.Y(n_1689)
);

AOI222xp33_ASAP7_75t_L g1690 ( 
.A1(n_1676),
.A2(n_1640),
.B1(n_1650),
.B2(n_1653),
.C1(n_1641),
.C2(n_1652),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1669),
.Y(n_1691)
);

AOI21xp33_ASAP7_75t_L g1692 ( 
.A1(n_1683),
.A2(n_1638),
.B(n_1652),
.Y(n_1692)
);

OR2x6_ASAP7_75t_L g1693 ( 
.A(n_1679),
.B(n_1638),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1683),
.A2(n_1638),
.B1(n_1634),
.B2(n_1595),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1669),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1664),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1678),
.B(n_1659),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1678),
.B(n_1634),
.Y(n_1698)
);

INVxp67_ASAP7_75t_L g1699 ( 
.A(n_1667),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_SL g1700 ( 
.A(n_1677),
.B(n_1657),
.Y(n_1700)
);

AOI222xp33_ASAP7_75t_L g1701 ( 
.A1(n_1676),
.A2(n_1651),
.B1(n_1610),
.B2(n_1663),
.C1(n_1649),
.C2(n_1588),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_SL g1702 ( 
.A1(n_1679),
.A2(n_1586),
.B1(n_1527),
.B2(n_1569),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1673),
.B(n_1626),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1665),
.B(n_1624),
.Y(n_1704)
);

NOR4xp25_ASAP7_75t_SL g1705 ( 
.A(n_1666),
.B(n_1629),
.C(n_1615),
.D(n_1644),
.Y(n_1705)
);

INVxp67_ASAP7_75t_SL g1706 ( 
.A(n_1672),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1677),
.B(n_1558),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_1681),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1679),
.A2(n_1638),
.B1(n_1579),
.B2(n_1658),
.Y(n_1709)
);

AND2x4_ASAP7_75t_SL g1710 ( 
.A(n_1679),
.B(n_1654),
.Y(n_1710)
);

AO21x2_ASAP7_75t_L g1711 ( 
.A1(n_1668),
.A2(n_1661),
.B(n_1662),
.Y(n_1711)
);

OA21x2_ASAP7_75t_L g1712 ( 
.A1(n_1675),
.A2(n_1639),
.B(n_1656),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1671),
.B(n_1687),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1679),
.A2(n_1638),
.B1(n_1537),
.B2(n_1637),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1673),
.B(n_1645),
.Y(n_1715)
);

INVx2_ASAP7_75t_SL g1716 ( 
.A(n_1671),
.Y(n_1716)
);

INVxp67_ASAP7_75t_L g1717 ( 
.A(n_1667),
.Y(n_1717)
);

NOR2x1_ASAP7_75t_R g1718 ( 
.A(n_1686),
.B(n_1615),
.Y(n_1718)
);

BUFx3_ASAP7_75t_L g1719 ( 
.A(n_1681),
.Y(n_1719)
);

INVx6_ASAP7_75t_L g1720 ( 
.A(n_1684),
.Y(n_1720)
);

OAI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1690),
.A2(n_1675),
.B(n_1637),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1696),
.Y(n_1722)
);

INVx3_ASAP7_75t_L g1723 ( 
.A(n_1713),
.Y(n_1723)
);

INVx3_ASAP7_75t_L g1724 ( 
.A(n_1713),
.Y(n_1724)
);

INVx2_ASAP7_75t_SL g1725 ( 
.A(n_1720),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1698),
.B(n_1686),
.Y(n_1726)
);

INVx2_ASAP7_75t_SL g1727 ( 
.A(n_1720),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1711),
.Y(n_1728)
);

HB1xp67_ASAP7_75t_L g1729 ( 
.A(n_1691),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1711),
.Y(n_1730)
);

BUFx2_ASAP7_75t_L g1731 ( 
.A(n_1716),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1698),
.B(n_1670),
.Y(n_1732)
);

INVxp67_ASAP7_75t_L g1733 ( 
.A(n_1706),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1695),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1703),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1720),
.B(n_1674),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1699),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1717),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1712),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1719),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1739),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1723),
.B(n_1704),
.Y(n_1742)
);

NAND2x1_ASAP7_75t_L g1743 ( 
.A(n_1723),
.B(n_1693),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1723),
.B(n_1724),
.Y(n_1744)
);

AND2x4_ASAP7_75t_L g1745 ( 
.A(n_1723),
.B(n_1710),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1739),
.Y(n_1746)
);

NOR2xp67_ASAP7_75t_L g1747 ( 
.A(n_1723),
.B(n_1671),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1737),
.B(n_1680),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1739),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1739),
.Y(n_1750)
);

INVxp67_ASAP7_75t_SL g1751 ( 
.A(n_1729),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1726),
.B(n_1718),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1722),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1730),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1730),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1724),
.B(n_1719),
.Y(n_1756)
);

INVxp67_ASAP7_75t_L g1757 ( 
.A(n_1726),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1737),
.B(n_1700),
.Y(n_1758)
);

NAND4xp25_ASAP7_75t_L g1759 ( 
.A(n_1721),
.B(n_1689),
.C(n_1701),
.D(n_1692),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1730),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1737),
.B(n_1700),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1732),
.B(n_1707),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1730),
.Y(n_1763)
);

INVx2_ASAP7_75t_SL g1764 ( 
.A(n_1725),
.Y(n_1764)
);

INVx1_ASAP7_75t_SL g1765 ( 
.A(n_1729),
.Y(n_1765)
);

AND3x2_ASAP7_75t_L g1766 ( 
.A(n_1733),
.B(n_1707),
.C(n_1685),
.Y(n_1766)
);

AND2x4_ASAP7_75t_L g1767 ( 
.A(n_1724),
.B(n_1710),
.Y(n_1767)
);

INVx1_ASAP7_75t_SL g1768 ( 
.A(n_1740),
.Y(n_1768)
);

AND3x2_ASAP7_75t_L g1769 ( 
.A(n_1733),
.B(n_1685),
.C(n_1672),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1738),
.B(n_1680),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1730),
.Y(n_1771)
);

BUFx6f_ASAP7_75t_L g1772 ( 
.A(n_1725),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1735),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1738),
.B(n_1715),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1738),
.B(n_1697),
.Y(n_1775)
);

NAND3xp33_ASAP7_75t_L g1776 ( 
.A(n_1721),
.B(n_1714),
.C(n_1694),
.Y(n_1776)
);

HB1xp67_ASAP7_75t_L g1777 ( 
.A(n_1735),
.Y(n_1777)
);

AND2x4_ASAP7_75t_L g1778 ( 
.A(n_1724),
.B(n_1693),
.Y(n_1778)
);

INVxp67_ASAP7_75t_L g1779 ( 
.A(n_1732),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1725),
.B(n_1693),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1773),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1777),
.Y(n_1782)
);

AND2x4_ASAP7_75t_L g1783 ( 
.A(n_1764),
.B(n_1725),
.Y(n_1783)
);

NAND2x1p5_ASAP7_75t_L g1784 ( 
.A(n_1743),
.B(n_1740),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1780),
.B(n_1740),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1757),
.B(n_1740),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1764),
.B(n_1727),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1753),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1775),
.B(n_1740),
.Y(n_1789)
);

INVxp67_ASAP7_75t_L g1790 ( 
.A(n_1751),
.Y(n_1790)
);

INVxp67_ASAP7_75t_L g1791 ( 
.A(n_1765),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1775),
.B(n_1734),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1779),
.B(n_1708),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1780),
.B(n_1736),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1780),
.B(n_1736),
.Y(n_1795)
);

INVx2_ASAP7_75t_SL g1796 ( 
.A(n_1772),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1762),
.B(n_1708),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1772),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1772),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1759),
.B(n_1670),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1774),
.B(n_1734),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1753),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1780),
.B(n_1736),
.Y(n_1803)
);

AOI211xp5_ASAP7_75t_L g1804 ( 
.A1(n_1759),
.A2(n_1721),
.B(n_1702),
.C(n_1709),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1774),
.B(n_1734),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_SL g1806 ( 
.A(n_1776),
.B(n_1688),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_L g1807 ( 
.A(n_1752),
.B(n_1561),
.Y(n_1807)
);

NOR2x1_ASAP7_75t_L g1808 ( 
.A(n_1765),
.B(n_1731),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1748),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1758),
.B(n_1687),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1776),
.B(n_1561),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1742),
.B(n_1736),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1758),
.B(n_1561),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1748),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1770),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1761),
.B(n_1770),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1791),
.B(n_1761),
.Y(n_1817)
);

BUFx2_ASAP7_75t_L g1818 ( 
.A(n_1808),
.Y(n_1818)
);

HB1xp67_ASAP7_75t_L g1819 ( 
.A(n_1791),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_L g1820 ( 
.A1(n_1806),
.A2(n_1693),
.B1(n_1778),
.B2(n_1714),
.Y(n_1820)
);

OAI21x1_ASAP7_75t_L g1821 ( 
.A1(n_1784),
.A2(n_1743),
.B(n_1728),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1790),
.B(n_1768),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1790),
.B(n_1768),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1788),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1802),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1785),
.B(n_1756),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1781),
.B(n_1766),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1796),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1801),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_L g1830 ( 
.A(n_1807),
.B(n_1778),
.Y(n_1830)
);

INVx2_ASAP7_75t_SL g1831 ( 
.A(n_1783),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1794),
.B(n_1756),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1805),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1809),
.Y(n_1834)
);

AND2x4_ASAP7_75t_L g1835 ( 
.A(n_1783),
.B(n_1747),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1795),
.B(n_1745),
.Y(n_1836)
);

INVx1_ASAP7_75t_SL g1837 ( 
.A(n_1783),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1787),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1803),
.B(n_1784),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1782),
.B(n_1722),
.Y(n_1840)
);

AOI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1806),
.A2(n_1778),
.B1(n_1679),
.B2(n_1745),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1816),
.B(n_1772),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1787),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_SL g1844 ( 
.A(n_1818),
.B(n_1804),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1819),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1822),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1836),
.B(n_1814),
.Y(n_1847)
);

AOI322xp5_ASAP7_75t_L g1848 ( 
.A1(n_1818),
.A2(n_1800),
.A3(n_1811),
.B1(n_1815),
.B2(n_1793),
.C1(n_1786),
.C2(n_1797),
.Y(n_1848)
);

OAI21xp33_ASAP7_75t_L g1849 ( 
.A1(n_1841),
.A2(n_1811),
.B(n_1813),
.Y(n_1849)
);

INVxp67_ASAP7_75t_SL g1850 ( 
.A(n_1831),
.Y(n_1850)
);

INVxp67_ASAP7_75t_SL g1851 ( 
.A(n_1831),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_SL g1852 ( 
.A(n_1837),
.B(n_1787),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1836),
.B(n_1796),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1822),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1823),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_L g1856 ( 
.A(n_1830),
.B(n_1807),
.Y(n_1856)
);

CKINVDCx16_ASAP7_75t_R g1857 ( 
.A(n_1817),
.Y(n_1857)
);

AOI322xp5_ASAP7_75t_L g1858 ( 
.A1(n_1820),
.A2(n_1827),
.A3(n_1823),
.B1(n_1834),
.B2(n_1837),
.C1(n_1829),
.C2(n_1833),
.Y(n_1858)
);

OAI221xp5_ASAP7_75t_L g1859 ( 
.A1(n_1827),
.A2(n_1813),
.B1(n_1789),
.B2(n_1792),
.C(n_1799),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1826),
.B(n_1798),
.Y(n_1860)
);

NAND2xp33_ASAP7_75t_L g1861 ( 
.A(n_1817),
.B(n_1559),
.Y(n_1861)
);

OAI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1821),
.A2(n_1799),
.B(n_1798),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1834),
.B(n_1812),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1824),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1857),
.B(n_1838),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1845),
.B(n_1829),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1853),
.B(n_1832),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1850),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1851),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1846),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1853),
.Y(n_1871)
);

AOI22xp33_ASAP7_75t_SL g1872 ( 
.A1(n_1859),
.A2(n_1839),
.B1(n_1832),
.B2(n_1826),
.Y(n_1872)
);

INVxp67_ASAP7_75t_L g1873 ( 
.A(n_1852),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1863),
.B(n_1842),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_L g1875 ( 
.A(n_1844),
.B(n_1833),
.Y(n_1875)
);

INVxp67_ASAP7_75t_SL g1876 ( 
.A(n_1852),
.Y(n_1876)
);

NOR2x1_ASAP7_75t_SL g1877 ( 
.A(n_1844),
.B(n_1842),
.Y(n_1877)
);

AOI221xp5_ASAP7_75t_L g1878 ( 
.A1(n_1876),
.A2(n_1875),
.B1(n_1873),
.B2(n_1866),
.C(n_1855),
.Y(n_1878)
);

NOR4xp25_ASAP7_75t_L g1879 ( 
.A(n_1875),
.B(n_1854),
.C(n_1864),
.D(n_1861),
.Y(n_1879)
);

O2A1O1Ixp33_ASAP7_75t_L g1880 ( 
.A1(n_1865),
.A2(n_1861),
.B(n_1849),
.C(n_1856),
.Y(n_1880)
);

OAI211xp5_ASAP7_75t_L g1881 ( 
.A1(n_1872),
.A2(n_1858),
.B(n_1848),
.C(n_1862),
.Y(n_1881)
);

NOR3xp33_ASAP7_75t_L g1882 ( 
.A(n_1868),
.B(n_1847),
.C(n_1860),
.Y(n_1882)
);

O2A1O1Ixp33_ASAP7_75t_L g1883 ( 
.A1(n_1869),
.A2(n_1828),
.B(n_1824),
.C(n_1825),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_L g1884 ( 
.A(n_1877),
.B(n_1847),
.Y(n_1884)
);

AOI221xp5_ASAP7_75t_L g1885 ( 
.A1(n_1866),
.A2(n_1860),
.B1(n_1825),
.B2(n_1843),
.C(n_1838),
.Y(n_1885)
);

NOR3xp33_ASAP7_75t_L g1886 ( 
.A(n_1870),
.B(n_1874),
.C(n_1871),
.Y(n_1886)
);

NOR2x1_ASAP7_75t_L g1887 ( 
.A(n_1871),
.B(n_1838),
.Y(n_1887)
);

AOI221xp5_ASAP7_75t_L g1888 ( 
.A1(n_1867),
.A2(n_1843),
.B1(n_1840),
.B2(n_1839),
.C(n_1835),
.Y(n_1888)
);

AOI22xp33_ASAP7_75t_L g1889 ( 
.A1(n_1878),
.A2(n_1843),
.B1(n_1835),
.B2(n_1778),
.Y(n_1889)
);

AOI321xp33_ASAP7_75t_L g1890 ( 
.A1(n_1881),
.A2(n_1840),
.A3(n_1835),
.B1(n_1771),
.B2(n_1754),
.C(n_1755),
.Y(n_1890)
);

OAI22xp33_ASAP7_75t_SL g1891 ( 
.A1(n_1884),
.A2(n_1835),
.B1(n_1727),
.B2(n_1728),
.Y(n_1891)
);

AOI22x1_ASAP7_75t_L g1892 ( 
.A1(n_1879),
.A2(n_1772),
.B1(n_1744),
.B2(n_1727),
.Y(n_1892)
);

OAI21xp5_ASAP7_75t_SL g1893 ( 
.A1(n_1880),
.A2(n_1882),
.B(n_1886),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1887),
.Y(n_1894)
);

INVx2_ASAP7_75t_SL g1895 ( 
.A(n_1883),
.Y(n_1895)
);

NAND3xp33_ASAP7_75t_L g1896 ( 
.A(n_1890),
.B(n_1885),
.C(n_1888),
.Y(n_1896)
);

HB1xp67_ASAP7_75t_L g1897 ( 
.A(n_1894),
.Y(n_1897)
);

HB1xp67_ASAP7_75t_L g1898 ( 
.A(n_1892),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1895),
.B(n_1769),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_SL g1900 ( 
.A(n_1891),
.B(n_1772),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1889),
.B(n_1742),
.Y(n_1901)
);

NOR3xp33_ASAP7_75t_L g1902 ( 
.A(n_1893),
.B(n_1821),
.C(n_1568),
.Y(n_1902)
);

OAI22xp5_ASAP7_75t_L g1903 ( 
.A1(n_1896),
.A2(n_1727),
.B1(n_1810),
.B2(n_1747),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_R g1904 ( 
.A(n_1897),
.B(n_1559),
.Y(n_1904)
);

OAI321xp33_ASAP7_75t_L g1905 ( 
.A1(n_1899),
.A2(n_1760),
.A3(n_1771),
.B1(n_1754),
.B2(n_1755),
.C(n_1763),
.Y(n_1905)
);

INVx2_ASAP7_75t_SL g1906 ( 
.A(n_1900),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_R g1907 ( 
.A(n_1898),
.B(n_1558),
.Y(n_1907)
);

XNOR2x1_ASAP7_75t_L g1908 ( 
.A(n_1901),
.B(n_1821),
.Y(n_1908)
);

NOR2x1_ASAP7_75t_L g1909 ( 
.A(n_1908),
.B(n_1902),
.Y(n_1909)
);

NAND2xp33_ASAP7_75t_R g1910 ( 
.A(n_1904),
.B(n_1705),
.Y(n_1910)
);

AOI322xp5_ASAP7_75t_L g1911 ( 
.A1(n_1906),
.A2(n_1728),
.A3(n_1771),
.B1(n_1763),
.B2(n_1760),
.C1(n_1755),
.C2(n_1754),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1909),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1912),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1913),
.Y(n_1914)
);

OAI21x1_ASAP7_75t_SL g1915 ( 
.A1(n_1913),
.A2(n_1907),
.B(n_1903),
.Y(n_1915)
);

OAI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1914),
.A2(n_1910),
.B1(n_1905),
.B2(n_1760),
.Y(n_1916)
);

AO22x2_ASAP7_75t_L g1917 ( 
.A1(n_1915),
.A2(n_1763),
.B1(n_1746),
.B2(n_1749),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1917),
.Y(n_1918)
);

AOI22xp5_ASAP7_75t_L g1919 ( 
.A1(n_1916),
.A2(n_1744),
.B1(n_1741),
.B2(n_1750),
.Y(n_1919)
);

AOI21xp33_ASAP7_75t_SL g1920 ( 
.A1(n_1918),
.A2(n_1911),
.B(n_1746),
.Y(n_1920)
);

OAI22xp5_ASAP7_75t_SL g1921 ( 
.A1(n_1920),
.A2(n_1919),
.B1(n_1566),
.B2(n_1616),
.Y(n_1921)
);

AOI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1921),
.A2(n_1746),
.B(n_1741),
.Y(n_1922)
);

AOI22xp5_ASAP7_75t_SL g1923 ( 
.A1(n_1922),
.A2(n_1566),
.B1(n_1616),
.B2(n_1767),
.Y(n_1923)
);

AOI22xp33_ASAP7_75t_L g1924 ( 
.A1(n_1923),
.A2(n_1741),
.B1(n_1749),
.B2(n_1750),
.Y(n_1924)
);

AOI211xp5_ASAP7_75t_L g1925 ( 
.A1(n_1924),
.A2(n_1750),
.B(n_1749),
.C(n_1728),
.Y(n_1925)
);


endmodule