module real_jpeg_7135_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_164;
wire n_48;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_222;
wire n_19;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_187;
wire n_75;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_202;
wire n_128;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_1),
.A2(n_163),
.B1(n_164),
.B2(n_167),
.Y(n_162)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_1),
.Y(n_167)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_3),
.A2(n_49),
.B1(n_61),
.B2(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_3),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_3),
.A2(n_93),
.B1(n_145),
.B2(n_147),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_3),
.A2(n_41),
.B1(n_93),
.B2(n_196),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_4),
.A2(n_21),
.B1(n_27),
.B2(n_28),
.Y(n_20)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_6),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_6),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_7),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_7),
.Y(n_160)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_9),
.A2(n_49),
.B1(n_97),
.B2(n_100),
.Y(n_96)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_9),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_9),
.A2(n_21),
.B1(n_100),
.B2(n_196),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_10),
.Y(n_79)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_10),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_11),
.A2(n_28),
.B1(n_41),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_11),
.A2(n_44),
.B1(n_127),
.B2(n_130),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_11),
.A2(n_44),
.B1(n_64),
.B2(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_12),
.B(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_12),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_12),
.A2(n_49),
.B1(n_123),
.B2(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_12),
.B(n_187),
.C(n_190),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_12),
.B(n_118),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_12),
.B(n_203),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_12),
.B(n_95),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_174),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_172),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_134),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_16),
.B(n_134),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_67),
.C(n_101),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_17),
.B(n_237),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_45),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_18),
.B(n_45),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_30),
.B(n_33),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_20),
.A2(n_34),
.B1(n_162),
.B2(n_168),
.Y(n_161)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx4_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_25),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_28),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_29),
.Y(n_192)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_31),
.A2(n_34),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_33),
.A2(n_222),
.B(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_40),
.Y(n_33)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_34),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_40),
.B(n_202),
.Y(n_201)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI32xp33_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_49),
.A3(n_51),
.B1(n_55),
.B2(n_60),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_47),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_48),
.Y(n_117)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_48),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_50),
.Y(n_120)
);

AO22x2_ASAP7_75t_L g118 ( 
.A1(n_51),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_118)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_59),
.Y(n_149)
);

NAND2xp33_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_66),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_67),
.A2(n_101),
.B1(n_102),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_67),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_92),
.B1(n_94),
.B2(n_96),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_68),
.A2(n_96),
.B(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_68),
.A2(n_138),
.B(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_69),
.B(n_139),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_83),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_73),
.B1(n_76),
.B2(n_80),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_82),
.Y(n_183)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_83),
.A2(n_92),
.B(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_86),
.B1(n_89),
.B2(n_91),
.Y(n_83)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_85),
.Y(n_189)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_88),
.Y(n_217)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_90),
.Y(n_166)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_95),
.B(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_122),
.B(n_125),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_103),
.B(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_118),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B1(n_111),
.B2(n_115),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_110),
.Y(n_157)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_SL g122 ( 
.A1(n_116),
.A2(n_123),
.B(n_124),
.Y(n_122)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_118),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_154),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_123),
.A2(n_200),
.B(n_201),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_133),
.Y(n_125)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_133),
.A2(n_144),
.B(n_150),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_142),
.B2(n_171),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_141),
.Y(n_136)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_152),
.Y(n_142)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_161),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_158),
.B2(n_159),
.Y(n_154)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_234),
.B(n_239),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_210),
.B(n_233),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_193),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_177),
.B(n_193),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_184),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_178),
.A2(n_184),
.B1(n_185),
.B2(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_178),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_204),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_194),
.B(n_205),
.C(n_209),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_200),
.B(n_201),
.Y(n_194)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_208),
.B2(n_209),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_226),
.B(n_232),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_220),
.B(n_225),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_219),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_218),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_224),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_224),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_222),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_230),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_236),
.Y(n_239)
);


endmodule