module fake_jpeg_27898_n_84 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_84);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_84;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_40),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_38),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_42),
.Y(n_55)
);

NOR3xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_13),
.C(n_27),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_1),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx6f_ASAP7_75t_SL g53 ( 
.A(n_45),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_37),
.B1(n_32),
.B2(n_31),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_46),
.A2(n_50),
.B1(n_51),
.B2(n_11),
.Y(n_57)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_3),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_36),
.B1(n_33),
.B2(n_37),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_30),
.B1(n_14),
.B2(n_16),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_43),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_52),
.B(n_56),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_60),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_55),
.A2(n_10),
.B1(n_26),
.B2(n_25),
.Y(n_59)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_50),
.A2(n_9),
.B1(n_24),
.B2(n_23),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_48),
.A2(n_29),
.B1(n_7),
.B2(n_8),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_63),
.Y(n_74)
);

O2A1O1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_6),
.B(n_21),
.C(n_18),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_66),
.B(n_68),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_1),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_22),
.Y(n_64)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_65),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_52),
.B(n_2),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_59),
.B1(n_62),
.B2(n_65),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_76),
.C(n_58),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_71),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

INVxp33_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

AOI21x1_ASAP7_75t_SL g81 ( 
.A1(n_80),
.A2(n_79),
.B(n_72),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_79),
.C(n_72),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_73),
.C(n_74),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_67),
.Y(n_84)
);


endmodule