module real_jpeg_29871_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_336, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_336;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_0),
.A2(n_31),
.B1(n_33),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_0),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_54),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_0),
.A2(n_54),
.B1(n_63),
.B2(n_65),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_0),
.A2(n_47),
.B1(n_48),
.B2(n_54),
.Y(n_134)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_1),
.Y(n_106)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_1),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_1),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_2),
.A2(n_35),
.B1(n_47),
.B2(n_48),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_2),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_2),
.A2(n_35),
.B1(n_63),
.B2(n_65),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_3),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_3),
.A2(n_31),
.B1(n_33),
.B2(n_152),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_3),
.A2(n_47),
.B1(n_48),
.B2(n_152),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_3),
.A2(n_63),
.B1(n_65),
.B2(n_152),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_4),
.A2(n_31),
.B1(n_33),
.B2(n_37),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_4),
.A2(n_37),
.B1(n_47),
.B2(n_48),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_4),
.A2(n_37),
.B1(n_63),
.B2(n_65),
.Y(n_140)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_6),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_6),
.B(n_30),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_6),
.B(n_33),
.Y(n_223)
);

AOI21xp33_ASAP7_75t_L g227 ( 
.A1(n_6),
.A2(n_33),
.B(n_223),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_6),
.A2(n_47),
.B1(n_48),
.B2(n_184),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_6),
.A2(n_60),
.B(n_63),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_6),
.B(n_88),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_6),
.A2(n_106),
.B1(n_129),
.B2(n_271),
.Y(n_273)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_8),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_8),
.A2(n_31),
.B1(n_33),
.B2(n_123),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_8),
.A2(n_47),
.B1(n_48),
.B2(n_123),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_8),
.A2(n_63),
.B1(n_65),
.B2(n_123),
.Y(n_258)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_10),
.A2(n_31),
.B1(n_33),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_10),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_10),
.A2(n_51),
.B1(n_63),
.B2(n_65),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_51),
.Y(n_125)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_12),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_12),
.A2(n_31),
.B1(n_33),
.B2(n_186),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_12),
.A2(n_47),
.B1(n_48),
.B2(n_186),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_12),
.A2(n_63),
.B1(n_65),
.B2(n_186),
.Y(n_271)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx11_ASAP7_75t_SL g64 ( 
.A(n_15),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_95),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_93),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_80),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_19),
.B(n_80),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_70),
.C(n_74),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_20),
.A2(n_21),
.B1(n_70),
.B2(n_322),
.Y(n_326)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_39),
.B1(n_40),
.B2(n_69),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_22),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_23),
.A2(n_122),
.B(n_124),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_23),
.A2(n_38),
.B1(n_122),
.B2(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_23),
.A2(n_38),
.B1(n_151),
.B2(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_24),
.B(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_24),
.A2(n_84),
.B(n_85),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_24),
.A2(n_85),
.B(n_125),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_24),
.A2(n_30),
.B1(n_183),
.B2(n_185),
.Y(n_182)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_26),
.B1(n_31),
.B2(n_33),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_25),
.B(n_33),
.Y(n_197)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

HAxp5_ASAP7_75t_SL g183 ( 
.A(n_27),
.B(n_184),
.CON(n_183),
.SN(n_183)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_29),
.A2(n_31),
.B1(n_183),
.B2(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_30),
.B(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_31),
.A2(n_33),
.B1(n_45),
.B2(n_49),
.Y(n_56)
);

AOI32xp33_ASAP7_75t_L g221 ( 
.A1(n_31),
.A2(n_47),
.A3(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_221)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_34),
.A2(n_38),
.B(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_36),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_38),
.B(n_73),
.Y(n_85)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_57),
.B2(n_68),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_42),
.B(n_57),
.C(n_69),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_52),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_43),
.A2(n_76),
.B(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_50),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_44),
.A2(n_55),
.B1(n_78),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_44),
.A2(n_55),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_44),
.A2(n_55),
.B1(n_180),
.B2(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_44),
.A2(n_55),
.B1(n_209),
.B2(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_44)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_45),
.Y(n_222)
);

NAND2xp33_ASAP7_75t_SL g224 ( 
.A(n_45),
.B(n_48),
.Y(n_224)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_48),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_48),
.A2(n_61),
.B(n_184),
.C(n_250),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_50),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_52),
.A2(n_88),
.B(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_57),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_57),
.A2(n_68),
.B1(n_75),
.B2(n_320),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_62),
.B(n_66),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_58),
.A2(n_62),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_58),
.A2(n_115),
.B(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_58),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_58),
.A2(n_66),
.B(n_133),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_58),
.A2(n_62),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_58),
.A2(n_158),
.B(n_231),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_58),
.A2(n_62),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_58),
.A2(n_62),
.B1(n_230),
.B2(n_248),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_65),
.Y(n_62)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_62),
.A2(n_114),
.B(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_62),
.B(n_184),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_63),
.Y(n_65)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_65),
.B(n_275),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_67),
.B(n_135),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_70),
.C(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_70),
.A2(n_319),
.B1(n_321),
.B2(n_322),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_70),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_74),
.B(n_326),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_75),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B(n_79),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_76),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_76),
.A2(n_79),
.B(n_89),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI321xp33_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_315),
.A3(n_327),
.B1(n_333),
.B2(n_334),
.C(n_336),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_169),
.B(n_314),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_153),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_98),
.B(n_153),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_126),
.C(n_137),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_99),
.A2(n_100),
.B1(n_126),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_116),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_101),
.B(n_118),
.C(n_120),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_113),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_102),
.B(n_113),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_109),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_103),
.A2(n_199),
.B(n_200),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_104),
.A2(n_112),
.B(n_142),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_104),
.A2(n_110),
.B1(n_262),
.B2(n_264),
.Y(n_261)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_106),
.A2(n_129),
.B1(n_263),
.B2(n_271),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_106),
.B(n_184),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_109),
.A2(n_129),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.Y(n_109)
);

INVx5_ASAP7_75t_SL g130 ( 
.A(n_110),
.Y(n_130)
);

INVx11_ASAP7_75t_L g200 ( 
.A(n_110),
.Y(n_200)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_112),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_119),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_126),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_132),
.B2(n_136),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_127),
.A2(n_128),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_132),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_L g324 ( 
.A1(n_128),
.A2(n_163),
.B(n_166),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B(n_131),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_129),
.A2(n_140),
.B(n_141),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_129),
.A2(n_140),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_132),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_134),
.B(n_147),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_137),
.B(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_148),
.C(n_149),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_138),
.B(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_145),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_145),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_304),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_148),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_167),
.B2(n_168),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_162),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_156),
.B(n_162),
.C(n_168),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_159),
.B(n_161),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_159),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_161),
.B(n_317),
.C(n_323),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_161),
.A2(n_317),
.B1(n_318),
.B2(n_332),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_161),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_167),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_308),
.B(n_313),
.Y(n_169)
);

O2A1O1Ixp33_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_213),
.B(n_294),
.C(n_307),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_201),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_172),
.B(n_201),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_187),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_174),
.B(n_175),
.C(n_187),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.C(n_182),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_182),
.B(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_185),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_195),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_189),
.B(n_193),
.C(n_195),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_198),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.C(n_207),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_202),
.A2(n_203),
.B1(n_289),
.B2(n_291),
.Y(n_288)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_290),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_207),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.C(n_212),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_212),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_293),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_286),
.B(n_292),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_241),
.B(n_285),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_232),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_217),
.B(n_232),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_225),
.C(n_228),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_218),
.A2(n_219),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_221),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_225),
.A2(n_226),
.B1(n_228),
.B2(n_229),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_237),
.B2(n_238),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_233),
.B(n_239),
.C(n_240),
.Y(n_287)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_279),
.B(n_284),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_259),
.B(n_278),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_251),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_244),
.B(n_251),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_249),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_245),
.A2(n_246),
.B1(n_249),
.B2(n_266),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_249),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_257),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_256),
.C(n_257),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_258),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_267),
.B(n_277),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_265),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_261),
.B(n_265),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_272),
.B(n_276),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_269),
.B(n_270),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_280),
.B(n_281),
.Y(n_284)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_287),
.B(n_288),
.Y(n_292)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_289),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_295),
.B(n_296),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_305),
.B2(n_306),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_301),
.B2(n_302),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_302),
.C(n_306),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_305),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_309),
.B(n_310),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_325),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_316),
.B(n_325),
.Y(n_334)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_319),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_323),
.A2(n_324),
.B1(n_330),
.B2(n_331),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_328),
.B(n_329),
.Y(n_333)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);


endmodule