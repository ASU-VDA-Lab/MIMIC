module fake_netlist_6_2889_n_1789 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1789);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1789;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_738;
wire n_189;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_122),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_91),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_51),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_138),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_15),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_41),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_5),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_89),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_87),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_83),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_28),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_71),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_17),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_49),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_53),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_22),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_11),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_20),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_64),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_51),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_133),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_65),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_46),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_121),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_98),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_96),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_17),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_146),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_6),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_28),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_26),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_72),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_136),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_50),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_110),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_63),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_41),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_115),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_117),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_56),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_38),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_103),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_49),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_130),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_128),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_18),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_15),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_39),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_19),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_4),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_73),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_139),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_132),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_23),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_151),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_88),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_134),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_38),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_32),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_119),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_35),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_62),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_40),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_34),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_23),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_45),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_106),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_47),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_126),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_60),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_107),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_34),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_104),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_77),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_59),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_21),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_69),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_36),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_111),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_48),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_66),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_0),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_58),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_10),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_21),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_112),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_57),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_79),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_45),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_14),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_12),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_36),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_154),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_70),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_95),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_114),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_109),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_39),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_6),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_44),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_40),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_155),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_80),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_105),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_24),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_13),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_92),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_12),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_26),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_24),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_152),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_149),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_68),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_46),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_76),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_148),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_116),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_124),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_7),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_75),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_100),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_30),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_113),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_43),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_125),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_129),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_118),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_85),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_101),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_43),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_84),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_81),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_123),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_22),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_32),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_10),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_3),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_150),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_50),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_29),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_127),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_143),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_30),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_1),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_35),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_14),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_52),
.Y(n_307)
);

BUFx10_ASAP7_75t_L g308 ( 
.A(n_16),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_82),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_208),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_240),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_289),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_203),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_240),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_225),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_188),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_217),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_197),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_290),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_157),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_201),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_290),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_209),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_214),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_223),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_236),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_238),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_245),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_259),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_260),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_268),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_269),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_188),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_157),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_274),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_177),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_282),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_295),
.Y(n_338)
);

INVxp33_ASAP7_75t_SL g339 ( 
.A(n_158),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_300),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_206),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_304),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_183),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_187),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_195),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_207),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_210),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_158),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_229),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_187),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_306),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_235),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_235),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_162),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_165),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_221),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_224),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_163),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_254),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_237),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_166),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_175),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_176),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_237),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_184),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_199),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_169),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_264),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_308),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_205),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_277),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_228),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_213),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_163),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_218),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g376 ( 
.A(n_301),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_218),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_244),
.Y(n_378)
);

BUFx10_ASAP7_75t_L g379 ( 
.A(n_256),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_220),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_230),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_231),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_239),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_222),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_360),
.B(n_256),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_316),
.Y(n_386)
);

INVx6_ASAP7_75t_L g387 ( 
.A(n_316),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_316),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_316),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_310),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_310),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_384),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_316),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_379),
.B(n_237),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_333),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_333),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_364),
.B(n_156),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_336),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_351),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_343),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_351),
.Y(n_401)
);

BUFx12f_ASAP7_75t_L g402 ( 
.A(n_313),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_323),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_345),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_323),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_324),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_352),
.B(n_283),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_333),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_324),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_379),
.B(n_283),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_353),
.B(n_283),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_320),
.B(n_179),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_325),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_354),
.B(n_355),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_333),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_383),
.B(n_179),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_333),
.Y(n_417)
);

AND2x2_ASAP7_75t_SL g418 ( 
.A(n_370),
.B(n_233),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_379),
.B(n_308),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_382),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_349),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_361),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_362),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_367),
.A2(n_173),
.B1(n_226),
.B2(n_242),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_325),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_326),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_381),
.B(n_233),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_348),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_363),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_317),
.B(n_339),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_326),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_334),
.B(n_219),
.Y(n_432)
);

INVx6_ASAP7_75t_L g433 ( 
.A(n_380),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_327),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_344),
.B(n_219),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_318),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_365),
.Y(n_437)
);

OR2x6_ASAP7_75t_L g438 ( 
.A(n_340),
.B(n_193),
.Y(n_438)
);

NOR2x1_ASAP7_75t_L g439 ( 
.A(n_366),
.B(n_241),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_373),
.B(n_156),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_327),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_328),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_313),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_328),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_329),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_329),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_330),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_350),
.B(n_159),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_330),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_311),
.B(n_159),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_331),
.Y(n_451)
);

INVx6_ASAP7_75t_L g452 ( 
.A(n_376),
.Y(n_452)
);

AND2x6_ASAP7_75t_L g453 ( 
.A(n_311),
.B(n_188),
.Y(n_453)
);

OR2x6_ASAP7_75t_L g454 ( 
.A(n_438),
.B(n_278),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_392),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_388),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_422),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_441),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_441),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_441),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_397),
.B(n_318),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_428),
.Y(n_462)
);

NAND2xp33_ASAP7_75t_L g463 ( 
.A(n_397),
.B(n_378),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_441),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_418),
.B(n_321),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_422),
.Y(n_466)
);

INVx8_ASAP7_75t_L g467 ( 
.A(n_453),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_412),
.B(n_312),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_441),
.Y(n_469)
);

BUFx8_ASAP7_75t_SL g470 ( 
.A(n_402),
.Y(n_470)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_444),
.Y(n_471)
);

NAND3xp33_ASAP7_75t_L g472 ( 
.A(n_412),
.B(n_342),
.C(n_315),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_398),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_422),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_444),
.Y(n_475)
);

NAND3xp33_ASAP7_75t_L g476 ( 
.A(n_412),
.B(n_314),
.C(n_331),
.Y(n_476)
);

NOR3xp33_ASAP7_75t_L g477 ( 
.A(n_424),
.B(n_369),
.C(n_341),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_422),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_444),
.Y(n_479)
);

NAND2xp33_ASAP7_75t_L g480 ( 
.A(n_448),
.B(n_378),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_418),
.A2(n_430),
.B1(n_448),
.B2(n_438),
.Y(n_481)
);

INVx8_ASAP7_75t_L g482 ( 
.A(n_453),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_422),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_444),
.Y(n_484)
);

AND2x6_ASAP7_75t_L g485 ( 
.A(n_432),
.B(n_188),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_444),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_388),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_423),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_444),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_444),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_418),
.B(n_321),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_445),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_445),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_445),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_418),
.B(n_341),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_445),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_445),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_445),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_388),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_388),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_445),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_388),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_430),
.B(n_346),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_428),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_446),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_385),
.B(n_346),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_446),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_419),
.Y(n_508)
);

OAI22xp33_ASAP7_75t_L g509 ( 
.A1(n_438),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_446),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_446),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_385),
.B(n_347),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_446),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_446),
.Y(n_514)
);

OAI21xp33_ASAP7_75t_SL g515 ( 
.A1(n_394),
.A2(n_322),
.B(n_319),
.Y(n_515)
);

NAND3xp33_ASAP7_75t_L g516 ( 
.A(n_432),
.B(n_335),
.C(n_332),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_432),
.B(n_319),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_435),
.B(n_347),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_435),
.B(n_322),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_446),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_420),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_435),
.B(n_358),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_394),
.B(n_356),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_388),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_388),
.Y(n_525)
);

NAND2xp33_ASAP7_75t_SL g526 ( 
.A(n_419),
.B(n_356),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_408),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_386),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_386),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_386),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_408),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_436),
.B(n_357),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_416),
.A2(n_188),
.B1(n_204),
.B2(n_332),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_408),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_420),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_443),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_420),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_408),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_408),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_410),
.B(n_357),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_410),
.B(n_372),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_453),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_398),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_400),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_416),
.A2(n_204),
.B1(n_335),
.B2(n_337),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_389),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_389),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_438),
.A2(n_372),
.B1(n_433),
.B2(n_440),
.Y(n_548)
);

AO21x2_ASAP7_75t_L g549 ( 
.A1(n_450),
.A2(n_262),
.B(n_246),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_408),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_389),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_395),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_395),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_443),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_395),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_396),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_429),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_440),
.B(n_359),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_423),
.Y(n_559)
);

INVx11_ASAP7_75t_L g560 ( 
.A(n_402),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_429),
.Y(n_561)
);

NAND2xp33_ASAP7_75t_L g562 ( 
.A(n_450),
.B(n_204),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_408),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_423),
.B(n_164),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_429),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_437),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_396),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_407),
.B(n_255),
.Y(n_568)
);

OAI22xp33_ASAP7_75t_L g569 ( 
.A1(n_438),
.A2(n_252),
.B1(n_232),
.B2(n_305),
.Y(n_569)
);

INVx5_ASAP7_75t_L g570 ( 
.A(n_453),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_437),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_407),
.B(n_271),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_433),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_438),
.B(n_368),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_433),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_392),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_407),
.B(n_286),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_437),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_451),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_411),
.B(n_196),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_451),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_451),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_403),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_400),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_452),
.B(n_371),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_453),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_396),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_417),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_452),
.B(n_358),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_403),
.Y(n_590)
);

INVxp67_ASAP7_75t_SL g591 ( 
.A(n_393),
.Y(n_591)
);

NAND2xp33_ASAP7_75t_L g592 ( 
.A(n_439),
.B(n_204),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_433),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_417),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_405),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_405),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_393),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_404),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_417),
.Y(n_599)
);

CKINVDCx6p67_ASAP7_75t_R g600 ( 
.A(n_402),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_424),
.A2(n_194),
.B1(n_186),
.B2(n_294),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_416),
.B(n_164),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_583),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_583),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_506),
.B(n_461),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_522),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_481),
.B(n_416),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_503),
.B(n_433),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_590),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_458),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_590),
.B(n_411),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_522),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_459),
.Y(n_613)
);

OR2x6_ASAP7_75t_L g614 ( 
.A(n_576),
.B(n_433),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_508),
.B(n_416),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_459),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_512),
.B(n_427),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_512),
.B(n_427),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_549),
.A2(n_411),
.B1(n_427),
.B2(n_299),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_517),
.Y(n_620)
);

AND2x6_ASAP7_75t_L g621 ( 
.A(n_457),
.B(n_267),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_460),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_465),
.A2(n_495),
.B1(n_491),
.B2(n_558),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_518),
.B(n_452),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_595),
.B(n_427),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_473),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_462),
.Y(n_627)
);

AND2x6_ASAP7_75t_L g628 ( 
.A(n_457),
.B(n_273),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_468),
.B(n_452),
.Y(n_629)
);

NOR2xp67_ASAP7_75t_L g630 ( 
.A(n_536),
.B(n_404),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_595),
.B(n_427),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_596),
.B(n_393),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_463),
.A2(n_480),
.B1(n_548),
.B2(n_526),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_542),
.B(n_276),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_462),
.B(n_421),
.Y(n_635)
);

NOR2xp67_ASAP7_75t_SL g636 ( 
.A(n_570),
.B(n_452),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_542),
.B(n_280),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_596),
.B(n_393),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_517),
.B(n_393),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_460),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_519),
.B(n_415),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_519),
.B(n_421),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_589),
.A2(n_452),
.B1(n_200),
.B2(n_198),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_504),
.B(n_406),
.Y(n_644)
);

BUFx5_ASAP7_75t_L g645 ( 
.A(n_466),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_464),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_549),
.A2(n_302),
.B1(n_307),
.B2(n_298),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_542),
.B(n_287),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_543),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_464),
.Y(n_650)
);

INVx8_ASAP7_75t_L g651 ( 
.A(n_454),
.Y(n_651)
);

CKINVDCx12_ASAP7_75t_R g652 ( 
.A(n_454),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_523),
.A2(n_541),
.B1(n_540),
.B2(n_568),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_554),
.B(n_414),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_572),
.B(n_577),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_469),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_488),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_580),
.B(n_414),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_515),
.A2(n_234),
.B1(n_309),
.B2(n_248),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_591),
.B(n_415),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_469),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_542),
.B(n_288),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_544),
.B(n_406),
.Y(n_663)
);

AO22x2_ASAP7_75t_L g664 ( 
.A1(n_477),
.A2(n_472),
.B1(n_601),
.B2(n_516),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_515),
.A2(n_202),
.B1(n_211),
.B2(n_212),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_488),
.B(n_168),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_488),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_485),
.B(n_415),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_559),
.B(n_168),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_559),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_485),
.B(n_415),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_SL g672 ( 
.A(n_600),
.B(n_171),
.Y(n_672)
);

A2O1A1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_516),
.A2(n_425),
.B(n_449),
.C(n_447),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_521),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_521),
.Y(n_675)
);

INVxp67_ASAP7_75t_L g676 ( 
.A(n_472),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_535),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_485),
.B(n_415),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_474),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_SL g680 ( 
.A1(n_455),
.A2(n_584),
.B1(n_598),
.B2(n_574),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_485),
.B(n_291),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_535),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_559),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_537),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_485),
.B(n_549),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_509),
.B(n_171),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_474),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_537),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_557),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_557),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_585),
.B(n_409),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_478),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_532),
.B(n_409),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_569),
.B(n_180),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_561),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_485),
.B(n_292),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_478),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_454),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_602),
.B(n_180),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_597),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_483),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_576),
.B(n_413),
.Y(n_702)
);

OR2x6_ASAP7_75t_L g703 ( 
.A(n_573),
.B(n_374),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_586),
.B(n_215),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_485),
.B(n_413),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_564),
.B(n_182),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_586),
.B(n_483),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_573),
.A2(n_275),
.B1(n_185),
.B2(n_192),
.Y(n_708)
);

INVx1_ASAP7_75t_SL g709 ( 
.A(n_584),
.Y(n_709)
);

OAI221xp5_ASAP7_75t_L g710 ( 
.A1(n_476),
.A2(n_434),
.B1(n_449),
.B2(n_447),
.C(n_442),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_586),
.B(n_216),
.Y(n_711)
);

NAND2xp33_ASAP7_75t_L g712 ( 
.A(n_575),
.B(n_227),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_561),
.Y(n_713)
);

BUFx5_ASAP7_75t_L g714 ( 
.A(n_484),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_597),
.B(n_565),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_597),
.B(n_425),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_565),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_467),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_566),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_586),
.B(n_243),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_566),
.B(n_426),
.Y(n_721)
);

INVx4_ASAP7_75t_L g722 ( 
.A(n_467),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_571),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_575),
.A2(n_247),
.B1(n_192),
.B2(n_182),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_571),
.Y(n_725)
);

NAND3xp33_ASAP7_75t_L g726 ( 
.A(n_476),
.B(n_281),
.C(n_185),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_578),
.B(n_426),
.Y(n_727)
);

AND2x4_ASAP7_75t_SL g728 ( 
.A(n_600),
.B(n_593),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_467),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_578),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_579),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_455),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_598),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_579),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_560),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_581),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_593),
.B(n_431),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_454),
.B(n_253),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_581),
.B(n_431),
.Y(n_739)
);

NOR2xp67_ASAP7_75t_L g740 ( 
.A(n_582),
.B(n_434),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_582),
.Y(n_741)
);

INVx3_ASAP7_75t_R g742 ( 
.A(n_470),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_531),
.B(n_442),
.Y(n_743)
);

NAND2x1p5_ASAP7_75t_L g744 ( 
.A(n_570),
.B(n_390),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_560),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_528),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_528),
.Y(n_747)
);

OAI21xp33_ASAP7_75t_L g748 ( 
.A1(n_601),
.A2(n_375),
.B(n_377),
.Y(n_748)
);

AND2x6_ASAP7_75t_L g749 ( 
.A(n_475),
.B(n_374),
.Y(n_749)
);

NAND3xp33_ASAP7_75t_L g750 ( 
.A(n_562),
.B(n_293),
.C(n_285),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_529),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_475),
.B(n_253),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_531),
.B(n_390),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_531),
.B(n_391),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_531),
.B(n_391),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_479),
.B(n_257),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_479),
.B(n_257),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_534),
.B(n_399),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_534),
.B(n_399),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_529),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_530),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_454),
.Y(n_762)
);

BUFx5_ASAP7_75t_L g763 ( 
.A(n_484),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_530),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_545),
.B(n_375),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_546),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_546),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_547),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_492),
.B(n_263),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_492),
.B(n_272),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_533),
.B(n_377),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_605),
.B(n_534),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_623),
.B(n_493),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_718),
.B(n_729),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_658),
.B(n_655),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_658),
.B(n_534),
.Y(n_776)
);

A2O1A1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_676),
.A2(n_337),
.B(n_338),
.C(n_305),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_627),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_642),
.B(n_308),
.Y(n_779)
);

NOR2x2_ASAP7_75t_L g780 ( 
.A(n_614),
.B(n_547),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_653),
.A2(n_505),
.B1(n_520),
.B2(n_513),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_691),
.B(n_538),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_676),
.B(n_486),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_629),
.B(n_538),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_629),
.B(n_538),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_679),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_687),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_692),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_624),
.B(n_538),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_610),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_613),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_607),
.A2(n_592),
.B1(n_261),
.B2(n_303),
.Y(n_792)
);

INVxp33_ASAP7_75t_L g793 ( 
.A(n_635),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_624),
.B(n_550),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_616),
.Y(n_795)
);

INVxp67_ASAP7_75t_L g796 ( 
.A(n_663),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_654),
.B(n_486),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_603),
.B(n_550),
.Y(n_798)
);

NAND2x1p5_ASAP7_75t_L g799 ( 
.A(n_718),
.B(n_570),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_626),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_702),
.Y(n_801)
);

CKINVDCx20_ASAP7_75t_R g802 ( 
.A(n_626),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_622),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_640),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_646),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_718),
.B(n_493),
.Y(n_806)
);

HB1xp67_ASAP7_75t_L g807 ( 
.A(n_606),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_604),
.B(n_550),
.Y(n_808)
);

AND2x6_ASAP7_75t_SL g809 ( 
.A(n_694),
.B(n_338),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_609),
.B(n_550),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_650),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_697),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_737),
.B(n_456),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_701),
.Y(n_814)
);

AND2x4_ASAP7_75t_SL g815 ( 
.A(n_614),
.B(n_497),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_656),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_718),
.B(n_497),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_661),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_611),
.B(n_608),
.Y(n_819)
);

HB1xp67_ASAP7_75t_L g820 ( 
.A(n_612),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_620),
.B(n_456),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_644),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_728),
.B(n_401),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_670),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_617),
.B(n_456),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_617),
.A2(n_511),
.B1(n_513),
.B2(n_489),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_713),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_618),
.B(n_489),
.Y(n_828)
);

OR2x2_ASAP7_75t_SL g829 ( 
.A(n_698),
.B(n_160),
.Y(n_829)
);

OR2x2_ASAP7_75t_L g830 ( 
.A(n_709),
.B(n_160),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_693),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_762),
.B(n_401),
.Y(n_832)
);

INVx4_ASAP7_75t_L g833 ( 
.A(n_729),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_618),
.B(n_499),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_698),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_745),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_717),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_639),
.B(n_499),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_641),
.B(n_499),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_633),
.A2(n_510),
.B1(n_511),
.B2(n_490),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_722),
.A2(n_467),
.B(n_482),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_733),
.B(n_161),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_670),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_615),
.A2(n_510),
.B1(n_520),
.B2(n_490),
.Y(n_844)
);

INVx4_ASAP7_75t_L g845 ( 
.A(n_729),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_647),
.B(n_500),
.Y(n_846)
);

INVx5_ASAP7_75t_L g847 ( 
.A(n_729),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_670),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_694),
.B(n_494),
.Y(n_849)
);

OR2x2_ASAP7_75t_L g850 ( 
.A(n_649),
.B(n_161),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_SL g851 ( 
.A1(n_732),
.A2(n_178),
.B1(n_167),
.B2(n_170),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_686),
.B(n_494),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_647),
.B(n_500),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_657),
.B(n_667),
.Y(n_854)
);

NOR3xp33_ASAP7_75t_SL g855 ( 
.A(n_686),
.B(n_174),
.C(n_167),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_670),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_683),
.B(n_500),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_700),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_645),
.B(n_498),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_762),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_645),
.B(n_498),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_719),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_730),
.Y(n_863)
);

NAND3xp33_ASAP7_75t_SL g864 ( 
.A(n_706),
.B(n_174),
.C(n_170),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_614),
.B(n_501),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_651),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_645),
.B(n_501),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_734),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_615),
.B(n_502),
.Y(n_869)
);

AND2x6_ASAP7_75t_L g870 ( 
.A(n_685),
.B(n_507),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_673),
.B(n_502),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_722),
.A2(n_467),
.B(n_482),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_673),
.B(n_502),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_703),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_732),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_666),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_746),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_666),
.B(n_524),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_645),
.B(n_507),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_645),
.B(n_514),
.Y(n_880)
);

INVx4_ASAP7_75t_L g881 ( 
.A(n_651),
.Y(n_881)
);

NOR2x2_ASAP7_75t_L g882 ( 
.A(n_703),
.B(n_551),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_699),
.B(n_505),
.Y(n_883)
);

BUFx4f_ASAP7_75t_L g884 ( 
.A(n_735),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_736),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_699),
.B(n_471),
.Y(n_886)
);

AND3x2_ASAP7_75t_SL g887 ( 
.A(n_664),
.B(n_172),
.C(n_178),
.Y(n_887)
);

AND2x6_ASAP7_75t_L g888 ( 
.A(n_771),
.B(n_514),
.Y(n_888)
);

CKINVDCx6p67_ASAP7_75t_R g889 ( 
.A(n_652),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_645),
.B(n_714),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_749),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_743),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_716),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_714),
.B(n_570),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_703),
.B(n_551),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_669),
.B(n_524),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_714),
.B(n_570),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_706),
.B(n_471),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_765),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_669),
.B(n_524),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_714),
.B(n_763),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_625),
.B(n_631),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_674),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_675),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_751),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_749),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_726),
.B(n_630),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_749),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_707),
.A2(n_482),
.B(n_471),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_760),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_664),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_677),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_619),
.B(n_527),
.Y(n_913)
);

AO22x1_ASAP7_75t_L g914 ( 
.A1(n_738),
.A2(n_297),
.B1(n_181),
.B2(n_189),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_664),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_682),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_738),
.B(n_471),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_684),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_688),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_619),
.B(n_527),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_761),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_740),
.B(n_527),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_752),
.B(n_552),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_749),
.Y(n_924)
);

BUFx8_ASAP7_75t_L g925 ( 
.A(n_742),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_689),
.Y(n_926)
);

NAND3xp33_ASAP7_75t_SL g927 ( 
.A(n_672),
.B(n_172),
.C(n_181),
.Y(n_927)
);

NAND2xp33_ASAP7_75t_SL g928 ( 
.A(n_708),
.B(n_281),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_690),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_680),
.B(n_189),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_651),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_748),
.B(n_190),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_764),
.Y(n_933)
);

INVx4_ASAP7_75t_L g934 ( 
.A(n_714),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_714),
.B(n_570),
.Y(n_935)
);

NOR2xp67_ASAP7_75t_L g936 ( 
.A(n_710),
.B(n_552),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_724),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_721),
.B(n_727),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_659),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_739),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_695),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_763),
.B(n_563),
.Y(n_942)
);

INVx4_ASAP7_75t_L g943 ( 
.A(n_763),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_763),
.B(n_563),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_607),
.A2(n_303),
.B(n_191),
.C(n_258),
.Y(n_945)
);

AND2x6_ASAP7_75t_SL g946 ( 
.A(n_681),
.B(n_190),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_752),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_723),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_621),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_725),
.Y(n_950)
);

INVxp67_ASAP7_75t_L g951 ( 
.A(n_756),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_731),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_768),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_763),
.B(n_496),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_763),
.B(n_563),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_741),
.B(n_553),
.Y(n_956)
);

INVx8_ASAP7_75t_L g957 ( 
.A(n_621),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_747),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_775),
.A2(n_665),
.B(n_705),
.C(n_648),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_822),
.B(n_756),
.Y(n_960)
);

BUFx12f_ASAP7_75t_L g961 ( 
.A(n_925),
.Y(n_961)
);

CKINVDCx20_ASAP7_75t_R g962 ( 
.A(n_802),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_822),
.B(n_757),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_940),
.B(n_757),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_940),
.B(n_769),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_902),
.A2(n_648),
.B(n_662),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_938),
.B(n_769),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_819),
.A2(n_637),
.B(n_662),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_938),
.B(n_770),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_827),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_846),
.A2(n_711),
.B(n_704),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_934),
.A2(n_637),
.B(n_634),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_876),
.B(n_770),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_SL g974 ( 
.A1(n_875),
.A2(n_270),
.B1(n_258),
.B2(n_261),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_945),
.A2(n_696),
.B(n_638),
.C(n_632),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_958),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_876),
.B(n_715),
.Y(n_977)
);

INVxp67_ASAP7_75t_SL g978 ( 
.A(n_824),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_866),
.Y(n_979)
);

INVxp67_ASAP7_75t_L g980 ( 
.A(n_801),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_934),
.A2(n_634),
.B(n_711),
.Y(n_981)
);

O2A1O1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_945),
.A2(n_754),
.B(n_753),
.C(n_755),
.Y(n_982)
);

OAI21x1_ASAP7_75t_L g983 ( 
.A1(n_942),
.A2(n_759),
.B(n_758),
.Y(n_983)
);

NAND2x1p5_ASAP7_75t_L g984 ( 
.A(n_847),
.B(n_707),
.Y(n_984)
);

BUFx8_ASAP7_75t_L g985 ( 
.A(n_778),
.Y(n_985)
);

BUFx6f_ASAP7_75t_SL g986 ( 
.A(n_907),
.Y(n_986)
);

AOI22x1_ASAP7_75t_L g987 ( 
.A1(n_892),
.A2(n_767),
.B1(n_766),
.B2(n_556),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_853),
.A2(n_720),
.B(n_660),
.Y(n_988)
);

INVx1_ASAP7_75t_SL g989 ( 
.A(n_800),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_793),
.B(n_643),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_796),
.B(n_191),
.Y(n_991)
);

CKINVDCx16_ASAP7_75t_R g992 ( 
.A(n_931),
.Y(n_992)
);

INVx2_ASAP7_75t_SL g993 ( 
.A(n_850),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_797),
.B(n_621),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_837),
.Y(n_995)
);

AOI21x1_ASAP7_75t_L g996 ( 
.A1(n_773),
.A2(n_668),
.B(n_671),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_793),
.B(n_712),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_797),
.B(n_621),
.Y(n_998)
);

NAND2xp33_ASAP7_75t_SL g999 ( 
.A(n_939),
.B(n_636),
.Y(n_999)
);

AND2x4_ASAP7_75t_SL g1000 ( 
.A(n_881),
.B(n_487),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_790),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_943),
.A2(n_496),
.B(n_678),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_943),
.A2(n_496),
.B(n_482),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_866),
.Y(n_1004)
);

INVx4_ASAP7_75t_L g1005 ( 
.A(n_866),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_784),
.A2(n_496),
.B(n_482),
.Y(n_1006)
);

INVx1_ASAP7_75t_SL g1007 ( 
.A(n_801),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_842),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_881),
.B(n_621),
.Y(n_1009)
);

OA21x2_ASAP7_75t_L g1010 ( 
.A1(n_789),
.A2(n_587),
.B(n_553),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_835),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_785),
.A2(n_794),
.B(n_776),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_852),
.A2(n_750),
.B1(n_744),
.B2(n_285),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_862),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_852),
.B(n_628),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_791),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_796),
.B(n_265),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_947),
.A2(n_951),
.B(n_849),
.C(n_883),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_SL g1019 ( 
.A1(n_898),
.A2(n_556),
.B(n_555),
.C(n_599),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_863),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_835),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_866),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_831),
.B(n_265),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_849),
.B(n_628),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_807),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_944),
.A2(n_744),
.B(n_587),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_878),
.A2(n_487),
.B(n_525),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_907),
.A2(n_628),
.B1(n_293),
.B2(n_594),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_SL g1029 ( 
.A1(n_898),
.A2(n_555),
.B(n_599),
.C(n_594),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_893),
.B(n_628),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_779),
.B(n_296),
.Y(n_1031)
);

HB1xp67_ASAP7_75t_L g1032 ( 
.A(n_807),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_832),
.B(n_628),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_868),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_899),
.B(n_539),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_915),
.A2(n_588),
.B(n_567),
.C(n_297),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_937),
.B(n_296),
.Y(n_1037)
);

O2A1O1Ixp5_ASAP7_75t_L g1038 ( 
.A1(n_773),
.A2(n_588),
.B(n_567),
.C(n_453),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_896),
.A2(n_539),
.B(n_525),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_951),
.A2(n_284),
.B(n_279),
.C(n_270),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_847),
.B(n_539),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_824),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_824),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_847),
.B(n_539),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_925),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_915),
.A2(n_266),
.B(n_279),
.C(n_284),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_882),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_911),
.A2(n_539),
.B1(n_525),
.B2(n_487),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_885),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_883),
.A2(n_266),
.B(n_525),
.C(n_487),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_847),
.B(n_525),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_795),
.Y(n_1052)
);

AOI221xp5_ASAP7_75t_L g1053 ( 
.A1(n_914),
.A2(n_864),
.B1(n_851),
.B2(n_930),
.C(n_932),
.Y(n_1053)
);

NOR2x1_ASAP7_75t_L g1054 ( 
.A(n_848),
.B(n_487),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_830),
.B(n_0),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_820),
.B(n_153),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_886),
.B(n_453),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_886),
.B(n_453),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_803),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_900),
.A2(n_387),
.B(n_453),
.Y(n_1060)
);

CKINVDCx20_ASAP7_75t_R g1061 ( 
.A(n_836),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_890),
.A2(n_387),
.B(n_453),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_804),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_805),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_890),
.A2(n_387),
.B(n_147),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_874),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_860),
.B(n_1),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_820),
.B(n_142),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_824),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_901),
.A2(n_387),
.B(n_141),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_889),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_832),
.B(n_135),
.Y(n_1072)
);

NOR3xp33_ASAP7_75t_SL g1073 ( 
.A(n_927),
.B(n_2),
.C(n_3),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_786),
.Y(n_1074)
);

INVx3_ASAP7_75t_L g1075 ( 
.A(n_843),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_860),
.Y(n_1076)
);

BUFx2_ASAP7_75t_L g1077 ( 
.A(n_874),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_917),
.A2(n_387),
.B1(n_131),
.B2(n_108),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_792),
.A2(n_387),
.B1(n_4),
.B2(n_5),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_783),
.B(n_917),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_787),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_783),
.B(n_2),
.Y(n_1082)
);

O2A1O1Ixp5_ASAP7_75t_L g1083 ( 
.A1(n_871),
.A2(n_102),
.B(n_99),
.C(n_97),
.Y(n_1083)
);

OAI22x1_ASAP7_75t_L g1084 ( 
.A1(n_887),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_811),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_855),
.B(n_8),
.Y(n_1086)
);

OAI33xp33_ASAP7_75t_L g1087 ( 
.A1(n_788),
.A2(n_9),
.A3(n_11),
.B1(n_13),
.B2(n_16),
.B3(n_18),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_828),
.A2(n_19),
.B(n_20),
.C(n_25),
.Y(n_1088)
);

AND2x6_ASAP7_75t_L g1089 ( 
.A(n_949),
.B(n_54),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_901),
.A2(n_78),
.B(n_93),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_809),
.B(n_25),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_777),
.A2(n_772),
.B(n_913),
.C(n_920),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_777),
.A2(n_27),
.B(n_29),
.C(n_31),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_816),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_855),
.B(n_27),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_843),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_818),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_812),
.Y(n_1098)
);

INVx4_ASAP7_75t_L g1099 ( 
.A(n_843),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_865),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_814),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_828),
.A2(n_31),
.B(n_33),
.C(n_37),
.Y(n_1102)
);

INVx2_ASAP7_75t_SL g1103 ( 
.A(n_823),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_865),
.B(n_55),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_877),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_SL g1106 ( 
.A1(n_873),
.A2(n_61),
.B(n_90),
.C(n_86),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_843),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1080),
.B(n_792),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_1026),
.A2(n_806),
.B(n_817),
.Y(n_1109)
);

O2A1O1Ixp5_ASAP7_75t_SL g1110 ( 
.A1(n_1082),
.A2(n_916),
.B(n_926),
.C(n_912),
.Y(n_1110)
);

AO21x2_ASAP7_75t_L g1111 ( 
.A1(n_1012),
.A2(n_840),
.B(n_806),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_985),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1055),
.A2(n_928),
.B1(n_888),
.B2(n_952),
.Y(n_1113)
);

BUFx10_ASAP7_75t_L g1114 ( 
.A(n_986),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_967),
.B(n_782),
.Y(n_1115)
);

CKINVDCx8_ASAP7_75t_R g1116 ( 
.A(n_992),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1031),
.B(n_823),
.Y(n_1117)
);

AO31x2_ASAP7_75t_L g1118 ( 
.A1(n_1012),
.A2(n_838),
.A3(n_839),
.B(n_834),
.Y(n_1118)
);

O2A1O1Ixp5_ASAP7_75t_L g1119 ( 
.A1(n_1015),
.A2(n_774),
.B(n_817),
.C(n_954),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_1061),
.Y(n_1120)
);

NOR2xp67_ASAP7_75t_L g1121 ( 
.A(n_1008),
.B(n_848),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_985),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_970),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_1027),
.A2(n_774),
.B(n_880),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_995),
.Y(n_1125)
);

AOI21x1_ASAP7_75t_SL g1126 ( 
.A1(n_1024),
.A2(n_854),
.B(n_922),
.Y(n_1126)
);

OA21x2_ASAP7_75t_L g1127 ( 
.A1(n_971),
.A2(n_781),
.B(n_810),
.Y(n_1127)
);

AO31x2_ASAP7_75t_L g1128 ( 
.A1(n_1050),
.A2(n_825),
.A3(n_955),
.B(n_869),
.Y(n_1128)
);

NAND2x1p5_ASAP7_75t_L g1129 ( 
.A(n_1005),
.B(n_833),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_1018),
.A2(n_948),
.B(n_903),
.C(n_919),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1027),
.A2(n_879),
.B(n_859),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_966),
.A2(n_872),
.B(n_841),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1014),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_SL g1134 ( 
.A(n_1005),
.B(n_884),
.Y(n_1134)
);

CKINVDCx11_ASAP7_75t_R g1135 ( 
.A(n_961),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_969),
.B(n_904),
.Y(n_1136)
);

HB1xp67_ASAP7_75t_L g1137 ( 
.A(n_1007),
.Y(n_1137)
);

OR2x2_ASAP7_75t_L g1138 ( 
.A(n_993),
.B(n_829),
.Y(n_1138)
);

OAI22x1_ASAP7_75t_L g1139 ( 
.A1(n_1091),
.A2(n_887),
.B1(n_895),
.B2(n_918),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_962),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_1053),
.B(n_884),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_1011),
.Y(n_1142)
);

OAI22x1_ASAP7_75t_L g1143 ( 
.A1(n_1037),
.A2(n_895),
.B1(n_929),
.B2(n_941),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1020),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1034),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_977),
.B(n_950),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_979),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_966),
.A2(n_981),
.B(n_968),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1039),
.A2(n_867),
.B(n_859),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1092),
.A2(n_936),
.B(n_826),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_973),
.B(n_888),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_960),
.B(n_905),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_SL g1153 ( 
.A1(n_1090),
.A2(n_808),
.B(n_798),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1039),
.A2(n_861),
.B(n_867),
.Y(n_1154)
);

OR2x6_ASAP7_75t_L g1155 ( 
.A(n_1072),
.B(n_957),
.Y(n_1155)
);

INVx6_ASAP7_75t_L g1156 ( 
.A(n_1071),
.Y(n_1156)
);

INVx1_ASAP7_75t_SL g1157 ( 
.A(n_1021),
.Y(n_1157)
);

OAI22x1_ASAP7_75t_L g1158 ( 
.A1(n_1067),
.A2(n_780),
.B1(n_858),
.B2(n_923),
.Y(n_1158)
);

CKINVDCx20_ASAP7_75t_R g1159 ( 
.A(n_1045),
.Y(n_1159)
);

INVx1_ASAP7_75t_SL g1160 ( 
.A(n_1025),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1049),
.Y(n_1161)
);

BUFx10_ASAP7_75t_L g1162 ( 
.A(n_986),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1079),
.A2(n_856),
.B1(n_813),
.B2(n_845),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_979),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_981),
.A2(n_954),
.B(n_833),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_990),
.B(n_946),
.Y(n_1166)
);

AO31x2_ASAP7_75t_L g1167 ( 
.A1(n_1006),
.A2(n_956),
.A3(n_857),
.B(n_909),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_963),
.B(n_953),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_972),
.A2(n_799),
.B(n_935),
.Y(n_1169)
);

INVx2_ASAP7_75t_SL g1170 ( 
.A(n_1025),
.Y(n_1170)
);

AND3x2_ASAP7_75t_L g1171 ( 
.A(n_1047),
.B(n_933),
.C(n_921),
.Y(n_1171)
);

INVx1_ASAP7_75t_SL g1172 ( 
.A(n_1032),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_979),
.Y(n_1173)
);

OR2x2_ASAP7_75t_L g1174 ( 
.A(n_964),
.B(n_910),
.Y(n_1174)
);

NAND2x1p5_ASAP7_75t_L g1175 ( 
.A(n_1004),
.B(n_856),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1092),
.A2(n_844),
.B(n_870),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_SL g1177 ( 
.A1(n_959),
.A2(n_1009),
.B(n_994),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_965),
.B(n_888),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_972),
.A2(n_988),
.B(n_1003),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_1032),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_SL g1181 ( 
.A1(n_1090),
.A2(n_821),
.B(n_870),
.Y(n_1181)
);

AOI221x1_ASAP7_75t_L g1182 ( 
.A1(n_1088),
.A2(n_924),
.B1(n_908),
.B2(n_906),
.C(n_856),
.Y(n_1182)
);

AOI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_997),
.A2(n_1086),
.B1(n_1095),
.B2(n_1072),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_1066),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1003),
.A2(n_894),
.B(n_935),
.Y(n_1185)
);

O2A1O1Ixp5_ASAP7_75t_L g1186 ( 
.A1(n_998),
.A2(n_879),
.B(n_861),
.C(n_880),
.Y(n_1186)
);

OA21x2_ASAP7_75t_L g1187 ( 
.A1(n_1038),
.A2(n_897),
.B(n_894),
.Y(n_1187)
);

OR2x6_ASAP7_75t_SL g1188 ( 
.A(n_976),
.B(n_815),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1100),
.B(n_888),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1006),
.A2(n_897),
.B(n_957),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_991),
.B(n_891),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_996),
.A2(n_924),
.B(n_906),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1038),
.A2(n_983),
.B(n_1060),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1100),
.B(n_870),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_980),
.Y(n_1195)
);

NOR2xp67_ASAP7_75t_L g1196 ( 
.A(n_1103),
.B(n_94),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1074),
.B(n_870),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1002),
.A2(n_1057),
.B(n_1058),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1017),
.B(n_1023),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1081),
.B(n_870),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1030),
.A2(n_74),
.B(n_67),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_SL g1202 ( 
.A1(n_1102),
.A2(n_1056),
.B(n_1068),
.C(n_1104),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1098),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1101),
.B(n_33),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_999),
.A2(n_37),
.B(n_42),
.Y(n_1205)
);

AO21x1_ASAP7_75t_L g1206 ( 
.A1(n_1093),
.A2(n_42),
.B(n_44),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_1033),
.B(n_47),
.Y(n_1207)
);

AOI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1060),
.A2(n_48),
.B(n_1010),
.Y(n_1208)
);

AOI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1010),
.A2(n_1070),
.B(n_1065),
.Y(n_1209)
);

NAND2x1p5_ASAP7_75t_L g1210 ( 
.A(n_1004),
.B(n_1022),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1077),
.Y(n_1211)
);

O2A1O1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1040),
.A2(n_1046),
.B(n_1093),
.C(n_980),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1076),
.B(n_1059),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_1076),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1001),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_987),
.A2(n_1062),
.B(n_1065),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1016),
.B(n_1097),
.Y(n_1217)
);

OR2x2_ASAP7_75t_L g1218 ( 
.A(n_989),
.B(n_1064),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_1004),
.Y(n_1219)
);

INVx5_ASAP7_75t_L g1220 ( 
.A(n_1042),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1036),
.A2(n_975),
.B(n_982),
.C(n_1046),
.Y(n_1221)
);

AO21x2_ASAP7_75t_L g1222 ( 
.A1(n_1019),
.A2(n_1029),
.B(n_1070),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1062),
.A2(n_975),
.B(n_982),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1052),
.B(n_1085),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1054),
.A2(n_984),
.B(n_1083),
.Y(n_1225)
);

OA22x2_ASAP7_75t_L g1226 ( 
.A1(n_1084),
.A2(n_974),
.B1(n_1028),
.B2(n_1048),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_978),
.A2(n_984),
.B1(n_1033),
.B2(n_1073),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1063),
.B(n_1105),
.Y(n_1228)
);

INVx4_ASAP7_75t_L g1229 ( 
.A(n_1022),
.Y(n_1229)
);

OA21x2_ASAP7_75t_L g1230 ( 
.A1(n_1083),
.A2(n_1078),
.B(n_1035),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_R g1231 ( 
.A(n_1022),
.B(n_1107),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1094),
.A2(n_1013),
.B1(n_1087),
.B2(n_1089),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_978),
.B(n_1036),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_SL g1234 ( 
.A(n_1089),
.B(n_1087),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1073),
.B(n_1107),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1041),
.A2(n_1044),
.B(n_1051),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1043),
.A2(n_1096),
.B(n_1075),
.Y(n_1237)
);

A2O1A1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1043),
.A2(n_1075),
.B(n_1096),
.C(n_1000),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1042),
.A2(n_1069),
.B1(n_1099),
.B2(n_1089),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1042),
.Y(n_1240)
);

O2A1O1Ixp5_ASAP7_75t_L g1241 ( 
.A1(n_1099),
.A2(n_1106),
.B(n_1089),
.C(n_1069),
.Y(n_1241)
);

AO31x2_ASAP7_75t_L g1242 ( 
.A1(n_1089),
.A2(n_1012),
.A3(n_1050),
.B(n_1018),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1069),
.A2(n_1026),
.B(n_1027),
.Y(n_1243)
);

NAND2x1p5_ASAP7_75t_L g1244 ( 
.A(n_1005),
.B(n_881),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1080),
.B(n_775),
.Y(n_1245)
);

AO31x2_ASAP7_75t_L g1246 ( 
.A1(n_1012),
.A2(n_1050),
.A3(n_1018),
.B(n_1080),
.Y(n_1246)
);

AOI22xp5_ASAP7_75t_SL g1247 ( 
.A1(n_1084),
.A2(n_605),
.B1(n_1091),
.B2(n_1055),
.Y(n_1247)
);

AO31x2_ASAP7_75t_L g1248 ( 
.A1(n_1012),
.A2(n_1050),
.A3(n_1018),
.B(n_1080),
.Y(n_1248)
);

NAND2x1p5_ASAP7_75t_L g1249 ( 
.A(n_1005),
.B(n_881),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1092),
.A2(n_1080),
.B(n_971),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_966),
.A2(n_943),
.B(n_934),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1080),
.A2(n_775),
.B1(n_605),
.B2(n_1018),
.Y(n_1252)
);

BUFx12f_ASAP7_75t_L g1253 ( 
.A(n_961),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1080),
.A2(n_605),
.B(n_775),
.C(n_623),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1243),
.A2(n_1132),
.B(n_1193),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1199),
.B(n_1152),
.Y(n_1256)
);

BUFx2_ASAP7_75t_L g1257 ( 
.A(n_1211),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1216),
.A2(n_1190),
.B(n_1208),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1109),
.A2(n_1223),
.B(n_1209),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1206),
.A2(n_1108),
.B1(n_1226),
.B2(n_1166),
.Y(n_1260)
);

INVxp67_ASAP7_75t_L g1261 ( 
.A(n_1137),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1123),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1148),
.A2(n_1124),
.B(n_1165),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1245),
.B(n_1146),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1125),
.Y(n_1265)
);

BUFx8_ASAP7_75t_L g1266 ( 
.A(n_1253),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1155),
.B(n_1207),
.Y(n_1267)
);

NAND2x1p5_ASAP7_75t_L g1268 ( 
.A(n_1220),
.B(n_1160),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1254),
.A2(n_1252),
.B(n_1221),
.Y(n_1269)
);

AO21x1_ASAP7_75t_L g1270 ( 
.A1(n_1252),
.A2(n_1234),
.B(n_1205),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_1142),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1133),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1168),
.B(n_1183),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1185),
.A2(n_1126),
.B(n_1169),
.Y(n_1274)
);

BUFx12f_ASAP7_75t_L g1275 ( 
.A(n_1135),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_SL g1276 ( 
.A(n_1120),
.B(n_1116),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1136),
.B(n_1117),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1144),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1145),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1161),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_1156),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1141),
.A2(n_1250),
.B1(n_1183),
.B2(n_1139),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1131),
.A2(n_1149),
.B(n_1154),
.Y(n_1283)
);

INVxp67_ASAP7_75t_L g1284 ( 
.A(n_1218),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1203),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1155),
.B(n_1207),
.Y(n_1286)
);

INVx3_ASAP7_75t_L g1287 ( 
.A(n_1237),
.Y(n_1287)
);

AO21x2_ASAP7_75t_L g1288 ( 
.A1(n_1150),
.A2(n_1181),
.B(n_1198),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1174),
.B(n_1191),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1192),
.A2(n_1225),
.B(n_1153),
.Y(n_1290)
);

AO21x2_ASAP7_75t_L g1291 ( 
.A1(n_1222),
.A2(n_1233),
.B(n_1177),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1110),
.A2(n_1119),
.B(n_1113),
.Y(n_1292)
);

AO21x2_ASAP7_75t_L g1293 ( 
.A1(n_1222),
.A2(n_1111),
.B(n_1130),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1234),
.A2(n_1143),
.B1(n_1158),
.B2(n_1115),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1228),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1215),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1228),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1118),
.Y(n_1298)
);

AOI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1155),
.A2(n_1227),
.B1(n_1138),
.B2(n_1202),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1157),
.B(n_1235),
.Y(n_1300)
);

NAND2x1p5_ASAP7_75t_L g1301 ( 
.A(n_1220),
.B(n_1160),
.Y(n_1301)
);

OAI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1113),
.A2(n_1134),
.B1(n_1204),
.B2(n_1188),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1186),
.A2(n_1241),
.B(n_1200),
.Y(n_1303)
);

INVx2_ASAP7_75t_SL g1304 ( 
.A(n_1220),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1197),
.A2(n_1236),
.B(n_1194),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1213),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1201),
.A2(n_1239),
.B(n_1182),
.Y(n_1307)
);

OAI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1115),
.A2(n_1212),
.B(n_1178),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1217),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1239),
.A2(n_1187),
.B(n_1151),
.Y(n_1310)
);

INVx3_ASAP7_75t_L g1311 ( 
.A(n_1242),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1187),
.A2(n_1151),
.B(n_1127),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_SL g1313 ( 
.A1(n_1227),
.A2(n_1232),
.B(n_1189),
.Y(n_1313)
);

AOI222xp33_ASAP7_75t_L g1314 ( 
.A1(n_1172),
.A2(n_1157),
.B1(n_1214),
.B2(n_1180),
.C1(n_1195),
.C2(n_1140),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1240),
.B(n_1238),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1118),
.Y(n_1316)
);

AO31x2_ASAP7_75t_L g1317 ( 
.A1(n_1163),
.A2(n_1167),
.A3(n_1118),
.B(n_1248),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1224),
.Y(n_1318)
);

NAND2x1p5_ASAP7_75t_L g1319 ( 
.A(n_1172),
.B(n_1170),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1219),
.B(n_1121),
.Y(n_1320)
);

O2A1O1Ixp33_ASAP7_75t_SL g1321 ( 
.A1(n_1163),
.A2(n_1247),
.B(n_1184),
.C(n_1242),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1242),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1246),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1247),
.A2(n_1230),
.B1(n_1114),
.B2(n_1162),
.Y(n_1324)
);

AOI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1134),
.A2(n_1196),
.B1(n_1159),
.B2(n_1171),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1244),
.B(n_1249),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1230),
.A2(n_1175),
.B(n_1244),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1175),
.A2(n_1249),
.B(n_1129),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1229),
.B(n_1156),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_SL g1330 ( 
.A1(n_1129),
.A2(n_1210),
.B(n_1164),
.Y(n_1330)
);

AO21x2_ASAP7_75t_L g1331 ( 
.A1(n_1167),
.A2(n_1248),
.B(n_1246),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_1114),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1162),
.A2(n_1112),
.B1(n_1122),
.B2(n_1147),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1147),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1246),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1167),
.A2(n_1128),
.B(n_1248),
.Y(n_1336)
);

OAI221xp5_ASAP7_75t_L g1337 ( 
.A1(n_1164),
.A2(n_605),
.B1(n_503),
.B2(n_1053),
.C(n_558),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1128),
.A2(n_1231),
.B(n_1173),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1173),
.Y(n_1339)
);

INVx2_ASAP7_75t_SL g1340 ( 
.A(n_1173),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1155),
.B(n_866),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1243),
.A2(n_1132),
.B(n_1193),
.Y(n_1342)
);

AND2x4_ASAP7_75t_L g1343 ( 
.A(n_1155),
.B(n_866),
.Y(n_1343)
);

CKINVDCx16_ASAP7_75t_R g1344 ( 
.A(n_1253),
.Y(n_1344)
);

AOI222xp33_ASAP7_75t_L g1345 ( 
.A1(n_1166),
.A2(n_424),
.B1(n_605),
.B2(n_1053),
.C1(n_1091),
.C2(n_1037),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1123),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1123),
.Y(n_1347)
);

AO31x2_ASAP7_75t_L g1348 ( 
.A1(n_1221),
.A2(n_1148),
.A3(n_1179),
.B(n_1182),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1206),
.A2(n_605),
.B1(n_1108),
.B2(n_1079),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1243),
.A2(n_1132),
.B(n_1193),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1254),
.A2(n_605),
.B(n_775),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1123),
.Y(n_1352)
);

BUFx4f_ASAP7_75t_SL g1353 ( 
.A(n_1253),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_1220),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1243),
.A2(n_1132),
.B(n_1193),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1123),
.Y(n_1356)
);

AO21x2_ASAP7_75t_L g1357 ( 
.A1(n_1179),
.A2(n_1148),
.B(n_1176),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1108),
.B(n_915),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1223),
.A2(n_1148),
.B(n_1193),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1243),
.A2(n_1132),
.B(n_1193),
.Y(n_1360)
);

INVx3_ASAP7_75t_SL g1361 ( 
.A(n_1120),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1243),
.A2(n_1132),
.B(n_1193),
.Y(n_1362)
);

O2A1O1Ixp33_ASAP7_75t_L g1363 ( 
.A1(n_1141),
.A2(n_605),
.B(n_503),
.C(n_1221),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_SL g1364 ( 
.A1(n_1206),
.A2(n_1212),
.B(n_1183),
.Y(n_1364)
);

INVx1_ASAP7_75t_SL g1365 ( 
.A(n_1157),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1123),
.Y(n_1366)
);

INVx2_ASAP7_75t_SL g1367 ( 
.A(n_1220),
.Y(n_1367)
);

BUFx3_ASAP7_75t_L g1368 ( 
.A(n_1156),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_SL g1369 ( 
.A1(n_1206),
.A2(n_1212),
.B(n_1183),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1123),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1243),
.A2(n_1132),
.B(n_1193),
.Y(n_1371)
);

OR2x2_ASAP7_75t_L g1372 ( 
.A(n_1157),
.B(n_1174),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1243),
.A2(n_1132),
.B(n_1193),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1243),
.A2(n_1132),
.B(n_1193),
.Y(n_1374)
);

OAI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1254),
.A2(n_605),
.B(n_775),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_1156),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1245),
.B(n_605),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1137),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1243),
.A2(n_1132),
.B(n_1193),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1123),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1243),
.A2(n_1132),
.B(n_1193),
.Y(n_1381)
);

NAND2x1p5_ASAP7_75t_L g1382 ( 
.A(n_1220),
.B(n_1160),
.Y(n_1382)
);

INVx1_ASAP7_75t_SL g1383 ( 
.A(n_1157),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1148),
.A2(n_1179),
.B(n_1251),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1243),
.A2(n_1132),
.B(n_1193),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1123),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1245),
.A2(n_605),
.B1(n_775),
.B2(n_1080),
.Y(n_1387)
);

INVx4_ASAP7_75t_L g1388 ( 
.A(n_1220),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1245),
.B(n_775),
.Y(n_1389)
);

CKINVDCx20_ASAP7_75t_R g1390 ( 
.A(n_1135),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1272),
.Y(n_1391)
);

O2A1O1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1363),
.A2(n_1337),
.B(n_1345),
.C(n_1351),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1260),
.A2(n_1377),
.B1(n_1389),
.B2(n_1264),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1378),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1260),
.A2(n_1377),
.B1(n_1349),
.B2(n_1282),
.Y(n_1395)
);

OA21x2_ASAP7_75t_L g1396 ( 
.A1(n_1292),
.A2(n_1336),
.B(n_1269),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1277),
.B(n_1284),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1349),
.A2(n_1282),
.B1(n_1387),
.B2(n_1300),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1375),
.A2(n_1384),
.B(n_1357),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1300),
.A2(n_1294),
.B1(n_1289),
.B2(n_1333),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1325),
.A2(n_1294),
.B1(n_1299),
.B2(n_1324),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1306),
.B(n_1372),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_1390),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1273),
.B(n_1358),
.Y(n_1404)
);

AOI221xp5_ASAP7_75t_L g1405 ( 
.A1(n_1364),
.A2(n_1369),
.B1(n_1321),
.B2(n_1270),
.C(n_1308),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_SL g1406 ( 
.A1(n_1354),
.A2(n_1388),
.B(n_1326),
.Y(n_1406)
);

O2A1O1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1302),
.A2(n_1321),
.B(n_1261),
.C(n_1324),
.Y(n_1407)
);

AOI21x1_ASAP7_75t_SL g1408 ( 
.A1(n_1315),
.A2(n_1341),
.B(n_1343),
.Y(n_1408)
);

O2A1O1Ixp5_ASAP7_75t_L g1409 ( 
.A1(n_1323),
.A2(n_1335),
.B(n_1322),
.C(n_1311),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1333),
.A2(n_1279),
.B1(n_1280),
.B2(n_1265),
.Y(n_1410)
);

OA21x2_ASAP7_75t_L g1411 ( 
.A1(n_1336),
.A2(n_1259),
.B(n_1274),
.Y(n_1411)
);

O2A1O1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1313),
.A2(n_1314),
.B(n_1365),
.C(n_1383),
.Y(n_1412)
);

INVx5_ASAP7_75t_L g1413 ( 
.A(n_1354),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_SL g1414 ( 
.A1(n_1354),
.A2(n_1388),
.B(n_1326),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1309),
.B(n_1318),
.Y(n_1415)
);

OA21x2_ASAP7_75t_L g1416 ( 
.A1(n_1259),
.A2(n_1274),
.B(n_1258),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1278),
.A2(n_1285),
.B1(n_1267),
.B2(n_1286),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_SL g1418 ( 
.A1(n_1390),
.A2(n_1344),
.B1(n_1361),
.B2(n_1275),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1273),
.B(n_1358),
.Y(n_1419)
);

O2A1O1Ixp5_ASAP7_75t_L g1420 ( 
.A1(n_1323),
.A2(n_1335),
.B(n_1311),
.C(n_1322),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1319),
.A2(n_1271),
.B1(n_1301),
.B2(n_1268),
.Y(n_1421)
);

O2A1O1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1332),
.A2(n_1366),
.B(n_1346),
.C(n_1386),
.Y(n_1422)
);

CKINVDCx16_ASAP7_75t_R g1423 ( 
.A(n_1275),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1295),
.B(n_1297),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1347),
.B(n_1380),
.Y(n_1425)
);

CKINVDCx16_ASAP7_75t_R g1426 ( 
.A(n_1276),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1296),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1262),
.A2(n_1370),
.B1(n_1352),
.B2(n_1356),
.Y(n_1428)
);

INVx3_ASAP7_75t_L g1429 ( 
.A(n_1354),
.Y(n_1429)
);

O2A1O1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1332),
.A2(n_1382),
.B(n_1301),
.C(n_1291),
.Y(n_1430)
);

BUFx6f_ASAP7_75t_L g1431 ( 
.A(n_1281),
.Y(n_1431)
);

O2A1O1Ixp5_ASAP7_75t_L g1432 ( 
.A1(n_1311),
.A2(n_1322),
.B(n_1316),
.C(n_1298),
.Y(n_1432)
);

INVx1_ASAP7_75t_SL g1433 ( 
.A(n_1382),
.Y(n_1433)
);

A2O1A1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1307),
.A2(n_1303),
.B(n_1338),
.C(n_1329),
.Y(n_1434)
);

O2A1O1Ixp5_ASAP7_75t_L g1435 ( 
.A1(n_1298),
.A2(n_1316),
.B(n_1287),
.C(n_1388),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1288),
.A2(n_1263),
.B(n_1293),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1257),
.A2(n_1320),
.B1(n_1361),
.B2(n_1329),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1334),
.B(n_1339),
.Y(n_1438)
);

CKINVDCx20_ASAP7_75t_R g1439 ( 
.A(n_1353),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1348),
.B(n_1305),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1293),
.A2(n_1307),
.B(n_1258),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1348),
.B(n_1305),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1328),
.B(n_1338),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1304),
.A2(n_1367),
.B1(n_1281),
.B2(n_1376),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1340),
.B(n_1348),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1348),
.B(n_1317),
.Y(n_1446)
);

OA21x2_ASAP7_75t_L g1447 ( 
.A1(n_1283),
.A2(n_1255),
.B(n_1385),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1310),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1304),
.B(n_1367),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1368),
.B(n_1376),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1368),
.B(n_1330),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1266),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1331),
.B(n_1317),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1312),
.B(n_1359),
.Y(n_1454)
);

CKINVDCx20_ASAP7_75t_R g1455 ( 
.A(n_1266),
.Y(n_1455)
);

O2A1O1Ixp33_ASAP7_75t_L g1456 ( 
.A1(n_1266),
.A2(n_1290),
.B(n_1327),
.C(n_1342),
.Y(n_1456)
);

OAI221xp5_ASAP7_75t_SL g1457 ( 
.A1(n_1327),
.A2(n_1290),
.B1(n_1342),
.B2(n_1350),
.C(n_1355),
.Y(n_1457)
);

OA21x2_ASAP7_75t_L g1458 ( 
.A1(n_1350),
.A2(n_1355),
.B(n_1360),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1362),
.A2(n_1381),
.B1(n_1373),
.B2(n_1374),
.Y(n_1459)
);

INVx1_ASAP7_75t_SL g1460 ( 
.A(n_1362),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1371),
.A2(n_1373),
.B1(n_1374),
.B2(n_1379),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1371),
.B(n_1379),
.Y(n_1462)
);

AOI21x1_ASAP7_75t_SL g1463 ( 
.A1(n_1381),
.A2(n_605),
.B(n_1086),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1267),
.B(n_1286),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1256),
.B(n_1273),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_SL g1466 ( 
.A1(n_1363),
.A2(n_1254),
.B(n_775),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1267),
.B(n_1286),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1260),
.A2(n_1080),
.B1(n_605),
.B2(n_1377),
.Y(n_1468)
);

NOR2xp67_ASAP7_75t_L g1469 ( 
.A(n_1284),
.B(n_1332),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1377),
.B(n_1264),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1260),
.A2(n_605),
.B1(n_775),
.B2(n_1337),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1256),
.B(n_1273),
.Y(n_1472)
);

A2O1A1Ixp33_ASAP7_75t_L g1473 ( 
.A1(n_1363),
.A2(n_605),
.B(n_1337),
.C(n_775),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1372),
.B(n_1289),
.Y(n_1474)
);

OA21x2_ASAP7_75t_L g1475 ( 
.A1(n_1292),
.A2(n_1336),
.B(n_1269),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1372),
.B(n_1289),
.Y(n_1476)
);

INVx2_ASAP7_75t_SL g1477 ( 
.A(n_1281),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1445),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1391),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1393),
.B(n_1470),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1448),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1443),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1453),
.B(n_1396),
.Y(n_1483)
);

AO21x2_ASAP7_75t_L g1484 ( 
.A1(n_1436),
.A2(n_1399),
.B(n_1441),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1393),
.B(n_1419),
.Y(n_1485)
);

INVx4_ASAP7_75t_L g1486 ( 
.A(n_1413),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1446),
.B(n_1440),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1442),
.B(n_1396),
.Y(n_1488)
);

INVx2_ASAP7_75t_SL g1489 ( 
.A(n_1443),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1424),
.B(n_1402),
.Y(n_1490)
);

INVx1_ASAP7_75t_SL g1491 ( 
.A(n_1433),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1475),
.B(n_1454),
.Y(n_1492)
);

OR2x6_ASAP7_75t_L g1493 ( 
.A(n_1456),
.B(n_1434),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1392),
.B(n_1400),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1411),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1473),
.A2(n_1471),
.B(n_1466),
.Y(n_1496)
);

AOI33xp33_ASAP7_75t_L g1497 ( 
.A1(n_1405),
.A2(n_1412),
.A3(n_1407),
.B1(n_1422),
.B2(n_1477),
.B3(n_1433),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1462),
.B(n_1460),
.Y(n_1498)
);

AO21x2_ASAP7_75t_L g1499 ( 
.A1(n_1459),
.A2(n_1461),
.B(n_1398),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1395),
.A2(n_1398),
.B1(n_1468),
.B2(n_1401),
.Y(n_1500)
);

AO21x2_ASAP7_75t_L g1501 ( 
.A1(n_1459),
.A2(n_1395),
.B(n_1468),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1416),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1404),
.B(n_1416),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1415),
.B(n_1394),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1474),
.B(n_1476),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1409),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1420),
.B(n_1432),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1447),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1465),
.B(n_1472),
.Y(n_1509)
);

OAI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1400),
.A2(n_1426),
.B1(n_1397),
.B2(n_1423),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1417),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1457),
.B(n_1447),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1428),
.B(n_1410),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1458),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1427),
.B(n_1435),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1428),
.Y(n_1516)
);

OA21x2_ASAP7_75t_L g1517 ( 
.A1(n_1425),
.A2(n_1417),
.B(n_1410),
.Y(n_1517)
);

AO21x2_ASAP7_75t_L g1518 ( 
.A1(n_1430),
.A2(n_1444),
.B(n_1463),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1438),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1444),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1421),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1449),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1464),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1437),
.B(n_1469),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1464),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1503),
.B(n_1451),
.Y(n_1526)
);

BUFx2_ASAP7_75t_L g1527 ( 
.A(n_1482),
.Y(n_1527)
);

AND2x4_ASAP7_75t_L g1528 ( 
.A(n_1482),
.B(n_1467),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1522),
.B(n_1450),
.Y(n_1529)
);

INVxp67_ASAP7_75t_L g1530 ( 
.A(n_1478),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1480),
.B(n_1429),
.Y(n_1531)
);

NAND2xp33_ASAP7_75t_SL g1532 ( 
.A(n_1497),
.B(n_1455),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1481),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1478),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1479),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1503),
.Y(n_1536)
);

AOI211xp5_ASAP7_75t_L g1537 ( 
.A1(n_1494),
.A2(n_1418),
.B(n_1414),
.C(n_1406),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1508),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1480),
.B(n_1413),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1479),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1505),
.B(n_1431),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1515),
.Y(n_1542)
);

AO21x2_ASAP7_75t_L g1543 ( 
.A1(n_1484),
.A2(n_1408),
.B(n_1413),
.Y(n_1543)
);

AOI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1500),
.A2(n_1403),
.B1(n_1452),
.B2(n_1431),
.Y(n_1544)
);

INVxp67_ASAP7_75t_L g1545 ( 
.A(n_1515),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1494),
.B(n_1439),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1498),
.B(n_1483),
.Y(n_1547)
);

NOR2x1_ASAP7_75t_L g1548 ( 
.A(n_1496),
.B(n_1518),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1498),
.B(n_1483),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1487),
.B(n_1506),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1516),
.B(n_1504),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1498),
.B(n_1483),
.Y(n_1552)
);

OAI221xp5_ASAP7_75t_L g1553 ( 
.A1(n_1532),
.A2(n_1496),
.B1(n_1500),
.B2(n_1493),
.C(n_1524),
.Y(n_1553)
);

NAND2xp33_ASAP7_75t_R g1554 ( 
.A(n_1531),
.B(n_1521),
.Y(n_1554)
);

OAI31xp33_ASAP7_75t_L g1555 ( 
.A1(n_1546),
.A2(n_1510),
.A3(n_1521),
.B(n_1513),
.Y(n_1555)
);

AOI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1537),
.A2(n_1510),
.B1(n_1521),
.B2(n_1501),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1531),
.B(n_1504),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1550),
.B(n_1487),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1538),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_SL g1560 ( 
.A1(n_1544),
.A2(n_1493),
.B1(n_1524),
.B2(n_1513),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1538),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1533),
.Y(n_1562)
);

OAI33xp33_ASAP7_75t_L g1563 ( 
.A1(n_1551),
.A2(n_1490),
.A3(n_1485),
.B1(n_1519),
.B2(n_1516),
.B3(n_1520),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1548),
.A2(n_1501),
.B1(n_1485),
.B2(n_1493),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1535),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1548),
.A2(n_1501),
.B1(n_1493),
.B2(n_1525),
.Y(n_1566)
);

OAI211xp5_ASAP7_75t_SL g1567 ( 
.A1(n_1544),
.A2(n_1497),
.B(n_1490),
.C(n_1520),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1550),
.B(n_1487),
.Y(n_1568)
);

NOR3xp33_ASAP7_75t_SL g1569 ( 
.A(n_1539),
.B(n_1506),
.C(n_1525),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1547),
.B(n_1489),
.Y(n_1570)
);

BUFx6f_ASAP7_75t_L g1571 ( 
.A(n_1539),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1540),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1542),
.B(n_1488),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1542),
.B(n_1488),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1533),
.Y(n_1575)
);

OAI221xp5_ASAP7_75t_L g1576 ( 
.A1(n_1537),
.A2(n_1493),
.B1(n_1491),
.B2(n_1489),
.C(n_1519),
.Y(n_1576)
);

AOI221xp5_ASAP7_75t_L g1577 ( 
.A1(n_1545),
.A2(n_1501),
.B1(n_1491),
.B2(n_1509),
.C(n_1511),
.Y(n_1577)
);

INVx1_ASAP7_75t_SL g1578 ( 
.A(n_1529),
.Y(n_1578)
);

AOI211xp5_ASAP7_75t_L g1579 ( 
.A1(n_1541),
.A2(n_1512),
.B(n_1507),
.C(n_1511),
.Y(n_1579)
);

OAI21xp33_ASAP7_75t_L g1580 ( 
.A1(n_1551),
.A2(n_1493),
.B(n_1492),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1526),
.A2(n_1501),
.B1(n_1493),
.B2(n_1523),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1547),
.B(n_1489),
.Y(n_1582)
);

BUFx6f_ASAP7_75t_L g1583 ( 
.A(n_1527),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_SL g1584 ( 
.A1(n_1543),
.A2(n_1499),
.B1(n_1518),
.B2(n_1517),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1549),
.B(n_1482),
.Y(n_1585)
);

AOI221xp5_ASAP7_75t_L g1586 ( 
.A1(n_1545),
.A2(n_1509),
.B1(n_1492),
.B2(n_1499),
.C(n_1507),
.Y(n_1586)
);

INVxp67_ASAP7_75t_L g1587 ( 
.A(n_1529),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1562),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1562),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1577),
.B(n_1530),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1555),
.B(n_1526),
.Y(n_1591)
);

INVx3_ASAP7_75t_L g1592 ( 
.A(n_1583),
.Y(n_1592)
);

BUFx6f_ASAP7_75t_L g1593 ( 
.A(n_1583),
.Y(n_1593)
);

INVx2_ASAP7_75t_SL g1594 ( 
.A(n_1583),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1575),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1559),
.Y(n_1596)
);

OAI21x1_ASAP7_75t_L g1597 ( 
.A1(n_1559),
.A2(n_1495),
.B(n_1502),
.Y(n_1597)
);

OR2x6_ASAP7_75t_L g1598 ( 
.A(n_1560),
.B(n_1486),
.Y(n_1598)
);

OAI21x1_ASAP7_75t_L g1599 ( 
.A1(n_1561),
.A2(n_1495),
.B(n_1502),
.Y(n_1599)
);

OAI21x1_ASAP7_75t_L g1600 ( 
.A1(n_1561),
.A2(n_1502),
.B(n_1514),
.Y(n_1600)
);

INVx1_ASAP7_75t_SL g1601 ( 
.A(n_1583),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1583),
.Y(n_1602)
);

INVx1_ASAP7_75t_SL g1603 ( 
.A(n_1558),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1575),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1557),
.B(n_1530),
.Y(n_1605)
);

AOI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1553),
.A2(n_1499),
.B(n_1543),
.Y(n_1606)
);

INVx5_ASAP7_75t_L g1607 ( 
.A(n_1571),
.Y(n_1607)
);

INVx4_ASAP7_75t_L g1608 ( 
.A(n_1571),
.Y(n_1608)
);

INVx2_ASAP7_75t_SL g1609 ( 
.A(n_1573),
.Y(n_1609)
);

INVxp67_ASAP7_75t_L g1610 ( 
.A(n_1571),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1571),
.B(n_1549),
.Y(n_1611)
);

NAND3xp33_ASAP7_75t_L g1612 ( 
.A(n_1556),
.B(n_1534),
.C(n_1512),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1558),
.B(n_1536),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1579),
.B(n_1528),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1568),
.B(n_1536),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1565),
.Y(n_1616)
);

BUFx3_ASAP7_75t_L g1617 ( 
.A(n_1571),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1570),
.B(n_1552),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1588),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1597),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1603),
.B(n_1585),
.Y(n_1621)
);

INVxp67_ASAP7_75t_SL g1622 ( 
.A(n_1614),
.Y(n_1622)
);

NAND4xp25_ASAP7_75t_SL g1623 ( 
.A(n_1612),
.B(n_1586),
.C(n_1564),
.D(n_1576),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1591),
.B(n_1569),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1588),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1589),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1589),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1595),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1590),
.B(n_1587),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1590),
.B(n_1568),
.Y(n_1630)
);

AOI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1612),
.A2(n_1567),
.B1(n_1554),
.B2(n_1566),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1602),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1595),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1603),
.B(n_1573),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1613),
.B(n_1574),
.Y(n_1635)
);

INVx2_ASAP7_75t_SL g1636 ( 
.A(n_1593),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1611),
.B(n_1585),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1604),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1611),
.B(n_1570),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1602),
.B(n_1582),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_SL g1641 ( 
.A(n_1605),
.B(n_1580),
.Y(n_1641)
);

NAND3xp33_ASAP7_75t_L g1642 ( 
.A(n_1606),
.B(n_1584),
.C(n_1581),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1616),
.Y(n_1643)
);

OAI21xp33_ASAP7_75t_L g1644 ( 
.A1(n_1606),
.A2(n_1507),
.B(n_1512),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1605),
.B(n_1552),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1610),
.B(n_1582),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1599),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1617),
.B(n_1578),
.Y(n_1648)
);

INVxp67_ASAP7_75t_L g1649 ( 
.A(n_1616),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1613),
.B(n_1609),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1599),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1599),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1609),
.B(n_1572),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1600),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1609),
.B(n_1534),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1617),
.B(n_1527),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1643),
.Y(n_1657)
);

OAI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1631),
.A2(n_1607),
.B(n_1594),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1619),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1640),
.B(n_1592),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1624),
.B(n_1618),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1619),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1650),
.B(n_1615),
.Y(n_1663)
);

AND2x4_ASAP7_75t_SL g1664 ( 
.A(n_1640),
.B(n_1598),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1625),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1632),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1632),
.B(n_1607),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1625),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1626),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1650),
.B(n_1615),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1631),
.B(n_1618),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1622),
.B(n_1601),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1637),
.B(n_1592),
.Y(n_1673)
);

OAI31xp33_ASAP7_75t_L g1674 ( 
.A1(n_1623),
.A2(n_1601),
.A3(n_1617),
.B(n_1594),
.Y(n_1674)
);

OR2x6_ASAP7_75t_L g1675 ( 
.A(n_1636),
.B(n_1598),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1626),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1636),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1629),
.B(n_1608),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1637),
.B(n_1592),
.Y(n_1679)
);

AND2x4_ASAP7_75t_L g1680 ( 
.A(n_1649),
.B(n_1607),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1656),
.B(n_1592),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1621),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1656),
.B(n_1594),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1627),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1630),
.B(n_1604),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1621),
.B(n_1607),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1630),
.B(n_1608),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1627),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1653),
.B(n_1596),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1628),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1628),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1683),
.B(n_1639),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1666),
.B(n_1682),
.Y(n_1693)
);

INVxp67_ASAP7_75t_L g1694 ( 
.A(n_1672),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1683),
.B(n_1681),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1668),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1674),
.B(n_1641),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1668),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1669),
.Y(n_1699)
);

INVxp67_ASAP7_75t_L g1700 ( 
.A(n_1678),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1663),
.B(n_1670),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1669),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1667),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1681),
.B(n_1639),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1660),
.B(n_1646),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1663),
.B(n_1653),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1661),
.B(n_1646),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1677),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_1667),
.Y(n_1709)
);

AOI22xp33_ASAP7_75t_L g1710 ( 
.A1(n_1658),
.A2(n_1642),
.B1(n_1644),
.B2(n_1598),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1671),
.B(n_1645),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1690),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1667),
.B(n_1633),
.Y(n_1713)
);

AND2x4_ASAP7_75t_L g1714 ( 
.A(n_1664),
.B(n_1633),
.Y(n_1714)
);

INVxp67_ASAP7_75t_L g1715 ( 
.A(n_1657),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1686),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1701),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1709),
.B(n_1657),
.Y(n_1718)
);

NOR2x1p5_ASAP7_75t_L g1719 ( 
.A(n_1693),
.B(n_1687),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1701),
.Y(n_1720)
);

OAI222xp33_ASAP7_75t_L g1721 ( 
.A1(n_1697),
.A2(n_1675),
.B1(n_1670),
.B2(n_1686),
.C1(n_1685),
.C2(n_1680),
.Y(n_1721)
);

NOR2xp67_ASAP7_75t_L g1722 ( 
.A(n_1714),
.B(n_1677),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1709),
.B(n_1673),
.Y(n_1723)
);

INVx3_ASAP7_75t_L g1724 ( 
.A(n_1714),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1703),
.B(n_1680),
.Y(n_1725)
);

OAI22xp33_ASAP7_75t_L g1726 ( 
.A1(n_1694),
.A2(n_1642),
.B1(n_1675),
.B2(n_1598),
.Y(n_1726)
);

AOI22xp33_ASAP7_75t_SL g1727 ( 
.A1(n_1711),
.A2(n_1695),
.B1(n_1715),
.B2(n_1700),
.Y(n_1727)
);

NOR4xp25_ASAP7_75t_L g1728 ( 
.A(n_1703),
.B(n_1644),
.C(n_1684),
.D(n_1691),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1708),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1696),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1695),
.Y(n_1731)
);

OAI221xp5_ASAP7_75t_L g1732 ( 
.A1(n_1710),
.A2(n_1675),
.B1(n_1598),
.B2(n_1662),
.C(n_1659),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1696),
.Y(n_1733)
);

AOI222xp33_ASAP7_75t_L g1734 ( 
.A1(n_1707),
.A2(n_1563),
.B1(n_1664),
.B2(n_1673),
.C1(n_1679),
.C2(n_1660),
.Y(n_1734)
);

AOI21x1_ASAP7_75t_L g1735 ( 
.A1(n_1714),
.A2(n_1680),
.B(n_1690),
.Y(n_1735)
);

OAI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1727),
.A2(n_1675),
.B1(n_1714),
.B2(n_1716),
.Y(n_1736)
);

AOI22xp33_ASAP7_75t_SL g1737 ( 
.A1(n_1732),
.A2(n_1692),
.B1(n_1705),
.B2(n_1704),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1727),
.B(n_1716),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1724),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1725),
.B(n_1692),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1731),
.B(n_1705),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1725),
.B(n_1704),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1717),
.Y(n_1743)
);

AOI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1734),
.A2(n_1679),
.B1(n_1713),
.B2(n_1598),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1720),
.B(n_1713),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1729),
.B(n_1713),
.Y(n_1746)
);

NOR3xp33_ASAP7_75t_L g1747 ( 
.A(n_1738),
.B(n_1721),
.C(n_1718),
.Y(n_1747)
);

NAND3xp33_ASAP7_75t_L g1748 ( 
.A(n_1736),
.B(n_1728),
.C(n_1724),
.Y(n_1748)
);

AOI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1736),
.A2(n_1721),
.B(n_1726),
.Y(n_1749)
);

NAND3xp33_ASAP7_75t_L g1750 ( 
.A(n_1744),
.B(n_1722),
.C(n_1723),
.Y(n_1750)
);

OAI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1737),
.A2(n_1732),
.B1(n_1719),
.B2(n_1706),
.Y(n_1751)
);

OAI211xp5_ASAP7_75t_L g1752 ( 
.A1(n_1746),
.A2(n_1735),
.B(n_1733),
.C(n_1730),
.Y(n_1752)
);

AOI222xp33_ASAP7_75t_L g1753 ( 
.A1(n_1743),
.A2(n_1712),
.B1(n_1698),
.B2(n_1702),
.C1(n_1699),
.C2(n_1713),
.Y(n_1753)
);

OAI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1740),
.A2(n_1706),
.B1(n_1607),
.B2(n_1685),
.Y(n_1754)
);

OAI221xp5_ASAP7_75t_L g1755 ( 
.A1(n_1742),
.A2(n_1712),
.B1(n_1702),
.B2(n_1699),
.C(n_1698),
.Y(n_1755)
);

NOR3xp33_ASAP7_75t_L g1756 ( 
.A(n_1739),
.B(n_1688),
.C(n_1676),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1753),
.Y(n_1757)
);

NOR2xp67_ASAP7_75t_L g1758 ( 
.A(n_1752),
.B(n_1745),
.Y(n_1758)
);

CKINVDCx20_ASAP7_75t_R g1759 ( 
.A(n_1751),
.Y(n_1759)
);

OA22x2_ASAP7_75t_L g1760 ( 
.A1(n_1754),
.A2(n_1741),
.B1(n_1665),
.B2(n_1608),
.Y(n_1760)
);

AOI221xp5_ASAP7_75t_L g1761 ( 
.A1(n_1747),
.A2(n_1608),
.B1(n_1689),
.B2(n_1593),
.C(n_1638),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1758),
.B(n_1750),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1757),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1761),
.B(n_1749),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1759),
.B(n_1748),
.Y(n_1765)
);

NOR2x1_ASAP7_75t_L g1766 ( 
.A(n_1760),
.B(n_1755),
.Y(n_1766)
);

NOR3xp33_ASAP7_75t_L g1767 ( 
.A(n_1761),
.B(n_1756),
.C(n_1689),
.Y(n_1767)
);

INVx3_ASAP7_75t_L g1768 ( 
.A(n_1762),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1765),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1763),
.B(n_1635),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1764),
.A2(n_1607),
.B1(n_1593),
.B2(n_1648),
.Y(n_1771)
);

AOI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1766),
.A2(n_1767),
.B(n_1634),
.Y(n_1772)
);

AOI211x1_ASAP7_75t_L g1773 ( 
.A1(n_1772),
.A2(n_1769),
.B(n_1771),
.C(n_1768),
.Y(n_1773)
);

AOI211xp5_ASAP7_75t_L g1774 ( 
.A1(n_1770),
.A2(n_1593),
.B(n_1648),
.C(n_1655),
.Y(n_1774)
);

NOR2x1_ASAP7_75t_L g1775 ( 
.A(n_1768),
.B(n_1638),
.Y(n_1775)
);

NOR2x1p5_ASAP7_75t_L g1776 ( 
.A(n_1773),
.B(n_1634),
.Y(n_1776)
);

NOR2x1_ASAP7_75t_L g1777 ( 
.A(n_1776),
.B(n_1775),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1777),
.Y(n_1778)
);

INVx1_ASAP7_75t_SL g1779 ( 
.A(n_1777),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1779),
.B(n_1774),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1778),
.B(n_1655),
.Y(n_1781)
);

AOI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1781),
.A2(n_1593),
.B1(n_1607),
.B2(n_1654),
.Y(n_1782)
);

AO22x2_ASAP7_75t_L g1783 ( 
.A1(n_1780),
.A2(n_1654),
.B1(n_1652),
.B2(n_1651),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1783),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1784),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1785),
.B(n_1782),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1786),
.A2(n_1593),
.B1(n_1654),
.B2(n_1652),
.Y(n_1787)
);

AOI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1787),
.A2(n_1652),
.B1(n_1620),
.B2(n_1651),
.Y(n_1788)
);

AOI211xp5_ASAP7_75t_L g1789 ( 
.A1(n_1788),
.A2(n_1651),
.B(n_1647),
.C(n_1620),
.Y(n_1789)
);


endmodule