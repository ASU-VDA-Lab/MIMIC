module fake_aes_6820_n_27 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_27);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_27;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
NAND2xp5_ASAP7_75t_L g12 ( .A(n_1), .B(n_6), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_9), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_10), .Y(n_14) );
HB1xp67_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
NOR2xp33_ASAP7_75t_R g16 ( .A(n_0), .B(n_11), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_8), .B(n_2), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_15), .Y(n_18) );
AOI21xp5_ASAP7_75t_L g19 ( .A1(n_12), .A2(n_4), .B(n_7), .Y(n_19) );
AO31x2_ASAP7_75t_L g20 ( .A1(n_18), .A2(n_12), .A3(n_17), .B(n_16), .Y(n_20) );
OR2x2_ASAP7_75t_L g21 ( .A(n_20), .B(n_0), .Y(n_21) );
OAI21xp33_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_17), .B(n_13), .Y(n_22) );
OAI21xp33_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_14), .B(n_19), .Y(n_23) );
HB1xp67_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
BUFx2_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
OAI22xp5_ASAP7_75t_SL g26 ( .A1(n_25), .A2(n_20), .B1(n_2), .B2(n_3), .Y(n_26) );
AOI22xp5_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_24), .B1(n_3), .B2(n_1), .Y(n_27) );
endmodule