module fake_aes_8749_n_34 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_34);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_34;
wire n_20;
wire n_23;
wire n_8;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_6), .Y(n_8) );
CKINVDCx5p33_ASAP7_75t_R g9 ( .A(n_7), .Y(n_9) );
CKINVDCx16_ASAP7_75t_R g10 ( .A(n_1), .Y(n_10) );
BUFx3_ASAP7_75t_L g11 ( .A(n_5), .Y(n_11) );
AND2x2_ASAP7_75t_L g12 ( .A(n_0), .B(n_2), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_2), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_10), .B(n_0), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_10), .B(n_1), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_11), .B(n_3), .Y(n_16) );
NOR2xp33_ASAP7_75t_L g17 ( .A(n_11), .B(n_3), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_14), .B(n_8), .Y(n_18) );
OR2x2_ASAP7_75t_L g19 ( .A(n_15), .B(n_13), .Y(n_19) );
INVx3_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
HB1xp67_ASAP7_75t_L g21 ( .A(n_17), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_20), .B(n_12), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_19), .Y(n_23) );
HB1xp67_ASAP7_75t_L g24 ( .A(n_20), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_23), .B(n_21), .Y(n_25) );
AOI22xp5_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_18), .B1(n_12), .B2(n_17), .Y(n_26) );
BUFx3_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_26), .B(n_22), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
XNOR2x1_ASAP7_75t_L g30 ( .A(n_27), .B(n_22), .Y(n_30) );
HB1xp67_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_29), .Y(n_32) );
AOI22xp5_ASAP7_75t_L g33 ( .A1(n_30), .A2(n_13), .B1(n_9), .B2(n_11), .Y(n_33) );
AOI22xp5_ASAP7_75t_L g34 ( .A1(n_32), .A2(n_4), .B1(n_31), .B2(n_33), .Y(n_34) );
endmodule