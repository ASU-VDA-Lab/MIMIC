module real_jpeg_20475_n_12 (n_5, n_4, n_8, n_0, n_280, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_280;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_276;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_255;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_0),
.A2(n_3),
.B1(n_18),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_0),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_0),
.A2(n_46),
.B1(n_47),
.B2(n_57),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_0),
.A2(n_25),
.B1(n_26),
.B2(n_57),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_0),
.A2(n_57),
.B1(n_72),
.B2(n_73),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_SL g164 ( 
.A1(n_0),
.A2(n_9),
.B(n_26),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_0),
.B(n_33),
.Y(n_178)
);

AOI21xp33_ASAP7_75t_L g193 ( 
.A1(n_0),
.A2(n_10),
.B(n_73),
.Y(n_193)
);

AOI21xp33_ASAP7_75t_SL g216 ( 
.A1(n_0),
.A2(n_47),
.B(n_48),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_1),
.A2(n_3),
.B1(n_18),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_31),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_1),
.A2(n_31),
.B1(n_46),
.B2(n_47),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_1),
.A2(n_31),
.B1(n_72),
.B2(n_73),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_2),
.A2(n_3),
.B1(n_18),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_2),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_61),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_2),
.A2(n_46),
.B1(n_47),
.B2(n_61),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_2),
.A2(n_61),
.B1(n_72),
.B2(n_73),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_3),
.A2(n_4),
.B1(n_17),
.B2(n_18),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

A2O1A1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_3),
.A2(n_22),
.B(n_57),
.C(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_4),
.A2(n_17),
.B1(n_25),
.B2(n_26),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_4),
.A2(n_17),
.B1(n_46),
.B2(n_47),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_4),
.A2(n_17),
.B1(n_72),
.B2(n_73),
.Y(n_88)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_5),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_5),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_6),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_9),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_70),
.Y(n_69)
);

INVx6_ASAP7_75t_SL g70 ( 
.A(n_10),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_10),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

BUFx3_ASAP7_75t_SL g47 ( 
.A(n_11),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_36),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_34),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_27),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_19),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_16),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_18),
.A2(n_21),
.B(n_23),
.C(n_24),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_21),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_19),
.B(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_24),
.Y(n_19)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_20),
.B(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_24),
.A2(n_30),
.B(n_54),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_25),
.A2(n_45),
.B(n_48),
.C(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_25),
.B(n_48),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g215 ( 
.A1(n_26),
.A2(n_49),
.B(n_57),
.C(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_28),
.B(n_38),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_32),
.A2(n_33),
.B1(n_60),
.B2(n_62),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_33),
.A2(n_55),
.B(n_60),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_75),
.B(n_278),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_39),
.B(n_276),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_39),
.B(n_276),
.Y(n_277)
);

FAx1_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_53),
.CI(n_58),
.CON(n_39),
.SN(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_44),
.B1(n_50),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_43),
.B(n_101),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_50),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_44),
.A2(n_100),
.B(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_45),
.A2(n_51),
.B1(n_99),
.B2(n_101),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_45),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_45),
.B(n_57),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_47),
.A2(n_57),
.B(n_70),
.C(n_193),
.Y(n_192)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_51),
.B(n_101),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_56),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_57),
.B(n_86),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_57),
.B(n_71),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.C(n_65),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_59),
.B(n_106),
.C(n_111),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_59),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_59),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_59),
.A2(n_98),
.B1(n_133),
.B2(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_59),
.B(n_160),
.C(n_161),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_59),
.A2(n_111),
.B1(n_133),
.B2(n_171),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_63),
.A2(n_65),
.B1(n_119),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_63),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_64),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_65),
.A2(n_119),
.B1(n_120),
.B2(n_123),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_65),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_74),
.Y(n_65)
);

INVxp33_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_67),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_68),
.A2(n_71),
.B1(n_74),
.B2(n_93),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_68),
.A2(n_71),
.B1(n_96),
.B2(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_71),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_71),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_72),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_72),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_73),
.B(n_86),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_275),
.B(n_277),
.Y(n_75)
);

OAI321xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_128),
.A3(n_139),
.B1(n_273),
.B2(n_274),
.C(n_280),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_113),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_78),
.B(n_113),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_97),
.C(n_104),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_79),
.B(n_97),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_91),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_89),
.B2(n_90),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_81),
.A2(n_82),
.B1(n_92),
.B2(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_92),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_82),
.A2(n_89),
.B(n_91),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_88),
.Y(n_82)
);

INVxp33_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_84),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_87),
.B1(n_88),
.B2(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_85),
.B(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_85),
.A2(n_86),
.B1(n_154),
.B2(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_86),
.A2(n_108),
.B(n_152),
.Y(n_151)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_86),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_89),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_92),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_95),
.A2(n_148),
.B(n_149),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_102),
.B(n_103),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_102),
.Y(n_103)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_98),
.B(n_177),
.C(n_179),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_98),
.A2(n_160),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_115),
.C(n_125),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_104),
.A2(n_105),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_106),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_107),
.A2(n_109),
.B1(n_208),
.B2(n_246),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_107),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_109),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_109),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_109),
.B(n_165),
.C(n_207),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_109),
.A2(n_208),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_109),
.B(n_226),
.C(n_231),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_111),
.B(n_116),
.C(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_111),
.A2(n_156),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_111),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_111),
.A2(n_146),
.B1(n_147),
.B2(n_171),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_111),
.B(n_147),
.C(n_214),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_113)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_124),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_116),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_116),
.A2(n_124),
.B1(n_132),
.B2(n_137),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_116),
.A2(n_124),
.B1(n_169),
.B2(n_172),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_116),
.A2(n_124),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_116),
.B(n_248),
.C(n_250),
.Y(n_265)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_123),
.C(n_124),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_120),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_124),
.B(n_137),
.C(n_138),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_129),
.B(n_130),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_138),
.Y(n_130)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_267),
.B(n_272),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_255),
.B(n_266),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_183),
.B(n_240),
.C(n_254),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_167),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_143),
.B(n_167),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_158),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_155),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_145),
.B(n_155),
.C(n_158),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_150),
.B2(n_151),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_146),
.A2(n_147),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_146),
.B(n_151),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_147),
.B(n_192),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_181),
.B(n_182),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_154),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_156),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_162),
.A2(n_163),
.B1(n_165),
.B2(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_199),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_165),
.A2(n_175),
.B1(n_205),
.B2(n_209),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_173),
.C(n_176),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_168),
.B(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_169),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_173),
.A2(n_174),
.B1(n_176),
.B2(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_176),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_190),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_239),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_233),
.B(n_238),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_223),
.B(n_232),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_211),
.B(n_222),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_202),
.B(n_210),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_194),
.B(n_201),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_198),
.B(n_200),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_204),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_205),
.Y(n_209)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_213),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_221),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_217),
.B1(n_218),
.B2(n_220),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_215),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_217),
.B(n_220),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_224),
.B(n_225),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_229),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_230),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_235),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_241),
.B(n_242),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_252),
.B2(n_253),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_247),
.C(n_253),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_252),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_256),
.B(n_257),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_265),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_263),
.C(n_265),
.Y(n_268)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_269),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);


endmodule