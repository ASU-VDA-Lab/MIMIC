module real_aes_6387_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_719;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g171 ( .A1(n_0), .A2(n_172), .B(n_173), .C(n_177), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_1), .B(n_166), .Y(n_179) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_2), .B(n_110), .C(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g439 ( .A(n_2), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_3), .B(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_4), .A2(n_160), .B(n_470), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_5), .A2(n_140), .B(n_157), .C(n_514), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_6), .A2(n_160), .B(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_7), .B(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_8), .B(n_166), .Y(n_476) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_9), .A2(n_132), .B(n_254), .Y(n_253) );
AOI222xp33_ASAP7_75t_L g445 ( .A1(n_10), .A2(n_446), .B1(n_715), .B2(n_718), .C1(n_722), .C2(n_723), .Y(n_445) );
AND2x6_ASAP7_75t_L g157 ( .A(n_11), .B(n_158), .Y(n_157) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_12), .A2(n_140), .B(n_157), .C(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g567 ( .A(n_13), .Y(n_567) );
INVx1_ASAP7_75t_L g107 ( .A(n_14), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_14), .B(n_40), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_15), .B(n_176), .Y(n_516) );
INVx1_ASAP7_75t_L g137 ( .A(n_16), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_17), .B(n_151), .Y(n_260) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_18), .A2(n_152), .B(n_525), .C(n_527), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_19), .B(n_166), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_20), .B(n_194), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g185 ( .A1(n_21), .A2(n_140), .B(n_186), .C(n_193), .Y(n_185) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_22), .A2(n_175), .B(n_228), .C(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_23), .B(n_176), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_24), .B(n_176), .Y(n_465) );
CKINVDCx16_ASAP7_75t_R g494 ( .A(n_25), .Y(n_494) );
INVx1_ASAP7_75t_L g464 ( .A(n_26), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_27), .A2(n_140), .B(n_193), .C(n_257), .Y(n_256) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_28), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_29), .Y(n_512) );
INVx1_ASAP7_75t_L g488 ( .A(n_30), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_31), .A2(n_160), .B(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g142 ( .A(n_32), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_33), .A2(n_155), .B(n_209), .C(n_210), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_34), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g472 ( .A1(n_35), .A2(n_175), .B(n_473), .C(n_475), .Y(n_472) );
INVxp67_ASAP7_75t_L g489 ( .A(n_36), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_37), .B(n_259), .Y(n_258) );
CKINVDCx14_ASAP7_75t_R g471 ( .A(n_38), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g462 ( .A1(n_39), .A2(n_140), .B(n_193), .C(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_40), .B(n_107), .Y(n_106) );
A2O1A1Ixp33_ASAP7_75t_L g564 ( .A1(n_41), .A2(n_177), .B(n_565), .C(n_566), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_42), .B(n_184), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g231 ( .A(n_43), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_44), .B(n_151), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_45), .B(n_160), .Y(n_255) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_46), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_47), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_48), .A2(n_155), .B(n_209), .C(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g174 ( .A(n_49), .Y(n_174) );
INVx1_ASAP7_75t_L g238 ( .A(n_50), .Y(n_238) );
INVx1_ASAP7_75t_L g532 ( .A(n_51), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_52), .B(n_160), .Y(n_235) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_53), .A2(n_71), .B1(n_123), .B2(n_124), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_53), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_54), .Y(n_198) );
CKINVDCx14_ASAP7_75t_R g563 ( .A(n_55), .Y(n_563) );
INVx1_ASAP7_75t_L g158 ( .A(n_56), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_57), .B(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_58), .B(n_166), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_59), .A2(n_147), .B(n_192), .C(n_249), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_60), .A2(n_70), .B1(n_716), .B2(n_717), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_60), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_61), .A2(n_102), .B1(n_114), .B2(n_728), .Y(n_101) );
INVx1_ASAP7_75t_L g136 ( .A(n_62), .Y(n_136) );
INVx1_ASAP7_75t_SL g474 ( .A(n_63), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_64), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_65), .B(n_151), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_66), .B(n_166), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_67), .B(n_152), .Y(n_225) );
INVx1_ASAP7_75t_L g497 ( .A(n_68), .Y(n_497) );
CKINVDCx16_ASAP7_75t_R g169 ( .A(n_69), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_70), .Y(n_717) );
INVx1_ASAP7_75t_L g124 ( .A(n_71), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_72), .B(n_188), .Y(n_187) );
A2O1A1Ixp33_ASAP7_75t_L g139 ( .A1(n_73), .A2(n_140), .B(n_145), .C(n_155), .Y(n_139) );
CKINVDCx16_ASAP7_75t_R g247 ( .A(n_74), .Y(n_247) );
INVx1_ASAP7_75t_L g113 ( .A(n_75), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_76), .A2(n_160), .B(n_562), .Y(n_561) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_77), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_78), .A2(n_160), .B(n_522), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_79), .A2(n_184), .B(n_484), .Y(n_483) );
CKINVDCx16_ASAP7_75t_R g461 ( .A(n_80), .Y(n_461) );
INVx1_ASAP7_75t_L g523 ( .A(n_81), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_82), .B(n_190), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_83), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_84), .A2(n_160), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g526 ( .A(n_85), .Y(n_526) );
INVx2_ASAP7_75t_L g134 ( .A(n_86), .Y(n_134) );
INVx1_ASAP7_75t_L g515 ( .A(n_87), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_88), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_89), .B(n_176), .Y(n_226) );
INVx2_ASAP7_75t_L g110 ( .A(n_90), .Y(n_110) );
OR2x2_ASAP7_75t_L g436 ( .A(n_90), .B(n_437), .Y(n_436) );
OR2x2_ASAP7_75t_L g450 ( .A(n_90), .B(n_438), .Y(n_450) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_91), .A2(n_140), .B(n_155), .C(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_92), .B(n_160), .Y(n_207) );
INVx1_ASAP7_75t_L g211 ( .A(n_93), .Y(n_211) );
INVxp67_ASAP7_75t_L g250 ( .A(n_94), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_95), .B(n_132), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_96), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g146 ( .A(n_97), .Y(n_146) );
INVx1_ASAP7_75t_L g221 ( .A(n_98), .Y(n_221) );
INVx2_ASAP7_75t_L g535 ( .A(n_99), .Y(n_535) );
AND2x2_ASAP7_75t_L g240 ( .A(n_100), .B(n_196), .Y(n_240) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_SL g728 ( .A(n_104), .Y(n_728) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_108), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g714 ( .A(n_110), .B(n_438), .Y(n_714) );
NOR2x2_ASAP7_75t_L g725 ( .A(n_110), .B(n_437), .Y(n_725) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
OA21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_120), .B(n_444), .Y(n_114) );
BUFx2_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_SL g727 ( .A(n_118), .Y(n_727) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI21xp5_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_435), .B(n_441), .Y(n_120) );
XNOR2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_125), .Y(n_121) );
INVx1_ASAP7_75t_L g447 ( .A(n_125), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_125), .A2(n_452), .B1(n_719), .B2(n_720), .Y(n_718) );
OR3x1_ASAP7_75t_L g125 ( .A(n_126), .B(n_343), .C(n_392), .Y(n_125) );
NAND5xp2_ASAP7_75t_L g126 ( .A(n_127), .B(n_277), .C(n_306), .D(n_314), .E(n_329), .Y(n_126) );
O2A1O1Ixp33_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_200), .B(n_216), .C(n_261), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_129), .B(n_180), .Y(n_128) );
AND2x2_ASAP7_75t_L g272 ( .A(n_129), .B(n_269), .Y(n_272) );
AND2x2_ASAP7_75t_L g305 ( .A(n_129), .B(n_181), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_129), .B(n_204), .Y(n_398) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_165), .Y(n_129) );
INVx2_ASAP7_75t_L g203 ( .A(n_130), .Y(n_203) );
BUFx2_ASAP7_75t_L g372 ( .A(n_130), .Y(n_372) );
AO21x2_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_138), .B(n_163), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_131), .B(n_164), .Y(n_163) );
INVx3_ASAP7_75t_L g166 ( .A(n_131), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_131), .B(n_215), .Y(n_214) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_131), .A2(n_220), .B(n_230), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_131), .B(n_467), .Y(n_466) );
AO21x2_ASAP7_75t_L g492 ( .A1(n_131), .A2(n_493), .B(n_500), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_131), .B(n_518), .Y(n_517) );
INVx4_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_132), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_132), .A2(n_255), .B(n_256), .Y(n_254) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g232 ( .A(n_133), .Y(n_232) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AND2x2_ASAP7_75t_SL g196 ( .A(n_134), .B(n_135), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_159), .Y(n_138) );
INVx5_ASAP7_75t_L g170 ( .A(n_140), .Y(n_170) );
AND2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_141), .Y(n_154) );
BUFx3_ASAP7_75t_L g178 ( .A(n_141), .Y(n_178) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g162 ( .A(n_142), .Y(n_162) );
INVx1_ASAP7_75t_L g229 ( .A(n_142), .Y(n_229) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_144), .Y(n_149) );
INVx3_ASAP7_75t_L g152 ( .A(n_144), .Y(n_152) );
AND2x2_ASAP7_75t_L g161 ( .A(n_144), .B(n_162), .Y(n_161) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_144), .Y(n_176) );
INVx1_ASAP7_75t_L g259 ( .A(n_144), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_150), .C(n_153), .Y(n_145) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
OAI22xp33_ASAP7_75t_L g487 ( .A1(n_148), .A2(n_151), .B1(n_488), .B2(n_489), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_148), .B(n_526), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_148), .B(n_535), .Y(n_534) );
INVx4_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g188 ( .A(n_149), .Y(n_188) );
INVx2_ASAP7_75t_L g172 ( .A(n_151), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_151), .B(n_250), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g463 ( .A1(n_151), .A2(n_191), .B(n_464), .C(n_465), .Y(n_463) );
INVx5_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_152), .B(n_567), .Y(n_566) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx3_ASAP7_75t_L g475 ( .A(n_154), .Y(n_475) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
O2A1O1Ixp33_ASAP7_75t_SL g168 ( .A1(n_156), .A2(n_169), .B(n_170), .C(n_171), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_L g246 ( .A1(n_156), .A2(n_170), .B(n_247), .C(n_248), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_156), .A2(n_170), .B(n_471), .C(n_472), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_SL g484 ( .A1(n_156), .A2(n_170), .B(n_485), .C(n_486), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_SL g522 ( .A1(n_156), .A2(n_170), .B(n_523), .C(n_524), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_SL g531 ( .A1(n_156), .A2(n_170), .B(n_532), .C(n_533), .Y(n_531) );
O2A1O1Ixp33_ASAP7_75t_SL g562 ( .A1(n_156), .A2(n_170), .B(n_563), .C(n_564), .Y(n_562) );
INVx4_ASAP7_75t_SL g156 ( .A(n_157), .Y(n_156) );
AND2x4_ASAP7_75t_L g160 ( .A(n_157), .B(n_161), .Y(n_160) );
BUFx3_ASAP7_75t_L g193 ( .A(n_157), .Y(n_193) );
NAND2x1p5_ASAP7_75t_L g222 ( .A(n_157), .B(n_161), .Y(n_222) );
BUFx2_ASAP7_75t_L g184 ( .A(n_160), .Y(n_184) );
INVx1_ASAP7_75t_L g192 ( .A(n_162), .Y(n_192) );
AND2x2_ASAP7_75t_L g180 ( .A(n_165), .B(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g270 ( .A(n_165), .Y(n_270) );
AND2x2_ASAP7_75t_L g356 ( .A(n_165), .B(n_269), .Y(n_356) );
AND2x2_ASAP7_75t_L g411 ( .A(n_165), .B(n_203), .Y(n_411) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_179), .Y(n_165) );
INVx2_ASAP7_75t_L g209 ( .A(n_170), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_175), .B(n_474), .Y(n_473) );
INVx4_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g565 ( .A(n_176), .Y(n_565) );
INVx2_ASAP7_75t_L g499 ( .A(n_177), .Y(n_499) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_178), .Y(n_213) );
INVx1_ASAP7_75t_L g527 ( .A(n_178), .Y(n_527) );
INVx1_ASAP7_75t_L g328 ( .A(n_180), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_180), .B(n_204), .Y(n_375) );
INVx5_ASAP7_75t_L g269 ( .A(n_181), .Y(n_269) );
AND2x4_ASAP7_75t_L g290 ( .A(n_181), .B(n_270), .Y(n_290) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_181), .Y(n_312) );
AND2x2_ASAP7_75t_L g387 ( .A(n_181), .B(n_372), .Y(n_387) );
AND2x2_ASAP7_75t_L g390 ( .A(n_181), .B(n_205), .Y(n_390) );
OR2x6_ASAP7_75t_L g181 ( .A(n_182), .B(n_197), .Y(n_181) );
AOI21xp5_ASAP7_75t_SL g182 ( .A1(n_183), .A2(n_185), .B(n_194), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_189), .B(n_191), .Y(n_186) );
INVx2_ASAP7_75t_L g190 ( .A(n_188), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g210 ( .A1(n_190), .A2(n_211), .B(n_212), .C(n_213), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_L g237 ( .A1(n_190), .A2(n_213), .B(n_238), .C(n_239), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g496 ( .A1(n_190), .A2(n_497), .B(n_498), .C(n_499), .Y(n_496) );
O2A1O1Ixp5_ASAP7_75t_L g514 ( .A1(n_190), .A2(n_499), .B(n_515), .C(n_516), .Y(n_514) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_192), .B(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_195), .B(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g199 ( .A(n_196), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_196), .A2(n_207), .B(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_196), .A2(n_235), .B(n_236), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g460 ( .A1(n_196), .A2(n_222), .B(n_461), .C(n_462), .Y(n_460) );
OA21x2_ASAP7_75t_L g560 ( .A1(n_196), .A2(n_561), .B(n_568), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
AO21x2_ASAP7_75t_L g510 ( .A1(n_199), .A2(n_511), .B(n_517), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_200), .B(n_270), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_200), .B(n_401), .Y(n_400) );
INVx2_ASAP7_75t_SL g200 ( .A(n_201), .Y(n_200) );
OR2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_204), .Y(n_201) );
AND2x2_ASAP7_75t_L g295 ( .A(n_202), .B(n_270), .Y(n_295) );
AND2x2_ASAP7_75t_L g313 ( .A(n_202), .B(n_205), .Y(n_313) );
INVx1_ASAP7_75t_L g333 ( .A(n_202), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_202), .B(n_269), .Y(n_378) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_202), .Y(n_420) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_203), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_204), .B(n_268), .Y(n_267) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_204), .Y(n_322) );
O2A1O1Ixp33_ASAP7_75t_L g325 ( .A1(n_204), .A2(n_265), .B(n_326), .C(n_328), .Y(n_325) );
AND2x2_ASAP7_75t_L g332 ( .A(n_204), .B(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g341 ( .A(n_204), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g345 ( .A(n_204), .B(n_269), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_204), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g360 ( .A(n_204), .B(n_270), .Y(n_360) );
AND2x2_ASAP7_75t_L g410 ( .A(n_204), .B(n_411), .Y(n_410) );
INVx5_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
BUFx2_ASAP7_75t_L g274 ( .A(n_205), .Y(n_274) );
AND2x2_ASAP7_75t_L g315 ( .A(n_205), .B(n_268), .Y(n_315) );
AND2x2_ASAP7_75t_L g327 ( .A(n_205), .B(n_302), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_205), .B(n_356), .Y(n_374) );
OR2x6_ASAP7_75t_L g205 ( .A(n_206), .B(n_214), .Y(n_205) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_241), .Y(n_216) );
INVx1_ASAP7_75t_L g263 ( .A(n_217), .Y(n_263) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_233), .Y(n_217) );
OR2x2_ASAP7_75t_L g265 ( .A(n_218), .B(n_233), .Y(n_265) );
NAND3xp33_ASAP7_75t_L g271 ( .A(n_218), .B(n_272), .C(n_273), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_218), .B(n_243), .Y(n_282) );
OR2x2_ASAP7_75t_L g297 ( .A(n_218), .B(n_285), .Y(n_297) );
AND2x2_ASAP7_75t_L g303 ( .A(n_218), .B(n_252), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_218), .B(n_434), .Y(n_433) );
INVx5_ASAP7_75t_SL g218 ( .A(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_219), .B(n_243), .Y(n_300) );
AND2x2_ASAP7_75t_L g339 ( .A(n_219), .B(n_253), .Y(n_339) );
NAND2xp5_ASAP7_75t_SL g367 ( .A(n_219), .B(n_252), .Y(n_367) );
OR2x2_ASAP7_75t_L g370 ( .A(n_219), .B(n_252), .Y(n_370) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_223), .Y(n_220) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_222), .A2(n_494), .B(n_495), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g511 ( .A1(n_222), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_227), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_227), .A2(n_258), .B(n_260), .Y(n_257) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
INVx2_ASAP7_75t_L g482 ( .A(n_232), .Y(n_482) );
INVx5_ASAP7_75t_SL g285 ( .A(n_233), .Y(n_285) );
OR2x2_ASAP7_75t_L g291 ( .A(n_233), .B(n_242), .Y(n_291) );
AND2x2_ASAP7_75t_L g307 ( .A(n_233), .B(n_308), .Y(n_307) );
AOI321xp33_ASAP7_75t_L g314 ( .A1(n_233), .A2(n_315), .A3(n_316), .B1(n_317), .B2(n_323), .C(n_325), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_233), .B(n_241), .Y(n_324) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_233), .Y(n_337) );
OR2x2_ASAP7_75t_L g384 ( .A(n_233), .B(n_282), .Y(n_384) );
AND2x2_ASAP7_75t_L g406 ( .A(n_233), .B(n_303), .Y(n_406) );
AND2x2_ASAP7_75t_L g425 ( .A(n_233), .B(n_243), .Y(n_425) );
OR2x6_ASAP7_75t_L g233 ( .A(n_234), .B(n_240), .Y(n_233) );
INVx1_ASAP7_75t_SL g241 ( .A(n_242), .Y(n_241) );
OR2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_252), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_243), .B(n_252), .Y(n_266) );
AND2x2_ASAP7_75t_L g275 ( .A(n_243), .B(n_276), .Y(n_275) );
INVx3_ASAP7_75t_L g302 ( .A(n_243), .Y(n_302) );
AND2x2_ASAP7_75t_L g308 ( .A(n_243), .B(n_303), .Y(n_308) );
INVxp67_ASAP7_75t_L g338 ( .A(n_243), .Y(n_338) );
OR2x2_ASAP7_75t_L g380 ( .A(n_243), .B(n_285), .Y(n_380) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_251), .Y(n_243) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_244), .A2(n_469), .B(n_476), .Y(n_468) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_244), .A2(n_521), .B(n_528), .Y(n_520) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_244), .A2(n_530), .B(n_536), .Y(n_529) );
OR2x2_ASAP7_75t_L g262 ( .A(n_252), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_SL g276 ( .A(n_252), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_252), .B(n_265), .Y(n_309) );
AND2x2_ASAP7_75t_L g358 ( .A(n_252), .B(n_302), .Y(n_358) );
AND2x2_ASAP7_75t_L g396 ( .A(n_252), .B(n_285), .Y(n_396) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_253), .B(n_285), .Y(n_284) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_264), .B(n_267), .C(n_271), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_262), .A2(n_264), .B1(n_389), .B2(n_391), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_264), .A2(n_287), .B1(n_342), .B2(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx1_ASAP7_75t_SL g416 ( .A(n_265), .Y(n_416) );
INVx1_ASAP7_75t_SL g316 ( .A(n_266), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_268), .B(n_288), .Y(n_318) );
AOI222xp33_ASAP7_75t_L g329 ( .A1(n_268), .A2(n_309), .B1(n_316), .B2(n_330), .C1(n_334), .C2(n_340), .Y(n_329) );
AND2x2_ASAP7_75t_L g419 ( .A(n_268), .B(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx2_ASAP7_75t_L g294 ( .A(n_269), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_269), .B(n_289), .Y(n_364) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_269), .Y(n_401) );
AND2x2_ASAP7_75t_L g404 ( .A(n_269), .B(n_313), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_269), .B(n_420), .Y(n_430) );
INVx1_ASAP7_75t_L g321 ( .A(n_270), .Y(n_321) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_270), .Y(n_349) );
O2A1O1Ixp33_ASAP7_75t_L g412 ( .A1(n_272), .A2(n_413), .B(n_414), .C(n_417), .Y(n_412) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
NAND3xp33_ASAP7_75t_L g335 ( .A(n_274), .B(n_336), .C(n_339), .Y(n_335) );
OR2x2_ASAP7_75t_L g363 ( .A(n_274), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_274), .B(n_290), .Y(n_391) );
OR2x2_ASAP7_75t_L g296 ( .A(n_276), .B(n_297), .Y(n_296) );
AOI211xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_280), .B(n_286), .C(n_298), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g407 ( .A(n_279), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g385 ( .A(n_280), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_281), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g299 ( .A(n_284), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_285), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g353 ( .A(n_285), .B(n_303), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_285), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_285), .B(n_302), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_291), .B1(n_292), .B2(n_296), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_288), .B(n_360), .Y(n_359) );
BUFx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_290), .B(n_332), .Y(n_331) );
OAI221xp5_ASAP7_75t_SL g354 ( .A1(n_291), .A2(n_355), .B1(n_357), .B2(n_359), .C(n_361), .Y(n_354) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AND2x2_ASAP7_75t_L g409 ( .A(n_294), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g422 ( .A(n_294), .B(n_411), .Y(n_422) );
INVx1_ASAP7_75t_L g342 ( .A(n_295), .Y(n_342) );
INVx1_ASAP7_75t_L g413 ( .A(n_296), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g402 ( .A1(n_297), .A2(n_380), .B(n_403), .Y(n_402) );
AOI21xp33_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_301), .B(n_304), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OAI21xp5_ASAP7_75t_SL g306 ( .A1(n_307), .A2(n_309), .B(n_310), .Y(n_306) );
INVx1_ASAP7_75t_L g346 ( .A(n_307), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_308), .A2(n_394), .B1(n_397), .B2(n_399), .C(n_402), .Y(n_393) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_316), .A2(n_406), .B1(n_407), .B2(n_409), .Y(n_405) );
NAND2xp5_ASAP7_75t_SL g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g382 ( .A(n_318), .Y(n_382) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NOR2xp67_ASAP7_75t_SL g320 ( .A(n_321), .B(n_322), .Y(n_320) );
AND2x2_ASAP7_75t_L g386 ( .A(n_322), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g351 ( .A(n_327), .Y(n_351) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_332), .B(n_356), .Y(n_408) );
INVxp67_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_338), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g424 ( .A(n_339), .B(n_425), .Y(n_424) );
AND2x4_ASAP7_75t_L g431 ( .A(n_339), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OAI211xp5_ASAP7_75t_SL g343 ( .A1(n_344), .A2(n_346), .B(n_347), .C(n_381), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AOI211xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_350), .B(n_354), .C(n_373), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_SL g434 ( .A(n_358), .Y(n_434) );
AND2x2_ASAP7_75t_L g371 ( .A(n_360), .B(n_372), .Y(n_371) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_365), .B1(n_369), .B2(n_371), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
OR2x2_ASAP7_75t_L g379 ( .A(n_367), .B(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g432 ( .A(n_368), .Y(n_432) );
INVxp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AOI31xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .A3(n_376), .B(n_379), .Y(n_373) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AOI211xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_383), .B(n_385), .C(n_388), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
CKINVDCx16_ASAP7_75t_R g389 ( .A(n_390), .Y(n_389) );
NAND5xp2_ASAP7_75t_L g392 ( .A(n_393), .B(n_405), .C(n_412), .D(n_426), .E(n_429), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_404), .A2(n_430), .B1(n_431), .B2(n_433), .Y(n_429) );
INVx1_ASAP7_75t_SL g428 ( .A(n_406), .Y(n_428) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AOI21xp33_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_421), .B(n_423), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_436), .Y(n_443) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
NAND3xp33_ASAP7_75t_L g444 ( .A(n_441), .B(n_445), .C(n_726), .Y(n_444) );
INVx1_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
OAI22xp5_ASAP7_75t_SL g446 ( .A1(n_447), .A2(n_448), .B1(n_451), .B2(n_714), .Y(n_446) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g719 ( .A(n_449), .Y(n_719) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OR3x1_ASAP7_75t_L g452 ( .A(n_453), .B(n_625), .C(n_672), .Y(n_452) );
NAND3xp33_ASAP7_75t_SL g453 ( .A(n_454), .B(n_571), .C(n_596), .Y(n_453) );
AOI221xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_509), .B1(n_537), .B2(n_540), .C(n_548), .Y(n_454) );
OAI21xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_477), .B(n_502), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_457), .B(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_457), .B(n_553), .Y(n_669) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_468), .Y(n_457) );
AND2x2_ASAP7_75t_L g539 ( .A(n_458), .B(n_508), .Y(n_539) );
AND2x2_ASAP7_75t_L g589 ( .A(n_458), .B(n_507), .Y(n_589) );
AND2x2_ASAP7_75t_L g610 ( .A(n_458), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g615 ( .A(n_458), .B(n_582), .Y(n_615) );
OR2x2_ASAP7_75t_L g623 ( .A(n_458), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g695 ( .A(n_458), .B(n_491), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_458), .B(n_644), .Y(n_709) );
INVx3_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g554 ( .A(n_459), .B(n_468), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_459), .B(n_491), .Y(n_555) );
AND2x4_ASAP7_75t_L g577 ( .A(n_459), .B(n_508), .Y(n_577) );
AND2x2_ASAP7_75t_L g607 ( .A(n_459), .B(n_479), .Y(n_607) );
AND2x2_ASAP7_75t_L g616 ( .A(n_459), .B(n_606), .Y(n_616) );
AND2x2_ASAP7_75t_L g632 ( .A(n_459), .B(n_492), .Y(n_632) );
OR2x2_ASAP7_75t_L g641 ( .A(n_459), .B(n_624), .Y(n_641) );
AND2x2_ASAP7_75t_L g647 ( .A(n_459), .B(n_582), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_459), .B(n_653), .Y(n_652) );
OR2x2_ASAP7_75t_L g661 ( .A(n_459), .B(n_504), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_459), .B(n_550), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_459), .B(n_611), .Y(n_700) );
OR2x6_ASAP7_75t_L g459 ( .A(n_460), .B(n_466), .Y(n_459) );
INVx2_ASAP7_75t_L g508 ( .A(n_468), .Y(n_508) );
AND2x2_ASAP7_75t_L g606 ( .A(n_468), .B(n_491), .Y(n_606) );
AND2x2_ASAP7_75t_L g611 ( .A(n_468), .B(n_492), .Y(n_611) );
INVx1_ASAP7_75t_L g667 ( .A(n_468), .Y(n_667) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g576 ( .A(n_478), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_491), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_479), .B(n_539), .Y(n_538) );
BUFx3_ASAP7_75t_L g553 ( .A(n_479), .Y(n_553) );
OR2x2_ASAP7_75t_L g624 ( .A(n_479), .B(n_491), .Y(n_624) );
OR2x2_ASAP7_75t_L g685 ( .A(n_479), .B(n_592), .Y(n_685) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_483), .B(n_490), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_481), .A2(n_505), .B(n_506), .Y(n_504) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g505 ( .A(n_483), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_490), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_491), .B(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g644 ( .A(n_491), .B(n_504), .Y(n_644) );
INVx2_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
BUFx2_ASAP7_75t_L g583 ( .A(n_492), .Y(n_583) );
INVx1_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_503), .A2(n_689), .B1(n_693), .B2(n_696), .C(n_697), .Y(n_688) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_507), .Y(n_503) );
INVx1_ASAP7_75t_SL g551 ( .A(n_504), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_504), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g683 ( .A(n_504), .B(n_539), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_507), .B(n_553), .Y(n_675) );
AND2x2_ASAP7_75t_L g582 ( .A(n_508), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_SL g586 ( .A(n_509), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_509), .B(n_592), .Y(n_622) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_519), .Y(n_509) );
AND2x2_ASAP7_75t_L g547 ( .A(n_510), .B(n_520), .Y(n_547) );
INVx4_ASAP7_75t_L g559 ( .A(n_510), .Y(n_559) );
BUFx3_ASAP7_75t_L g602 ( .A(n_510), .Y(n_602) );
AND3x2_ASAP7_75t_L g617 ( .A(n_510), .B(n_618), .C(n_619), .Y(n_617) );
AND2x2_ASAP7_75t_L g699 ( .A(n_519), .B(n_613), .Y(n_699) );
AND2x2_ASAP7_75t_L g707 ( .A(n_519), .B(n_592), .Y(n_707) );
INVx1_ASAP7_75t_SL g712 ( .A(n_519), .Y(n_712) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_529), .Y(n_519) );
INVx1_ASAP7_75t_SL g570 ( .A(n_520), .Y(n_570) );
AND2x2_ASAP7_75t_L g593 ( .A(n_520), .B(n_559), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_520), .B(n_543), .Y(n_595) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_520), .Y(n_635) );
OR2x2_ASAP7_75t_L g640 ( .A(n_520), .B(n_559), .Y(n_640) );
INVx2_ASAP7_75t_L g545 ( .A(n_529), .Y(n_545) );
AND2x2_ASAP7_75t_L g580 ( .A(n_529), .B(n_560), .Y(n_580) );
OR2x2_ASAP7_75t_L g600 ( .A(n_529), .B(n_560), .Y(n_600) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_529), .Y(n_620) );
INVx1_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
AOI21xp33_ASAP7_75t_L g670 ( .A1(n_538), .A2(n_579), .B(n_671), .Y(n_670) );
AOI322xp5_ASAP7_75t_L g706 ( .A1(n_540), .A2(n_550), .A3(n_577), .B1(n_707), .B2(n_708), .C1(n_710), .C2(n_713), .Y(n_706) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_546), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_542), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_543), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g569 ( .A(n_544), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g637 ( .A(n_545), .B(n_559), .Y(n_637) );
AND2x2_ASAP7_75t_L g704 ( .A(n_545), .B(n_560), .Y(n_704) );
INVx1_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g645 ( .A(n_547), .B(n_599), .Y(n_645) );
AOI31xp33_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_552), .A3(n_555), .B(n_556), .Y(n_548) );
AND2x2_ASAP7_75t_L g604 ( .A(n_550), .B(n_582), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_550), .B(n_574), .Y(n_686) );
AND2x2_ASAP7_75t_L g705 ( .A(n_550), .B(n_610), .Y(n_705) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_553), .B(n_582), .Y(n_594) );
NAND2x1p5_ASAP7_75t_L g628 ( .A(n_553), .B(n_611), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_553), .B(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_553), .B(n_695), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_554), .B(n_611), .Y(n_643) );
INVx1_ASAP7_75t_L g687 ( .A(n_554), .Y(n_687) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_569), .Y(n_557) );
INVxp67_ASAP7_75t_L g639 ( .A(n_558), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_559), .B(n_570), .Y(n_575) );
INVx1_ASAP7_75t_L g681 ( .A(n_559), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_559), .B(n_658), .Y(n_692) );
BUFx3_ASAP7_75t_L g592 ( .A(n_560), .Y(n_592) );
AND2x2_ASAP7_75t_L g618 ( .A(n_560), .B(n_570), .Y(n_618) );
INVx2_ASAP7_75t_L g658 ( .A(n_560), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_569), .B(n_691), .Y(n_690) );
AOI211xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_576), .B(n_578), .C(n_587), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AOI21xp33_ASAP7_75t_L g621 ( .A1(n_573), .A2(n_622), .B(n_623), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_574), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_574), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g654 ( .A(n_575), .B(n_600), .Y(n_654) );
INVx3_ASAP7_75t_L g585 ( .A(n_577), .Y(n_585) );
OAI22xp5_ASAP7_75t_SL g578 ( .A1(n_579), .A2(n_581), .B1(n_584), .B2(n_586), .Y(n_578) );
OAI21xp5_ASAP7_75t_SL g603 ( .A1(n_580), .A2(n_604), .B(n_605), .Y(n_603) );
AND2x2_ASAP7_75t_L g629 ( .A(n_580), .B(n_593), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_580), .B(n_681), .Y(n_680) );
INVxp67_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g584 ( .A(n_583), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g653 ( .A(n_583), .Y(n_653) );
OAI21xp5_ASAP7_75t_SL g597 ( .A1(n_584), .A2(n_598), .B(n_603), .Y(n_597) );
OAI22xp33_ASAP7_75t_SL g587 ( .A1(n_588), .A2(n_590), .B1(n_594), .B2(n_595), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_589), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVx1_ASAP7_75t_L g613 ( .A(n_592), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_592), .B(n_635), .Y(n_634) );
NOR3xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_608), .C(n_621), .Y(n_596) );
OAI22xp5_ASAP7_75t_SL g663 ( .A1(n_598), .A2(n_664), .B1(n_668), .B2(n_669), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_599), .B(n_601), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g668 ( .A(n_600), .B(n_601), .Y(n_668) );
AND2x2_ASAP7_75t_L g676 ( .A(n_601), .B(n_657), .Y(n_676) );
CKINVDCx16_ASAP7_75t_R g601 ( .A(n_602), .Y(n_601) );
O2A1O1Ixp33_ASAP7_75t_SL g684 ( .A1(n_602), .A2(n_685), .B(n_686), .C(n_687), .Y(n_684) );
OR2x2_ASAP7_75t_L g711 ( .A(n_602), .B(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
OAI21xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_612), .B(n_614), .Y(n_608) );
INVx1_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
O2A1O1Ixp33_ASAP7_75t_L g646 ( .A1(n_610), .A2(n_647), .B(n_648), .C(n_651), .Y(n_646) );
OAI21xp33_ASAP7_75t_SL g614 ( .A1(n_615), .A2(n_616), .B(n_617), .Y(n_614) );
AND2x2_ASAP7_75t_L g679 ( .A(n_618), .B(n_637), .Y(n_679) );
INVxp67_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g657 ( .A(n_620), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g662 ( .A(n_622), .Y(n_662) );
NAND3xp33_ASAP7_75t_SL g625 ( .A(n_626), .B(n_646), .C(n_659), .Y(n_625) );
AOI211xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_629), .B(n_630), .C(n_638), .Y(n_626) );
INVx1_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
INVx1_ASAP7_75t_L g696 ( .A(n_633), .Y(n_696) );
OR2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
INVx1_ASAP7_75t_L g656 ( .A(n_635), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_635), .B(n_704), .Y(n_703) );
INVxp67_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
A2O1A1Ixp33_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_640), .B(n_641), .C(n_642), .Y(n_638) );
INVx2_ASAP7_75t_SL g650 ( .A(n_640), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_641), .A2(n_652), .B1(n_654), .B2(n_655), .Y(n_651) );
OAI21xp33_ASAP7_75t_SL g642 ( .A1(n_643), .A2(n_644), .B(n_645), .Y(n_642) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
AOI211xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_662), .B(n_663), .C(n_670), .Y(n_659) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
INVxp33_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g713 ( .A(n_667), .Y(n_713) );
NAND4xp25_ASAP7_75t_L g672 ( .A(n_673), .B(n_688), .C(n_701), .D(n_706), .Y(n_672) );
AOI211xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_676), .B(n_677), .C(n_684), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AOI21xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_680), .B(n_682), .Y(n_677) );
AOI21xp33_ASAP7_75t_L g697 ( .A1(n_678), .A2(n_698), .B(n_700), .Y(n_697) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_685), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_705), .Y(n_701) );
INVxp67_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g721 ( .A(n_714), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_715), .Y(n_722) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
INVx3_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
endmodule