module fake_ibex_766_n_979 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_163, n_26, n_188, n_114, n_34, n_97, n_102, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_979);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_163;
input n_26;
input n_188;
input n_114;
input n_34;
input n_97;
input n_102;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_979;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_328;
wire n_372;
wire n_341;
wire n_293;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_947;
wire n_972;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_909;
wire n_545;
wire n_862;
wire n_583;
wire n_887;
wire n_957;
wire n_678;
wire n_663;
wire n_969;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_698;
wire n_375;
wire n_280;
wire n_340;
wire n_317;
wire n_708;
wire n_901;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_270;
wire n_383;
wire n_346;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_243;
wire n_497;
wire n_287;
wire n_711;
wire n_228;
wire n_671;
wire n_876;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_928;
wire n_655;
wire n_333;
wire n_898;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_732;
wire n_673;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_490;
wire n_407;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_858;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_960;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_648;
wire n_571;
wire n_472;
wire n_209;
wire n_229;
wire n_589;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_949;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_354;
wire n_392;
wire n_206;
wire n_630;
wire n_516;
wire n_567;
wire n_548;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_200;
wire n_506;
wire n_444;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_320;
wire n_285;
wire n_379;
wire n_247;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_440;
wire n_268;
wire n_955;
wire n_385;
wire n_342;
wire n_233;
wire n_414;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_450;
wire n_302;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_897;
wire n_889;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_890;
wire n_816;
wire n_912;
wire n_921;
wire n_874;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_202;
wire n_298;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVx2_ASAP7_75t_L g193 ( 
.A(n_43),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_167),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_117),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_45),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_185),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_172),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_146),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_142),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_55),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_138),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_134),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_0),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_150),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_118),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_135),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_98),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_162),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_61),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_183),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_123),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_57),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_63),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_84),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_110),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_179),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_93),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_25),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_99),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_182),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_5),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_33),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_171),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_36),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_21),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_39),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_86),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_20),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_119),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_37),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_158),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_153),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_51),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_112),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_26),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_36),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_124),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_24),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_94),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_136),
.B(n_107),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_1),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_9),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_26),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_69),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_96),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_178),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_42),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_187),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_66),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_77),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_44),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_180),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_85),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_64),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_163),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_58),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_181),
.Y(n_259)
);

BUFx5_ASAP7_75t_L g260 ( 
.A(n_79),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_131),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_106),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_105),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_137),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_165),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_177),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_49),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_111),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_65),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_97),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_149),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_62),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_161),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_35),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_145),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_60),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_154),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_54),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_78),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_70),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_2),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_141),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_102),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_40),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_87),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_160),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_116),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_4),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_80),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_113),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_52),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_164),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_175),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_56),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_53),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_68),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_14),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_0),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_39),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_29),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_100),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_132),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_71),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_81),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_2),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_152),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_156),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_174),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_46),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_101),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_6),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_59),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_191),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_121),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_126),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_115),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_74),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_108),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_83),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_249),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_305),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_205),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_210),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_307),
.Y(n_324)
);

OA21x2_ASAP7_75t_L g325 ( 
.A1(n_193),
.A2(n_92),
.B(n_190),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_307),
.Y(n_326)
);

AND2x2_ASAP7_75t_R g327 ( 
.A(n_220),
.B(n_1),
.Y(n_327)
);

BUFx8_ASAP7_75t_L g328 ( 
.A(n_254),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_260),
.Y(n_329)
);

INVxp33_ASAP7_75t_SL g330 ( 
.A(n_239),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_205),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_204),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_271),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_279),
.B(n_3),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_308),
.Y(n_335)
);

AND2x4_ASAP7_75t_L g336 ( 
.A(n_226),
.B(n_300),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_295),
.Y(n_337)
);

AND2x6_ASAP7_75t_L g338 ( 
.A(n_199),
.B(n_41),
.Y(n_338)
);

AND2x6_ASAP7_75t_L g339 ( 
.A(n_199),
.B(n_309),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_205),
.Y(n_340)
);

AND2x4_ASAP7_75t_L g341 ( 
.A(n_300),
.B(n_3),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_260),
.Y(n_342)
);

OA21x2_ASAP7_75t_L g343 ( 
.A1(n_193),
.A2(n_95),
.B(n_189),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_307),
.Y(n_344)
);

AND2x4_ASAP7_75t_L g345 ( 
.A(n_223),
.B(n_4),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_205),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_298),
.B(n_5),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_224),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_284),
.Y(n_349)
);

AND2x4_ASAP7_75t_L g350 ( 
.A(n_227),
.B(n_6),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_260),
.Y(n_351)
);

OAI21x1_ASAP7_75t_L g352 ( 
.A1(n_196),
.A2(n_234),
.B(n_215),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_236),
.B(n_7),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_230),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_260),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_260),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_309),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_270),
.B(n_7),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_260),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_284),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_243),
.Y(n_361)
);

OAI22xp33_ASAP7_75t_L g362 ( 
.A1(n_220),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_362)
);

BUFx8_ASAP7_75t_L g363 ( 
.A(n_277),
.Y(n_363)
);

OAI21x1_ASAP7_75t_L g364 ( 
.A1(n_196),
.A2(n_103),
.B(n_186),
.Y(n_364)
);

BUFx12f_ASAP7_75t_L g365 ( 
.A(n_204),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_288),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_299),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_311),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_284),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_291),
.B(n_276),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_262),
.Y(n_371)
);

BUFx8_ASAP7_75t_L g372 ( 
.A(n_284),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_215),
.B(n_8),
.Y(n_373)
);

CKINVDCx11_ASAP7_75t_R g374 ( 
.A(n_238),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_234),
.B(n_10),
.Y(n_375)
);

INVx6_ASAP7_75t_L g376 ( 
.A(n_316),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_250),
.B(n_11),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_250),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_195),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_297),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_197),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_272),
.Y(n_382)
);

BUFx8_ASAP7_75t_SL g383 ( 
.A(n_238),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_272),
.B(n_11),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_275),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_275),
.B(n_12),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_278),
.B(n_12),
.Y(n_387)
);

BUFx8_ASAP7_75t_L g388 ( 
.A(n_201),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_278),
.B(n_13),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_262),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_301),
.B(n_312),
.Y(n_391)
);

OAI21x1_ASAP7_75t_L g392 ( 
.A1(n_301),
.A2(n_109),
.B(n_184),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_312),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_314),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_240),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_202),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_341),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_341),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_352),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_377),
.B(n_387),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_377),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_387),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_332),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_382),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_389),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_389),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_324),
.B(n_203),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_339),
.Y(n_408)
);

INVx2_ASAP7_75t_SL g409 ( 
.A(n_332),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_321),
.Y(n_410)
);

BUFx6f_ASAP7_75t_SL g411 ( 
.A(n_345),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_391),
.B(n_207),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_321),
.B(n_253),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_345),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_339),
.Y(n_415)
);

INVx5_ASAP7_75t_L g416 ( 
.A(n_338),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_334),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_320),
.B(n_253),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_320),
.B(n_380),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_372),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_350),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_329),
.B(n_209),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_350),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_385),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g425 ( 
.A(n_324),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_322),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_385),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_336),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_385),
.Y(n_429)
);

AND2x6_ASAP7_75t_L g430 ( 
.A(n_344),
.B(n_213),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_385),
.Y(n_431)
);

OAI22xp33_ASAP7_75t_L g432 ( 
.A1(n_390),
.A2(n_240),
.B1(n_314),
.B2(n_228),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_393),
.Y(n_433)
);

AO21x2_ASAP7_75t_L g434 ( 
.A1(n_364),
.A2(n_221),
.B(n_218),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_344),
.B(n_225),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_365),
.Y(n_436)
);

BUFx10_ASAP7_75t_L g437 ( 
.A(n_323),
.Y(n_437)
);

OAI22xp33_ASAP7_75t_L g438 ( 
.A1(n_394),
.A2(n_245),
.B1(n_274),
.B2(n_281),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_370),
.B(n_198),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_378),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g441 ( 
.A(n_333),
.B(n_232),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_393),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_393),
.Y(n_443)
);

NAND2xp33_ASAP7_75t_L g444 ( 
.A(n_338),
.B(n_339),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_371),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_378),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_348),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_335),
.B(n_237),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_342),
.B(n_233),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_347),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_393),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_354),
.Y(n_452)
);

INVx5_ASAP7_75t_L g453 ( 
.A(n_338),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_370),
.B(n_198),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_351),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_361),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_355),
.B(n_256),
.Y(n_457)
);

NAND2xp33_ASAP7_75t_L g458 ( 
.A(n_338),
.B(n_208),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_366),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_367),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_337),
.B(n_200),
.Y(n_461)
);

NAND2xp33_ASAP7_75t_R g462 ( 
.A(n_330),
.B(n_244),
.Y(n_462)
);

INVx4_ASAP7_75t_L g463 ( 
.A(n_338),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_330),
.B(n_200),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_356),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_359),
.B(n_257),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_L g467 ( 
.A(n_339),
.B(n_306),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_368),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_379),
.A2(n_396),
.B1(n_381),
.B2(n_375),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_357),
.B(n_258),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_339),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_373),
.Y(n_472)
);

AO21x2_ASAP7_75t_L g473 ( 
.A1(n_392),
.A2(n_269),
.B(n_261),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_375),
.Y(n_474)
);

BUFx6f_ASAP7_75t_SL g475 ( 
.A(n_326),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_363),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_363),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_322),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_372),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_384),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_331),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_376),
.B(n_273),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_331),
.Y(n_483)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_376),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_376),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_384),
.B(n_285),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_386),
.B(n_286),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_353),
.B(n_310),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_358),
.B(n_310),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_386),
.Y(n_490)
);

NAND2xp33_ASAP7_75t_L g491 ( 
.A(n_334),
.B(n_313),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_349),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_340),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_340),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_328),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_388),
.B(n_290),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_388),
.B(n_304),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_463),
.B(n_194),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_439),
.B(n_328),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_413),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_410),
.B(n_394),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_403),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_417),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_408),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_416),
.B(n_206),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_472),
.Y(n_506)
);

NOR3xp33_ASAP7_75t_L g507 ( 
.A(n_432),
.B(n_362),
.C(n_374),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_462),
.Y(n_508)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_419),
.B(n_362),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_474),
.B(n_325),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_480),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_416),
.B(n_211),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_490),
.Y(n_513)
);

OAI22xp33_ASAP7_75t_L g514 ( 
.A1(n_462),
.A2(n_395),
.B1(n_327),
.B2(n_325),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_454),
.B(n_212),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_469),
.B(n_343),
.Y(n_516)
);

NOR2xp67_ASAP7_75t_L g517 ( 
.A(n_495),
.B(n_16),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_469),
.B(n_343),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_447),
.B(n_452),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_408),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_450),
.B(n_418),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_440),
.Y(n_522)
);

NAND3xp33_ASAP7_75t_L g523 ( 
.A(n_491),
.B(n_343),
.C(n_216),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_456),
.B(n_214),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_464),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_414),
.A2(n_219),
.B1(n_251),
.B2(n_267),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_459),
.B(n_217),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_460),
.B(n_222),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_446),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_416),
.B(n_229),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_409),
.B(n_374),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_468),
.B(n_231),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_425),
.B(n_235),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_421),
.A2(n_242),
.B1(n_349),
.B2(n_369),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_420),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_420),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_401),
.B(n_241),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_479),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_461),
.A2(n_283),
.B1(n_247),
.B2(n_248),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_453),
.B(n_246),
.Y(n_540)
);

NOR2xp67_ASAP7_75t_L g541 ( 
.A(n_476),
.B(n_17),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_477),
.B(n_395),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_402),
.B(n_252),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_428),
.B(n_255),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_488),
.B(n_259),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_405),
.B(n_263),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_453),
.B(n_264),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_484),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_397),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_404),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_441),
.B(n_383),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_406),
.B(n_423),
.Y(n_552)
);

INVxp33_ASAP7_75t_L g553 ( 
.A(n_436),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_489),
.B(n_265),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_453),
.B(n_266),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_415),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_486),
.B(n_487),
.Y(n_557)
);

BUFx5_ASAP7_75t_L g558 ( 
.A(n_471),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_486),
.B(n_268),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_411),
.B(n_448),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_487),
.B(n_398),
.Y(n_561)
);

O2A1O1Ixp33_ASAP7_75t_L g562 ( 
.A1(n_400),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_437),
.Y(n_563)
);

BUFx8_ASAP7_75t_L g564 ( 
.A(n_475),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_496),
.B(n_280),
.Y(n_565)
);

CKINVDCx11_ASAP7_75t_R g566 ( 
.A(n_437),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_496),
.B(n_282),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_497),
.B(n_287),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_491),
.A2(n_411),
.B1(n_438),
.B2(n_497),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_407),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_445),
.A2(n_383),
.B1(n_319),
.B2(n_318),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_435),
.B(n_289),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_412),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_412),
.B(n_292),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_435),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_485),
.B(n_293),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_430),
.B(n_470),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_430),
.B(n_294),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_506),
.B(n_511),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_510),
.A2(n_444),
.B(n_458),
.Y(n_580)
);

AND2x2_ASAP7_75t_SL g581 ( 
.A(n_507),
.B(n_458),
.Y(n_581)
);

O2A1O1Ixp33_ASAP7_75t_L g582 ( 
.A1(n_509),
.A2(n_422),
.B(n_466),
.C(n_449),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_513),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_570),
.B(n_482),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_510),
.A2(n_444),
.B(n_467),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_503),
.B(n_482),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_525),
.B(n_422),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g588 ( 
.A1(n_516),
.A2(n_399),
.B(n_434),
.Y(n_588)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_518),
.A2(n_434),
.B(n_473),
.Y(n_589)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_518),
.A2(n_473),
.B(n_449),
.Y(n_590)
);

A2O1A1Ixp33_ASAP7_75t_L g591 ( 
.A1(n_575),
.A2(n_457),
.B(n_466),
.C(n_465),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_519),
.A2(n_465),
.B(n_455),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_563),
.B(n_455),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_519),
.B(n_296),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_501),
.A2(n_475),
.B1(n_303),
.B2(n_315),
.Y(n_595)
);

AO21x2_ASAP7_75t_L g596 ( 
.A1(n_523),
.A2(n_442),
.B(n_424),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_514),
.A2(n_302),
.B1(n_317),
.B2(n_349),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_574),
.B(n_18),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_574),
.B(n_19),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_557),
.A2(n_443),
.B1(n_451),
.B2(n_442),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_502),
.B(n_21),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_561),
.A2(n_433),
.B(n_427),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_L g603 ( 
.A1(n_552),
.A2(n_451),
.B1(n_429),
.B2(n_431),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_561),
.A2(n_433),
.B(n_429),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_549),
.B(n_22),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_504),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_535),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_524),
.A2(n_494),
.B(n_493),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_527),
.A2(n_494),
.B(n_478),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_552),
.A2(n_360),
.B1(n_369),
.B2(n_346),
.Y(n_610)
);

OAI321xp33_ASAP7_75t_L g611 ( 
.A1(n_562),
.A2(n_369),
.A3(n_360),
.B1(n_569),
.B2(n_521),
.C(n_346),
.Y(n_611)
);

A2O1A1Ixp33_ASAP7_75t_L g612 ( 
.A1(n_515),
.A2(n_360),
.B(n_369),
.C(n_492),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_527),
.A2(n_483),
.B(n_481),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_500),
.B(n_531),
.Y(n_614)
);

OAI321xp33_ASAP7_75t_L g615 ( 
.A1(n_562),
.A2(n_360),
.A3(n_346),
.B1(n_340),
.B2(n_478),
.C(n_426),
.Y(n_615)
);

INVx1_ASAP7_75t_SL g616 ( 
.A(n_566),
.Y(n_616)
);

AND2x2_ASAP7_75t_SL g617 ( 
.A(n_542),
.B(n_22),
.Y(n_617)
);

O2A1O1Ixp33_ASAP7_75t_L g618 ( 
.A1(n_508),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_618)
);

OAI21xp33_ASAP7_75t_L g619 ( 
.A1(n_499),
.A2(n_543),
.B(n_537),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_522),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_528),
.B(n_532),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_560),
.B(n_23),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_528),
.B(n_27),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_529),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_573),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_546),
.B(n_27),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_551),
.B(n_28),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_534),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_628)
);

CKINVDCx8_ASAP7_75t_R g629 ( 
.A(n_564),
.Y(n_629)
);

AND3x2_ASAP7_75t_L g630 ( 
.A(n_564),
.B(n_30),
.C(n_31),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_545),
.B(n_32),
.Y(n_631)
);

A2O1A1Ixp33_ASAP7_75t_L g632 ( 
.A1(n_554),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_632)
);

BUFx12f_ASAP7_75t_L g633 ( 
.A(n_536),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_577),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_571),
.B(n_38),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_559),
.A2(n_498),
.B(n_572),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_539),
.B(n_526),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_L g638 ( 
.A1(n_578),
.A2(n_122),
.B(n_176),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_544),
.B(n_38),
.Y(n_639)
);

OAI321xp33_ASAP7_75t_L g640 ( 
.A1(n_578),
.A2(n_565),
.A3(n_568),
.B1(n_567),
.B2(n_533),
.C(n_576),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_505),
.A2(n_120),
.B(n_47),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_512),
.A2(n_125),
.B(n_48),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_530),
.A2(n_127),
.B(n_50),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_553),
.B(n_40),
.Y(n_644)
);

OR2x6_ASAP7_75t_L g645 ( 
.A(n_538),
.B(n_67),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_548),
.A2(n_72),
.B1(n_73),
.B2(n_75),
.Y(n_646)
);

BUFx8_ASAP7_75t_L g647 ( 
.A(n_517),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_548),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_L g649 ( 
.A1(n_550),
.A2(n_76),
.B(n_82),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_540),
.A2(n_88),
.B(n_89),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_541),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_547),
.A2(n_90),
.B(n_91),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_555),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_520),
.B(n_192),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_520),
.B(n_104),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_579),
.B(n_556),
.Y(n_656)
);

NOR2x1_ASAP7_75t_SL g657 ( 
.A(n_645),
.B(n_621),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_583),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_614),
.Y(n_659)
);

INVx6_ASAP7_75t_L g660 ( 
.A(n_633),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_624),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_645),
.Y(n_662)
);

AO21x1_ASAP7_75t_L g663 ( 
.A1(n_638),
.A2(n_649),
.B(n_646),
.Y(n_663)
);

INVx1_ASAP7_75t_SL g664 ( 
.A(n_593),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_L g665 ( 
.A1(n_591),
.A2(n_558),
.B(n_114),
.Y(n_665)
);

AO21x2_ASAP7_75t_L g666 ( 
.A1(n_638),
.A2(n_558),
.B(n_128),
.Y(n_666)
);

NOR2xp67_ASAP7_75t_L g667 ( 
.A(n_627),
.B(n_129),
.Y(n_667)
);

OAI21x1_ASAP7_75t_L g668 ( 
.A1(n_654),
.A2(n_130),
.B(n_133),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_625),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_620),
.Y(n_670)
);

OAI21x1_ASAP7_75t_L g671 ( 
.A1(n_655),
.A2(n_139),
.B(n_140),
.Y(n_671)
);

INVx3_ASAP7_75t_SL g672 ( 
.A(n_616),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_592),
.A2(n_143),
.B(n_144),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_617),
.B(n_147),
.Y(n_674)
);

AOI21xp33_ASAP7_75t_L g675 ( 
.A1(n_595),
.A2(n_148),
.B(n_151),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g676 ( 
.A1(n_582),
.A2(n_155),
.B(n_157),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_645),
.B(n_159),
.Y(n_677)
);

INVx1_ASAP7_75t_SL g678 ( 
.A(n_593),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_581),
.B(n_168),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_644),
.B(n_169),
.Y(n_680)
);

OAI21x1_ASAP7_75t_SL g681 ( 
.A1(n_623),
.A2(n_170),
.B(n_173),
.Y(n_681)
);

INVx1_ASAP7_75t_SL g682 ( 
.A(n_607),
.Y(n_682)
);

NOR4xp25_ASAP7_75t_L g683 ( 
.A(n_618),
.B(n_632),
.C(n_634),
.D(n_611),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_651),
.B(n_598),
.Y(n_684)
);

BUFx12f_ASAP7_75t_L g685 ( 
.A(n_647),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_587),
.B(n_594),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_599),
.B(n_586),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_636),
.A2(n_604),
.B(n_602),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_597),
.B(n_601),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_622),
.B(n_605),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_L g691 ( 
.A1(n_626),
.A2(n_631),
.B1(n_639),
.B2(n_628),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_608),
.A2(n_613),
.B(n_609),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_647),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_596),
.A2(n_640),
.B(n_600),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_640),
.B(n_606),
.Y(n_695)
);

AOI21xp33_ASAP7_75t_L g696 ( 
.A1(n_653),
.A2(n_648),
.B(n_603),
.Y(n_696)
);

AOI211x1_ASAP7_75t_L g697 ( 
.A1(n_635),
.A2(n_652),
.B(n_642),
.C(n_641),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_630),
.B(n_606),
.Y(n_698)
);

AO31x2_ASAP7_75t_L g699 ( 
.A1(n_612),
.A2(n_610),
.A3(n_650),
.B(n_643),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_606),
.Y(n_700)
);

OAI21x1_ASAP7_75t_L g701 ( 
.A1(n_615),
.A2(n_611),
.B(n_629),
.Y(n_701)
);

OAI21xp5_ASAP7_75t_L g702 ( 
.A1(n_615),
.A2(n_580),
.B(n_590),
.Y(n_702)
);

CKINVDCx6p67_ASAP7_75t_R g703 ( 
.A(n_633),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_579),
.B(n_417),
.Y(n_704)
);

AND2x6_ASAP7_75t_L g705 ( 
.A(n_579),
.B(n_506),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_617),
.A2(n_371),
.B1(n_507),
.B2(n_502),
.Y(n_706)
);

O2A1O1Ixp5_ASAP7_75t_L g707 ( 
.A1(n_589),
.A2(n_631),
.B(n_639),
.C(n_580),
.Y(n_707)
);

AOI21xp33_ASAP7_75t_L g708 ( 
.A1(n_619),
.A2(n_462),
.B(n_499),
.Y(n_708)
);

INVx5_ASAP7_75t_L g709 ( 
.A(n_645),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_606),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_617),
.B(n_563),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_583),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_579),
.B(n_417),
.Y(n_713)
);

INVx4_ASAP7_75t_L g714 ( 
.A(n_633),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_637),
.B(n_501),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_579),
.A2(n_570),
.B1(n_584),
.B2(n_511),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_L g717 ( 
.A1(n_588),
.A2(n_444),
.B(n_510),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_579),
.B(n_417),
.Y(n_718)
);

AND2x6_ASAP7_75t_L g719 ( 
.A(n_579),
.B(n_506),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_588),
.A2(n_444),
.B(n_510),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_583),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_579),
.A2(n_570),
.B1(n_584),
.B2(n_511),
.Y(n_722)
);

INVxp67_ASAP7_75t_SL g723 ( 
.A(n_579),
.Y(n_723)
);

OA21x2_ASAP7_75t_L g724 ( 
.A1(n_589),
.A2(n_588),
.B(n_590),
.Y(n_724)
);

NOR2x1_ASAP7_75t_L g725 ( 
.A(n_616),
.B(n_645),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_588),
.A2(n_444),
.B(n_510),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_637),
.B(n_501),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_579),
.B(n_506),
.Y(n_728)
);

OAI21x1_ASAP7_75t_SL g729 ( 
.A1(n_621),
.A2(n_638),
.B(n_649),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_579),
.B(n_417),
.Y(n_730)
);

OAI21xp5_ASAP7_75t_L g731 ( 
.A1(n_580),
.A2(n_590),
.B(n_585),
.Y(n_731)
);

OAI21xp5_ASAP7_75t_L g732 ( 
.A1(n_580),
.A2(n_590),
.B(n_585),
.Y(n_732)
);

OAI21xp33_ASAP7_75t_L g733 ( 
.A1(n_621),
.A2(n_450),
.B(n_521),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_633),
.Y(n_734)
);

INVx1_ASAP7_75t_SL g735 ( 
.A(n_614),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_614),
.B(n_410),
.Y(n_736)
);

O2A1O1Ixp33_ASAP7_75t_L g737 ( 
.A1(n_621),
.A2(n_514),
.B(n_438),
.C(n_632),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_614),
.B(n_410),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_579),
.B(n_417),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_606),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_L g741 ( 
.A1(n_579),
.A2(n_570),
.B1(n_584),
.B2(n_511),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_579),
.B(n_417),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_658),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_692),
.A2(n_729),
.B(n_688),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_661),
.Y(n_745)
);

OR2x2_ASAP7_75t_SL g746 ( 
.A(n_660),
.B(n_698),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_710),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_SL g748 ( 
.A1(n_657),
.A2(n_677),
.B1(n_709),
.B2(n_719),
.Y(n_748)
);

AO31x2_ASAP7_75t_L g749 ( 
.A1(n_663),
.A2(n_726),
.A3(n_720),
.B(n_717),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_728),
.B(n_735),
.Y(n_750)
);

INVx4_ASAP7_75t_L g751 ( 
.A(n_709),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_711),
.A2(n_716),
.B1(n_741),
.B2(n_722),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_660),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_685),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_723),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_SL g756 ( 
.A1(n_677),
.A2(n_657),
.B(n_676),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_732),
.A2(n_707),
.B(n_724),
.Y(n_757)
);

AOI222xp33_ASAP7_75t_L g758 ( 
.A1(n_733),
.A2(n_659),
.B1(n_674),
.B2(n_728),
.C1(n_686),
.C2(n_687),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_706),
.B(n_736),
.Y(n_759)
);

OAI21xp5_ASAP7_75t_L g760 ( 
.A1(n_737),
.A2(n_683),
.B(n_665),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_709),
.A2(n_690),
.B1(n_725),
.B2(n_721),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_658),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_703),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_738),
.B(n_742),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_670),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_705),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_704),
.B(n_730),
.Y(n_767)
);

OAI21x1_ASAP7_75t_SL g768 ( 
.A1(n_681),
.A2(n_673),
.B(n_679),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_712),
.Y(n_769)
);

OA21x2_ASAP7_75t_L g770 ( 
.A1(n_701),
.A2(n_668),
.B(n_671),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_672),
.Y(n_771)
);

BUFx2_ASAP7_75t_L g772 ( 
.A(n_705),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_712),
.Y(n_773)
);

AO21x2_ASAP7_75t_L g774 ( 
.A1(n_666),
.A2(n_675),
.B(n_667),
.Y(n_774)
);

OA21x2_ASAP7_75t_L g775 ( 
.A1(n_700),
.A2(n_669),
.B(n_708),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_719),
.B(n_713),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_689),
.A2(n_684),
.B(n_680),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_718),
.B(n_739),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_714),
.Y(n_779)
);

CKINVDCx20_ASAP7_75t_R g780 ( 
.A(n_714),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_664),
.B(n_678),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_734),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_719),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_693),
.Y(n_784)
);

OAI21x1_ASAP7_75t_L g785 ( 
.A1(n_710),
.A2(n_740),
.B(n_697),
.Y(n_785)
);

OAI21xp5_ASAP7_75t_L g786 ( 
.A1(n_696),
.A2(n_656),
.B(n_682),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_L g787 ( 
.A1(n_699),
.A2(n_590),
.B(n_580),
.Y(n_787)
);

NAND2x1p5_ASAP7_75t_L g788 ( 
.A(n_740),
.B(n_699),
.Y(n_788)
);

NOR2xp67_ASAP7_75t_SL g789 ( 
.A(n_685),
.B(n_629),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_685),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_705),
.Y(n_791)
);

OR2x6_ASAP7_75t_L g792 ( 
.A(n_677),
.B(n_645),
.Y(n_792)
);

INVx1_ASAP7_75t_SL g793 ( 
.A(n_705),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_SL g794 ( 
.A(n_709),
.B(n_677),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_658),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_715),
.A2(n_507),
.B1(n_727),
.B2(n_617),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_709),
.B(n_705),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_728),
.B(n_417),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_715),
.B(n_727),
.Y(n_799)
);

INVx2_ASAP7_75t_R g800 ( 
.A(n_709),
.Y(n_800)
);

O2A1O1Ixp5_ASAP7_75t_L g801 ( 
.A1(n_695),
.A2(n_663),
.B(n_732),
.C(n_731),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_661),
.Y(n_802)
);

AO21x2_ASAP7_75t_L g803 ( 
.A1(n_702),
.A2(n_694),
.B(n_731),
.Y(n_803)
);

BUFx2_ASAP7_75t_L g804 ( 
.A(n_705),
.Y(n_804)
);

NAND2x1p5_ASAP7_75t_L g805 ( 
.A(n_709),
.B(n_677),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_715),
.B(n_727),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_707),
.A2(n_590),
.B(n_580),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_685),
.Y(n_808)
);

AO31x2_ASAP7_75t_L g809 ( 
.A1(n_663),
.A2(n_694),
.A3(n_589),
.B(n_717),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_658),
.Y(n_810)
);

NAND2x1p5_ASAP7_75t_L g811 ( 
.A(n_709),
.B(n_677),
.Y(n_811)
);

AO32x2_ASAP7_75t_L g812 ( 
.A1(n_662),
.A2(n_634),
.A3(n_628),
.B1(n_691),
.B2(n_716),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_715),
.A2(n_507),
.B1(n_727),
.B2(n_617),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_750),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_745),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_792),
.B(n_797),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_792),
.A2(n_813),
.B1(n_796),
.B2(n_811),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_743),
.B(n_762),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_765),
.B(n_773),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_792),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_802),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_764),
.B(n_799),
.Y(n_822)
);

AO31x2_ASAP7_75t_L g823 ( 
.A1(n_744),
.A2(n_757),
.A3(n_777),
.B(n_761),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_764),
.B(n_759),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_805),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_769),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_813),
.A2(n_796),
.B1(n_806),
.B2(n_758),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_795),
.B(n_810),
.Y(n_828)
);

BUFx2_ASAP7_75t_L g829 ( 
.A(n_805),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_811),
.B(n_755),
.Y(n_830)
);

INVx1_ASAP7_75t_SL g831 ( 
.A(n_780),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_777),
.A2(n_752),
.B(n_758),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_766),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_785),
.Y(n_834)
);

NAND2x1_ASAP7_75t_L g835 ( 
.A(n_756),
.B(n_768),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_755),
.B(n_776),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_798),
.Y(n_837)
);

BUFx2_ASAP7_75t_L g838 ( 
.A(n_772),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_781),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_776),
.B(n_778),
.Y(n_840)
);

BUFx4f_ASAP7_75t_SL g841 ( 
.A(n_780),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_767),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_788),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_783),
.B(n_791),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_748),
.B(n_804),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_759),
.B(n_784),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_747),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_794),
.A2(n_748),
.B1(n_786),
.B2(n_800),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_746),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_760),
.B(n_791),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_751),
.Y(n_851)
);

OR2x2_ASAP7_75t_L g852 ( 
.A(n_793),
.B(n_760),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_782),
.Y(n_853)
);

AO21x2_ASAP7_75t_L g854 ( 
.A1(n_744),
.A2(n_807),
.B(n_787),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_812),
.B(n_803),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_784),
.Y(n_856)
);

OAI21x1_ASAP7_75t_L g857 ( 
.A1(n_807),
.A2(n_787),
.B(n_801),
.Y(n_857)
);

HB1xp67_ASAP7_75t_L g858 ( 
.A(n_771),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_779),
.A2(n_753),
.B1(n_763),
.B2(n_775),
.Y(n_859)
);

BUFx2_ASAP7_75t_L g860 ( 
.A(n_838),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_815),
.Y(n_861)
);

BUFx2_ASAP7_75t_SL g862 ( 
.A(n_825),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_821),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_821),
.Y(n_864)
);

INVx5_ASAP7_75t_L g865 ( 
.A(n_847),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_850),
.B(n_818),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_826),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_850),
.B(n_809),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_814),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_818),
.B(n_809),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_832),
.B(n_809),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_819),
.B(n_809),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_819),
.B(n_828),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_842),
.B(n_779),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_855),
.B(n_749),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_836),
.B(n_749),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_855),
.B(n_812),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_839),
.Y(n_878)
);

BUFx2_ASAP7_75t_SL g879 ( 
.A(n_825),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_840),
.B(n_770),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_824),
.B(n_789),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_827),
.B(n_763),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_830),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_840),
.B(n_774),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_880),
.B(n_843),
.Y(n_885)
);

INVxp67_ASAP7_75t_SL g886 ( 
.A(n_869),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_861),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_868),
.B(n_854),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_868),
.B(n_854),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_866),
.B(n_854),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_866),
.B(n_857),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_861),
.Y(n_892)
);

OR2x2_ASAP7_75t_L g893 ( 
.A(n_876),
.B(n_852),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_873),
.B(n_822),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_870),
.B(n_823),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_875),
.B(n_834),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_870),
.B(n_872),
.Y(n_897)
);

AOI211xp5_ASAP7_75t_L g898 ( 
.A1(n_882),
.A2(n_817),
.B(n_846),
.C(n_849),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_878),
.B(n_883),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_872),
.B(n_823),
.Y(n_900)
);

OR2x2_ASAP7_75t_L g901 ( 
.A(n_876),
.B(n_852),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_865),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_897),
.B(n_863),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_897),
.B(n_864),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_887),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_890),
.B(n_884),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_887),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_886),
.B(n_864),
.Y(n_908)
);

OR2x2_ASAP7_75t_L g909 ( 
.A(n_893),
.B(n_871),
.Y(n_909)
);

NAND2x1_ASAP7_75t_L g910 ( 
.A(n_902),
.B(n_860),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_892),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_890),
.B(n_884),
.Y(n_912)
);

AND2x4_ASAP7_75t_SL g913 ( 
.A(n_902),
.B(n_816),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_894),
.B(n_867),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_891),
.B(n_877),
.Y(n_915)
);

INVx4_ASAP7_75t_L g916 ( 
.A(n_885),
.Y(n_916)
);

OR2x2_ASAP7_75t_L g917 ( 
.A(n_909),
.B(n_893),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_908),
.Y(n_918)
);

NAND2xp67_ASAP7_75t_L g919 ( 
.A(n_913),
.B(n_899),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_915),
.B(n_891),
.Y(n_920)
);

AND2x2_ASAP7_75t_SL g921 ( 
.A(n_916),
.B(n_860),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_905),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_910),
.Y(n_923)
);

OR2x2_ASAP7_75t_L g924 ( 
.A(n_909),
.B(n_901),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_907),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_911),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_914),
.B(n_881),
.Y(n_927)
);

NAND2xp33_ASAP7_75t_L g928 ( 
.A(n_903),
.B(n_848),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_916),
.Y(n_929)
);

AOI22xp5_ASAP7_75t_L g930 ( 
.A1(n_928),
.A2(n_898),
.B1(n_913),
.B2(n_910),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_929),
.Y(n_931)
);

OAI31xp33_ASAP7_75t_L g932 ( 
.A1(n_923),
.A2(n_831),
.A3(n_859),
.B(n_845),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_929),
.Y(n_933)
);

OAI22xp33_ASAP7_75t_L g934 ( 
.A1(n_929),
.A2(n_916),
.B1(n_904),
.B2(n_835),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_917),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_918),
.B(n_906),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_927),
.B(n_912),
.Y(n_937)
);

AOI322xp5_ASAP7_75t_L g938 ( 
.A1(n_921),
.A2(n_915),
.A3(n_912),
.B1(n_900),
.B2(n_895),
.C1(n_889),
.C2(n_888),
.Y(n_938)
);

BUFx2_ASAP7_75t_L g939 ( 
.A(n_921),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_917),
.B(n_896),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_922),
.Y(n_941)
);

NOR3xp33_ASAP7_75t_L g942 ( 
.A(n_930),
.B(n_856),
.C(n_853),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_930),
.A2(n_928),
.B1(n_898),
.B2(n_924),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_935),
.B(n_924),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_941),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_938),
.B(n_920),
.Y(n_946)
);

INVxp33_ASAP7_75t_L g947 ( 
.A(n_939),
.Y(n_947)
);

OAI211xp5_ASAP7_75t_SL g948 ( 
.A1(n_943),
.A2(n_932),
.B(n_938),
.C(n_934),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_942),
.A2(n_933),
.B(n_931),
.Y(n_949)
);

O2A1O1Ixp5_ASAP7_75t_L g950 ( 
.A1(n_947),
.A2(n_936),
.B(n_937),
.C(n_940),
.Y(n_950)
);

NOR3x1_ASAP7_75t_L g951 ( 
.A(n_948),
.B(n_946),
.C(n_856),
.Y(n_951)
);

INVx1_ASAP7_75t_SL g952 ( 
.A(n_949),
.Y(n_952)
);

OR2x2_ASAP7_75t_L g953 ( 
.A(n_952),
.B(n_944),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_951),
.B(n_950),
.Y(n_954)
);

NOR2x1_ASAP7_75t_L g955 ( 
.A(n_953),
.B(n_841),
.Y(n_955)
);

INVx1_ASAP7_75t_SL g956 ( 
.A(n_954),
.Y(n_956)
);

NOR2x1_ASAP7_75t_L g957 ( 
.A(n_956),
.B(n_754),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_955),
.B(n_945),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_957),
.A2(n_790),
.B1(n_808),
.B2(n_858),
.Y(n_959)
);

BUFx2_ASAP7_75t_L g960 ( 
.A(n_958),
.Y(n_960)
);

OAI22x1_ASAP7_75t_SL g961 ( 
.A1(n_957),
.A2(n_851),
.B1(n_919),
.B2(n_874),
.Y(n_961)
);

INVx4_ASAP7_75t_L g962 ( 
.A(n_960),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_959),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_961),
.B(n_940),
.Y(n_964)
);

INVx1_ASAP7_75t_SL g965 ( 
.A(n_959),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_959),
.Y(n_966)
);

OAI22xp33_ASAP7_75t_L g967 ( 
.A1(n_962),
.A2(n_820),
.B1(n_829),
.B2(n_835),
.Y(n_967)
);

AND2x4_ASAP7_75t_SL g968 ( 
.A(n_966),
.B(n_816),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_963),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_965),
.A2(n_829),
.B(n_816),
.Y(n_970)
);

AO21x1_ASAP7_75t_L g971 ( 
.A1(n_964),
.A2(n_926),
.B(n_925),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_962),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_972),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_SL g974 ( 
.A1(n_970),
.A2(n_820),
.B(n_837),
.Y(n_974)
);

AO221x1_ASAP7_75t_L g975 ( 
.A1(n_967),
.A2(n_969),
.B1(n_968),
.B2(n_971),
.C(n_833),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_973),
.A2(n_862),
.B1(n_879),
.B2(n_844),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_976),
.B(n_975),
.Y(n_977)
);

OR2x6_ASAP7_75t_L g978 ( 
.A(n_977),
.B(n_974),
.Y(n_978)
);

AOI22xp33_ASAP7_75t_L g979 ( 
.A1(n_978),
.A2(n_862),
.B1(n_879),
.B2(n_920),
.Y(n_979)
);


endmodule