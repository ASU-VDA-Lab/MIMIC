module fake_jpeg_3559_n_427 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_427);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_427;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_5),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_4),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_55),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_16),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_58),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_60),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_15),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_61),
.B(n_63),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_18),
.B(n_14),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_62),
.B(n_67),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_12),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_66),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_12),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

BUFx4f_ASAP7_75t_SL g154 ( 
.A(n_68),
.Y(n_154)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_70),
.Y(n_166)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_72),
.Y(n_159)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_16),
.Y(n_73)
);

CKINVDCx9p33_ASAP7_75t_R g170 ( 
.A(n_73),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_20),
.B(n_14),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_74),
.B(n_78),
.Y(n_130)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_16),
.Y(n_75)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_75),
.Y(n_151)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_16),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_85),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_20),
.B(n_0),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_79),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_80),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_17),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_82),
.B(n_98),
.Y(n_155)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_84),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_30),
.B(n_0),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_30),
.B(n_32),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_87),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_46),
.B(n_0),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

BUFx10_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_89),
.Y(n_173)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_17),
.Y(n_91)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_91),
.Y(n_157)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_92),
.Y(n_174)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_93),
.Y(n_176)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_17),
.Y(n_94)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_94),
.Y(n_177)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_95),
.Y(n_165)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_96),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_32),
.B(n_53),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_102),
.Y(n_118)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_99),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_100),
.Y(n_138)
);

HAxp5_ASAP7_75t_SL g101 ( 
.A(n_52),
.B(n_1),
.CON(n_101),
.SN(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_101),
.A2(n_54),
.B(n_21),
.C(n_31),
.Y(n_139)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_104),
.Y(n_135)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_38),
.Y(n_104)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx11_ASAP7_75t_L g161 ( 
.A(n_105),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_108),
.Y(n_140)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_107),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_38),
.B(n_1),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_111),
.Y(n_145)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

INVx11_ASAP7_75t_L g168 ( 
.A(n_110),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_44),
.B(n_1),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_111),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_112),
.B(n_121),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_78),
.A2(n_31),
.B1(n_45),
.B2(n_42),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_116),
.A2(n_131),
.B1(n_134),
.B2(n_137),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_44),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_57),
.A2(n_52),
.B1(n_53),
.B2(n_47),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_123),
.A2(n_24),
.B1(n_8),
.B2(n_9),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_63),
.A2(n_47),
.B1(n_43),
.B2(n_33),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g228 ( 
.A1(n_125),
.A2(n_126),
.B1(n_161),
.B2(n_159),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_67),
.A2(n_36),
.B1(n_45),
.B2(n_42),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_86),
.B(n_26),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_133),
.B(n_147),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_59),
.A2(n_37),
.B1(n_36),
.B2(n_35),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_82),
.A2(n_50),
.B1(n_26),
.B2(n_43),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_97),
.A2(n_54),
.B1(n_37),
.B2(n_35),
.Y(n_137)
);

AOI21xp33_ASAP7_75t_L g187 ( 
.A1(n_139),
.A2(n_130),
.B(n_133),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_65),
.A2(n_79),
.B1(n_68),
.B2(n_80),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_143),
.A2(n_154),
.B1(n_173),
.B2(n_120),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_61),
.B(n_29),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_58),
.A2(n_33),
.B1(n_19),
.B2(n_27),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_148),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_73),
.B(n_29),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_149),
.B(n_156),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_75),
.B(n_21),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_69),
.B(n_27),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_158),
.B(n_164),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_81),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_89),
.A2(n_23),
.B1(n_19),
.B2(n_24),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_167),
.A2(n_171),
.B1(n_128),
.B2(n_154),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_99),
.A2(n_23),
.B1(n_24),
.B2(n_5),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_112),
.B(n_100),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_179),
.B(n_187),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_101),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_180),
.B(n_181),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_1),
.Y(n_181)
);

O2A1O1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_139),
.A2(n_24),
.B(n_7),
.C(n_8),
.Y(n_182)
);

A2O1A1Ixp33_ASAP7_75t_L g238 ( 
.A1(n_182),
.A2(n_192),
.B(n_218),
.C(n_180),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_183),
.A2(n_207),
.B1(n_219),
.B2(n_221),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_125),
.A2(n_4),
.B1(n_24),
.B2(n_140),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_184),
.A2(n_232),
.B1(n_196),
.B2(n_190),
.Y(n_269)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_127),
.Y(n_185)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_185),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_145),
.A2(n_4),
.B1(n_150),
.B2(n_121),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_186),
.A2(n_204),
.B(n_181),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_170),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_188),
.B(n_195),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_118),
.B(n_135),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_189),
.B(n_209),
.Y(n_254)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_132),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_190),
.Y(n_263)
);

BUFx8_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

INVx5_ASAP7_75t_SL g248 ( 
.A(n_191),
.Y(n_248)
);

A2O1A1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_117),
.A2(n_146),
.B(n_113),
.C(n_155),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_122),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_193),
.Y(n_247)
);

AND2x2_ASAP7_75t_SL g194 ( 
.A(n_157),
.B(n_169),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_194),
.B(n_196),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_153),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_132),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_142),
.B(n_165),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_214),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_141),
.B(n_152),
.C(n_177),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_199),
.B(n_211),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_144),
.A2(n_175),
.B1(n_162),
.B2(n_115),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_201),
.A2(n_208),
.B1(n_217),
.B2(n_191),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_151),
.B(n_141),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_202),
.Y(n_261)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_124),
.Y(n_203)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

OR2x2_ASAP7_75t_SL g204 ( 
.A(n_152),
.B(n_177),
.Y(n_204)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_122),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g244 ( 
.A(n_206),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_123),
.A2(n_119),
.B1(n_124),
.B2(n_129),
.Y(n_207)
);

AOI22x1_ASAP7_75t_L g208 ( 
.A1(n_143),
.A2(n_115),
.B1(n_162),
.B2(n_175),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_114),
.B(n_138),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_119),
.Y(n_210)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_176),
.C(n_151),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_129),
.Y(n_213)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_213),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_172),
.B(n_176),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_174),
.Y(n_215)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_128),
.Y(n_216)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_216),
.Y(n_273)
);

O2A1O1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_126),
.A2(n_154),
.B(n_166),
.C(n_160),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_174),
.Y(n_220)
);

INVxp33_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_160),
.A2(n_163),
.B1(n_166),
.B2(n_120),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_163),
.B(n_173),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_222),
.B(n_202),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_168),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_226),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_168),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_126),
.Y(n_227)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_228),
.B(n_231),
.Y(n_272)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_126),
.Y(n_229)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_229),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_159),
.Y(n_230)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_230),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_161),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_162),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_179),
.A2(n_200),
.B1(n_178),
.B2(n_217),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_234),
.A2(n_227),
.B1(n_216),
.B2(n_230),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_237),
.B(n_238),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_207),
.A2(n_183),
.B1(n_212),
.B2(n_200),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_242),
.A2(n_245),
.B1(n_260),
.B2(n_266),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_180),
.A2(n_178),
.B1(n_208),
.B2(n_189),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_197),
.B(n_192),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_249),
.B(n_264),
.C(n_274),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_250),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_186),
.A2(n_182),
.B1(n_225),
.B2(n_209),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_255),
.A2(n_268),
.B1(n_235),
.B2(n_272),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_205),
.A2(n_181),
.B(n_204),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_257),
.B(n_258),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_228),
.A2(n_194),
.B(n_202),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_208),
.A2(n_221),
.B1(n_228),
.B2(n_199),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_262),
.B(n_251),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_228),
.A2(n_194),
.B(n_224),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_211),
.A2(n_210),
.B1(n_222),
.B2(n_232),
.Y(n_266)
);

FAx1_ASAP7_75t_SL g267 ( 
.A(n_218),
.B(n_191),
.CI(n_222),
.CON(n_267),
.SN(n_267)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_258),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_269),
.A2(n_270),
.B1(n_261),
.B2(n_236),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_203),
.A2(n_213),
.B1(n_206),
.B2(n_193),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_253),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_275),
.B(n_287),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_220),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_278),
.B(n_298),
.Y(n_321)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_241),
.Y(n_279)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_279),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_280),
.A2(n_287),
.B1(n_289),
.B2(n_276),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_242),
.A2(n_234),
.B1(n_272),
.B2(n_260),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_281),
.A2(n_299),
.B1(n_301),
.B2(n_244),
.Y(n_313)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_240),
.Y(n_282)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_282),
.Y(n_330)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_283),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_284),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_285),
.A2(n_277),
.B1(n_303),
.B2(n_305),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_254),
.B(n_233),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_286),
.B(n_307),
.Y(n_312)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_261),
.Y(n_287)
);

OAI211xp5_ASAP7_75t_L g288 ( 
.A1(n_235),
.A2(n_245),
.B(n_257),
.C(n_238),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_288),
.B(n_289),
.Y(n_319)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_246),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_290),
.B(n_294),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_239),
.B(n_249),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_291),
.B(n_296),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_292),
.A2(n_293),
.B(n_294),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_266),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_251),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_259),
.B(n_252),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_243),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_297),
.B(n_306),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_264),
.B(n_268),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_236),
.A2(n_268),
.B1(n_274),
.B2(n_250),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_295),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_241),
.A2(n_267),
.B1(n_256),
.B2(n_247),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_246),
.B(n_256),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_302),
.B(n_305),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_244),
.Y(n_304)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_304),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_267),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_271),
.B(n_273),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_263),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_308),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_281),
.A2(n_263),
.B1(n_248),
.B2(n_244),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_310),
.A2(n_323),
.B1(n_327),
.B2(n_304),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_313),
.A2(n_320),
.B1(n_326),
.B2(n_308),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_277),
.A2(n_248),
.B(n_244),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_314),
.A2(n_326),
.B(n_331),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_316),
.A2(n_323),
.B1(n_314),
.B2(n_310),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_317),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_277),
.A2(n_292),
.B1(n_299),
.B2(n_298),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_293),
.A2(n_278),
.B1(n_295),
.B2(n_290),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_324),
.B(n_331),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_293),
.A2(n_290),
.B(n_301),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_294),
.A2(n_300),
.B1(n_280),
.B2(n_302),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_279),
.B(n_283),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_328),
.B(n_332),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_282),
.B(n_307),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_328),
.Y(n_334)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_334),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_335),
.Y(n_362)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_332),
.Y(n_336)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_336),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_337),
.A2(n_340),
.B1(n_344),
.B2(n_346),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_338),
.B(n_349),
.C(n_344),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_318),
.Y(n_339)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_339),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_313),
.A2(n_320),
.B1(n_321),
.B2(n_319),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_329),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_341),
.B(n_351),
.Y(n_360)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_333),
.Y(n_342)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_342),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_322),
.B(n_318),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_343),
.B(n_345),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_316),
.A2(n_319),
.B1(n_321),
.B2(n_327),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_322),
.B(n_329),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_347),
.A2(n_309),
.B(n_346),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_312),
.B(n_315),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_312),
.B(n_315),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_352),
.B(n_353),
.Y(n_363)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_333),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_325),
.B(n_317),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_354),
.B(n_330),
.Y(n_364)
);

OA21x2_ASAP7_75t_L g355 ( 
.A1(n_330),
.A2(n_309),
.B(n_325),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_355),
.B(n_350),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_311),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_359),
.B(n_364),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_338),
.B(n_324),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_361),
.B(n_369),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_366),
.B(n_368),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_339),
.B(n_354),
.Y(n_367)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_367),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_343),
.B(n_340),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_372),
.B(n_335),
.C(n_355),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_347),
.A2(n_337),
.B(n_340),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_373),
.B(n_355),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_360),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_376),
.B(n_378),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_377),
.B(n_380),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_362),
.A2(n_337),
.B1(n_350),
.B2(n_336),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_362),
.A2(n_350),
.B1(n_334),
.B2(n_345),
.Y(n_380)
);

A2O1A1Ixp33_ASAP7_75t_SL g390 ( 
.A1(n_381),
.A2(n_374),
.B(n_386),
.C(n_378),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_370),
.A2(n_351),
.B1(n_352),
.B2(n_348),
.Y(n_383)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_383),
.Y(n_393)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_360),
.Y(n_384)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_384),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_370),
.A2(n_355),
.B1(n_348),
.B2(n_353),
.Y(n_385)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_385),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_373),
.A2(n_342),
.B1(n_355),
.B2(n_368),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_386),
.B(n_387),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_372),
.A2(n_366),
.B1(n_356),
.B2(n_357),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_382),
.Y(n_389)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_389),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_390),
.A2(n_397),
.B1(n_385),
.B2(n_374),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_375),
.B(n_361),
.C(n_369),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_396),
.B(n_375),
.C(n_365),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_374),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_381),
.A2(n_356),
.B(n_357),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_398),
.A2(n_365),
.B(n_363),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_399),
.B(n_400),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_396),
.B(n_377),
.C(n_387),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_SL g410 ( 
.A1(n_401),
.A2(n_390),
.B1(n_388),
.B2(n_394),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_391),
.B(n_380),
.C(n_379),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_402),
.B(n_404),
.Y(n_409)
);

AOI21x1_ASAP7_75t_SL g408 ( 
.A1(n_403),
.A2(n_398),
.B(n_363),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_391),
.B(n_383),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_392),
.B(n_388),
.Y(n_406)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_406),
.Y(n_413)
);

OAI21xp33_ASAP7_75t_SL g407 ( 
.A1(n_406),
.A2(n_395),
.B(n_393),
.Y(n_407)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_407),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_408),
.A2(n_402),
.B(n_358),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_410),
.A2(n_404),
.B1(n_413),
.B2(n_400),
.Y(n_417)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_405),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_412),
.B(n_371),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_414),
.A2(n_417),
.B1(n_390),
.B2(n_371),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_416),
.B(n_418),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_411),
.B(n_399),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_414),
.A2(n_410),
.B1(n_409),
.B2(n_407),
.Y(n_419)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_419),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_420),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_422),
.A2(n_421),
.B(n_420),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_424),
.B(n_423),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_425),
.B(n_415),
.Y(n_426)
);

BUFx24_ASAP7_75t_SL g427 ( 
.A(n_426),
.Y(n_427)
);


endmodule