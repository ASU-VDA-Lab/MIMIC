module fake_ariane_3073_n_1884 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1884);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1884;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1769;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_186),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_150),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_77),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_160),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_79),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_8),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_137),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_112),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_157),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_128),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_12),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_188),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_129),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_51),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g205 ( 
.A(n_38),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_74),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_16),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_122),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_176),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_23),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_149),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_116),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_94),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_169),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_88),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_105),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_25),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

INVxp67_ASAP7_75t_SL g219 ( 
.A(n_46),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_138),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_90),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_68),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_104),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_56),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_184),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_162),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_168),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_108),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_113),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_0),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_161),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_45),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_182),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_120),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_67),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_93),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_78),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_38),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_25),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_139),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_42),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_174),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_158),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_19),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_82),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_36),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_115),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_66),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_170),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_64),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_69),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_27),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_111),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_32),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_89),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_52),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_41),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_81),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_136),
.Y(n_259)
);

BUFx10_ASAP7_75t_L g260 ( 
.A(n_86),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_62),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_1),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_187),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_42),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_106),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_164),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_15),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_62),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_103),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_75),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_9),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_178),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_132),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_180),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_144),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_34),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_33),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_101),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_97),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_151),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_14),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_20),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_84),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_147),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_172),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_9),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_109),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_119),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_146),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_131),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_24),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_121),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_145),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_142),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_71),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_1),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_91),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_171),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_185),
.Y(n_299)
);

BUFx10_ASAP7_75t_L g300 ( 
.A(n_33),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_167),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_117),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_102),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_73),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g305 ( 
.A(n_16),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_20),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_166),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_51),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_46),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_165),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_54),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_59),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_28),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_3),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_13),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_130),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_7),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_179),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_7),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_2),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_58),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_17),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_54),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_50),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_76),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_177),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_63),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_87),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_13),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_14),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_32),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_40),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_27),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_85),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_6),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_127),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_154),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_183),
.Y(n_338)
);

BUFx10_ASAP7_75t_L g339 ( 
.A(n_148),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_133),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_24),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_3),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_28),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_80),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_29),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_100),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_15),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_110),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_163),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_95),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_118),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_10),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_18),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_4),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_12),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_55),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_53),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_65),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_35),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_99),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_181),
.Y(n_361)
);

BUFx10_ASAP7_75t_L g362 ( 
.A(n_17),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_18),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_125),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_141),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_21),
.Y(n_366)
);

BUFx10_ASAP7_75t_L g367 ( 
.A(n_45),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_114),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_36),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_55),
.Y(n_370)
);

BUFx10_ASAP7_75t_L g371 ( 
.A(n_53),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_135),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_6),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_156),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_37),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_70),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_47),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_152),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_22),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_10),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_34),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_59),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_57),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_155),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_19),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_315),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_201),
.Y(n_387)
);

INVxp33_ASAP7_75t_SL g388 ( 
.A(n_363),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_315),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_273),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_315),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_274),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_200),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_314),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_238),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_286),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_267),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_241),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_286),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_286),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_244),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_286),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_281),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_342),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_373),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_279),
.B(n_2),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_267),
.B(n_4),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_254),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_256),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_257),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_261),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_194),
.B(n_5),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_262),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_205),
.B(n_5),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_276),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_205),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_222),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_277),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_282),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_291),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_286),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_245),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_264),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_221),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_264),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_308),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_333),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_311),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_333),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_312),
.Y(n_430)
);

NOR2xp67_ASAP7_75t_L g431 ( 
.A(n_306),
.B(n_8),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_354),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_195),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_293),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_317),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_354),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_195),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_379),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_202),
.B(n_211),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_323),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_297),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_376),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_260),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_324),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_379),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_381),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_381),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_327),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_260),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_218),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_260),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_339),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_229),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_329),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_330),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g456 ( 
.A(n_207),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_216),
.B(n_11),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_221),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_229),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_339),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_339),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_204),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_331),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_205),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_223),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_204),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_223),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_348),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_217),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_348),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_231),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_231),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_210),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_R g474 ( 
.A(n_235),
.B(n_126),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_300),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_316),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_316),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_300),
.Y(n_478)
);

INVxp67_ASAP7_75t_SL g479 ( 
.A(n_224),
.Y(n_479)
);

INVxp33_ASAP7_75t_SL g480 ( 
.A(n_217),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_300),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_239),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_332),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_340),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_340),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_346),
.Y(n_486)
);

AND2x6_ASAP7_75t_L g487 ( 
.A(n_468),
.B(n_346),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_468),
.B(n_220),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_393),
.B(n_230),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_386),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_397),
.B(n_305),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_386),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_390),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_392),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_417),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_396),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_387),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_389),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_389),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_422),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_434),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_391),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_421),
.Y(n_503)
);

AND2x2_ASAP7_75t_SL g504 ( 
.A(n_414),
.B(n_460),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_460),
.B(n_190),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_424),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_424),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_403),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_441),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_R g510 ( 
.A(n_395),
.B(n_237),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_399),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_404),
.Y(n_512)
);

NAND2xp33_ASAP7_75t_L g513 ( 
.A(n_398),
.B(n_385),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_424),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_442),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_458),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_401),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_456),
.B(n_305),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_R g519 ( 
.A(n_408),
.B(n_247),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_458),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_409),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_468),
.B(n_236),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_421),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_410),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_411),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_399),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_413),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_400),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_414),
.B(n_263),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_415),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_442),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_400),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_402),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_465),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_473),
.B(n_305),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_443),
.B(n_230),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_402),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_479),
.B(n_362),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_418),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_449),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_450),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_419),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_433),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_450),
.Y(n_544)
);

AND2x6_ASAP7_75t_L g545 ( 
.A(n_453),
.B(n_215),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_453),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_459),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_471),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_471),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_472),
.B(n_263),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_472),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_439),
.B(n_240),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_476),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_420),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_476),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_426),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_R g557 ( 
.A(n_428),
.B(n_248),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_477),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_430),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_435),
.Y(n_560)
);

OR2x6_ASAP7_75t_L g561 ( 
.A(n_406),
.B(n_309),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_526),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_561),
.A2(n_552),
.B1(n_505),
.B2(n_543),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_491),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_561),
.A2(n_480),
.B1(n_388),
.B2(n_444),
.Y(n_565)
);

INVxp67_ASAP7_75t_SL g566 ( 
.A(n_488),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_528),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_529),
.B(n_440),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_490),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_492),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_498),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_529),
.B(n_475),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_499),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_510),
.B(n_448),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_528),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_532),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_491),
.B(n_454),
.Y(n_577)
);

AND3x4_ASAP7_75t_L g578 ( 
.A(n_529),
.B(n_431),
.C(n_475),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_511),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_518),
.B(n_455),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_532),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_533),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_526),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_529),
.B(n_482),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_493),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_511),
.Y(n_586)
);

NAND2x1p5_ASAP7_75t_L g587 ( 
.A(n_504),
.B(n_299),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_526),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_506),
.Y(n_589)
);

NAND2xp33_ASAP7_75t_L g590 ( 
.A(n_519),
.B(n_463),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_561),
.A2(n_457),
.B1(n_412),
.B2(n_405),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_507),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_544),
.Y(n_593)
);

BUFx4f_ASAP7_75t_L g594 ( 
.A(n_487),
.Y(n_594)
);

AO22x2_ASAP7_75t_L g595 ( 
.A1(n_518),
.A2(n_416),
.B1(n_478),
.B2(n_464),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_535),
.B(n_483),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_526),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_561),
.A2(n_550),
.B1(n_504),
.B2(n_538),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_533),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_514),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_537),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_535),
.B(n_467),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_537),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_508),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_538),
.B(n_513),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_L g606 ( 
.A(n_557),
.B(n_215),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_502),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_561),
.A2(n_394),
.B1(n_407),
.B2(n_437),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_516),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_493),
.Y(n_610)
);

INVx5_ASAP7_75t_L g611 ( 
.A(n_545),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_504),
.B(n_462),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_487),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_522),
.B(n_470),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_526),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_487),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_550),
.A2(n_466),
.B1(n_469),
.B2(n_431),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_517),
.B(n_190),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_520),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_544),
.Y(n_620)
);

BUFx10_ASAP7_75t_L g621 ( 
.A(n_517),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_544),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_487),
.Y(n_623)
);

AND2x6_ASAP7_75t_L g624 ( 
.A(n_553),
.B(n_215),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_548),
.A2(n_271),
.B1(n_246),
.B2(n_252),
.Y(n_625)
);

OR2x6_ASAP7_75t_L g626 ( 
.A(n_521),
.B(n_423),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_541),
.B(n_423),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_496),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_544),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_525),
.B(n_451),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_546),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_549),
.A2(n_356),
.B1(n_268),
.B2(n_296),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_546),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_546),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_546),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_546),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_541),
.B(n_484),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_551),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_551),
.A2(n_320),
.B1(n_353),
.B2(n_375),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_551),
.A2(n_366),
.B1(n_313),
.B2(n_321),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_521),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_541),
.B(n_485),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_553),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_551),
.Y(n_644)
);

INVx1_ASAP7_75t_SL g645 ( 
.A(n_512),
.Y(n_645)
);

BUFx8_ASAP7_75t_SL g646 ( 
.A(n_515),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_551),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_523),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_555),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_531),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_524),
.A2(n_347),
.B1(n_369),
.B2(n_359),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_555),
.B(n_485),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_534),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_547),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_494),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_523),
.Y(n_656)
);

INVx4_ASAP7_75t_L g657 ( 
.A(n_487),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_523),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_524),
.B(n_527),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_489),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_487),
.A2(n_380),
.B1(n_352),
.B2(n_322),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_527),
.B(n_191),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_555),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_523),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_547),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_523),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_489),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_558),
.B(n_486),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_530),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_530),
.B(n_191),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_503),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_539),
.B(n_452),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_558),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_SL g674 ( 
.A(n_539),
.B(n_542),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_494),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_542),
.B(n_461),
.Y(n_676)
);

INVx4_ASAP7_75t_L g677 ( 
.A(n_545),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_545),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_503),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_SL g680 ( 
.A1(n_536),
.A2(n_481),
.B1(n_357),
.B2(n_355),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_554),
.B(n_192),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_554),
.B(n_556),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_503),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_545),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_545),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_545),
.A2(n_486),
.B1(n_319),
.B2(n_219),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_556),
.B(n_425),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_545),
.Y(n_688)
);

AO22x2_ASAP7_75t_L g689 ( 
.A1(n_534),
.A2(n_345),
.B1(n_299),
.B2(n_365),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_559),
.B(n_232),
.Y(n_690)
);

NOR2x1p5_ASAP7_75t_L g691 ( 
.A(n_559),
.B(n_232),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_560),
.B(n_425),
.Y(n_692)
);

OR2x6_ASAP7_75t_L g693 ( 
.A(n_495),
.B(n_427),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_495),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_497),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_497),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_500),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_500),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_501),
.B(n_192),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_641),
.B(n_501),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_566),
.B(n_605),
.Y(n_701)
);

NOR3xp33_ASAP7_75t_L g702 ( 
.A(n_563),
.B(n_347),
.C(n_343),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_564),
.B(n_335),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_564),
.B(n_341),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_580),
.B(n_343),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_669),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_614),
.B(n_509),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_584),
.B(n_272),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_596),
.A2(n_234),
.B1(n_198),
.B2(n_214),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_584),
.B(n_302),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_626),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_593),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_577),
.B(n_193),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_584),
.B(n_193),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_627),
.B(n_196),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_579),
.Y(n_716)
);

NAND3xp33_ASAP7_75t_L g717 ( 
.A(n_659),
.B(n_357),
.C(n_355),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_626),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_579),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_593),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_586),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_641),
.B(n_196),
.Y(n_722)
);

OR2x6_ASAP7_75t_L g723 ( 
.A(n_693),
.B(n_429),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_586),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_654),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_598),
.A2(n_360),
.B1(n_197),
.B2(n_198),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_626),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_568),
.B(n_359),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_665),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_665),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_578),
.A2(n_362),
.B1(n_367),
.B2(n_371),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_627),
.B(n_197),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_602),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_687),
.B(n_199),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_687),
.B(n_199),
.Y(n_735)
);

HB1xp67_ASAP7_75t_L g736 ( 
.A(n_626),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_692),
.B(n_509),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_578),
.A2(n_214),
.B1(n_203),
.B2(n_206),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_587),
.B(n_369),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_587),
.B(n_370),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_569),
.B(n_208),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_587),
.B(n_572),
.Y(n_742)
);

NAND3xp33_ASAP7_75t_L g743 ( 
.A(n_674),
.B(n_377),
.C(n_370),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_565),
.B(n_208),
.Y(n_744)
);

OR2x6_ASAP7_75t_L g745 ( 
.A(n_693),
.B(n_429),
.Y(n_745)
);

O2A1O1Ixp33_ASAP7_75t_L g746 ( 
.A1(n_643),
.A2(n_432),
.B(n_447),
.C(n_446),
.Y(n_746)
);

INVxp67_ASAP7_75t_L g747 ( 
.A(n_604),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_572),
.B(n_209),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_649),
.B(n_209),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_663),
.B(n_570),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_669),
.B(n_212),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_571),
.B(n_212),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_573),
.B(n_213),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_673),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_690),
.B(n_536),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_620),
.A2(n_255),
.B(n_337),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_693),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_683),
.Y(n_758)
);

NAND3xp33_ASAP7_75t_L g759 ( 
.A(n_590),
.B(n_382),
.C(n_377),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_593),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_589),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_690),
.B(n_540),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_618),
.B(n_382),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_607),
.B(n_225),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_612),
.A2(n_227),
.B1(n_226),
.B2(n_344),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_662),
.B(n_383),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_621),
.B(n_362),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_621),
.B(n_227),
.Y(n_768)
);

AO221x1_ASAP7_75t_L g769 ( 
.A1(n_689),
.A2(n_215),
.B1(n_303),
.B2(n_325),
.C(n_307),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_693),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_694),
.Y(n_771)
);

AND2x2_ASAP7_75t_SL g772 ( 
.A(n_606),
.B(n_242),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_670),
.B(n_383),
.Y(n_773)
);

OR2x6_ASAP7_75t_L g774 ( 
.A(n_697),
.B(n_432),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_621),
.B(n_228),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_592),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_612),
.B(n_233),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_574),
.B(n_233),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_585),
.B(n_344),
.Y(n_779)
);

A2O1A1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_591),
.A2(n_258),
.B(n_292),
.C(n_310),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_585),
.B(n_351),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_592),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_600),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_600),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_668),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_681),
.B(n_367),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_609),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_619),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_610),
.B(n_358),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_619),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_593),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_671),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_699),
.B(n_367),
.Y(n_793)
);

OR2x6_ASAP7_75t_L g794 ( 
.A(n_697),
.B(n_436),
.Y(n_794)
);

NAND2x1p5_ASAP7_75t_L g795 ( 
.A(n_613),
.B(n_243),
.Y(n_795)
);

BUFx8_ASAP7_75t_L g796 ( 
.A(n_650),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_638),
.B(n_371),
.Y(n_797)
);

INVx4_ASAP7_75t_L g798 ( 
.A(n_613),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_683),
.Y(n_799)
);

BUFx8_ASAP7_75t_L g800 ( 
.A(n_650),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_610),
.B(n_361),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_590),
.A2(n_606),
.B1(n_595),
.B2(n_608),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_646),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_628),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_637),
.B(n_361),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_671),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_655),
.B(n_675),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_628),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_655),
.B(n_364),
.Y(n_809)
);

OAI22xp33_ASAP7_75t_L g810 ( 
.A1(n_675),
.A2(n_447),
.B1(n_446),
.B2(n_445),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_638),
.B(n_371),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_697),
.B(n_364),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_697),
.B(n_368),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_679),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_697),
.B(n_368),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_694),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_653),
.B(n_374),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_642),
.B(n_652),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_679),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_617),
.B(n_384),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_647),
.B(n_384),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_683),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_682),
.B(n_474),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_595),
.A2(n_265),
.B1(n_266),
.B2(n_250),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_647),
.B(n_280),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_645),
.Y(n_826)
);

INVxp67_ASAP7_75t_L g827 ( 
.A(n_672),
.Y(n_827)
);

NOR2xp67_ASAP7_75t_L g828 ( 
.A(n_676),
.B(n_436),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_696),
.B(n_249),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_647),
.B(n_284),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_567),
.B(n_251),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_575),
.B(n_253),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_689),
.A2(n_445),
.B1(n_438),
.B2(n_378),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_689),
.A2(n_438),
.B1(n_372),
.B2(n_350),
.Y(n_834)
);

OR2x2_ASAP7_75t_L g835 ( 
.A(n_696),
.B(n_11),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_695),
.B(n_630),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_691),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_695),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_576),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_576),
.B(n_259),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_581),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_581),
.B(n_269),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_651),
.B(n_270),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_582),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_701),
.B(n_595),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_818),
.A2(n_636),
.B(n_620),
.Y(n_846)
);

O2A1O1Ixp5_ASAP7_75t_L g847 ( 
.A1(n_705),
.A2(n_615),
.B(n_562),
.C(n_597),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_798),
.A2(n_636),
.B(n_622),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_712),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_798),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_705),
.B(n_595),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_750),
.A2(n_622),
.B(n_629),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_706),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_733),
.B(n_698),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_733),
.B(n_646),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_716),
.A2(n_644),
.B(n_629),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_785),
.B(n_689),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_719),
.A2(n_594),
.B(n_633),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_721),
.A2(n_594),
.B(n_633),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_723),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_827),
.B(n_680),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_724),
.A2(n_594),
.B(n_635),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_758),
.A2(n_822),
.B(n_799),
.Y(n_863)
);

O2A1O1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_827),
.A2(n_836),
.B(n_780),
.C(n_702),
.Y(n_864)
);

OAI321xp33_ASAP7_75t_L g865 ( 
.A1(n_824),
.A2(n_625),
.A3(n_632),
.B1(n_640),
.B2(n_639),
.C(n_661),
.Y(n_865)
);

OAI21xp5_ASAP7_75t_L g866 ( 
.A1(n_725),
.A2(n_635),
.B(n_634),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_742),
.B(n_728),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_707),
.B(n_660),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_747),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_761),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_729),
.A2(n_631),
.B(n_588),
.Y(n_871)
);

NAND2xp33_ASAP7_75t_SL g872 ( 
.A(n_838),
.B(n_711),
.Y(n_872)
);

O2A1O1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_702),
.A2(n_597),
.B(n_588),
.C(n_615),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_747),
.B(n_660),
.Y(n_874)
);

OAI321xp33_ASAP7_75t_L g875 ( 
.A1(n_834),
.A2(n_686),
.A3(n_349),
.B1(n_287),
.B2(n_294),
.C(n_336),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_737),
.B(n_667),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_742),
.B(n_728),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_700),
.B(n_755),
.Y(n_878)
);

OAI21xp5_ASAP7_75t_L g879 ( 
.A1(n_730),
.A2(n_631),
.B(n_562),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_821),
.A2(n_597),
.B(n_583),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_708),
.B(n_582),
.Y(n_881)
);

HB1xp67_ASAP7_75t_L g882 ( 
.A(n_723),
.Y(n_882)
);

O2A1O1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_810),
.A2(n_583),
.B(n_599),
.C(n_601),
.Y(n_883)
);

BUFx12f_ASAP7_75t_L g884 ( 
.A(n_796),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_710),
.B(n_599),
.Y(n_885)
);

AOI21x1_ASAP7_75t_L g886 ( 
.A1(n_841),
.A2(n_658),
.B(n_648),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_776),
.A2(n_783),
.B1(n_784),
.B2(n_782),
.Y(n_887)
);

OAI321xp33_ASAP7_75t_L g888 ( 
.A1(n_834),
.A2(n_601),
.A3(n_603),
.B1(n_215),
.B2(n_303),
.C(n_666),
.Y(n_888)
);

BUFx12f_ASAP7_75t_L g889 ( 
.A(n_796),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_754),
.A2(n_664),
.B(n_666),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_712),
.Y(n_891)
);

OAI21xp33_ASAP7_75t_L g892 ( 
.A1(n_709),
.A2(n_603),
.B(n_683),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_718),
.B(n_613),
.Y(n_893)
);

NAND2x1p5_ASAP7_75t_L g894 ( 
.A(n_727),
.B(n_616),
.Y(n_894)
);

NOR2x1p5_ASAP7_75t_SL g895 ( 
.A(n_792),
.B(n_806),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_826),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_800),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_715),
.B(n_683),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_749),
.A2(n_732),
.B(n_814),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_819),
.A2(n_805),
.B(n_741),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_712),
.Y(n_901)
);

O2A1O1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_810),
.A2(n_684),
.B(n_685),
.C(n_678),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_712),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_720),
.Y(n_904)
);

O2A1O1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_734),
.A2(n_684),
.B(n_678),
.C(n_23),
.Y(n_905)
);

O2A1O1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_735),
.A2(n_678),
.B(n_22),
.C(n_26),
.Y(n_906)
);

AO22x1_ASAP7_75t_L g907 ( 
.A1(n_800),
.A2(n_667),
.B1(n_624),
.B2(n_688),
.Y(n_907)
);

AND2x6_ASAP7_75t_L g908 ( 
.A(n_802),
.B(n_688),
.Y(n_908)
);

INVx11_ASAP7_75t_L g909 ( 
.A(n_803),
.Y(n_909)
);

INVxp67_ASAP7_75t_SL g910 ( 
.A(n_736),
.Y(n_910)
);

A2O1A1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_739),
.A2(n_656),
.B(n_688),
.C(n_304),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_SL g912 ( 
.A(n_772),
.B(n_623),
.Y(n_912)
);

A2O1A1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_739),
.A2(n_656),
.B(n_688),
.C(n_318),
.Y(n_913)
);

NAND2x1_ASAP7_75t_L g914 ( 
.A(n_720),
.B(n_657),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_713),
.A2(n_656),
.B(n_677),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_752),
.A2(n_298),
.B(n_278),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_723),
.B(n_21),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_763),
.A2(n_26),
.B(n_29),
.C(n_30),
.Y(n_918)
);

BUFx4f_ASAP7_75t_L g919 ( 
.A(n_745),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_740),
.B(n_828),
.Y(n_920)
);

NAND3xp33_ASAP7_75t_L g921 ( 
.A(n_763),
.B(n_275),
.C(n_283),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_740),
.B(n_703),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_L g923 ( 
.A1(n_825),
.A2(n_624),
.B(n_611),
.Y(n_923)
);

AOI21x1_ASAP7_75t_L g924 ( 
.A1(n_839),
.A2(n_624),
.B(n_303),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_757),
.B(n_285),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_745),
.Y(n_926)
);

AND2x2_ASAP7_75t_SL g927 ( 
.A(n_772),
.B(n_731),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_703),
.B(n_624),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_704),
.B(n_624),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_704),
.B(n_288),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_714),
.B(n_289),
.Y(n_931)
);

NOR3xp33_ASAP7_75t_L g932 ( 
.A(n_807),
.B(n_290),
.C(n_295),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_771),
.B(n_301),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_753),
.A2(n_338),
.B(n_334),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_726),
.A2(n_328),
.B1(n_326),
.B2(n_611),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_816),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_764),
.A2(n_611),
.B(n_83),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_745),
.B(n_30),
.Y(n_938)
);

AND2x6_ASAP7_75t_L g939 ( 
.A(n_720),
.B(n_72),
.Y(n_939)
);

NOR2x1p5_ASAP7_75t_L g940 ( 
.A(n_762),
.B(n_31),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_817),
.B(n_31),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_787),
.B(n_37),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_788),
.B(n_39),
.Y(n_943)
);

INVxp67_ASAP7_75t_L g944 ( 
.A(n_767),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_770),
.B(n_39),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_765),
.B(n_40),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_774),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_774),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_790),
.B(n_41),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_777),
.B(n_43),
.Y(n_950)
);

O2A1O1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_766),
.A2(n_43),
.B(n_44),
.C(n_47),
.Y(n_951)
);

O2A1O1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_766),
.A2(n_773),
.B(n_748),
.C(n_809),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_797),
.B(n_44),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_738),
.B(n_48),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_773),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_955)
);

A2O1A1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_786),
.A2(n_49),
.B(n_52),
.C(n_56),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_L g957 ( 
.A1(n_795),
.A2(n_57),
.B1(n_58),
.B2(n_60),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_720),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_797),
.B(n_60),
.Y(n_959)
);

INVx1_ASAP7_75t_SL g960 ( 
.A(n_774),
.Y(n_960)
);

INVx4_ASAP7_75t_L g961 ( 
.A(n_794),
.Y(n_961)
);

BUFx2_ASAP7_75t_L g962 ( 
.A(n_794),
.Y(n_962)
);

OAI21xp33_ASAP7_75t_L g963 ( 
.A1(n_786),
.A2(n_61),
.B(n_63),
.Y(n_963)
);

INVxp67_ASAP7_75t_SL g964 ( 
.A(n_760),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_744),
.B(n_61),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_825),
.A2(n_92),
.B(n_96),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_L g967 ( 
.A1(n_795),
.A2(n_794),
.B1(n_731),
.B2(n_760),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_793),
.A2(n_98),
.B1(n_107),
.B2(n_123),
.Y(n_968)
);

OAI21xp5_ASAP7_75t_L g969 ( 
.A1(n_830),
.A2(n_124),
.B(n_134),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_779),
.B(n_189),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_829),
.A2(n_140),
.B(n_143),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_781),
.A2(n_153),
.B(n_159),
.C(n_801),
.Y(n_972)
);

O2A1O1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_789),
.A2(n_722),
.B(n_843),
.C(n_751),
.Y(n_973)
);

O2A1O1Ixp33_ASAP7_75t_SL g974 ( 
.A1(n_823),
.A2(n_775),
.B(n_768),
.C(n_813),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_811),
.B(n_793),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_831),
.A2(n_842),
.B(n_840),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_832),
.A2(n_760),
.B(n_791),
.Y(n_977)
);

OAI21xp33_ASAP7_75t_L g978 ( 
.A1(n_717),
.A2(n_743),
.B(n_835),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_811),
.A2(n_815),
.B1(n_812),
.B2(n_759),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_830),
.A2(n_756),
.B(n_746),
.C(n_833),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_760),
.A2(n_791),
.B(n_804),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_791),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_833),
.B(n_820),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_808),
.B(n_791),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_778),
.B(n_837),
.Y(n_985)
);

CKINVDCx6p67_ASAP7_75t_R g986 ( 
.A(n_769),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_818),
.A2(n_701),
.B(n_798),
.Y(n_987)
);

O2A1O1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_705),
.A2(n_733),
.B(n_827),
.C(n_563),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_701),
.B(n_705),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_711),
.B(n_641),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_701),
.B(n_705),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_701),
.B(n_705),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_733),
.B(n_827),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_826),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_701),
.B(n_705),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_705),
.A2(n_733),
.B(n_827),
.C(n_563),
.Y(n_996)
);

NOR2x1p5_ASAP7_75t_SL g997 ( 
.A(n_716),
.B(n_719),
.Y(n_997)
);

AO21x1_ASAP7_75t_L g998 ( 
.A1(n_702),
.A2(n_701),
.B(n_705),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_705),
.A2(n_605),
.B(n_702),
.C(n_739),
.Y(n_999)
);

O2A1O1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_705),
.A2(n_733),
.B(n_827),
.C(n_563),
.Y(n_1000)
);

OR2x6_ASAP7_75t_L g1001 ( 
.A(n_723),
.B(n_745),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_712),
.Y(n_1002)
);

BUFx4f_ASAP7_75t_L g1003 ( 
.A(n_723),
.Y(n_1003)
);

AOI21x1_ASAP7_75t_L g1004 ( 
.A1(n_841),
.A2(n_844),
.B(n_586),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_SL g1005 ( 
.A(n_927),
.B(n_912),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_999),
.A2(n_987),
.B(n_989),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_993),
.B(n_867),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_991),
.B(n_992),
.Y(n_1008)
);

BUFx2_ASAP7_75t_L g1009 ( 
.A(n_869),
.Y(n_1009)
);

OAI22x1_ASAP7_75t_L g1010 ( 
.A1(n_861),
.A2(n_940),
.B1(n_868),
.B2(n_946),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_877),
.B(n_922),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_854),
.B(n_988),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_894),
.Y(n_1013)
);

OAI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_847),
.A2(n_846),
.B(n_858),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_870),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_981),
.A2(n_859),
.B(n_858),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_975),
.B(n_996),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_1000),
.B(n_876),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_983),
.B(n_845),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_L g1020 ( 
.A1(n_859),
.A2(n_862),
.B(n_879),
.Y(n_1020)
);

O2A1O1Ixp5_ASAP7_75t_L g1021 ( 
.A1(n_998),
.A2(n_941),
.B(n_953),
.C(n_959),
.Y(n_1021)
);

AOI21x1_ASAP7_75t_L g1022 ( 
.A1(n_900),
.A2(n_899),
.B(n_928),
.Y(n_1022)
);

OR2x2_ASAP7_75t_L g1023 ( 
.A(n_878),
.B(n_874),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_887),
.B(n_908),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_1001),
.Y(n_1025)
);

AO21x2_ASAP7_75t_L g1026 ( 
.A1(n_871),
.A2(n_913),
.B(n_911),
.Y(n_1026)
);

INVx1_ASAP7_75t_SL g1027 ( 
.A(n_960),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_919),
.B(n_1003),
.Y(n_1028)
);

AOI21x1_ASAP7_75t_L g1029 ( 
.A1(n_929),
.A2(n_898),
.B(n_880),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_851),
.B(n_910),
.Y(n_1030)
);

AOI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_963),
.A2(n_950),
.B1(n_954),
.B2(n_857),
.Y(n_1031)
);

OR2x6_ASAP7_75t_L g1032 ( 
.A(n_1001),
.B(n_897),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_890),
.A2(n_856),
.B(n_863),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_866),
.A2(n_852),
.B(n_980),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_883),
.A2(n_873),
.B(n_864),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_1001),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_848),
.A2(n_937),
.B(n_924),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_919),
.B(n_1003),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_966),
.A2(n_969),
.B(n_952),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_905),
.A2(n_915),
.B(n_906),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_908),
.B(n_881),
.Y(n_1041)
);

AO31x2_ASAP7_75t_L g1042 ( 
.A1(n_920),
.A2(n_885),
.A3(n_984),
.B(n_967),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_930),
.A2(n_892),
.B(n_974),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_973),
.A2(n_888),
.B(n_850),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_853),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_SL g1046 ( 
.A1(n_972),
.A2(n_918),
.B(n_951),
.Y(n_1046)
);

AO21x2_ASAP7_75t_L g1047 ( 
.A1(n_888),
.A2(n_923),
.B(n_979),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_894),
.Y(n_1048)
);

OR2x2_ASAP7_75t_L g1049 ( 
.A(n_855),
.B(n_896),
.Y(n_1049)
);

AOI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_965),
.A2(n_944),
.B1(n_960),
.B2(n_926),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_849),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_936),
.B(n_961),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_860),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_849),
.Y(n_1054)
);

HB1xp67_ASAP7_75t_L g1055 ( 
.A(n_882),
.Y(n_1055)
);

AOI21x1_ASAP7_75t_SL g1056 ( 
.A1(n_942),
.A2(n_943),
.B(n_949),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_849),
.Y(n_1057)
);

INVx3_ASAP7_75t_SL g1058 ( 
.A(n_994),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_SL g1059 ( 
.A1(n_961),
.A2(n_971),
.B(n_968),
.Y(n_1059)
);

BUFx4f_ASAP7_75t_L g1060 ( 
.A(n_884),
.Y(n_1060)
);

NAND2x1_ASAP7_75t_L g1061 ( 
.A(n_850),
.B(n_982),
.Y(n_1061)
);

AO21x1_ASAP7_75t_L g1062 ( 
.A1(n_970),
.A2(n_957),
.B(n_955),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_904),
.B(n_982),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_904),
.A2(n_914),
.B(n_902),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_931),
.A2(n_964),
.B(n_934),
.Y(n_1065)
);

NAND2x1_ASAP7_75t_L g1066 ( 
.A(n_891),
.B(n_1002),
.Y(n_1066)
);

AOI21x1_ASAP7_75t_L g1067 ( 
.A1(n_893),
.A2(n_916),
.B(n_921),
.Y(n_1067)
);

NAND2x1p5_ASAP7_75t_L g1068 ( 
.A(n_962),
.B(n_1002),
.Y(n_1068)
);

AOI21x1_ASAP7_75t_L g1069 ( 
.A1(n_933),
.A2(n_947),
.B(n_948),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_978),
.B(n_1002),
.Y(n_1070)
);

AND2x2_ASAP7_75t_SL g1071 ( 
.A(n_917),
.B(n_938),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_990),
.A2(n_945),
.B(n_895),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_891),
.A2(n_903),
.B(n_958),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_901),
.B(n_958),
.Y(n_1074)
);

NAND2x1_ASAP7_75t_L g1075 ( 
.A(n_901),
.B(n_958),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_901),
.A2(n_903),
.B(n_872),
.Y(n_1076)
);

AOI21x1_ASAP7_75t_L g1077 ( 
.A1(n_935),
.A2(n_997),
.B(n_907),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_903),
.B(n_932),
.Y(n_1078)
);

A2O1A1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_956),
.A2(n_985),
.B(n_925),
.C(n_875),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_889),
.B(n_986),
.Y(n_1080)
);

OAI21xp33_ASAP7_75t_L g1081 ( 
.A1(n_875),
.A2(n_865),
.B(n_909),
.Y(n_1081)
);

NOR2x1_ASAP7_75t_SL g1082 ( 
.A(n_939),
.B(n_1001),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_939),
.B(n_878),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_939),
.B(n_1001),
.Y(n_1084)
);

AOI21x1_ASAP7_75t_L g1085 ( 
.A1(n_886),
.A2(n_1004),
.B(n_977),
.Y(n_1085)
);

BUFx2_ASAP7_75t_L g1086 ( 
.A(n_869),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_989),
.B(n_991),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_999),
.A2(n_987),
.B(n_989),
.Y(n_1088)
);

AO31x2_ASAP7_75t_L g1089 ( 
.A1(n_998),
.A2(n_976),
.A3(n_899),
.B(n_900),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_999),
.A2(n_988),
.B(n_1000),
.C(n_996),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_999),
.A2(n_987),
.B(n_989),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_989),
.A2(n_991),
.B1(n_995),
.B2(n_992),
.Y(n_1092)
);

AOI21x1_ASAP7_75t_L g1093 ( 
.A1(n_886),
.A2(n_1004),
.B(n_977),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_989),
.B(n_991),
.Y(n_1094)
);

AO21x1_ASAP7_75t_L g1095 ( 
.A1(n_922),
.A2(n_975),
.B(n_989),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_989),
.B(n_991),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_878),
.B(n_755),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_989),
.B(n_991),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_878),
.B(n_755),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_1001),
.B(n_926),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_870),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_870),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_989),
.B(n_991),
.Y(n_1103)
);

A2O1A1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_999),
.A2(n_988),
.B(n_1000),
.C(n_996),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_989),
.B(n_991),
.Y(n_1105)
);

AO31x2_ASAP7_75t_L g1106 ( 
.A1(n_998),
.A2(n_976),
.A3(n_899),
.B(n_900),
.Y(n_1106)
);

INVx5_ASAP7_75t_L g1107 ( 
.A(n_1001),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_999),
.A2(n_988),
.B(n_1000),
.C(n_996),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_1001),
.B(n_926),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_999),
.A2(n_987),
.B(n_989),
.Y(n_1110)
);

AOI221xp5_ASAP7_75t_L g1111 ( 
.A1(n_861),
.A2(n_563),
.B1(n_868),
.B2(n_705),
.C(n_676),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_894),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_993),
.B(n_989),
.Y(n_1113)
);

NAND3xp33_ASAP7_75t_SL g1114 ( 
.A(n_988),
.B(n_610),
.C(n_585),
.Y(n_1114)
);

AO31x2_ASAP7_75t_L g1115 ( 
.A1(n_998),
.A2(n_976),
.A3(n_899),
.B(n_900),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_993),
.B(n_989),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_999),
.A2(n_987),
.B(n_989),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_999),
.A2(n_987),
.B(n_989),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_989),
.B(n_991),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_869),
.Y(n_1120)
);

INVxp67_ASAP7_75t_L g1121 ( 
.A(n_869),
.Y(n_1121)
);

INVx3_ASAP7_75t_L g1122 ( 
.A(n_894),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_999),
.A2(n_988),
.B(n_1000),
.C(n_996),
.Y(n_1123)
);

HB1xp67_ASAP7_75t_L g1124 ( 
.A(n_869),
.Y(n_1124)
);

OAI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_999),
.A2(n_987),
.B(n_989),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_989),
.B(n_991),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_993),
.B(n_641),
.Y(n_1127)
);

O2A1O1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_999),
.A2(n_996),
.B(n_1000),
.C(n_988),
.Y(n_1128)
);

AO31x2_ASAP7_75t_L g1129 ( 
.A1(n_998),
.A2(n_976),
.A3(n_899),
.B(n_900),
.Y(n_1129)
);

AOI221x1_ASAP7_75t_L g1130 ( 
.A1(n_999),
.A2(n_963),
.B1(n_702),
.B2(n_975),
.C(n_922),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_989),
.B(n_991),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_869),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_993),
.B(n_989),
.Y(n_1133)
);

AOI21x1_ASAP7_75t_SL g1134 ( 
.A1(n_941),
.A2(n_991),
.B(n_989),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_1107),
.B(n_1028),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1092),
.A2(n_1012),
.B1(n_1119),
.B2(n_1126),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_SL g1137 ( 
.A1(n_1018),
.A2(n_1010),
.B1(n_1116),
.B2(n_1113),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1015),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1097),
.B(n_1099),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_1107),
.Y(n_1140)
);

BUFx5_ASAP7_75t_L g1141 ( 
.A(n_1084),
.Y(n_1141)
);

O2A1O1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_1111),
.A2(n_1092),
.B(n_1133),
.C(n_1104),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1101),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1008),
.A2(n_1105),
.B1(n_1126),
.B2(n_1119),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_SL g1145 ( 
.A(n_1071),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1008),
.B(n_1087),
.Y(n_1146)
);

INVx3_ASAP7_75t_L g1147 ( 
.A(n_1084),
.Y(n_1147)
);

NAND3xp33_ASAP7_75t_L g1148 ( 
.A(n_1130),
.B(n_1108),
.C(n_1090),
.Y(n_1148)
);

NAND2x1p5_ASAP7_75t_L g1149 ( 
.A(n_1107),
.B(n_1038),
.Y(n_1149)
);

O2A1O1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_1123),
.A2(n_1007),
.B(n_1131),
.C(n_1087),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_1060),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_1124),
.Y(n_1152)
);

INVx2_ASAP7_75t_SL g1153 ( 
.A(n_1060),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_1094),
.B(n_1096),
.Y(n_1154)
);

INVx1_ASAP7_75t_SL g1155 ( 
.A(n_1009),
.Y(n_1155)
);

INVx2_ASAP7_75t_SL g1156 ( 
.A(n_1045),
.Y(n_1156)
);

BUFx2_ASAP7_75t_SL g1157 ( 
.A(n_1086),
.Y(n_1157)
);

NAND2x1p5_ASAP7_75t_L g1158 ( 
.A(n_1107),
.B(n_1036),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_1120),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1094),
.A2(n_1131),
.B1(n_1105),
.B2(n_1103),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_1132),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1023),
.B(n_1121),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1096),
.A2(n_1098),
.B1(n_1103),
.B2(n_1017),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1006),
.A2(n_1091),
.B(n_1088),
.Y(n_1164)
);

OR2x2_ASAP7_75t_L g1165 ( 
.A(n_1098),
.B(n_1027),
.Y(n_1165)
);

OR2x6_ASAP7_75t_L g1166 ( 
.A(n_1032),
.B(n_1036),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1053),
.B(n_1055),
.Y(n_1167)
);

HB1xp67_ASAP7_75t_L g1168 ( 
.A(n_1070),
.Y(n_1168)
);

OR2x6_ASAP7_75t_L g1169 ( 
.A(n_1032),
.B(n_1036),
.Y(n_1169)
);

INVx2_ASAP7_75t_SL g1170 ( 
.A(n_1058),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_SL g1171 ( 
.A1(n_1079),
.A2(n_1082),
.B(n_1047),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1102),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1032),
.B(n_1027),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_1017),
.B(n_1081),
.Y(n_1174)
);

OR2x6_ASAP7_75t_L g1175 ( 
.A(n_1100),
.B(n_1109),
.Y(n_1175)
);

OA22x2_ASAP7_75t_L g1176 ( 
.A1(n_1050),
.A2(n_1080),
.B1(n_1109),
.B2(n_1100),
.Y(n_1176)
);

INVx4_ASAP7_75t_L g1177 ( 
.A(n_1051),
.Y(n_1177)
);

AO21x1_ASAP7_75t_L g1178 ( 
.A1(n_1005),
.A2(n_1043),
.B(n_1024),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_1068),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1127),
.B(n_1083),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1011),
.B(n_1019),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1024),
.A2(n_1128),
.B1(n_1006),
.B2(n_1110),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1019),
.B(n_1095),
.Y(n_1183)
);

INVx6_ASAP7_75t_L g1184 ( 
.A(n_1049),
.Y(n_1184)
);

OR2x6_ASAP7_75t_L g1185 ( 
.A(n_1025),
.B(n_1068),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_1070),
.Y(n_1186)
);

INVx2_ASAP7_75t_SL g1187 ( 
.A(n_1052),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1030),
.B(n_1005),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_1051),
.Y(n_1189)
);

AOI21xp33_ASAP7_75t_L g1190 ( 
.A1(n_1062),
.A2(n_1047),
.B(n_1046),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_1051),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1069),
.Y(n_1192)
);

BUFx3_ASAP7_75t_L g1193 ( 
.A(n_1054),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1078),
.B(n_1031),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_1078),
.Y(n_1195)
);

OAI22xp33_ASAP7_75t_L g1196 ( 
.A1(n_1114),
.A2(n_1110),
.B1(n_1118),
.B2(n_1088),
.Y(n_1196)
);

A2O1A1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1021),
.A2(n_1044),
.B(n_1117),
.C(n_1091),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1117),
.A2(n_1125),
.B(n_1118),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1035),
.A2(n_1125),
.B(n_1034),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_1054),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1041),
.B(n_1063),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1041),
.B(n_1063),
.Y(n_1202)
);

INVx1_ASAP7_75t_SL g1203 ( 
.A(n_1074),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_1013),
.B(n_1122),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1048),
.B(n_1112),
.Y(n_1205)
);

OR2x2_ASAP7_75t_L g1206 ( 
.A(n_1074),
.B(n_1042),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1054),
.B(n_1057),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1040),
.A2(n_1014),
.B1(n_1061),
.B2(n_1065),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1072),
.Y(n_1209)
);

OR2x2_ASAP7_75t_L g1210 ( 
.A(n_1042),
.B(n_1057),
.Y(n_1210)
);

NAND2xp33_ASAP7_75t_L g1211 ( 
.A(n_1057),
.B(n_1040),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1076),
.B(n_1073),
.Y(n_1212)
);

OR2x6_ASAP7_75t_L g1213 ( 
.A(n_1066),
.B(n_1075),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_1064),
.Y(n_1214)
);

OAI22x1_ASAP7_75t_L g1215 ( 
.A1(n_1077),
.A2(n_1067),
.B1(n_1022),
.B2(n_1093),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_1016),
.B(n_1033),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1134),
.A2(n_1029),
.B1(n_1056),
.B2(n_1059),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1089),
.B(n_1129),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1089),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1020),
.A2(n_1037),
.B(n_1026),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1106),
.B(n_1115),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1106),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1115),
.A2(n_1129),
.B(n_1085),
.Y(n_1223)
);

INVx6_ASAP7_75t_L g1224 ( 
.A(n_1107),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1113),
.B(n_1116),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1113),
.B(n_1116),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1092),
.B(n_1008),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_1107),
.Y(n_1228)
);

O2A1O1Ixp5_ASAP7_75t_SL g1229 ( 
.A1(n_1006),
.A2(n_1091),
.B(n_1110),
.C(n_1088),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1097),
.B(n_1099),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1015),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1113),
.B(n_1116),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_1045),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1113),
.B(n_1116),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_1124),
.Y(n_1235)
);

AOI221x1_ASAP7_75t_L g1236 ( 
.A1(n_1039),
.A2(n_999),
.B1(n_1081),
.B2(n_702),
.C(n_963),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1015),
.Y(n_1237)
);

INVx4_ASAP7_75t_L g1238 ( 
.A(n_1060),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1097),
.B(n_1099),
.Y(n_1239)
);

INVx2_ASAP7_75t_SL g1240 ( 
.A(n_1060),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1107),
.B(n_1028),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1107),
.B(n_1028),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1092),
.B(n_1008),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1092),
.B(n_1008),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1092),
.B(n_1008),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1009),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1092),
.A2(n_1012),
.B1(n_989),
.B2(n_992),
.Y(n_1247)
);

BUFx10_ASAP7_75t_L g1248 ( 
.A(n_1018),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1107),
.B(n_1028),
.Y(n_1249)
);

INVxp67_ASAP7_75t_L g1250 ( 
.A(n_1124),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1092),
.B(n_1008),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1015),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_1107),
.B(n_1028),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1015),
.Y(n_1254)
);

AOI21xp33_ASAP7_75t_SL g1255 ( 
.A1(n_1012),
.A2(n_610),
.B(n_585),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1107),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1081),
.A2(n_927),
.B1(n_1111),
.B2(n_868),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1015),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1097),
.B(n_1099),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1097),
.B(n_1099),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1081),
.A2(n_927),
.B1(n_1111),
.B2(n_868),
.Y(n_1261)
);

OR2x2_ASAP7_75t_L g1262 ( 
.A(n_1023),
.B(n_1113),
.Y(n_1262)
);

BUFx10_ASAP7_75t_L g1263 ( 
.A(n_1018),
.Y(n_1263)
);

OR2x2_ASAP7_75t_SL g1264 ( 
.A(n_1023),
.B(n_876),
.Y(n_1264)
);

OAI21xp33_ASAP7_75t_L g1265 ( 
.A1(n_1012),
.A2(n_991),
.B(n_989),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_1107),
.Y(n_1266)
);

AOI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1111),
.A2(n_927),
.B1(n_1012),
.B2(n_861),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1045),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1097),
.B(n_1099),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_SL g1270 ( 
.A1(n_1267),
.A2(n_1137),
.B1(n_1261),
.B2(n_1257),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1221),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1233),
.Y(n_1272)
);

AO21x2_ASAP7_75t_L g1273 ( 
.A1(n_1220),
.A2(n_1190),
.B(n_1223),
.Y(n_1273)
);

INVx3_ASAP7_75t_L g1274 ( 
.A(n_1221),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1147),
.B(n_1135),
.Y(n_1275)
);

INVx11_ASAP7_75t_L g1276 ( 
.A(n_1238),
.Y(n_1276)
);

BUFx8_ASAP7_75t_L g1277 ( 
.A(n_1145),
.Y(n_1277)
);

INVx1_ASAP7_75t_SL g1278 ( 
.A(n_1184),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1267),
.A2(n_1137),
.B1(n_1145),
.B2(n_1194),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1143),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1172),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1247),
.A2(n_1142),
.B1(n_1265),
.B2(n_1136),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1247),
.A2(n_1265),
.B1(n_1176),
.B2(n_1136),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1152),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1231),
.Y(n_1285)
);

INVx3_ASAP7_75t_L g1286 ( 
.A(n_1219),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1237),
.Y(n_1287)
);

INVx4_ASAP7_75t_L g1288 ( 
.A(n_1177),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1252),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1174),
.A2(n_1248),
.B1(n_1263),
.B2(n_1154),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1254),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1258),
.Y(n_1292)
);

INVx2_ASAP7_75t_SL g1293 ( 
.A(n_1173),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1209),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_SL g1295 ( 
.A1(n_1248),
.A2(n_1263),
.B1(n_1148),
.B2(n_1163),
.Y(n_1295)
);

AO21x1_ASAP7_75t_SL g1296 ( 
.A1(n_1199),
.A2(n_1190),
.B(n_1218),
.Y(n_1296)
);

BUFx4f_ASAP7_75t_SL g1297 ( 
.A(n_1153),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1165),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1199),
.B(n_1227),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1227),
.B(n_1243),
.Y(n_1300)
);

AOI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1144),
.A2(n_1160),
.B1(n_1163),
.B2(n_1269),
.Y(n_1301)
);

AOI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1215),
.A2(n_1217),
.B(n_1208),
.Y(n_1302)
);

INVx3_ASAP7_75t_L g1303 ( 
.A(n_1216),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_1184),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_SL g1305 ( 
.A1(n_1148),
.A2(n_1243),
.B1(n_1251),
.B2(n_1245),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1188),
.A2(n_1260),
.B1(n_1139),
.B2(n_1230),
.Y(n_1306)
);

BUFx3_ASAP7_75t_L g1307 ( 
.A(n_1268),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1168),
.Y(n_1308)
);

INVx3_ASAP7_75t_L g1309 ( 
.A(n_1216),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1217),
.A2(n_1229),
.B(n_1198),
.Y(n_1310)
);

INVx6_ASAP7_75t_L g1311 ( 
.A(n_1141),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1164),
.A2(n_1214),
.B(n_1212),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1225),
.B(n_1226),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1222),
.Y(n_1314)
);

INVx2_ASAP7_75t_SL g1315 ( 
.A(n_1210),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1186),
.Y(n_1316)
);

AO21x2_ASAP7_75t_L g1317 ( 
.A1(n_1183),
.A2(n_1171),
.B(n_1197),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1188),
.A2(n_1239),
.B1(n_1259),
.B2(n_1144),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_1140),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1160),
.A2(n_1244),
.B1(n_1245),
.B2(n_1251),
.Y(n_1320)
);

AOI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1236),
.A2(n_1182),
.B(n_1178),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1214),
.Y(n_1322)
);

BUFx2_ASAP7_75t_SL g1323 ( 
.A(n_1240),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1206),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1235),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1201),
.Y(n_1326)
);

INVxp67_ASAP7_75t_SL g1327 ( 
.A(n_1202),
.Y(n_1327)
);

HB1xp67_ASAP7_75t_L g1328 ( 
.A(n_1167),
.Y(n_1328)
);

CKINVDCx20_ASAP7_75t_R g1329 ( 
.A(n_1151),
.Y(n_1329)
);

OAI21xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1146),
.A2(n_1181),
.B(n_1234),
.Y(n_1330)
);

OAI22xp33_ASAP7_75t_SL g1331 ( 
.A1(n_1146),
.A2(n_1232),
.B1(n_1262),
.B2(n_1195),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1157),
.Y(n_1332)
);

INVx1_ASAP7_75t_SL g1333 ( 
.A(n_1155),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_1196),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_1264),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_1246),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_SL g1337 ( 
.A1(n_1180),
.A2(n_1147),
.B1(n_1141),
.B2(n_1253),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1192),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1203),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1189),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1155),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1200),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_1193),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1150),
.B(n_1162),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1185),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1250),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1175),
.B(n_1161),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1175),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1156),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1187),
.A2(n_1159),
.B1(n_1169),
.B2(n_1166),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1213),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1175),
.B(n_1166),
.Y(n_1352)
);

AO21x1_ASAP7_75t_L g1353 ( 
.A1(n_1211),
.A2(n_1205),
.B(n_1207),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1141),
.B(n_1191),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1191),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1170),
.Y(n_1356)
);

OAI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1255),
.A2(n_1185),
.B1(n_1149),
.B2(n_1228),
.Y(n_1357)
);

INVx2_ASAP7_75t_SL g1358 ( 
.A(n_1224),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1241),
.B(n_1249),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1179),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1149),
.Y(n_1361)
);

INVx4_ASAP7_75t_L g1362 ( 
.A(n_1140),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1158),
.Y(n_1363)
);

BUFx6f_ASAP7_75t_L g1364 ( 
.A(n_1228),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1256),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1256),
.Y(n_1366)
);

BUFx4_ASAP7_75t_SL g1367 ( 
.A(n_1204),
.Y(n_1367)
);

INVx4_ASAP7_75t_L g1368 ( 
.A(n_1256),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1242),
.A2(n_927),
.B1(n_1111),
.B2(n_1267),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1266),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1266),
.A2(n_1267),
.B1(n_1111),
.B2(n_1012),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1266),
.Y(n_1372)
);

AO21x1_ASAP7_75t_SL g1373 ( 
.A1(n_1199),
.A2(n_1190),
.B(n_1218),
.Y(n_1373)
);

BUFx12f_ASAP7_75t_L g1374 ( 
.A(n_1151),
.Y(n_1374)
);

OR2x6_ASAP7_75t_L g1375 ( 
.A(n_1171),
.B(n_1084),
.Y(n_1375)
);

OAI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1267),
.A2(n_1111),
.B1(n_1005),
.B2(n_802),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1138),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1138),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1199),
.B(n_1227),
.Y(n_1379)
);

CKINVDCx6p67_ASAP7_75t_R g1380 ( 
.A(n_1238),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1247),
.A2(n_1039),
.B(n_1164),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1154),
.B(n_1136),
.Y(n_1382)
);

CKINVDCx20_ASAP7_75t_R g1383 ( 
.A(n_1151),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1152),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_SL g1385 ( 
.A1(n_1137),
.A2(n_927),
.B1(n_1005),
.B2(n_689),
.Y(n_1385)
);

BUFx12f_ASAP7_75t_L g1386 ( 
.A(n_1151),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1138),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1138),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1138),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1320),
.B(n_1300),
.Y(n_1390)
);

INVxp67_ASAP7_75t_L g1391 ( 
.A(n_1296),
.Y(n_1391)
);

AO21x2_ASAP7_75t_L g1392 ( 
.A1(n_1381),
.A2(n_1321),
.B(n_1376),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1300),
.B(n_1299),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1324),
.B(n_1299),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1284),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1314),
.Y(n_1396)
);

BUFx2_ASAP7_75t_L g1397 ( 
.A(n_1303),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1379),
.B(n_1296),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1379),
.B(n_1373),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1325),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1382),
.B(n_1327),
.Y(n_1401)
);

BUFx8_ASAP7_75t_SL g1402 ( 
.A(n_1329),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1338),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1373),
.B(n_1334),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1303),
.Y(n_1405)
);

INVx3_ASAP7_75t_L g1406 ( 
.A(n_1303),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1384),
.Y(n_1407)
);

INVx5_ASAP7_75t_L g1408 ( 
.A(n_1375),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1324),
.B(n_1271),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1334),
.B(n_1271),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1305),
.B(n_1330),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1310),
.A2(n_1302),
.B(n_1312),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1341),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1271),
.B(n_1274),
.Y(n_1414)
);

OA21x2_ASAP7_75t_L g1415 ( 
.A1(n_1283),
.A2(n_1353),
.B(n_1294),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1317),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1317),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1294),
.Y(n_1418)
);

OA21x2_ASAP7_75t_L g1419 ( 
.A1(n_1353),
.A2(n_1322),
.B(n_1282),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1326),
.B(n_1301),
.Y(n_1420)
);

INVx1_ASAP7_75t_SL g1421 ( 
.A(n_1333),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1328),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1274),
.B(n_1309),
.Y(n_1423)
);

INVx3_ASAP7_75t_L g1424 ( 
.A(n_1309),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1389),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1317),
.Y(n_1426)
);

INVx8_ASAP7_75t_L g1427 ( 
.A(n_1375),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1309),
.Y(n_1428)
);

INVxp67_ASAP7_75t_L g1429 ( 
.A(n_1346),
.Y(n_1429)
);

INVx2_ASAP7_75t_SL g1430 ( 
.A(n_1311),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1280),
.B(n_1281),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1371),
.A2(n_1273),
.B(n_1270),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1315),
.B(n_1308),
.Y(n_1433)
);

INVx1_ASAP7_75t_SL g1434 ( 
.A(n_1347),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1340),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1388),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1285),
.Y(n_1437)
);

AO21x1_ASAP7_75t_L g1438 ( 
.A1(n_1344),
.A2(n_1331),
.B(n_1387),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1287),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1289),
.B(n_1291),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1292),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1342),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1377),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1378),
.B(n_1318),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1273),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1306),
.B(n_1315),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1286),
.Y(n_1447)
);

BUFx6f_ASAP7_75t_L g1448 ( 
.A(n_1311),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1293),
.B(n_1322),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1339),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1316),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1293),
.B(n_1298),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1313),
.B(n_1295),
.Y(n_1453)
);

OA21x2_ASAP7_75t_L g1454 ( 
.A1(n_1369),
.A2(n_1279),
.B(n_1348),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1355),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1290),
.B(n_1351),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1354),
.B(n_1347),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1345),
.B(n_1336),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1349),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1385),
.B(n_1361),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1272),
.B(n_1307),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1272),
.B(n_1307),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1361),
.B(n_1345),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1349),
.B(n_1375),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1336),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1375),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1360),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1352),
.B(n_1304),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1343),
.Y(n_1469)
);

INVx1_ASAP7_75t_SL g1470 ( 
.A(n_1370),
.Y(n_1470)
);

BUFx4f_ASAP7_75t_L g1471 ( 
.A(n_1319),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1288),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1365),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1393),
.B(n_1356),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1401),
.B(n_1357),
.Y(n_1475)
);

BUFx12f_ASAP7_75t_L g1476 ( 
.A(n_1458),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1401),
.B(n_1332),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1396),
.Y(n_1478)
);

INVx3_ASAP7_75t_SL g1479 ( 
.A(n_1419),
.Y(n_1479)
);

NOR2xp33_ASAP7_75t_L g1480 ( 
.A(n_1402),
.B(n_1332),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1393),
.B(n_1356),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1403),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1394),
.B(n_1278),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1403),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1398),
.B(n_1275),
.Y(n_1485)
);

AO21x2_ASAP7_75t_L g1486 ( 
.A1(n_1432),
.A2(n_1350),
.B(n_1363),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1418),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1390),
.B(n_1343),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1398),
.B(n_1399),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1390),
.B(n_1366),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1420),
.B(n_1319),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1420),
.B(n_1319),
.Y(n_1492)
);

BUFx3_ASAP7_75t_L g1493 ( 
.A(n_1397),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1399),
.B(n_1275),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1425),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_L g1496 ( 
.A(n_1448),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1411),
.B(n_1364),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1433),
.B(n_1372),
.Y(n_1498)
);

NAND3xp33_ASAP7_75t_L g1499 ( 
.A(n_1432),
.B(n_1277),
.C(n_1288),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1425),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1457),
.B(n_1404),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1457),
.B(n_1275),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1418),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1419),
.Y(n_1504)
);

INVx4_ASAP7_75t_L g1505 ( 
.A(n_1472),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1411),
.B(n_1364),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1433),
.B(n_1358),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1419),
.Y(n_1508)
);

BUFx4f_ASAP7_75t_L g1509 ( 
.A(n_1427),
.Y(n_1509)
);

AND2x4_ASAP7_75t_L g1510 ( 
.A(n_1408),
.B(n_1362),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1404),
.B(n_1337),
.Y(n_1511)
);

INVxp67_ASAP7_75t_SL g1512 ( 
.A(n_1419),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1449),
.B(n_1359),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1449),
.B(n_1359),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1395),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_1397),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1410),
.B(n_1359),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1410),
.B(n_1423),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1423),
.B(n_1362),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1413),
.B(n_1364),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1391),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1422),
.B(n_1400),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1423),
.B(n_1368),
.Y(n_1523)
);

INVxp67_ASAP7_75t_L g1524 ( 
.A(n_1455),
.Y(n_1524)
);

OAI211xp5_ASAP7_75t_L g1525 ( 
.A1(n_1453),
.A2(n_1335),
.B(n_1383),
.C(n_1329),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1414),
.B(n_1335),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1407),
.B(n_1358),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1436),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1515),
.B(n_1429),
.Y(n_1529)
);

OA21x2_ASAP7_75t_L g1530 ( 
.A1(n_1512),
.A2(n_1445),
.B(n_1412),
.Y(n_1530)
);

NAND3xp33_ASAP7_75t_L g1531 ( 
.A(n_1504),
.B(n_1467),
.C(n_1456),
.Y(n_1531)
);

OAI21xp5_ASAP7_75t_SL g1532 ( 
.A1(n_1525),
.A2(n_1391),
.B(n_1464),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1501),
.B(n_1405),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1515),
.B(n_1421),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1524),
.B(n_1421),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1501),
.B(n_1405),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1524),
.B(n_1435),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1522),
.B(n_1442),
.Y(n_1538)
);

OAI21xp33_ASAP7_75t_L g1539 ( 
.A1(n_1512),
.A2(n_1451),
.B(n_1439),
.Y(n_1539)
);

OA21x2_ASAP7_75t_L g1540 ( 
.A1(n_1504),
.A2(n_1445),
.B(n_1412),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1522),
.B(n_1431),
.Y(n_1541)
);

OAI21xp33_ASAP7_75t_L g1542 ( 
.A1(n_1508),
.A2(n_1451),
.B(n_1439),
.Y(n_1542)
);

NAND3xp33_ASAP7_75t_L g1543 ( 
.A(n_1508),
.B(n_1456),
.C(n_1415),
.Y(n_1543)
);

OAI221xp5_ASAP7_75t_L g1544 ( 
.A1(n_1479),
.A2(n_1415),
.B1(n_1444),
.B2(n_1441),
.C(n_1443),
.Y(n_1544)
);

OAI221xp5_ASAP7_75t_L g1545 ( 
.A1(n_1479),
.A2(n_1415),
.B1(n_1444),
.B2(n_1441),
.C(n_1443),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1488),
.B(n_1431),
.Y(n_1546)
);

OAI221xp5_ASAP7_75t_L g1547 ( 
.A1(n_1479),
.A2(n_1415),
.B1(n_1437),
.B2(n_1468),
.C(n_1463),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1477),
.B(n_1469),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1489),
.B(n_1406),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1499),
.A2(n_1458),
.B1(n_1465),
.B2(n_1459),
.Y(n_1550)
);

OA21x2_ASAP7_75t_L g1551 ( 
.A1(n_1475),
.A2(n_1445),
.B(n_1412),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1488),
.B(n_1440),
.Y(n_1552)
);

NAND3xp33_ASAP7_75t_L g1553 ( 
.A(n_1497),
.B(n_1437),
.C(n_1450),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1490),
.B(n_1440),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1487),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1489),
.B(n_1406),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1490),
.B(n_1392),
.Y(n_1557)
);

AOI21xp33_ASAP7_75t_L g1558 ( 
.A1(n_1475),
.A2(n_1438),
.B(n_1392),
.Y(n_1558)
);

NAND3xp33_ASAP7_75t_L g1559 ( 
.A(n_1497),
.B(n_1450),
.C(n_1463),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1486),
.A2(n_1438),
.B1(n_1454),
.B2(n_1392),
.Y(n_1560)
);

NAND3xp33_ASAP7_75t_L g1561 ( 
.A(n_1506),
.B(n_1450),
.C(n_1473),
.Y(n_1561)
);

OAI21xp5_ASAP7_75t_SL g1562 ( 
.A1(n_1525),
.A2(n_1464),
.B(n_1461),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1477),
.B(n_1506),
.Y(n_1563)
);

OAI221xp5_ASAP7_75t_L g1564 ( 
.A1(n_1499),
.A2(n_1468),
.B1(n_1460),
.B2(n_1434),
.C(n_1470),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1478),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1478),
.Y(n_1566)
);

NAND3xp33_ASAP7_75t_L g1567 ( 
.A(n_1491),
.B(n_1473),
.C(n_1447),
.Y(n_1567)
);

NAND3xp33_ASAP7_75t_L g1568 ( 
.A(n_1491),
.B(n_1447),
.C(n_1416),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1518),
.B(n_1406),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1487),
.Y(n_1570)
);

NAND3xp33_ASAP7_75t_L g1571 ( 
.A(n_1492),
.B(n_1447),
.C(n_1416),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1474),
.B(n_1392),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1518),
.B(n_1474),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1481),
.B(n_1406),
.Y(n_1574)
);

NAND3xp33_ASAP7_75t_L g1575 ( 
.A(n_1503),
.B(n_1417),
.C(n_1426),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1481),
.B(n_1424),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1502),
.B(n_1424),
.Y(n_1577)
);

OAI21xp33_ASAP7_75t_SL g1578 ( 
.A1(n_1485),
.A2(n_1461),
.B(n_1462),
.Y(n_1578)
);

OAI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1476),
.A2(n_1471),
.B1(n_1460),
.B2(n_1424),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1507),
.B(n_1462),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_SL g1581 ( 
.A(n_1505),
.B(n_1448),
.Y(n_1581)
);

AND2x2_ASAP7_75t_SL g1582 ( 
.A(n_1509),
.B(n_1466),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1507),
.B(n_1434),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1520),
.B(n_1470),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1502),
.B(n_1424),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1503),
.B(n_1409),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1517),
.B(n_1428),
.Y(n_1587)
);

NAND3xp33_ASAP7_75t_L g1588 ( 
.A(n_1520),
.B(n_1417),
.C(n_1426),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1517),
.B(n_1428),
.Y(n_1589)
);

OAI21xp5_ASAP7_75t_SL g1590 ( 
.A1(n_1511),
.A2(n_1480),
.B(n_1521),
.Y(n_1590)
);

AOI211xp5_ASAP7_75t_L g1591 ( 
.A1(n_1511),
.A2(n_1446),
.B(n_1452),
.C(n_1430),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1527),
.B(n_1452),
.Y(n_1592)
);

INVx2_ASAP7_75t_SL g1593 ( 
.A(n_1570),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1573),
.B(n_1485),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1555),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1586),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1590),
.B(n_1476),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1540),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1540),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1563),
.B(n_1476),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1586),
.Y(n_1601)
);

INVx4_ASAP7_75t_L g1602 ( 
.A(n_1530),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1573),
.B(n_1494),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1533),
.B(n_1494),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1553),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1540),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1565),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1533),
.B(n_1521),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1557),
.B(n_1482),
.Y(n_1609)
);

AND2x4_ASAP7_75t_SL g1610 ( 
.A(n_1577),
.B(n_1510),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1536),
.B(n_1549),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1572),
.B(n_1482),
.Y(n_1612)
);

AND2x4_ASAP7_75t_L g1613 ( 
.A(n_1581),
.B(n_1493),
.Y(n_1613)
);

INVxp67_ASAP7_75t_SL g1614 ( 
.A(n_1531),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1536),
.B(n_1513),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1541),
.B(n_1538),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1534),
.Y(n_1617)
);

CKINVDCx20_ASAP7_75t_R g1618 ( 
.A(n_1580),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1542),
.B(n_1484),
.Y(n_1619)
);

NAND2x1p5_ASAP7_75t_L g1620 ( 
.A(n_1582),
.B(n_1408),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1581),
.B(n_1493),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1549),
.B(n_1513),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1554),
.B(n_1498),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1565),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1556),
.B(n_1514),
.Y(n_1625)
);

BUFx2_ASAP7_75t_L g1626 ( 
.A(n_1578),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1566),
.Y(n_1627)
);

INVxp67_ASAP7_75t_L g1628 ( 
.A(n_1547),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1539),
.B(n_1484),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1546),
.B(n_1498),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1561),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1556),
.B(n_1514),
.Y(n_1632)
);

INVxp67_ASAP7_75t_SL g1633 ( 
.A(n_1551),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1552),
.B(n_1527),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1569),
.B(n_1493),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1567),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1569),
.B(n_1516),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1577),
.B(n_1516),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1585),
.B(n_1516),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1585),
.B(n_1505),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1587),
.B(n_1526),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1587),
.B(n_1526),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1559),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1537),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1619),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1617),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1626),
.B(n_1589),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1619),
.Y(n_1648)
);

NAND2x1p5_ASAP7_75t_L g1649 ( 
.A(n_1626),
.B(n_1582),
.Y(n_1649)
);

NAND2x1p5_ASAP7_75t_L g1650 ( 
.A(n_1613),
.B(n_1509),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1629),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1595),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1617),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1600),
.B(n_1548),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1643),
.B(n_1529),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1610),
.B(n_1574),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1595),
.Y(n_1657)
);

NAND2x1p5_ASAP7_75t_L g1658 ( 
.A(n_1613),
.B(n_1509),
.Y(n_1658)
);

INVx2_ASAP7_75t_SL g1659 ( 
.A(n_1610),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1610),
.B(n_1574),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1596),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1643),
.B(n_1548),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1605),
.B(n_1592),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1629),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1605),
.B(n_1583),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1634),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1594),
.B(n_1576),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1628),
.A2(n_1558),
.B(n_1545),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1594),
.B(n_1576),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1636),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1636),
.B(n_1535),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1631),
.B(n_1584),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1598),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1631),
.B(n_1495),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1596),
.B(n_1601),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1603),
.B(n_1519),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1634),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1644),
.Y(n_1678)
);

INVxp67_ASAP7_75t_SL g1679 ( 
.A(n_1633),
.Y(n_1679)
);

NAND3xp33_ASAP7_75t_L g1680 ( 
.A(n_1628),
.B(n_1543),
.C(n_1544),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1644),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1603),
.B(n_1519),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1611),
.B(n_1523),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1598),
.Y(n_1684)
);

OR2x6_ASAP7_75t_L g1685 ( 
.A(n_1620),
.B(n_1427),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1623),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1623),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1630),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1662),
.B(n_1614),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1674),
.Y(n_1690)
);

INVx2_ASAP7_75t_SL g1691 ( 
.A(n_1649),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_L g1692 ( 
.A(n_1654),
.B(n_1600),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1647),
.B(n_1614),
.Y(n_1693)
);

HB1xp67_ASAP7_75t_L g1694 ( 
.A(n_1670),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1652),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1646),
.B(n_1593),
.Y(n_1696)
);

AOI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1680),
.A2(n_1560),
.B1(n_1564),
.B2(n_1633),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1652),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1647),
.B(n_1615),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1671),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1653),
.B(n_1593),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1657),
.Y(n_1702)
);

NOR2x1_ASAP7_75t_L g1703 ( 
.A(n_1671),
.B(n_1597),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1673),
.Y(n_1704)
);

NOR2x2_ASAP7_75t_L g1705 ( 
.A(n_1685),
.B(n_1597),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1675),
.B(n_1612),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1657),
.Y(n_1707)
);

INVxp67_ASAP7_75t_SL g1708 ( 
.A(n_1649),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1673),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1647),
.B(n_1615),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1686),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1687),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1649),
.B(n_1615),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1688),
.Y(n_1714)
);

OAI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1668),
.A2(n_1618),
.B1(n_1560),
.B2(n_1591),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1675),
.B(n_1612),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1663),
.B(n_1609),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1659),
.B(n_1604),
.Y(n_1718)
);

OAI21xp5_ASAP7_75t_L g1719 ( 
.A1(n_1679),
.A2(n_1609),
.B(n_1602),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1655),
.B(n_1593),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1663),
.B(n_1616),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1645),
.B(n_1601),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1659),
.B(n_1604),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1648),
.B(n_1616),
.Y(n_1724)
);

NAND2xp67_ASAP7_75t_SL g1725 ( 
.A(n_1656),
.B(n_1608),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1666),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1667),
.B(n_1641),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1661),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1677),
.Y(n_1729)
);

OAI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1650),
.A2(n_1532),
.B1(n_1562),
.B2(n_1630),
.Y(n_1730)
);

OAI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1672),
.A2(n_1664),
.B(n_1651),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1665),
.B(n_1661),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1684),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1678),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1721),
.B(n_1665),
.Y(n_1735)
);

INVx1_ASAP7_75t_SL g1736 ( 
.A(n_1705),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1700),
.B(n_1681),
.Y(n_1737)
);

INVx1_ASAP7_75t_SL g1738 ( 
.A(n_1705),
.Y(n_1738)
);

AND2x4_ASAP7_75t_L g1739 ( 
.A(n_1699),
.B(n_1667),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1699),
.B(n_1669),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1728),
.Y(n_1741)
);

INVx1_ASAP7_75t_SL g1742 ( 
.A(n_1693),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1721),
.B(n_1669),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1728),
.Y(n_1744)
);

INVx1_ASAP7_75t_SL g1745 ( 
.A(n_1693),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1695),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1698),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1710),
.B(n_1676),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1732),
.B(n_1684),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1702),
.Y(n_1750)
);

INVxp67_ASAP7_75t_L g1751 ( 
.A(n_1694),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1710),
.B(n_1713),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1707),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1713),
.B(n_1676),
.Y(n_1754)
);

AND2x4_ASAP7_75t_L g1755 ( 
.A(n_1727),
.B(n_1656),
.Y(n_1755)
);

CKINVDCx16_ASAP7_75t_R g1756 ( 
.A(n_1692),
.Y(n_1756)
);

AOI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1715),
.A2(n_1602),
.B1(n_1685),
.B2(n_1486),
.Y(n_1757)
);

HB1xp67_ASAP7_75t_L g1758 ( 
.A(n_1734),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1704),
.Y(n_1759)
);

INVxp33_ASAP7_75t_SL g1760 ( 
.A(n_1730),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1734),
.Y(n_1761)
);

NOR2x1p5_ASAP7_75t_L g1762 ( 
.A(n_1708),
.B(n_1374),
.Y(n_1762)
);

OAI21x1_ASAP7_75t_L g1763 ( 
.A1(n_1719),
.A2(n_1658),
.B(n_1650),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1732),
.B(n_1717),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1727),
.B(n_1682),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1711),
.Y(n_1766)
);

NAND2x1p5_ASAP7_75t_L g1767 ( 
.A(n_1691),
.B(n_1471),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1697),
.A2(n_1602),
.B1(n_1685),
.B2(n_1486),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_SL g1769 ( 
.A1(n_1689),
.A2(n_1602),
.B1(n_1606),
.B2(n_1599),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1718),
.B(n_1682),
.Y(n_1770)
);

INVx1_ASAP7_75t_SL g1771 ( 
.A(n_1703),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1712),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1758),
.Y(n_1773)
);

AOI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1757),
.A2(n_1691),
.B1(n_1726),
.B2(n_1714),
.Y(n_1774)
);

CKINVDCx16_ASAP7_75t_R g1775 ( 
.A(n_1756),
.Y(n_1775)
);

OAI222xp33_ASAP7_75t_L g1776 ( 
.A1(n_1736),
.A2(n_1717),
.B1(n_1704),
.B2(n_1733),
.C1(n_1709),
.C2(n_1729),
.Y(n_1776)
);

OAI211xp5_ASAP7_75t_L g1777 ( 
.A1(n_1771),
.A2(n_1696),
.B(n_1701),
.C(n_1720),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1742),
.B(n_1690),
.Y(n_1778)
);

OA211x2_ASAP7_75t_L g1779 ( 
.A1(n_1751),
.A2(n_1731),
.B(n_1725),
.C(n_1724),
.Y(n_1779)
);

NOR2x1_ASAP7_75t_L g1780 ( 
.A(n_1762),
.B(n_1725),
.Y(n_1780)
);

INVxp67_ASAP7_75t_L g1781 ( 
.A(n_1738),
.Y(n_1781)
);

AOI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1760),
.A2(n_1733),
.B1(n_1709),
.B2(n_1722),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1752),
.B(n_1718),
.Y(n_1783)
);

INVxp67_ASAP7_75t_L g1784 ( 
.A(n_1766),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1741),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1741),
.Y(n_1786)
);

OAI221xp5_ASAP7_75t_L g1787 ( 
.A1(n_1768),
.A2(n_1599),
.B1(n_1606),
.B2(n_1598),
.C(n_1706),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1735),
.B(n_1706),
.Y(n_1788)
);

AOI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1760),
.A2(n_1685),
.B1(n_1606),
.B2(n_1599),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1752),
.B(n_1723),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1744),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1745),
.A2(n_1550),
.B1(n_1723),
.B2(n_1650),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1739),
.Y(n_1793)
);

OAI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1769),
.A2(n_1735),
.B1(n_1764),
.B2(n_1743),
.Y(n_1794)
);

AOI22xp5_ASAP7_75t_L g1795 ( 
.A1(n_1759),
.A2(n_1658),
.B1(n_1486),
.B2(n_1551),
.Y(n_1795)
);

OAI21xp33_ASAP7_75t_L g1796 ( 
.A1(n_1737),
.A2(n_1716),
.B(n_1658),
.Y(n_1796)
);

O2A1O1Ixp33_ASAP7_75t_L g1797 ( 
.A1(n_1772),
.A2(n_1716),
.B(n_1579),
.C(n_1383),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1744),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1746),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1764),
.B(n_1683),
.Y(n_1800)
);

BUFx4f_ASAP7_75t_SL g1801 ( 
.A(n_1775),
.Y(n_1801)
);

INVx1_ASAP7_75t_SL g1802 ( 
.A(n_1793),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1800),
.B(n_1743),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1782),
.B(n_1765),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1781),
.B(n_1765),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1783),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1785),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1790),
.B(n_1770),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1788),
.B(n_1770),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1786),
.Y(n_1810)
);

OAI221xp5_ASAP7_75t_L g1811 ( 
.A1(n_1794),
.A2(n_1749),
.B1(n_1767),
.B2(n_1772),
.C(n_1759),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1791),
.Y(n_1812)
);

AOI221xp5_ASAP7_75t_L g1813 ( 
.A1(n_1776),
.A2(n_1761),
.B1(n_1746),
.B2(n_1750),
.C(n_1747),
.Y(n_1813)
);

NAND2x1_ASAP7_75t_L g1814 ( 
.A(n_1780),
.B(n_1755),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1800),
.B(n_1748),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1788),
.B(n_1740),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1784),
.B(n_1740),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1798),
.Y(n_1818)
);

NOR2x1_ASAP7_75t_L g1819 ( 
.A(n_1773),
.B(n_1747),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1792),
.B(n_1748),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1799),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1808),
.B(n_1778),
.Y(n_1822)
);

NOR2xp33_ASAP7_75t_SL g1823 ( 
.A(n_1801),
.B(n_1374),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_L g1824 ( 
.A(n_1801),
.B(n_1777),
.Y(n_1824)
);

A2O1A1Ixp33_ASAP7_75t_SL g1825 ( 
.A1(n_1811),
.A2(n_1794),
.B(n_1779),
.C(n_1787),
.Y(n_1825)
);

AOI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1813),
.A2(n_1774),
.B1(n_1795),
.B2(n_1820),
.Y(n_1826)
);

AOI221xp5_ASAP7_75t_L g1827 ( 
.A1(n_1804),
.A2(n_1789),
.B1(n_1796),
.B2(n_1797),
.C(n_1750),
.Y(n_1827)
);

OAI211xp5_ASAP7_75t_SL g1828 ( 
.A1(n_1819),
.A2(n_1753),
.B(n_1749),
.C(n_1763),
.Y(n_1828)
);

AOI21xp5_ASAP7_75t_L g1829 ( 
.A1(n_1814),
.A2(n_1755),
.B(n_1739),
.Y(n_1829)
);

AOI211xp5_ASAP7_75t_L g1830 ( 
.A1(n_1802),
.A2(n_1763),
.B(n_1754),
.C(n_1755),
.Y(n_1830)
);

AOI311xp33_ASAP7_75t_L g1831 ( 
.A1(n_1816),
.A2(n_1739),
.A3(n_1754),
.B(n_1767),
.C(n_1495),
.Y(n_1831)
);

NOR4xp25_ASAP7_75t_L g1832 ( 
.A(n_1805),
.B(n_1608),
.C(n_1660),
.D(n_1641),
.Y(n_1832)
);

NOR3xp33_ASAP7_75t_L g1833 ( 
.A(n_1809),
.B(n_1386),
.C(n_1568),
.Y(n_1833)
);

NAND2x1_ASAP7_75t_L g1834 ( 
.A(n_1806),
.B(n_1660),
.Y(n_1834)
);

AND3x1_ASAP7_75t_L g1835 ( 
.A(n_1823),
.B(n_1806),
.C(n_1817),
.Y(n_1835)
);

OAI322xp33_ASAP7_75t_L g1836 ( 
.A1(n_1824),
.A2(n_1821),
.A3(n_1807),
.B1(n_1818),
.B2(n_1810),
.C1(n_1812),
.C2(n_1803),
.Y(n_1836)
);

AOI31xp33_ASAP7_75t_L g1837 ( 
.A1(n_1822),
.A2(n_1820),
.A3(n_1808),
.B(n_1815),
.Y(n_1837)
);

NAND4xp75_ASAP7_75t_L g1838 ( 
.A(n_1829),
.B(n_1815),
.C(n_1386),
.D(n_1297),
.Y(n_1838)
);

HB1xp67_ASAP7_75t_L g1839 ( 
.A(n_1834),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1832),
.B(n_1767),
.Y(n_1840)
);

NOR3xp33_ASAP7_75t_L g1841 ( 
.A(n_1828),
.B(n_1571),
.C(n_1575),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1827),
.Y(n_1842)
);

OAI211xp5_ASAP7_75t_L g1843 ( 
.A1(n_1825),
.A2(n_1276),
.B(n_1642),
.C(n_1683),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1830),
.Y(n_1844)
);

NAND4xp25_ASAP7_75t_L g1845 ( 
.A(n_1831),
.B(n_1613),
.C(n_1621),
.D(n_1640),
.Y(n_1845)
);

INVxp67_ASAP7_75t_L g1846 ( 
.A(n_1826),
.Y(n_1846)
);

NAND3xp33_ASAP7_75t_SL g1847 ( 
.A(n_1843),
.B(n_1833),
.C(n_1620),
.Y(n_1847)
);

NAND3xp33_ASAP7_75t_L g1848 ( 
.A(n_1842),
.B(n_1835),
.C(n_1844),
.Y(n_1848)
);

A2O1A1Ixp33_ASAP7_75t_L g1849 ( 
.A1(n_1843),
.A2(n_1323),
.B(n_1613),
.C(n_1621),
.Y(n_1849)
);

NAND3xp33_ASAP7_75t_L g1850 ( 
.A(n_1846),
.B(n_1277),
.C(n_1621),
.Y(n_1850)
);

HB1xp67_ASAP7_75t_L g1851 ( 
.A(n_1839),
.Y(n_1851)
);

HB1xp67_ASAP7_75t_L g1852 ( 
.A(n_1840),
.Y(n_1852)
);

AOI221xp5_ASAP7_75t_L g1853 ( 
.A1(n_1841),
.A2(n_1588),
.B1(n_1607),
.B2(n_1624),
.C(n_1627),
.Y(n_1853)
);

NAND4xp25_ASAP7_75t_L g1854 ( 
.A(n_1845),
.B(n_1621),
.C(n_1276),
.D(n_1640),
.Y(n_1854)
);

AOI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1848),
.A2(n_1838),
.B1(n_1837),
.B2(n_1836),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1851),
.Y(n_1856)
);

NOR2x1_ASAP7_75t_L g1857 ( 
.A(n_1850),
.B(n_1642),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1852),
.Y(n_1858)
);

NOR2x1_ASAP7_75t_L g1859 ( 
.A(n_1847),
.B(n_1640),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1854),
.Y(n_1860)
);

AOI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1849),
.A2(n_1277),
.B1(n_1380),
.B2(n_1551),
.Y(n_1861)
);

AOI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1853),
.A2(n_1380),
.B1(n_1530),
.B2(n_1483),
.Y(n_1862)
);

OR2x6_ASAP7_75t_L g1863 ( 
.A(n_1856),
.B(n_1367),
.Y(n_1863)
);

INVx5_ASAP7_75t_L g1864 ( 
.A(n_1858),
.Y(n_1864)
);

NAND3x1_ASAP7_75t_L g1865 ( 
.A(n_1855),
.B(n_1611),
.C(n_1635),
.Y(n_1865)
);

INVxp67_ASAP7_75t_SL g1866 ( 
.A(n_1860),
.Y(n_1866)
);

NOR2x1_ASAP7_75t_L g1867 ( 
.A(n_1859),
.B(n_1640),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1857),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1864),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1863),
.Y(n_1870)
);

HB1xp67_ASAP7_75t_L g1871 ( 
.A(n_1868),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1866),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1871),
.Y(n_1873)
);

OAI22x1_ASAP7_75t_L g1874 ( 
.A1(n_1872),
.A2(n_1861),
.B1(n_1867),
.B2(n_1862),
.Y(n_1874)
);

NOR2x1p5_ASAP7_75t_L g1875 ( 
.A(n_1873),
.B(n_1869),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1875),
.Y(n_1876)
);

OAI22xp33_ASAP7_75t_SL g1877 ( 
.A1(n_1875),
.A2(n_1871),
.B1(n_1870),
.B2(n_1874),
.Y(n_1877)
);

AOI21xp33_ASAP7_75t_L g1878 ( 
.A1(n_1877),
.A2(n_1865),
.B(n_1483),
.Y(n_1878)
);

OAI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1876),
.A2(n_1625),
.B1(n_1622),
.B2(n_1632),
.Y(n_1879)
);

OAI21x1_ASAP7_75t_L g1880 ( 
.A1(n_1879),
.A2(n_1625),
.B(n_1622),
.Y(n_1880)
);

INVxp67_ASAP7_75t_L g1881 ( 
.A(n_1880),
.Y(n_1881)
);

AOI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1881),
.A2(n_1878),
.B1(n_1632),
.B2(n_1288),
.Y(n_1882)
);

OAI221xp5_ASAP7_75t_R g1883 ( 
.A1(n_1882),
.A2(n_1635),
.B1(n_1637),
.B2(n_1638),
.C(n_1639),
.Y(n_1883)
);

AOI211xp5_ASAP7_75t_L g1884 ( 
.A1(n_1883),
.A2(n_1496),
.B(n_1500),
.C(n_1528),
.Y(n_1884)
);


endmodule