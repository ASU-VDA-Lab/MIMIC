module fake_netlist_6_2964_n_2352 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_507, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_396, n_495, n_350, n_78, n_84, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_468, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_466, n_506, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_153, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_493, n_397, n_155, n_109, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_363, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_483, n_102, n_204, n_482, n_474, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_33, n_477, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_487, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2352);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_507;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_468;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_493;
input n_397;
input n_155;
input n_109;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_33;
input n_477;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2352;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2291;
wire n_830;
wire n_2299;
wire n_873;
wire n_1371;
wire n_1285;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_539;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_2190;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2207;
wire n_1970;
wire n_608;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_792;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2193;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_2178;
wire n_950;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_644;
wire n_682;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_1492;
wire n_987;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_2231;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_811;
wire n_683;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_1053;
wire n_1681;
wire n_520;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2204;
wire n_1520;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_2278;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2052;
wire n_1847;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_1997;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_2310;
wire n_584;
wire n_2141;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1949;
wire n_545;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_646;
wire n_528;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_1283;
wire n_918;
wire n_748;
wire n_1114;
wire n_1848;
wire n_1147;
wire n_763;
wire n_1785;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_2287;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_924;
wire n_1582;
wire n_2318;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_1218;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_985;
wire n_2233;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1996;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_1025;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_72),
.Y(n_511)
);

BUFx10_ASAP7_75t_L g512 ( 
.A(n_321),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_141),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_209),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_21),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_62),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_255),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_235),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_407),
.Y(n_519)
);

BUFx10_ASAP7_75t_L g520 ( 
.A(n_32),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_67),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_421),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_452),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_241),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_146),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_231),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_149),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_25),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_25),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_448),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_135),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_492),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_397),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_110),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_55),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_311),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g537 ( 
.A(n_301),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_263),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_332),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_338),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_498),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_476),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_28),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_245),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_70),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_386),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_491),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_90),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_164),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_139),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_285),
.Y(n_551)
);

CKINVDCx14_ASAP7_75t_R g552 ( 
.A(n_162),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_12),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_482),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_406),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_97),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_246),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_468),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_270),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_211),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_53),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_371),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_73),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_178),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_484),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_42),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_226),
.Y(n_567)
);

BUFx10_ASAP7_75t_L g568 ( 
.A(n_114),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_210),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_249),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_345),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_200),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_429),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_8),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_161),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_107),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_404),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_199),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_419),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_292),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_447),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_40),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_453),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_480),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_68),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_39),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_194),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_359),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_222),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_462),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_116),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_394),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_418),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_14),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_165),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_3),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_6),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_256),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_505),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_490),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_305),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_165),
.Y(n_602)
);

BUFx8_ASAP7_75t_SL g603 ( 
.A(n_6),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_496),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_401),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_218),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_38),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_104),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_5),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_494),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_178),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_70),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_76),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_336),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_368),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_247),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_486),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_495),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_322),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_97),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_472),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_84),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_113),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_140),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_225),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_502),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_112),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_160),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_16),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_243),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_10),
.Y(n_631)
);

CKINVDCx16_ASAP7_75t_R g632 ( 
.A(n_199),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_59),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_14),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_434),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_341),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_228),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_300),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_215),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_445),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_148),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_55),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_500),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_280),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_48),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_446),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_351),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_230),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_149),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_478),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_349),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_483),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_81),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_348),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_45),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_61),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_343),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_81),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_479),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_26),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_402),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_493),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_475),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_499),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_485),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_323),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_156),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_370),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_372),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_275),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_130),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_175),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_15),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_410),
.Y(n_674)
);

BUFx5_ASAP7_75t_L g675 ( 
.A(n_125),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_327),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_157),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_293),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_106),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_488),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_145),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_405),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_399),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_391),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_27),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_320),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_127),
.Y(n_687)
);

CKINVDCx20_ASAP7_75t_R g688 ( 
.A(n_57),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_437),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_150),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_354),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_20),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_473),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_501),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_274),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_340),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_315),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_87),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_460),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_179),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_68),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_101),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_115),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_48),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_358),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_400),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_90),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_489),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_94),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_229),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_481),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_0),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_176),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_82),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_383),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_251),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_389),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_75),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_497),
.Y(n_719)
);

INVx1_ASAP7_75t_SL g720 ( 
.A(n_33),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_303),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_356),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_45),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_330),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_395),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_487),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_195),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_102),
.Y(n_728)
);

INVxp67_ASAP7_75t_SL g729 ( 
.A(n_684),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_675),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_675),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_675),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_523),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_675),
.Y(n_734)
);

CKINVDCx16_ASAP7_75t_R g735 ( 
.A(n_632),
.Y(n_735)
);

INVxp67_ASAP7_75t_SL g736 ( 
.A(n_555),
.Y(n_736)
);

INVxp67_ASAP7_75t_SL g737 ( 
.A(n_559),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_603),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_675),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_675),
.Y(n_740)
);

INVxp67_ASAP7_75t_SL g741 ( 
.A(n_598),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_675),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_709),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_603),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_709),
.Y(n_745)
);

INVxp33_ASAP7_75t_SL g746 ( 
.A(n_511),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_514),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_627),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_517),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_519),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_514),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_516),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_514),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_514),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_513),
.Y(n_755)
);

INVxp33_ASAP7_75t_L g756 ( 
.A(n_560),
.Y(n_756)
);

BUFx2_ASAP7_75t_L g757 ( 
.A(n_552),
.Y(n_757)
);

CKINVDCx16_ASAP7_75t_R g758 ( 
.A(n_552),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_526),
.Y(n_759)
);

INVxp67_ASAP7_75t_SL g760 ( 
.A(n_659),
.Y(n_760)
);

INVxp33_ASAP7_75t_L g761 ( 
.A(n_560),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_520),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_515),
.Y(n_763)
);

CKINVDCx20_ASAP7_75t_R g764 ( 
.A(n_627),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_527),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_528),
.Y(n_766)
);

INVxp67_ASAP7_75t_SL g767 ( 
.A(n_554),
.Y(n_767)
);

INVxp33_ASAP7_75t_L g768 ( 
.A(n_572),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_529),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_534),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_549),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_521),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_550),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_530),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_679),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_556),
.Y(n_776)
);

CKINVDCx14_ASAP7_75t_R g777 ( 
.A(n_512),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_532),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_569),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_582),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_585),
.Y(n_781)
);

BUFx2_ASAP7_75t_L g782 ( 
.A(n_525),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_586),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_587),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_607),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_533),
.Y(n_786)
);

INVxp33_ASAP7_75t_SL g787 ( 
.A(n_531),
.Y(n_787)
);

INVxp67_ASAP7_75t_SL g788 ( 
.A(n_554),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_613),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_536),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_540),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_541),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_535),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_620),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_622),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_544),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_628),
.Y(n_797)
);

INVxp33_ASAP7_75t_SL g798 ( 
.A(n_543),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_679),
.Y(n_799)
);

INVxp33_ASAP7_75t_SL g800 ( 
.A(n_545),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_631),
.Y(n_801)
);

CKINVDCx14_ASAP7_75t_R g802 ( 
.A(n_512),
.Y(n_802)
);

INVxp67_ASAP7_75t_L g803 ( 
.A(n_520),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_633),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_641),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_687),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_653),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_656),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_660),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_572),
.Y(n_810)
);

INVxp67_ASAP7_75t_SL g811 ( 
.A(n_518),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_690),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_523),
.Y(n_813)
);

INVxp33_ASAP7_75t_L g814 ( 
.A(n_642),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_548),
.Y(n_815)
);

INVxp33_ASAP7_75t_SL g816 ( 
.A(n_561),
.Y(n_816)
);

INVxp67_ASAP7_75t_SL g817 ( 
.A(n_522),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_700),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_701),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_703),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_524),
.B(n_1),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_704),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_520),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_712),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_811),
.B(n_542),
.Y(n_825)
);

OA21x2_ASAP7_75t_L g826 ( 
.A1(n_730),
.A2(n_558),
.B(n_542),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_733),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_733),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_733),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_733),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_813),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_749),
.Y(n_832)
);

BUFx8_ASAP7_75t_SL g833 ( 
.A(n_738),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_817),
.B(n_558),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_751),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_813),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_735),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_751),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_736),
.A2(n_686),
.B1(n_661),
.B2(n_565),
.Y(n_839)
);

CKINVDCx16_ASAP7_75t_R g840 ( 
.A(n_758),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_747),
.Y(n_841)
);

INVx5_ASAP7_75t_L g842 ( 
.A(n_813),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_813),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_752),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_753),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_750),
.B(n_588),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_732),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_767),
.B(n_788),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_759),
.B(n_588),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_774),
.B(n_668),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_732),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_754),
.Y(n_852)
);

INVx5_ASAP7_75t_L g853 ( 
.A(n_810),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_731),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_734),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_772),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_739),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_L g858 ( 
.A1(n_737),
.A2(n_566),
.B1(n_574),
.B2(n_564),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_778),
.B(n_668),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_740),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_810),
.Y(n_861)
);

CKINVDCx14_ASAP7_75t_R g862 ( 
.A(n_777),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_742),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_786),
.B(n_717),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_755),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_763),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_765),
.Y(n_867)
);

OA21x2_ASAP7_75t_L g868 ( 
.A1(n_821),
.A2(n_717),
.B(n_551),
.Y(n_868)
);

NAND2xp33_ASAP7_75t_L g869 ( 
.A(n_756),
.B(n_642),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_766),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_769),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_743),
.B(n_538),
.Y(n_872)
);

OA21x2_ASAP7_75t_L g873 ( 
.A1(n_770),
.A2(n_567),
.B(n_557),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_771),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_773),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_776),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_779),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_790),
.B(n_570),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_780),
.Y(n_879)
);

OAI22x1_ASAP7_75t_R g880 ( 
.A1(n_738),
.A2(n_688),
.B1(n_687),
.B2(n_563),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_745),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_791),
.B(n_571),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_781),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_783),
.Y(n_884)
);

OAI22x1_ASAP7_75t_R g885 ( 
.A1(n_748),
.A2(n_688),
.B1(n_727),
.B2(n_575),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_793),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_792),
.B(n_573),
.Y(n_887)
);

HB1xp67_ASAP7_75t_L g888 ( 
.A(n_815),
.Y(n_888)
);

INVx5_ASAP7_75t_L g889 ( 
.A(n_757),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_863),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_863),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_836),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_836),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_855),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_855),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_857),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_861),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_836),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_857),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_860),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_861),
.Y(n_901)
);

CKINVDCx6p67_ASAP7_75t_R g902 ( 
.A(n_840),
.Y(n_902)
);

OA21x2_ASAP7_75t_L g903 ( 
.A1(n_860),
.A2(n_604),
.B(n_584),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_854),
.B(n_729),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_861),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_881),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_881),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_854),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_836),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_854),
.Y(n_910)
);

INVxp67_ASAP7_75t_L g911 ( 
.A(n_844),
.Y(n_911)
);

OR2x2_ASAP7_75t_L g912 ( 
.A(n_858),
.B(n_782),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_865),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_861),
.Y(n_914)
);

CKINVDCx20_ASAP7_75t_R g915 ( 
.A(n_837),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_848),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_836),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_865),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_843),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_861),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_843),
.Y(n_921)
);

INVx4_ASAP7_75t_L g922 ( 
.A(n_848),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_847),
.B(n_741),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_848),
.B(n_784),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_872),
.B(n_785),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_847),
.B(n_760),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_871),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_851),
.B(n_796),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_856),
.A2(n_787),
.B1(n_816),
.B2(n_798),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_871),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_883),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_883),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_829),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_843),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_839),
.A2(n_720),
.B1(n_594),
.B2(n_756),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_874),
.Y(n_936)
);

INVx1_ASAP7_75t_SL g937 ( 
.A(n_833),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_874),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_874),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_829),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_829),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_827),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_827),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_862),
.B(n_777),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_856),
.A2(n_888),
.B1(n_886),
.B2(n_787),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_851),
.B(n_610),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_872),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_874),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_868),
.B(n_615),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_874),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_876),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_872),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_876),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_876),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_828),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_868),
.B(n_617),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_868),
.B(n_826),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_843),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_876),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_832),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_825),
.B(n_523),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_832),
.A2(n_768),
.B1(n_814),
.B2(n_761),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_826),
.B(n_873),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_876),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_843),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_867),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_867),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_867),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_835),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_852),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_889),
.B(n_789),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_828),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_830),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_826),
.B(n_873),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_830),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_831),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_852),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_969),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_894),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_906),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_922),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_913),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_L g983 ( 
.A1(n_916),
.A2(n_834),
.B1(n_825),
.B2(n_873),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_928),
.B(n_746),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_918),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_927),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_922),
.B(n_846),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_962),
.B(n_889),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_907),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_962),
.B(n_802),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_902),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_916),
.B(n_924),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_930),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_890),
.B(n_849),
.Y(n_994)
);

BUFx3_ASAP7_75t_L g995 ( 
.A(n_925),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_931),
.Y(n_996)
);

AND2x6_ASAP7_75t_L g997 ( 
.A(n_957),
.B(n_523),
.Y(n_997)
);

AND2x2_ASAP7_75t_SL g998 ( 
.A(n_912),
.B(n_944),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_924),
.B(n_889),
.Y(n_999)
);

INVxp33_ASAP7_75t_L g1000 ( 
.A(n_945),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_895),
.Y(n_1001)
);

INVxp67_ASAP7_75t_L g1002 ( 
.A(n_929),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_932),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_966),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_961),
.A2(n_834),
.B1(n_825),
.B2(n_869),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_891),
.B(n_850),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_967),
.Y(n_1007)
);

INVx5_ASAP7_75t_L g1008 ( 
.A(n_970),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_968),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_904),
.B(n_859),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_961),
.A2(n_834),
.B1(n_869),
.B2(n_686),
.Y(n_1011)
);

BUFx3_ASAP7_75t_L g1012 ( 
.A(n_925),
.Y(n_1012)
);

INVx2_ASAP7_75t_SL g1013 ( 
.A(n_928),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_947),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_896),
.Y(n_1015)
);

INVx1_ASAP7_75t_SL g1016 ( 
.A(n_915),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_SL g1017 ( 
.A1(n_915),
.A2(n_748),
.B1(n_775),
.B2(n_764),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_942),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_949),
.B(n_864),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_904),
.B(n_878),
.Y(n_1020)
);

INVx1_ASAP7_75t_SL g1021 ( 
.A(n_960),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_949),
.A2(n_887),
.B1(n_882),
.B2(n_816),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_947),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_952),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_923),
.B(n_926),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_971),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_892),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_952),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_937),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_908),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_910),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_892),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_923),
.B(n_889),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_971),
.B(n_800),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_911),
.B(n_802),
.Y(n_1035)
);

INVx5_ASAP7_75t_L g1036 ( 
.A(n_970),
.Y(n_1036)
);

INVx4_ASAP7_75t_L g1037 ( 
.A(n_970),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_926),
.B(n_831),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_911),
.B(n_744),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_935),
.A2(n_661),
.B1(n_707),
.B2(n_553),
.Y(n_1040)
);

OR2x2_ASAP7_75t_L g1041 ( 
.A(n_935),
.B(n_762),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_899),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_956),
.A2(n_637),
.B1(n_646),
.B2(n_625),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_900),
.Y(n_1044)
);

INVx4_ASAP7_75t_L g1045 ( 
.A(n_970),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_943),
.Y(n_1046)
);

NOR2x1p5_ASAP7_75t_L g1047 ( 
.A(n_956),
.B(n_576),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_957),
.B(n_841),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_936),
.B(n_866),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_955),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_938),
.B(n_866),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_939),
.B(n_803),
.Y(n_1052)
);

INVx1_ASAP7_75t_SL g1053 ( 
.A(n_946),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_948),
.B(n_539),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_972),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_973),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_975),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_976),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_950),
.B(n_823),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_903),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_946),
.Y(n_1061)
);

BUFx4f_ASAP7_75t_L g1062 ( 
.A(n_903),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_963),
.A2(n_665),
.B1(n_670),
.B2(n_664),
.Y(n_1063)
);

BUFx4f_ASAP7_75t_L g1064 ( 
.A(n_903),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_933),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_940),
.Y(n_1066)
);

AO22x2_ASAP7_75t_L g1067 ( 
.A1(n_963),
.A2(n_885),
.B1(n_880),
.B2(n_707),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_951),
.B(n_852),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_953),
.B(n_590),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_941),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_909),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_954),
.B(n_764),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_974),
.B(n_841),
.Y(n_1073)
);

CKINVDCx20_ASAP7_75t_R g1074 ( 
.A(n_959),
.Y(n_1074)
);

AND2x2_ASAP7_75t_SL g1075 ( 
.A(n_974),
.B(n_676),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_914),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_964),
.B(n_593),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_914),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_909),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_897),
.B(n_852),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_901),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_905),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_920),
.B(n_852),
.Y(n_1083)
);

INVx5_ASAP7_75t_L g1084 ( 
.A(n_892),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_977),
.B(n_695),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_SL g1086 ( 
.A(n_977),
.B(n_600),
.Y(n_1086)
);

INVx1_ASAP7_75t_SL g1087 ( 
.A(n_921),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_921),
.Y(n_1088)
);

CKINVDCx20_ASAP7_75t_R g1089 ( 
.A(n_958),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_958),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_892),
.B(n_775),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_893),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_893),
.B(n_799),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_893),
.Y(n_1094)
);

BUFx10_ASAP7_75t_L g1095 ( 
.A(n_893),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_898),
.Y(n_1096)
);

OR2x2_ASAP7_75t_L g1097 ( 
.A(n_898),
.B(n_761),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_898),
.B(n_799),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_898),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_917),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_917),
.B(n_845),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_917),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_917),
.B(n_697),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_965),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_965),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_919),
.B(n_934),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_965),
.Y(n_1107)
);

INVx4_ASAP7_75t_L g1108 ( 
.A(n_919),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_965),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_919),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_919),
.B(n_806),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_934),
.Y(n_1112)
);

INVx5_ASAP7_75t_L g1113 ( 
.A(n_934),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_913),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_1013),
.B(n_601),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_982),
.Y(n_1116)
);

BUFx5_ASAP7_75t_L g1117 ( 
.A(n_1060),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1049),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1020),
.B(n_711),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1010),
.B(n_725),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_1019),
.A2(n_726),
.B(n_537),
.C(n_635),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_984),
.B(n_716),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_1000),
.B(n_806),
.Y(n_1123)
);

NOR3xp33_ASAP7_75t_L g1124 ( 
.A(n_1017),
.B(n_822),
.C(n_820),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_992),
.B(n_870),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_1089),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_1025),
.A2(n_875),
.B(n_879),
.C(n_877),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_985),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1053),
.B(n_845),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_1053),
.B(n_546),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_1022),
.B(n_547),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_1002),
.B(n_833),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1061),
.B(n_562),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_994),
.B(n_577),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_1075),
.A2(n_512),
.B1(n_879),
.B2(n_877),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_1011),
.A2(n_1005),
.B(n_1006),
.C(n_1063),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_1086),
.B(n_579),
.Y(n_1137)
);

NAND2xp33_ASAP7_75t_SL g1138 ( 
.A(n_1047),
.B(n_580),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_986),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_993),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_1041),
.B(n_988),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1049),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1014),
.B(n_884),
.Y(n_1143)
);

AOI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1005),
.A2(n_583),
.B1(n_589),
.B2(n_581),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_1086),
.B(n_592),
.Y(n_1145)
);

INVx2_ASAP7_75t_SL g1146 ( 
.A(n_1097),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_1072),
.B(n_578),
.Y(n_1147)
);

INVx4_ASAP7_75t_L g1148 ( 
.A(n_995),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_1026),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_1011),
.B(n_599),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_987),
.B(n_605),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1051),
.Y(n_1152)
);

AOI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_983),
.A2(n_614),
.B1(n_616),
.B2(n_606),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_981),
.B(n_618),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_996),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1003),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1082),
.B(n_619),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1051),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1082),
.B(n_621),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1114),
.B(n_1033),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_990),
.B(n_591),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_979),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1023),
.B(n_884),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_1043),
.A2(n_630),
.B1(n_636),
.B2(n_626),
.Y(n_1164)
);

INVxp33_ASAP7_75t_L g1165 ( 
.A(n_1017),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1048),
.B(n_638),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1024),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1048),
.B(n_640),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1001),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1015),
.Y(n_1170)
);

INVx2_ASAP7_75t_SL g1171 ( 
.A(n_980),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1012),
.B(n_643),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1028),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_SL g1174 ( 
.A(n_991),
.Y(n_1174)
);

NOR2xp67_ASAP7_75t_L g1175 ( 
.A(n_1042),
.B(n_217),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1044),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_978),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_989),
.B(n_1074),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_998),
.B(n_644),
.Y(n_1179)
);

NOR2x1p5_ASAP7_75t_L g1180 ( 
.A(n_1029),
.B(n_595),
.Y(n_1180)
);

INVx2_ASAP7_75t_SL g1181 ( 
.A(n_1016),
.Y(n_1181)
);

NAND3xp33_ASAP7_75t_L g1182 ( 
.A(n_1004),
.B(n_648),
.C(n_647),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_1016),
.Y(n_1183)
);

INVxp67_ASAP7_75t_L g1184 ( 
.A(n_1091),
.Y(n_1184)
);

OR2x2_ASAP7_75t_L g1185 ( 
.A(n_1021),
.B(n_794),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1076),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_1027),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1021),
.B(n_568),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1039),
.B(n_596),
.Y(n_1189)
);

BUFx2_ASAP7_75t_L g1190 ( 
.A(n_1093),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1054),
.B(n_597),
.Y(n_1191)
);

INVxp67_ASAP7_75t_L g1192 ( 
.A(n_1098),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1007),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1038),
.B(n_650),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1073),
.B(n_651),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1073),
.B(n_652),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1035),
.B(n_568),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1008),
.B(n_654),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1087),
.B(n_657),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1009),
.A2(n_663),
.B1(n_666),
.B2(n_662),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1078),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1030),
.Y(n_1202)
);

INVxp67_ASAP7_75t_L g1203 ( 
.A(n_1111),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_1069),
.B(n_602),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_1008),
.B(n_669),
.Y(n_1205)
);

INVx2_ASAP7_75t_SL g1206 ( 
.A(n_1034),
.Y(n_1206)
);

INVxp67_ASAP7_75t_L g1207 ( 
.A(n_1052),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1077),
.B(n_608),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1031),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1087),
.B(n_674),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1059),
.B(n_568),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_997),
.B(n_678),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1101),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_997),
.B(n_680),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_1008),
.B(n_682),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_997),
.B(n_683),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_997),
.B(n_689),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1101),
.B(n_691),
.Y(n_1218)
);

INVx2_ASAP7_75t_SL g1219 ( 
.A(n_1065),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_1036),
.B(n_1084),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_1036),
.B(n_693),
.Y(n_1221)
);

NAND2xp33_ASAP7_75t_L g1222 ( 
.A(n_1027),
.B(n_694),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1050),
.Y(n_1223)
);

INVx8_ASAP7_75t_L g1224 ( 
.A(n_1027),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_999),
.B(n_609),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1018),
.B(n_696),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1046),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1040),
.B(n_611),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_1036),
.B(n_699),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1040),
.B(n_612),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_1084),
.B(n_705),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1056),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1057),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1058),
.Y(n_1234)
);

INVxp67_ASAP7_75t_L g1235 ( 
.A(n_1067),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1018),
.B(n_706),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1055),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1055),
.B(n_708),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1066),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1071),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1070),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_1081),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1079),
.B(n_710),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1032),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1032),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_1085),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1037),
.B(n_715),
.Y(n_1247)
);

CKINVDCx20_ASAP7_75t_R g1248 ( 
.A(n_1103),
.Y(n_1248)
);

AO22x2_ASAP7_75t_L g1249 ( 
.A1(n_1067),
.A2(n_797),
.B1(n_801),
.B2(n_795),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1088),
.Y(n_1250)
);

O2A1O1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1090),
.A2(n_838),
.B(n_835),
.C(n_805),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1062),
.A2(n_721),
.B1(n_722),
.B2(n_719),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1045),
.B(n_724),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1045),
.B(n_838),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1094),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1109),
.B(n_804),
.Y(n_1256)
);

INVx2_ASAP7_75t_SL g1257 ( 
.A(n_1064),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1112),
.B(n_623),
.Y(n_1258)
);

O2A1O1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1092),
.A2(n_1096),
.B(n_1104),
.C(n_1100),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1105),
.Y(n_1260)
);

INVx5_ASAP7_75t_L g1261 ( 
.A(n_1095),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1113),
.B(n_842),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1084),
.A2(n_842),
.B(n_853),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_SL g1264 ( 
.A(n_1099),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1102),
.Y(n_1265)
);

INVx3_ASAP7_75t_L g1266 ( 
.A(n_1032),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1107),
.Y(n_1267)
);

AOI22x1_ASAP7_75t_SL g1268 ( 
.A1(n_1110),
.A2(n_629),
.B1(n_634),
.B2(n_624),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1108),
.B(n_639),
.Y(n_1269)
);

NAND2xp33_ASAP7_75t_L g1270 ( 
.A(n_1113),
.B(n_645),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_SL g1271 ( 
.A(n_1113),
.B(n_842),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1106),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_1095),
.Y(n_1273)
);

INVxp33_ASAP7_75t_L g1274 ( 
.A(n_1080),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1083),
.Y(n_1275)
);

O2A1O1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1068),
.A2(n_808),
.B(n_809),
.C(n_807),
.Y(n_1276)
);

NOR3xp33_ASAP7_75t_L g1277 ( 
.A(n_1108),
.B(n_818),
.C(n_812),
.Y(n_1277)
);

AO22x1_ASAP7_75t_L g1278 ( 
.A1(n_1000),
.A2(n_655),
.B1(n_658),
.B2(n_649),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_982),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1075),
.A2(n_824),
.B1(n_819),
.B2(n_671),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1020),
.B(n_667),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1020),
.B(n_672),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1020),
.B(n_673),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_SL g1284 ( 
.A(n_1013),
.B(n_842),
.Y(n_1284)
);

NAND2xp33_ASAP7_75t_L g1285 ( 
.A(n_1019),
.B(n_677),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1020),
.B(n_681),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_982),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_1013),
.B(n_842),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_982),
.Y(n_1289)
);

INVxp67_ASAP7_75t_L g1290 ( 
.A(n_1072),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_SL g1291 ( 
.A(n_1013),
.B(n_685),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1020),
.B(n_692),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_982),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1020),
.B(n_698),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1020),
.B(n_702),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_982),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_982),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_981),
.A2(n_853),
.B(n_714),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_982),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1020),
.B(n_713),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1020),
.B(n_718),
.Y(n_1301)
);

INVxp67_ASAP7_75t_L g1302 ( 
.A(n_1072),
.Y(n_1302)
);

NAND2xp33_ASAP7_75t_L g1303 ( 
.A(n_1019),
.B(n_723),
.Y(n_1303)
);

CKINVDCx20_ASAP7_75t_R g1304 ( 
.A(n_991),
.Y(n_1304)
);

NOR2xp67_ASAP7_75t_L g1305 ( 
.A(n_981),
.B(n_219),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1049),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1020),
.B(n_728),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_982),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_982),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1020),
.B(n_853),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_1181),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1118),
.Y(n_1312)
);

AOI211xp5_ASAP7_75t_L g1313 ( 
.A1(n_1228),
.A2(n_3),
.B(n_1),
.C(n_2),
.Y(n_1313)
);

INVx2_ASAP7_75t_SL g1314 ( 
.A(n_1178),
.Y(n_1314)
);

OAI221xp5_ASAP7_75t_L g1315 ( 
.A1(n_1230),
.A2(n_5),
.B1(n_2),
.B2(n_4),
.C(n_7),
.Y(n_1315)
);

BUFx2_ASAP7_75t_L g1316 ( 
.A(n_1183),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1281),
.B(n_4),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1116),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1290),
.B(n_1302),
.Y(n_1319)
);

INVx4_ASAP7_75t_L g1320 ( 
.A(n_1261),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1189),
.A2(n_853),
.B1(n_221),
.B2(n_223),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_SL g1322 ( 
.A(n_1246),
.B(n_853),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_SL g1323 ( 
.A(n_1184),
.B(n_220),
.Y(n_1323)
);

BUFx8_ASAP7_75t_L g1324 ( 
.A(n_1174),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1282),
.B(n_7),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1149),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_SL g1327 ( 
.A1(n_1147),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1150),
.A2(n_12),
.B1(n_9),
.B2(n_11),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1283),
.B(n_11),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1286),
.B(n_13),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1142),
.Y(n_1331)
);

AND2x4_ASAP7_75t_SL g1332 ( 
.A(n_1178),
.B(n_224),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1128),
.Y(n_1333)
);

BUFx4f_ASAP7_75t_L g1334 ( 
.A(n_1149),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1139),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1305),
.A2(n_232),
.B(n_227),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1152),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1192),
.B(n_233),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1211),
.B(n_13),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1136),
.A2(n_236),
.B(n_234),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1140),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1155),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1292),
.B(n_15),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1294),
.B(n_16),
.Y(n_1344)
);

NAND2x1p5_ASAP7_75t_L g1345 ( 
.A(n_1261),
.B(n_237),
.Y(n_1345)
);

BUFx3_ASAP7_75t_L g1346 ( 
.A(n_1126),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1141),
.A2(n_239),
.B1(n_240),
.B2(n_238),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1158),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1156),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1279),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_1304),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1287),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1295),
.B(n_17),
.Y(n_1353)
);

OAI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1213),
.A2(n_1160),
.B(n_1166),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1306),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1289),
.Y(n_1356)
);

INVx2_ASAP7_75t_SL g1357 ( 
.A(n_1185),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1300),
.B(n_17),
.Y(n_1358)
);

INVx2_ASAP7_75t_SL g1359 ( 
.A(n_1188),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1301),
.B(n_1307),
.Y(n_1360)
);

A2O1A1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1191),
.A2(n_20),
.B(n_18),
.C(n_19),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_SL g1362 ( 
.A(n_1203),
.B(n_242),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_1149),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1134),
.B(n_18),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_SL g1365 ( 
.A(n_1261),
.B(n_244),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1273),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1122),
.A2(n_1285),
.B1(n_1303),
.B2(n_1208),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1293),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1296),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1146),
.B(n_248),
.Y(n_1370)
);

INVx2_ASAP7_75t_SL g1371 ( 
.A(n_1171),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_1187),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1201),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1256),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1207),
.B(n_19),
.Y(n_1375)
);

INVx5_ASAP7_75t_L g1376 ( 
.A(n_1224),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1310),
.A2(n_252),
.B(n_250),
.Y(n_1377)
);

INVx5_ASAP7_75t_L g1378 ( 
.A(n_1224),
.Y(n_1378)
);

INVx3_ASAP7_75t_L g1379 ( 
.A(n_1265),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_1174),
.Y(n_1380)
);

AND2x2_ASAP7_75t_SL g1381 ( 
.A(n_1190),
.B(n_1204),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1186),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1187),
.Y(n_1383)
);

BUFx2_ASAP7_75t_L g1384 ( 
.A(n_1187),
.Y(n_1384)
);

NOR2x1p5_ASAP7_75t_L g1385 ( 
.A(n_1148),
.B(n_1167),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1297),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1125),
.B(n_1197),
.Y(n_1387)
);

INVx5_ASAP7_75t_L g1388 ( 
.A(n_1224),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1148),
.B(n_253),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1144),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1119),
.B(n_22),
.Y(n_1391)
);

OR2x6_ASAP7_75t_L g1392 ( 
.A(n_1206),
.B(n_23),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1299),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1161),
.B(n_24),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_1248),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1168),
.B(n_24),
.Y(n_1396)
);

INVx5_ASAP7_75t_L g1397 ( 
.A(n_1244),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_R g1398 ( 
.A(n_1138),
.B(n_254),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1195),
.B(n_26),
.Y(n_1399)
);

NAND2x1p5_ASAP7_75t_L g1400 ( 
.A(n_1244),
.B(n_257),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1173),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1209),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_1244),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1120),
.A2(n_259),
.B1(n_260),
.B2(n_258),
.Y(n_1404)
);

OAI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1196),
.A2(n_262),
.B(n_261),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1308),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_1245),
.Y(n_1407)
);

NAND2x1p5_ASAP7_75t_L g1408 ( 
.A(n_1245),
.B(n_1266),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1309),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1153),
.A2(n_265),
.B1(n_266),
.B2(n_264),
.Y(n_1410)
);

BUFx2_ASAP7_75t_SL g1411 ( 
.A(n_1264),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1129),
.B(n_27),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1133),
.B(n_28),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1143),
.Y(n_1414)
);

BUFx6f_ASAP7_75t_L g1415 ( 
.A(n_1245),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1272),
.B(n_29),
.Y(n_1416)
);

OAI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1144),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1163),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1151),
.B(n_30),
.Y(n_1419)
);

BUFx6f_ASAP7_75t_L g1420 ( 
.A(n_1242),
.Y(n_1420)
);

O2A1O1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1121),
.A2(n_33),
.B(n_31),
.C(n_32),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1157),
.B(n_267),
.Y(n_1422)
);

BUFx12f_ASAP7_75t_L g1423 ( 
.A(n_1180),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1176),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_SL g1425 ( 
.A(n_1159),
.B(n_268),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1193),
.B(n_34),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1202),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1232),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1260),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1275),
.B(n_34),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1264),
.Y(n_1431)
);

NAND3xp33_ASAP7_75t_L g1432 ( 
.A(n_1123),
.B(n_35),
.C(n_36),
.Y(n_1432)
);

NAND2xp33_ASAP7_75t_L g1433 ( 
.A(n_1117),
.B(n_269),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1223),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1115),
.B(n_35),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1239),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1241),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1233),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1165),
.B(n_36),
.Y(n_1439)
);

AND2x4_ASAP7_75t_L g1440 ( 
.A(n_1177),
.B(n_271),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1194),
.B(n_37),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1235),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1154),
.A2(n_273),
.B(n_272),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_SL g1444 ( 
.A(n_1199),
.B(n_276),
.Y(n_1444)
);

OR2x6_ASAP7_75t_L g1445 ( 
.A(n_1219),
.B(n_37),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1162),
.B(n_277),
.Y(n_1446)
);

INVx3_ASAP7_75t_L g1447 ( 
.A(n_1169),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1130),
.B(n_1258),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_1170),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_L g1450 ( 
.A(n_1234),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1227),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1267),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1240),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1274),
.B(n_38),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1131),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_1455)
);

CKINVDCx20_ASAP7_75t_R g1456 ( 
.A(n_1268),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1237),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1172),
.B(n_278),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1255),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1124),
.B(n_41),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1210),
.B(n_42),
.Y(n_1461)
);

INVx1_ASAP7_75t_SL g1462 ( 
.A(n_1291),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1266),
.Y(n_1463)
);

INVx2_ASAP7_75t_SL g1464 ( 
.A(n_1249),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_1257),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1225),
.B(n_43),
.Y(n_1466)
);

BUFx6f_ASAP7_75t_L g1467 ( 
.A(n_1250),
.Y(n_1467)
);

AND2x2_ASAP7_75t_SL g1468 ( 
.A(n_1132),
.B(n_43),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1269),
.B(n_44),
.Y(n_1469)
);

OAI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1153),
.A2(n_281),
.B(n_279),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1117),
.Y(n_1471)
);

AOI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1179),
.A2(n_283),
.B1(n_284),
.B2(n_282),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1137),
.A2(n_47),
.B1(n_44),
.B2(n_46),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1127),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1251),
.Y(n_1475)
);

NAND2xp33_ASAP7_75t_L g1476 ( 
.A(n_1117),
.B(n_286),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1145),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1254),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1276),
.Y(n_1479)
);

AO22x1_ASAP7_75t_L g1480 ( 
.A1(n_1277),
.A2(n_49),
.B1(n_46),
.B2(n_47),
.Y(n_1480)
);

AND2x6_ASAP7_75t_L g1481 ( 
.A(n_1218),
.B(n_287),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1259),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1117),
.B(n_1280),
.Y(n_1483)
);

NAND2x1p5_ASAP7_75t_L g1484 ( 
.A(n_1220),
.B(n_288),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_1278),
.Y(n_1485)
);

INVxp67_ASAP7_75t_L g1486 ( 
.A(n_1249),
.Y(n_1486)
);

BUFx2_ASAP7_75t_L g1487 ( 
.A(n_1117),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1226),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1284),
.B(n_289),
.Y(n_1489)
);

INVxp67_ASAP7_75t_SL g1490 ( 
.A(n_1175),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1135),
.B(n_49),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1236),
.Y(n_1492)
);

XOR2x2_ASAP7_75t_SL g1493 ( 
.A(n_1252),
.B(n_50),
.Y(n_1493)
);

INVx2_ASAP7_75t_SL g1494 ( 
.A(n_1238),
.Y(n_1494)
);

INVx3_ASAP7_75t_L g1495 ( 
.A(n_1243),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1252),
.B(n_50),
.Y(n_1496)
);

NAND2xp33_ASAP7_75t_SL g1497 ( 
.A(n_1288),
.B(n_51),
.Y(n_1497)
);

CKINVDCx20_ASAP7_75t_R g1498 ( 
.A(n_1200),
.Y(n_1498)
);

INVx1_ASAP7_75t_SL g1499 ( 
.A(n_1200),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1247),
.B(n_51),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1212),
.B(n_52),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1175),
.Y(n_1502)
);

NAND3xp33_ASAP7_75t_SL g1503 ( 
.A(n_1182),
.B(n_53),
.C(n_54),
.Y(n_1503)
);

INVx2_ASAP7_75t_SL g1504 ( 
.A(n_1182),
.Y(n_1504)
);

INVx1_ASAP7_75t_SL g1505 ( 
.A(n_1222),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1253),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_SL g1507 ( 
.A(n_1214),
.B(n_290),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1216),
.B(n_54),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1262),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1217),
.B(n_56),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1164),
.B(n_56),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1271),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1270),
.B(n_1198),
.Y(n_1513)
);

INVx3_ASAP7_75t_L g1514 ( 
.A(n_1205),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1334),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1318),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_1366),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1387),
.B(n_1215),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1316),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1360),
.B(n_1221),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1414),
.B(n_1229),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1333),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1418),
.B(n_1231),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1335),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1341),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1427),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1478),
.B(n_1298),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_SL g1528 ( 
.A(n_1357),
.B(n_1263),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1316),
.Y(n_1529)
);

BUFx2_ASAP7_75t_L g1530 ( 
.A(n_1311),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1442),
.Y(n_1531)
);

INVx3_ASAP7_75t_L g1532 ( 
.A(n_1376),
.Y(n_1532)
);

OR2x6_ASAP7_75t_L g1533 ( 
.A(n_1411),
.B(n_291),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1499),
.B(n_57),
.Y(n_1534)
);

INVx3_ASAP7_75t_L g1535 ( 
.A(n_1376),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1374),
.B(n_58),
.Y(n_1536)
);

INVx5_ASAP7_75t_L g1537 ( 
.A(n_1376),
.Y(n_1537)
);

INVxp67_ASAP7_75t_L g1538 ( 
.A(n_1319),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1342),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1349),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1381),
.B(n_58),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1354),
.B(n_59),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1498),
.B(n_60),
.Y(n_1543)
);

BUFx6f_ASAP7_75t_L g1544 ( 
.A(n_1372),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1468),
.B(n_60),
.Y(n_1545)
);

BUFx2_ASAP7_75t_L g1546 ( 
.A(n_1395),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1350),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1492),
.B(n_61),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1352),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1506),
.B(n_62),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1359),
.B(n_1314),
.Y(n_1551)
);

BUFx6f_ASAP7_75t_L g1552 ( 
.A(n_1372),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1394),
.B(n_63),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1356),
.Y(n_1554)
);

OAI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1367),
.A2(n_1490),
.B1(n_1483),
.B2(n_1448),
.Y(n_1555)
);

AOI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1485),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_1556)
);

OR2x6_ASAP7_75t_L g1557 ( 
.A(n_1320),
.B(n_1326),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1368),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1488),
.B(n_64),
.Y(n_1559)
);

BUFx3_ASAP7_75t_L g1560 ( 
.A(n_1326),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1462),
.B(n_65),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1369),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1339),
.B(n_66),
.Y(n_1563)
);

A2O1A1Ixp33_ASAP7_75t_L g1564 ( 
.A1(n_1470),
.A2(n_69),
.B(n_66),
.C(n_67),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1386),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1393),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1406),
.Y(n_1567)
);

INVx4_ASAP7_75t_L g1568 ( 
.A(n_1378),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1378),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1409),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_1324),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1363),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1424),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1493),
.B(n_69),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1434),
.Y(n_1575)
);

INVx5_ASAP7_75t_L g1576 ( 
.A(n_1378),
.Y(n_1576)
);

BUFx6f_ASAP7_75t_L g1577 ( 
.A(n_1372),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1436),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1363),
.Y(n_1579)
);

INVx3_ASAP7_75t_L g1580 ( 
.A(n_1388),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1437),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1412),
.B(n_71),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1402),
.Y(n_1583)
);

NOR2x2_ASAP7_75t_L g1584 ( 
.A(n_1392),
.B(n_71),
.Y(n_1584)
);

A2O1A1Ixp33_ASAP7_75t_L g1585 ( 
.A1(n_1469),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1452),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1494),
.B(n_74),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1451),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1373),
.Y(n_1589)
);

A2O1A1Ixp33_ASAP7_75t_L g1590 ( 
.A1(n_1466),
.A2(n_77),
.B(n_75),
.C(n_76),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1428),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_1351),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1487),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1429),
.Y(n_1594)
);

BUFx6f_ASAP7_75t_L g1595 ( 
.A(n_1403),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1438),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1382),
.Y(n_1597)
);

INVx2_ASAP7_75t_SL g1598 ( 
.A(n_1420),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1495),
.B(n_77),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1312),
.Y(n_1600)
);

INVxp67_ASAP7_75t_L g1601 ( 
.A(n_1420),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1317),
.B(n_78),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1331),
.Y(n_1603)
);

NAND2x1p5_ASAP7_75t_L g1604 ( 
.A(n_1388),
.B(n_294),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1487),
.Y(n_1605)
);

BUFx2_ASAP7_75t_L g1606 ( 
.A(n_1346),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1401),
.Y(n_1607)
);

BUFx3_ASAP7_75t_L g1608 ( 
.A(n_1379),
.Y(n_1608)
);

AOI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1458),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1496),
.A2(n_82),
.B1(n_79),
.B2(n_80),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1325),
.B(n_83),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1384),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1457),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1375),
.B(n_83),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1459),
.Y(n_1615)
);

INVx3_ASAP7_75t_L g1616 ( 
.A(n_1388),
.Y(n_1616)
);

BUFx3_ASAP7_75t_L g1617 ( 
.A(n_1324),
.Y(n_1617)
);

BUFx6f_ASAP7_75t_L g1618 ( 
.A(n_1403),
.Y(n_1618)
);

BUFx2_ASAP7_75t_L g1619 ( 
.A(n_1384),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1439),
.B(n_84),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1329),
.B(n_85),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1337),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1348),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1435),
.B(n_85),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1474),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1482),
.Y(n_1626)
);

AND3x1_ASAP7_75t_SL g1627 ( 
.A(n_1315),
.B(n_1385),
.C(n_1313),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1355),
.Y(n_1628)
);

INVx3_ASAP7_75t_L g1629 ( 
.A(n_1463),
.Y(n_1629)
);

BUFx6f_ASAP7_75t_L g1630 ( 
.A(n_1403),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_1423),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1511),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1486),
.B(n_86),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1453),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1447),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1463),
.Y(n_1636)
);

BUFx6f_ASAP7_75t_L g1637 ( 
.A(n_1407),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1332),
.B(n_88),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1330),
.B(n_1343),
.Y(n_1639)
);

BUFx6f_ASAP7_75t_L g1640 ( 
.A(n_1407),
.Y(n_1640)
);

BUFx6f_ASAP7_75t_L g1641 ( 
.A(n_1407),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1449),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1450),
.Y(n_1643)
);

BUFx2_ASAP7_75t_L g1644 ( 
.A(n_1464),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1465),
.B(n_295),
.Y(n_1645)
);

BUFx6f_ASAP7_75t_L g1646 ( 
.A(n_1383),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1344),
.B(n_89),
.Y(n_1647)
);

INVx3_ASAP7_75t_L g1648 ( 
.A(n_1467),
.Y(n_1648)
);

INVx5_ASAP7_75t_L g1649 ( 
.A(n_1397),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1353),
.B(n_89),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1358),
.B(n_91),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1450),
.Y(n_1652)
);

AOI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1433),
.A2(n_297),
.B(n_296),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1491),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1465),
.B(n_510),
.Y(n_1655)
);

A2O1A1Ixp33_ASAP7_75t_L g1656 ( 
.A1(n_1364),
.A2(n_94),
.B(n_92),
.C(n_93),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1465),
.B(n_509),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1396),
.B(n_95),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1467),
.Y(n_1659)
);

INVxp33_ASAP7_75t_L g1660 ( 
.A(n_1431),
.Y(n_1660)
);

NAND2x1p5_ASAP7_75t_L g1661 ( 
.A(n_1397),
.B(n_298),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1477),
.B(n_95),
.Y(n_1662)
);

INVx3_ASAP7_75t_L g1663 ( 
.A(n_1467),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1460),
.B(n_96),
.Y(n_1664)
);

INVx3_ASAP7_75t_L g1665 ( 
.A(n_1440),
.Y(n_1665)
);

BUFx3_ASAP7_75t_L g1666 ( 
.A(n_1371),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1399),
.B(n_96),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1471),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1390),
.A2(n_1510),
.B1(n_1508),
.B2(n_1503),
.Y(n_1669)
);

BUFx2_ASAP7_75t_L g1670 ( 
.A(n_1370),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1461),
.B(n_98),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1408),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1391),
.B(n_98),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1454),
.B(n_99),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1413),
.B(n_1441),
.Y(n_1675)
);

BUFx2_ASAP7_75t_L g1676 ( 
.A(n_1370),
.Y(n_1676)
);

BUFx10_ASAP7_75t_L g1677 ( 
.A(n_1380),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1475),
.Y(n_1678)
);

AOI22x1_ASAP7_75t_L g1679 ( 
.A1(n_1340),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1477),
.B(n_100),
.Y(n_1680)
);

BUFx2_ASAP7_75t_L g1681 ( 
.A(n_1383),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1440),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1509),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1512),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1416),
.Y(n_1685)
);

NOR2x1_ASAP7_75t_L g1686 ( 
.A(n_1513),
.B(n_1432),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1502),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1426),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1430),
.B(n_103),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1419),
.B(n_105),
.Y(n_1690)
);

INVx3_ASAP7_75t_L g1691 ( 
.A(n_1446),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1504),
.B(n_105),
.Y(n_1692)
);

BUFx2_ASAP7_75t_L g1693 ( 
.A(n_1415),
.Y(n_1693)
);

CKINVDCx6p67_ASAP7_75t_R g1694 ( 
.A(n_1445),
.Y(n_1694)
);

AND2x2_ASAP7_75t_SL g1695 ( 
.A(n_1476),
.B(n_106),
.Y(n_1695)
);

BUFx2_ASAP7_75t_L g1696 ( 
.A(n_1415),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1446),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1392),
.B(n_107),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1514),
.B(n_108),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1397),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1505),
.B(n_108),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1389),
.B(n_299),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_SL g1703 ( 
.A(n_1389),
.B(n_109),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1688),
.B(n_1500),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1516),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1516),
.Y(n_1706)
);

INVx2_ASAP7_75t_SL g1707 ( 
.A(n_1517),
.Y(n_1707)
);

AOI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1527),
.A2(n_1405),
.B(n_1444),
.Y(n_1708)
);

OAI21x1_ASAP7_75t_L g1709 ( 
.A1(n_1626),
.A2(n_1377),
.B(n_1336),
.Y(n_1709)
);

AOI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1555),
.A2(n_1675),
.B(n_1639),
.Y(n_1710)
);

OAI21x1_ASAP7_75t_L g1711 ( 
.A1(n_1625),
.A2(n_1443),
.B(n_1507),
.Y(n_1711)
);

INVx2_ASAP7_75t_SL g1712 ( 
.A(n_1608),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1670),
.B(n_1489),
.Y(n_1713)
);

OAI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1669),
.A2(n_1479),
.B(n_1501),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1685),
.B(n_1327),
.Y(n_1715)
);

AO21x1_ASAP7_75t_L g1716 ( 
.A1(n_1542),
.A2(n_1421),
.B(n_1417),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1538),
.B(n_1520),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1647),
.B(n_1455),
.Y(n_1718)
);

O2A1O1Ixp5_ASAP7_75t_L g1719 ( 
.A1(n_1564),
.A2(n_1410),
.B(n_1425),
.C(n_1422),
.Y(n_1719)
);

OAI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1686),
.A2(n_1361),
.B(n_1472),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1650),
.B(n_1328),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1522),
.Y(n_1722)
);

OAI21x1_ASAP7_75t_L g1723 ( 
.A1(n_1625),
.A2(n_1404),
.B(n_1400),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1620),
.B(n_1445),
.Y(n_1724)
);

AOI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1653),
.A2(n_1338),
.B(n_1323),
.Y(n_1725)
);

AOI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1695),
.A2(n_1362),
.B(n_1365),
.Y(n_1726)
);

BUFx2_ASAP7_75t_L g1727 ( 
.A(n_1519),
.Y(n_1727)
);

NOR2x1_ASAP7_75t_L g1728 ( 
.A(n_1568),
.B(n_1322),
.Y(n_1728)
);

INVx2_ASAP7_75t_SL g1729 ( 
.A(n_1560),
.Y(n_1729)
);

OAI21x1_ASAP7_75t_L g1730 ( 
.A1(n_1678),
.A2(n_1679),
.B(n_1668),
.Y(n_1730)
);

AO31x2_ASAP7_75t_L g1731 ( 
.A1(n_1593),
.A2(n_1347),
.A3(n_1481),
.B(n_1321),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1559),
.B(n_1473),
.Y(n_1732)
);

OAI21x1_ASAP7_75t_L g1733 ( 
.A1(n_1679),
.A2(n_1484),
.B(n_1345),
.Y(n_1733)
);

BUFx6f_ASAP7_75t_L g1734 ( 
.A(n_1649),
.Y(n_1734)
);

INVx4_ASAP7_75t_L g1735 ( 
.A(n_1649),
.Y(n_1735)
);

AOI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1665),
.A2(n_1691),
.B(n_1682),
.Y(n_1736)
);

AOI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1665),
.A2(n_1497),
.B(n_1480),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1664),
.B(n_1398),
.Y(n_1738)
);

NAND3x1_ASAP7_75t_L g1739 ( 
.A(n_1556),
.B(n_1456),
.C(n_109),
.Y(n_1739)
);

OAI21x1_ASAP7_75t_L g1740 ( 
.A1(n_1668),
.A2(n_1481),
.B(n_304),
.Y(n_1740)
);

INVxp67_ASAP7_75t_L g1741 ( 
.A(n_1594),
.Y(n_1741)
);

CKINVDCx11_ASAP7_75t_R g1742 ( 
.A(n_1677),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1518),
.B(n_1481),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1676),
.B(n_302),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_SL g1745 ( 
.A(n_1691),
.B(n_110),
.Y(n_1745)
);

INVx3_ASAP7_75t_L g1746 ( 
.A(n_1649),
.Y(n_1746)
);

OAI21x1_ASAP7_75t_L g1747 ( 
.A1(n_1528),
.A2(n_307),
.B(n_306),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1529),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1607),
.B(n_111),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1624),
.B(n_111),
.Y(n_1750)
);

A2O1A1Ixp33_ASAP7_75t_L g1751 ( 
.A1(n_1614),
.A2(n_114),
.B(n_112),
.C(n_113),
.Y(n_1751)
);

NAND2x1p5_ASAP7_75t_L g1752 ( 
.A(n_1537),
.B(n_308),
.Y(n_1752)
);

OA21x2_ASAP7_75t_L g1753 ( 
.A1(n_1593),
.A2(n_1605),
.B(n_1582),
.Y(n_1753)
);

INVx5_ASAP7_75t_L g1754 ( 
.A(n_1537),
.Y(n_1754)
);

INVx3_ASAP7_75t_L g1755 ( 
.A(n_1666),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_SL g1756 ( 
.A(n_1571),
.B(n_309),
.Y(n_1756)
);

A2O1A1Ixp33_ASAP7_75t_L g1757 ( 
.A1(n_1602),
.A2(n_117),
.B(n_115),
.C(n_116),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1549),
.Y(n_1758)
);

AOI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1682),
.A2(n_508),
.B(n_312),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1541),
.B(n_117),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1522),
.Y(n_1761)
);

OAI21x1_ASAP7_75t_SL g1762 ( 
.A1(n_1692),
.A2(n_118),
.B(n_119),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1524),
.Y(n_1763)
);

OA22x2_ASAP7_75t_L g1764 ( 
.A1(n_1574),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_1764)
);

BUFx2_ASAP7_75t_L g1765 ( 
.A(n_1612),
.Y(n_1765)
);

AND2x4_ASAP7_75t_L g1766 ( 
.A(n_1643),
.B(n_310),
.Y(n_1766)
);

INVx3_ASAP7_75t_L g1767 ( 
.A(n_1648),
.Y(n_1767)
);

AOI21xp33_ASAP7_75t_L g1768 ( 
.A1(n_1667),
.A2(n_120),
.B(n_121),
.Y(n_1768)
);

INVx3_ASAP7_75t_SL g1769 ( 
.A(n_1694),
.Y(n_1769)
);

OAI21x1_ASAP7_75t_L g1770 ( 
.A1(n_1697),
.A2(n_314),
.B(n_313),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1548),
.B(n_121),
.Y(n_1771)
);

AOI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1697),
.A2(n_507),
.B(n_317),
.Y(n_1772)
);

OAI21x1_ASAP7_75t_L g1773 ( 
.A1(n_1605),
.A2(n_318),
.B(n_316),
.Y(n_1773)
);

AO31x2_ASAP7_75t_L g1774 ( 
.A1(n_1585),
.A2(n_1656),
.A3(n_1590),
.B(n_1621),
.Y(n_1774)
);

AO21x1_ASAP7_75t_L g1775 ( 
.A1(n_1671),
.A2(n_122),
.B(n_123),
.Y(n_1775)
);

INVx3_ASAP7_75t_L g1776 ( 
.A(n_1648),
.Y(n_1776)
);

OA22x2_ASAP7_75t_L g1777 ( 
.A1(n_1609),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1550),
.B(n_124),
.Y(n_1778)
);

NAND2x1p5_ASAP7_75t_L g1779 ( 
.A(n_1537),
.B(n_319),
.Y(n_1779)
);

AOI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1702),
.A2(n_1690),
.B(n_1611),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1689),
.B(n_1702),
.Y(n_1781)
);

OAI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1521),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_1782)
);

OAI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1523),
.A2(n_129),
.B1(n_126),
.B2(n_128),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_SL g1784 ( 
.A(n_1534),
.B(n_128),
.Y(n_1784)
);

AOI21x1_ASAP7_75t_L g1785 ( 
.A1(n_1673),
.A2(n_325),
.B(n_324),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1674),
.B(n_129),
.Y(n_1786)
);

OAI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1553),
.A2(n_130),
.B(n_131),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1558),
.Y(n_1788)
);

OAI22x1_ASAP7_75t_L g1789 ( 
.A1(n_1545),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.Y(n_1789)
);

INVx1_ASAP7_75t_SL g1790 ( 
.A(n_1530),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1525),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_SL g1792 ( 
.A(n_1599),
.B(n_132),
.Y(n_1792)
);

OAI21x1_ASAP7_75t_L g1793 ( 
.A1(n_1547),
.A2(n_328),
.B(n_326),
.Y(n_1793)
);

OAI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1658),
.A2(n_1651),
.B(n_1632),
.Y(n_1794)
);

AO32x2_ASAP7_75t_L g1795 ( 
.A1(n_1687),
.A2(n_133),
.A3(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_1795)
);

NAND3xp33_ASAP7_75t_L g1796 ( 
.A(n_1610),
.B(n_134),
.C(n_136),
.Y(n_1796)
);

NAND2x1p5_ASAP7_75t_L g1797 ( 
.A(n_1576),
.B(n_329),
.Y(n_1797)
);

BUFx2_ASAP7_75t_L g1798 ( 
.A(n_1619),
.Y(n_1798)
);

AOI21x1_ASAP7_75t_L g1799 ( 
.A1(n_1547),
.A2(n_333),
.B(n_331),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1565),
.Y(n_1800)
);

OAI21x1_ASAP7_75t_L g1801 ( 
.A1(n_1565),
.A2(n_1581),
.B(n_1575),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1575),
.Y(n_1802)
);

AOI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1703),
.A2(n_335),
.B(n_334),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1581),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1526),
.B(n_1562),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1566),
.Y(n_1806)
);

BUFx2_ASAP7_75t_L g1807 ( 
.A(n_1606),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1567),
.Y(n_1808)
);

INVx3_ASAP7_75t_L g1809 ( 
.A(n_1572),
.Y(n_1809)
);

A2O1A1Ixp33_ASAP7_75t_L g1810 ( 
.A1(n_1699),
.A2(n_139),
.B(n_137),
.C(n_138),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1570),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1563),
.B(n_137),
.Y(n_1812)
);

AOI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1683),
.A2(n_339),
.B(n_337),
.Y(n_1813)
);

NAND2x1_ASAP7_75t_L g1814 ( 
.A(n_1568),
.B(n_342),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1573),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1578),
.B(n_138),
.Y(n_1816)
);

INVx6_ASAP7_75t_L g1817 ( 
.A(n_1677),
.Y(n_1817)
);

INVx3_ASAP7_75t_L g1818 ( 
.A(n_1557),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1583),
.B(n_140),
.Y(n_1819)
);

AOI21xp5_ASAP7_75t_L g1820 ( 
.A1(n_1684),
.A2(n_506),
.B(n_346),
.Y(n_1820)
);

OAI21x1_ASAP7_75t_L g1821 ( 
.A1(n_1634),
.A2(n_1615),
.B(n_1613),
.Y(n_1821)
);

AOI21x1_ASAP7_75t_L g1822 ( 
.A1(n_1644),
.A2(n_347),
.B(n_344),
.Y(n_1822)
);

NAND3xp33_ASAP7_75t_SL g1823 ( 
.A(n_1543),
.B(n_141),
.C(n_142),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1536),
.B(n_142),
.Y(n_1824)
);

OAI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1654),
.A2(n_143),
.B(n_144),
.Y(n_1825)
);

AOI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1576),
.A2(n_504),
.B(n_350),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1638),
.B(n_143),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_1546),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1588),
.B(n_1591),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1539),
.Y(n_1830)
);

OAI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1587),
.A2(n_144),
.B(n_145),
.Y(n_1831)
);

OAI21x1_ASAP7_75t_L g1832 ( 
.A1(n_1634),
.A2(n_1554),
.B(n_1540),
.Y(n_1832)
);

AOI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1576),
.A2(n_353),
.B(n_352),
.Y(n_1833)
);

AOI211x1_ASAP7_75t_L g1834 ( 
.A1(n_1662),
.A2(n_148),
.B(n_146),
.C(n_147),
.Y(n_1834)
);

AND3x2_ASAP7_75t_L g1835 ( 
.A(n_1561),
.B(n_147),
.C(n_150),
.Y(n_1835)
);

INVx2_ASAP7_75t_SL g1836 ( 
.A(n_1598),
.Y(n_1836)
);

A2O1A1Ixp33_ASAP7_75t_L g1837 ( 
.A1(n_1680),
.A2(n_153),
.B(n_151),
.C(n_152),
.Y(n_1837)
);

NAND2x1_ASAP7_75t_L g1838 ( 
.A(n_1532),
.B(n_355),
.Y(n_1838)
);

AO21x1_ASAP7_75t_L g1839 ( 
.A1(n_1701),
.A2(n_151),
.B(n_152),
.Y(n_1839)
);

OAI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1589),
.A2(n_1551),
.B(n_1628),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1586),
.Y(n_1841)
);

AOI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1627),
.A2(n_155),
.B1(n_153),
.B2(n_154),
.Y(n_1842)
);

OAI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1531),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_1843)
);

A2O1A1Ixp33_ASAP7_75t_L g1844 ( 
.A1(n_1633),
.A2(n_159),
.B(n_157),
.C(n_158),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_SL g1845 ( 
.A(n_1592),
.B(n_158),
.Y(n_1845)
);

OAI21x1_ASAP7_75t_L g1846 ( 
.A1(n_1663),
.A2(n_360),
.B(n_357),
.Y(n_1846)
);

OAI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1635),
.A2(n_161),
.B1(n_159),
.B2(n_160),
.Y(n_1847)
);

INVxp67_ASAP7_75t_SL g1848 ( 
.A(n_1663),
.Y(n_1848)
);

OA21x2_ASAP7_75t_L g1849 ( 
.A1(n_1596),
.A2(n_1597),
.B(n_1600),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1603),
.Y(n_1850)
);

OAI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1642),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.Y(n_1851)
);

NOR2x1_ASAP7_75t_SL g1852 ( 
.A(n_1533),
.B(n_361),
.Y(n_1852)
);

OAI21x1_ASAP7_75t_L g1853 ( 
.A1(n_1661),
.A2(n_363),
.B(n_362),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1660),
.B(n_364),
.Y(n_1854)
);

INVxp67_ASAP7_75t_SL g1855 ( 
.A(n_1622),
.Y(n_1855)
);

OA21x2_ASAP7_75t_L g1856 ( 
.A1(n_1623),
.A2(n_366),
.B(n_365),
.Y(n_1856)
);

NOR2xp67_ASAP7_75t_L g1857 ( 
.A(n_1652),
.B(n_367),
.Y(n_1857)
);

AOI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1604),
.A2(n_503),
.B(n_373),
.Y(n_1858)
);

OAI21x1_ASAP7_75t_L g1859 ( 
.A1(n_1535),
.A2(n_1580),
.B(n_1569),
.Y(n_1859)
);

AOI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1645),
.A2(n_163),
.B1(n_166),
.B2(n_167),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1698),
.B(n_166),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1659),
.B(n_167),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_1742),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1710),
.B(n_1645),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1705),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1704),
.B(n_1780),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1748),
.B(n_1579),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1758),
.Y(n_1868)
);

AOI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1721),
.A2(n_1533),
.B1(n_1657),
.B2(n_1655),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_L g1870 ( 
.A(n_1717),
.B(n_1601),
.Y(n_1870)
);

OAI22xp5_ASAP7_75t_L g1871 ( 
.A1(n_1718),
.A2(n_1732),
.B1(n_1715),
.B2(n_1781),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1788),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1806),
.Y(n_1873)
);

BUFx6f_ASAP7_75t_L g1874 ( 
.A(n_1734),
.Y(n_1874)
);

AND2x4_ASAP7_75t_L g1875 ( 
.A(n_1713),
.B(n_1535),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1706),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1760),
.B(n_1655),
.Y(n_1877)
);

BUFx2_ASAP7_75t_L g1878 ( 
.A(n_1765),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_1828),
.Y(n_1879)
);

AOI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1708),
.A2(n_1657),
.B(n_1580),
.Y(n_1880)
);

CKINVDCx20_ASAP7_75t_R g1881 ( 
.A(n_1807),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1714),
.B(n_1672),
.Y(n_1882)
);

AND2x4_ASAP7_75t_L g1883 ( 
.A(n_1713),
.B(n_1569),
.Y(n_1883)
);

OAI21x1_ASAP7_75t_L g1884 ( 
.A1(n_1709),
.A2(n_1616),
.B(n_1629),
.Y(n_1884)
);

O2A1O1Ixp33_ASAP7_75t_L g1885 ( 
.A1(n_1751),
.A2(n_1515),
.B(n_1700),
.C(n_1557),
.Y(n_1885)
);

INVx1_ASAP7_75t_SL g1886 ( 
.A(n_1790),
.Y(n_1886)
);

INVx3_ASAP7_75t_L g1887 ( 
.A(n_1734),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1722),
.Y(n_1888)
);

AOI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1725),
.A2(n_1616),
.B(n_1552),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1724),
.B(n_1750),
.Y(n_1890)
);

AND2x4_ASAP7_75t_L g1891 ( 
.A(n_1727),
.B(n_1681),
.Y(n_1891)
);

INVx2_ASAP7_75t_SL g1892 ( 
.A(n_1817),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1761),
.Y(n_1893)
);

AOI22xp33_ASAP7_75t_L g1894 ( 
.A1(n_1823),
.A2(n_1796),
.B1(n_1825),
.B2(n_1787),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1832),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1794),
.B(n_1696),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1763),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1741),
.B(n_1693),
.Y(n_1898)
);

INVx1_ASAP7_75t_SL g1899 ( 
.A(n_1798),
.Y(n_1899)
);

INVx3_ASAP7_75t_L g1900 ( 
.A(n_1734),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1812),
.B(n_1738),
.Y(n_1901)
);

AOI21xp5_ASAP7_75t_L g1902 ( 
.A1(n_1720),
.A2(n_1552),
.B(n_1544),
.Y(n_1902)
);

AOI22xp33_ASAP7_75t_L g1903 ( 
.A1(n_1831),
.A2(n_1617),
.B1(n_1631),
.B2(n_1629),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1855),
.B(n_1636),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1801),
.Y(n_1905)
);

OAI21xp33_ASAP7_75t_L g1906 ( 
.A1(n_1842),
.A2(n_1636),
.B(n_1584),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1840),
.B(n_1544),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1791),
.Y(n_1908)
);

OR2x6_ASAP7_75t_L g1909 ( 
.A(n_1817),
.B(n_1544),
.Y(n_1909)
);

OAI22xp5_ASAP7_75t_L g1910 ( 
.A1(n_1739),
.A2(n_1646),
.B1(n_1641),
.B2(n_1640),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1800),
.Y(n_1911)
);

CKINVDCx11_ASAP7_75t_R g1912 ( 
.A(n_1769),
.Y(n_1912)
);

NAND2x1p5_ASAP7_75t_L g1913 ( 
.A(n_1754),
.B(n_1552),
.Y(n_1913)
);

NOR4xp25_ASAP7_75t_L g1914 ( 
.A(n_1844),
.B(n_168),
.C(n_169),
.D(n_170),
.Y(n_1914)
);

NOR2xp67_ASAP7_75t_L g1915 ( 
.A(n_1755),
.B(n_1646),
.Y(n_1915)
);

INVx5_ASAP7_75t_L g1916 ( 
.A(n_1754),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1861),
.B(n_1577),
.Y(n_1917)
);

AND2x4_ASAP7_75t_L g1918 ( 
.A(n_1848),
.B(n_1577),
.Y(n_1918)
);

NOR2x1_ASAP7_75t_SL g1919 ( 
.A(n_1754),
.B(n_1577),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1805),
.B(n_1595),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_1707),
.Y(n_1921)
);

O2A1O1Ixp5_ASAP7_75t_SL g1922 ( 
.A1(n_1768),
.A2(n_168),
.B(n_169),
.C(n_170),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1802),
.Y(n_1923)
);

AOI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1719),
.A2(n_1618),
.B(n_1595),
.Y(n_1924)
);

BUFx6f_ASAP7_75t_L g1925 ( 
.A(n_1712),
.Y(n_1925)
);

AND2x4_ASAP7_75t_L g1926 ( 
.A(n_1818),
.B(n_1595),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1804),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1827),
.B(n_1618),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1850),
.B(n_1618),
.Y(n_1929)
);

INVx1_ASAP7_75t_SL g1930 ( 
.A(n_1809),
.Y(n_1930)
);

OAI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1743),
.A2(n_1646),
.B1(n_1641),
.B2(n_1640),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1830),
.Y(n_1932)
);

A2O1A1Ixp33_ASAP7_75t_L g1933 ( 
.A1(n_1726),
.A2(n_1641),
.B(n_1640),
.C(n_1637),
.Y(n_1933)
);

OAI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1860),
.A2(n_1637),
.B1(n_1630),
.B2(n_173),
.Y(n_1934)
);

AND2x4_ASAP7_75t_L g1935 ( 
.A(n_1744),
.B(n_1746),
.Y(n_1935)
);

BUFx2_ASAP7_75t_L g1936 ( 
.A(n_1746),
.Y(n_1936)
);

BUFx3_ASAP7_75t_L g1937 ( 
.A(n_1729),
.Y(n_1937)
);

O2A1O1Ixp33_ASAP7_75t_L g1938 ( 
.A1(n_1810),
.A2(n_171),
.B(n_172),
.C(n_173),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1808),
.B(n_1630),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_SL g1940 ( 
.A(n_1756),
.B(n_369),
.Y(n_1940)
);

BUFx2_ASAP7_75t_L g1941 ( 
.A(n_1767),
.Y(n_1941)
);

BUFx2_ASAP7_75t_L g1942 ( 
.A(n_1767),
.Y(n_1942)
);

OAI22xp5_ASAP7_75t_L g1943 ( 
.A1(n_1777),
.A2(n_171),
.B1(n_172),
.B2(n_174),
.Y(n_1943)
);

INVx3_ASAP7_75t_L g1944 ( 
.A(n_1776),
.Y(n_1944)
);

OR2x2_ASAP7_75t_L g1945 ( 
.A(n_1753),
.B(n_174),
.Y(n_1945)
);

OA21x2_ASAP7_75t_L g1946 ( 
.A1(n_1730),
.A2(n_175),
.B(n_176),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1764),
.B(n_374),
.Y(n_1947)
);

AOI21xp5_ASAP7_75t_L g1948 ( 
.A1(n_1711),
.A2(n_376),
.B(n_375),
.Y(n_1948)
);

OAI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1737),
.A2(n_177),
.B(n_179),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1841),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1786),
.B(n_377),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1836),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1753),
.Y(n_1953)
);

NOR2xp67_ASAP7_75t_L g1954 ( 
.A(n_1811),
.B(n_378),
.Y(n_1954)
);

HB1xp67_ASAP7_75t_L g1955 ( 
.A(n_1821),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1815),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1829),
.B(n_1771),
.Y(n_1957)
);

AND2x4_ASAP7_75t_L g1958 ( 
.A(n_1744),
.B(n_1859),
.Y(n_1958)
);

AOI21xp5_ASAP7_75t_L g1959 ( 
.A1(n_1733),
.A2(n_380),
.B(n_379),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1862),
.B(n_1792),
.Y(n_1960)
);

OAI22xp5_ASAP7_75t_L g1961 ( 
.A1(n_1778),
.A2(n_177),
.B1(n_180),
.B2(n_181),
.Y(n_1961)
);

O2A1O1Ixp33_ASAP7_75t_L g1962 ( 
.A1(n_1837),
.A2(n_180),
.B(n_181),
.C(n_182),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1824),
.B(n_182),
.Y(n_1963)
);

HB1xp67_ASAP7_75t_L g1964 ( 
.A(n_1849),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_SL g1965 ( 
.A(n_1728),
.B(n_381),
.Y(n_1965)
);

OAI22xp5_ASAP7_75t_L g1966 ( 
.A1(n_1894),
.A2(n_1757),
.B1(n_1784),
.B2(n_1783),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1917),
.B(n_1749),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1865),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1866),
.B(n_1839),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1928),
.B(n_1854),
.Y(n_1970)
);

INVx1_ASAP7_75t_SL g1971 ( 
.A(n_1881),
.Y(n_1971)
);

NOR2x1_ASAP7_75t_L g1972 ( 
.A(n_1945),
.B(n_1735),
.Y(n_1972)
);

AOI21xp5_ASAP7_75t_L g1973 ( 
.A1(n_1864),
.A2(n_1716),
.B(n_1813),
.Y(n_1973)
);

AOI21xp5_ASAP7_75t_SL g1974 ( 
.A1(n_1938),
.A2(n_1852),
.B(n_1779),
.Y(n_1974)
);

A2O1A1Ixp33_ASAP7_75t_SL g1975 ( 
.A1(n_1949),
.A2(n_1782),
.B(n_1833),
.C(n_1826),
.Y(n_1975)
);

NOR2x2_ASAP7_75t_L g1976 ( 
.A(n_1909),
.B(n_1835),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1890),
.B(n_1776),
.Y(n_1977)
);

HB1xp67_ASAP7_75t_L g1978 ( 
.A(n_1964),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1871),
.B(n_1775),
.Y(n_1979)
);

AND2x4_ASAP7_75t_L g1980 ( 
.A(n_1958),
.B(n_1932),
.Y(n_1980)
);

AND2x4_ASAP7_75t_L g1981 ( 
.A(n_1958),
.B(n_1735),
.Y(n_1981)
);

A2O1A1Ixp33_ASAP7_75t_L g1982 ( 
.A1(n_1962),
.A2(n_1803),
.B(n_1772),
.C(n_1759),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1957),
.B(n_1834),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1877),
.B(n_1789),
.Y(n_1984)
);

BUFx2_ASAP7_75t_L g1985 ( 
.A(n_1878),
.Y(n_1985)
);

HB1xp67_ASAP7_75t_L g1986 ( 
.A(n_1953),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1901),
.B(n_1731),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1876),
.Y(n_1988)
);

O2A1O1Ixp5_ASAP7_75t_L g1989 ( 
.A1(n_1948),
.A2(n_1799),
.B(n_1822),
.C(n_1785),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1956),
.Y(n_1990)
);

CKINVDCx6p67_ASAP7_75t_R g1991 ( 
.A(n_1912),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1899),
.B(n_1816),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1907),
.B(n_1731),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1950),
.Y(n_1994)
);

INVxp67_ASAP7_75t_L g1995 ( 
.A(n_1955),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1888),
.Y(n_1996)
);

O2A1O1Ixp5_ASAP7_75t_L g1997 ( 
.A1(n_1959),
.A2(n_1880),
.B(n_1943),
.C(n_1924),
.Y(n_1997)
);

BUFx6f_ASAP7_75t_L g1998 ( 
.A(n_1925),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1936),
.B(n_1731),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1882),
.B(n_1774),
.Y(n_2000)
);

BUFx3_ASAP7_75t_L g2001 ( 
.A(n_1874),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1893),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1960),
.B(n_1766),
.Y(n_2003)
);

BUFx3_ASAP7_75t_L g2004 ( 
.A(n_1874),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1891),
.B(n_1766),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1896),
.B(n_1774),
.Y(n_2006)
);

OAI22xp5_ASAP7_75t_L g2007 ( 
.A1(n_1869),
.A2(n_1845),
.B1(n_1843),
.B2(n_1745),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1868),
.B(n_1774),
.Y(n_2008)
);

OA21x2_ASAP7_75t_L g2009 ( 
.A1(n_1905),
.A2(n_1723),
.B(n_1773),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1891),
.B(n_1849),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1872),
.B(n_1819),
.Y(n_2011)
);

INVxp67_ASAP7_75t_SL g2012 ( 
.A(n_1895),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1897),
.Y(n_2013)
);

OAI22xp5_ASAP7_75t_L g2014 ( 
.A1(n_1903),
.A2(n_1847),
.B1(n_1851),
.B2(n_1857),
.Y(n_2014)
);

NOR2xp67_ASAP7_75t_L g2015 ( 
.A(n_1892),
.B(n_1820),
.Y(n_2015)
);

OR2x2_ASAP7_75t_L g2016 ( 
.A(n_1908),
.B(n_1736),
.Y(n_2016)
);

A2O1A1Ixp33_ASAP7_75t_L g2017 ( 
.A1(n_1940),
.A2(n_1858),
.B(n_1740),
.C(n_1793),
.Y(n_2017)
);

OR2x2_ASAP7_75t_L g2018 ( 
.A(n_1911),
.B(n_1856),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1873),
.B(n_1762),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1941),
.B(n_1770),
.Y(n_2020)
);

O2A1O1Ixp33_ASAP7_75t_L g2021 ( 
.A1(n_1961),
.A2(n_1838),
.B(n_1814),
.C(n_1797),
.Y(n_2021)
);

OAI22xp5_ASAP7_75t_L g2022 ( 
.A1(n_1934),
.A2(n_1752),
.B1(n_1838),
.B2(n_1814),
.Y(n_2022)
);

BUFx6f_ASAP7_75t_L g2023 ( 
.A(n_1925),
.Y(n_2023)
);

NOR2xp33_ASAP7_75t_L g2024 ( 
.A(n_1885),
.B(n_1856),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1923),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1986),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_2000),
.B(n_1927),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1986),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1978),
.Y(n_2029)
);

OAI21xp5_ASAP7_75t_L g2030 ( 
.A1(n_1997),
.A2(n_1914),
.B(n_1922),
.Y(n_2030)
);

AO21x2_ASAP7_75t_L g2031 ( 
.A1(n_1973),
.A2(n_1933),
.B(n_1889),
.Y(n_2031)
);

INVx5_ASAP7_75t_L g2032 ( 
.A(n_1981),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1978),
.Y(n_2033)
);

AO21x2_ASAP7_75t_L g2034 ( 
.A1(n_1979),
.A2(n_1884),
.B(n_1902),
.Y(n_2034)
);

BUFx2_ASAP7_75t_L g2035 ( 
.A(n_1980),
.Y(n_2035)
);

OA21x2_ASAP7_75t_L g2036 ( 
.A1(n_1997),
.A2(n_1989),
.B(n_2024),
.Y(n_2036)
);

HB1xp67_ASAP7_75t_L g2037 ( 
.A(n_1972),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1968),
.Y(n_2038)
);

HB1xp67_ASAP7_75t_L g2039 ( 
.A(n_2010),
.Y(n_2039)
);

INVx5_ASAP7_75t_L g2040 ( 
.A(n_1981),
.Y(n_2040)
);

OR2x2_ASAP7_75t_L g2041 ( 
.A(n_1995),
.B(n_2012),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1993),
.B(n_1946),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1996),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1988),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_2002),
.Y(n_2045)
);

INVx1_ASAP7_75t_SL g2046 ( 
.A(n_1980),
.Y(n_2046)
);

INVx3_ASAP7_75t_L g2047 ( 
.A(n_2009),
.Y(n_2047)
);

HB1xp67_ASAP7_75t_L g2048 ( 
.A(n_1985),
.Y(n_2048)
);

INVxp33_ASAP7_75t_L g2049 ( 
.A(n_1970),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1994),
.Y(n_2050)
);

NOR2xp33_ASAP7_75t_L g2051 ( 
.A(n_1971),
.B(n_1886),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1987),
.B(n_1942),
.Y(n_2052)
);

BUFx2_ASAP7_75t_L g2053 ( 
.A(n_1995),
.Y(n_2053)
);

HB1xp67_ASAP7_75t_L g2054 ( 
.A(n_2016),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2013),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_2025),
.Y(n_2056)
);

INVx3_ASAP7_75t_L g2057 ( 
.A(n_2009),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1990),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_2018),
.Y(n_2059)
);

HB1xp67_ASAP7_75t_L g2060 ( 
.A(n_2012),
.Y(n_2060)
);

NAND2x1_ASAP7_75t_L g2061 ( 
.A(n_2053),
.B(n_2024),
.Y(n_2061)
);

AND2x4_ASAP7_75t_L g2062 ( 
.A(n_2032),
.B(n_2020),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2038),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_2039),
.B(n_1999),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_2035),
.B(n_1967),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_2035),
.B(n_1984),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2038),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_2046),
.B(n_2006),
.Y(n_2068)
);

OAI211xp5_ASAP7_75t_SL g2069 ( 
.A1(n_2030),
.A2(n_1963),
.B(n_1992),
.C(n_1969),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_2046),
.B(n_2052),
.Y(n_2070)
);

BUFx2_ASAP7_75t_L g2071 ( 
.A(n_2054),
.Y(n_2071)
);

AOI22xp5_ASAP7_75t_L g2072 ( 
.A1(n_2031),
.A2(n_1966),
.B1(n_2022),
.B2(n_2007),
.Y(n_2072)
);

OR2x2_ASAP7_75t_L g2073 ( 
.A(n_2059),
.B(n_2008),
.Y(n_2073)
);

OAI222xp33_ASAP7_75t_L g2074 ( 
.A1(n_2048),
.A2(n_1983),
.B1(n_2014),
.B2(n_2019),
.C1(n_2003),
.C2(n_2011),
.Y(n_2074)
);

AND2x4_ASAP7_75t_L g2075 ( 
.A(n_2032),
.B(n_2001),
.Y(n_2075)
);

CKINVDCx5p33_ASAP7_75t_R g2076 ( 
.A(n_2051),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2044),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_2052),
.B(n_1977),
.Y(n_2078)
);

OR2x2_ASAP7_75t_L g2079 ( 
.A(n_2059),
.B(n_2009),
.Y(n_2079)
);

INVx3_ASAP7_75t_L g2080 ( 
.A(n_2026),
.Y(n_2080)
);

OAI222xp33_ASAP7_75t_L g2081 ( 
.A1(n_2042),
.A2(n_1947),
.B1(n_2021),
.B2(n_2005),
.C1(n_1867),
.C2(n_1931),
.Y(n_2081)
);

BUFx2_ASAP7_75t_L g2082 ( 
.A(n_2037),
.Y(n_2082)
);

INVx2_ASAP7_75t_L g2083 ( 
.A(n_2080),
.Y(n_2083)
);

OR2x2_ASAP7_75t_L g2084 ( 
.A(n_2071),
.B(n_2059),
.Y(n_2084)
);

HB1xp67_ASAP7_75t_L g2085 ( 
.A(n_2080),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_2080),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_2063),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2067),
.Y(n_2088)
);

HB1xp67_ASAP7_75t_L g2089 ( 
.A(n_2073),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2077),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2073),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2088),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_2083),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_2091),
.B(n_2082),
.Y(n_2094)
);

AND2x4_ASAP7_75t_L g2095 ( 
.A(n_2087),
.B(n_2075),
.Y(n_2095)
);

INVx5_ASAP7_75t_L g2096 ( 
.A(n_2086),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2090),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2092),
.Y(n_2098)
);

OAI22xp5_ASAP7_75t_L g2099 ( 
.A1(n_2094),
.A2(n_2072),
.B1(n_2076),
.B2(n_2061),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_2095),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2097),
.Y(n_2101)
);

AOI22xp5_ASAP7_75t_L g2102 ( 
.A1(n_2094),
.A2(n_2069),
.B1(n_1906),
.B2(n_2036),
.Y(n_2102)
);

BUFx3_ASAP7_75t_L g2103 ( 
.A(n_2095),
.Y(n_2103)
);

INVx2_ASAP7_75t_SL g2104 ( 
.A(n_2096),
.Y(n_2104)
);

INVx2_ASAP7_75t_SL g2105 ( 
.A(n_2096),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2093),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2093),
.Y(n_2107)
);

OR2x2_ASAP7_75t_L g2108 ( 
.A(n_2100),
.B(n_2084),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2098),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2102),
.B(n_2095),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_2103),
.B(n_2066),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2102),
.B(n_2089),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_2101),
.B(n_2089),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_2104),
.B(n_2066),
.Y(n_2114)
);

NOR2xp33_ASAP7_75t_L g2115 ( 
.A(n_2099),
.B(n_1991),
.Y(n_2115)
);

OR2x2_ASAP7_75t_L g2116 ( 
.A(n_2106),
.B(n_2065),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2107),
.Y(n_2117)
);

OR2x2_ASAP7_75t_L g2118 ( 
.A(n_2099),
.B(n_2065),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2117),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_2111),
.B(n_2105),
.Y(n_2120)
);

NAND2x1_ASAP7_75t_L g2121 ( 
.A(n_2114),
.B(n_2075),
.Y(n_2121)
);

HB1xp67_ASAP7_75t_L g2122 ( 
.A(n_2113),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_2108),
.Y(n_2123)
);

CKINVDCx16_ASAP7_75t_R g2124 ( 
.A(n_2115),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2109),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_2113),
.B(n_2085),
.Y(n_2126)
);

INVx1_ASAP7_75t_SL g2127 ( 
.A(n_2120),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2122),
.Y(n_2128)
);

INVx1_ASAP7_75t_SL g2129 ( 
.A(n_2124),
.Y(n_2129)
);

OAI31xp33_ASAP7_75t_L g2130 ( 
.A1(n_2123),
.A2(n_2112),
.A3(n_2110),
.B(n_2118),
.Y(n_2130)
);

INVx3_ASAP7_75t_L g2131 ( 
.A(n_2129),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2128),
.Y(n_2132)
);

INVx1_ASAP7_75t_SL g2133 ( 
.A(n_2127),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2128),
.Y(n_2134)
);

INVxp67_ASAP7_75t_L g2135 ( 
.A(n_2131),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2131),
.B(n_2133),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_2132),
.Y(n_2137)
);

NOR3xp33_ASAP7_75t_L g2138 ( 
.A(n_2134),
.B(n_2125),
.C(n_2119),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_2131),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2136),
.Y(n_2140)
);

OR2x2_ASAP7_75t_L g2141 ( 
.A(n_2139),
.B(n_2130),
.Y(n_2141)
);

CKINVDCx5p33_ASAP7_75t_R g2142 ( 
.A(n_2135),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_2137),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_2138),
.B(n_2121),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2136),
.B(n_2116),
.Y(n_2145)
);

INVxp67_ASAP7_75t_L g2146 ( 
.A(n_2136),
.Y(n_2146)
);

NAND4xp25_ASAP7_75t_L g2147 ( 
.A(n_2136),
.B(n_2126),
.C(n_1870),
.D(n_1937),
.Y(n_2147)
);

HB1xp67_ASAP7_75t_L g2148 ( 
.A(n_2136),
.Y(n_2148)
);

INVx3_ASAP7_75t_L g2149 ( 
.A(n_2139),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_2148),
.B(n_2126),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2145),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_2149),
.B(n_2076),
.Y(n_2152)
);

OAI32xp33_ASAP7_75t_L g2153 ( 
.A1(n_2141),
.A2(n_1863),
.A3(n_2085),
.B1(n_1879),
.B2(n_1921),
.Y(n_2153)
);

OAI22xp5_ASAP7_75t_L g2154 ( 
.A1(n_2146),
.A2(n_2096),
.B1(n_1952),
.B2(n_2075),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_2149),
.Y(n_2155)
);

XOR2x2_ASAP7_75t_L g2156 ( 
.A(n_2140),
.B(n_1930),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_2144),
.B(n_2096),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2142),
.Y(n_2158)
);

OAI21xp5_ASAP7_75t_L g2159 ( 
.A1(n_2143),
.A2(n_2074),
.B(n_1898),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_2147),
.Y(n_2160)
);

XOR2xp5_ASAP7_75t_L g2161 ( 
.A(n_2147),
.B(n_1925),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_SL g2162 ( 
.A(n_2148),
.B(n_1998),
.Y(n_2162)
);

AOI22xp33_ASAP7_75t_L g2163 ( 
.A1(n_2151),
.A2(n_2036),
.B1(n_2030),
.B2(n_2023),
.Y(n_2163)
);

NAND4xp25_ASAP7_75t_L g2164 ( 
.A(n_2152),
.B(n_2158),
.C(n_2157),
.D(n_2153),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2150),
.B(n_2070),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_2155),
.B(n_2070),
.Y(n_2166)
);

AND3x1_ASAP7_75t_L g2167 ( 
.A(n_2160),
.B(n_1951),
.C(n_1976),
.Y(n_2167)
);

NOR2x1_ASAP7_75t_L g2168 ( 
.A(n_2158),
.B(n_1909),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2156),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_2161),
.B(n_2068),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_2162),
.B(n_2154),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_SL g2172 ( 
.A(n_2159),
.B(n_1998),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2150),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2150),
.Y(n_2174)
);

NOR2xp33_ASAP7_75t_L g2175 ( 
.A(n_2151),
.B(n_1998),
.Y(n_2175)
);

AOI21xp5_ASAP7_75t_L g2176 ( 
.A1(n_2171),
.A2(n_1975),
.B(n_1974),
.Y(n_2176)
);

NOR2xp67_ASAP7_75t_L g2177 ( 
.A(n_2173),
.B(n_183),
.Y(n_2177)
);

NAND3xp33_ASAP7_75t_L g2178 ( 
.A(n_2174),
.B(n_2164),
.C(n_2169),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_2167),
.B(n_2078),
.Y(n_2179)
);

NOR3xp33_ASAP7_75t_L g2180 ( 
.A(n_2175),
.B(n_1910),
.C(n_1915),
.Y(n_2180)
);

OR2x2_ASAP7_75t_L g2181 ( 
.A(n_2165),
.B(n_2049),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_SL g2182 ( 
.A(n_2168),
.B(n_1998),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_2166),
.B(n_2036),
.Y(n_2183)
);

NAND5xp2_ASAP7_75t_L g2184 ( 
.A(n_2170),
.B(n_2021),
.C(n_1913),
.D(n_1982),
.E(n_2017),
.Y(n_2184)
);

AOI21xp33_ASAP7_75t_L g2185 ( 
.A1(n_2172),
.A2(n_183),
.B(n_184),
.Y(n_2185)
);

NAND4xp25_ASAP7_75t_L g2186 ( 
.A(n_2163),
.B(n_2015),
.C(n_1954),
.D(n_1975),
.Y(n_2186)
);

NOR2x1_ASAP7_75t_L g2187 ( 
.A(n_2173),
.B(n_184),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2187),
.Y(n_2188)
);

OAI32xp33_ASAP7_75t_L g2189 ( 
.A1(n_2178),
.A2(n_1887),
.A3(n_1900),
.B1(n_2001),
.B2(n_2004),
.Y(n_2189)
);

NOR3xp33_ASAP7_75t_L g2190 ( 
.A(n_2185),
.B(n_2081),
.C(n_1965),
.Y(n_2190)
);

NOR3xp33_ASAP7_75t_L g2191 ( 
.A(n_2177),
.B(n_1900),
.C(n_1887),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_2179),
.B(n_185),
.Y(n_2192)
);

NOR2xp33_ASAP7_75t_L g2193 ( 
.A(n_2181),
.B(n_185),
.Y(n_2193)
);

XOR2x2_ASAP7_75t_L g2194 ( 
.A(n_2182),
.B(n_186),
.Y(n_2194)
);

NOR3xp33_ASAP7_75t_L g2195 ( 
.A(n_2176),
.B(n_1853),
.C(n_1982),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_2183),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2180),
.B(n_186),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_2186),
.Y(n_2198)
);

NOR3xp33_ASAP7_75t_L g2199 ( 
.A(n_2184),
.B(n_187),
.C(n_188),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_2177),
.B(n_187),
.Y(n_2200)
);

OAI21xp33_ASAP7_75t_L g2201 ( 
.A1(n_2178),
.A2(n_2023),
.B(n_2068),
.Y(n_2201)
);

NOR2x1_ASAP7_75t_L g2202 ( 
.A(n_2187),
.B(n_188),
.Y(n_2202)
);

HB1xp67_ASAP7_75t_L g2203 ( 
.A(n_2177),
.Y(n_2203)
);

NAND3xp33_ASAP7_75t_L g2204 ( 
.A(n_2202),
.B(n_1916),
.C(n_189),
.Y(n_2204)
);

NOR2x1_ASAP7_75t_L g2205 ( 
.A(n_2188),
.B(n_189),
.Y(n_2205)
);

INVxp67_ASAP7_75t_L g2206 ( 
.A(n_2203),
.Y(n_2206)
);

NOR2xp67_ASAP7_75t_SL g2207 ( 
.A(n_2200),
.B(n_2023),
.Y(n_2207)
);

NOR2x1_ASAP7_75t_L g2208 ( 
.A(n_2192),
.B(n_190),
.Y(n_2208)
);

NOR3x1_ASAP7_75t_L g2209 ( 
.A(n_2197),
.B(n_190),
.C(n_191),
.Y(n_2209)
);

OAI31xp33_ASAP7_75t_L g2210 ( 
.A1(n_2201),
.A2(n_2062),
.A3(n_193),
.B(n_191),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2191),
.B(n_192),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2193),
.B(n_192),
.Y(n_2212)
);

NAND4xp75_ASAP7_75t_L g2213 ( 
.A(n_2196),
.B(n_196),
.C(n_193),
.D(n_194),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2194),
.Y(n_2214)
);

NOR3xp33_ASAP7_75t_L g2215 ( 
.A(n_2198),
.B(n_196),
.C(n_197),
.Y(n_2215)
);

NAND3xp33_ASAP7_75t_L g2216 ( 
.A(n_2199),
.B(n_1916),
.C(n_197),
.Y(n_2216)
);

INVxp67_ASAP7_75t_SL g2217 ( 
.A(n_2190),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_2189),
.B(n_2078),
.Y(n_2218)
);

NOR2x1_ASAP7_75t_L g2219 ( 
.A(n_2195),
.B(n_198),
.Y(n_2219)
);

NOR2x1_ASAP7_75t_L g2220 ( 
.A(n_2202),
.B(n_198),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2202),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2202),
.Y(n_2222)
);

NOR2xp67_ASAP7_75t_L g2223 ( 
.A(n_2188),
.B(n_200),
.Y(n_2223)
);

OAI211xp5_ASAP7_75t_L g2224 ( 
.A1(n_2202),
.A2(n_1916),
.B(n_202),
.C(n_203),
.Y(n_2224)
);

NAND3x2_ASAP7_75t_L g2225 ( 
.A(n_2188),
.B(n_2053),
.C(n_201),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2203),
.B(n_201),
.Y(n_2226)
);

AND2x4_ASAP7_75t_L g2227 ( 
.A(n_2202),
.B(n_2023),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2202),
.Y(n_2228)
);

NAND2x1p5_ASAP7_75t_L g2229 ( 
.A(n_2202),
.B(n_1874),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2220),
.Y(n_2230)
);

OAI21xp5_ASAP7_75t_L g2231 ( 
.A1(n_2206),
.A2(n_1846),
.B(n_1747),
.Y(n_2231)
);

INVx1_ASAP7_75t_SL g2232 ( 
.A(n_2227),
.Y(n_2232)
);

AND2x2_ASAP7_75t_L g2233 ( 
.A(n_2218),
.B(n_2064),
.Y(n_2233)
);

NOR3xp33_ASAP7_75t_L g2234 ( 
.A(n_2226),
.B(n_202),
.C(n_203),
.Y(n_2234)
);

NAND2xp33_ASAP7_75t_R g2235 ( 
.A(n_2221),
.B(n_204),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2223),
.B(n_204),
.Y(n_2236)
);

NOR3x1_ASAP7_75t_L g2237 ( 
.A(n_2216),
.B(n_205),
.C(n_206),
.Y(n_2237)
);

OR2x2_ASAP7_75t_L g2238 ( 
.A(n_2229),
.B(n_205),
.Y(n_2238)
);

OR2x2_ASAP7_75t_L g2239 ( 
.A(n_2222),
.B(n_206),
.Y(n_2239)
);

NOR2x1_ASAP7_75t_L g2240 ( 
.A(n_2205),
.B(n_207),
.Y(n_2240)
);

OAI21xp33_ASAP7_75t_L g2241 ( 
.A1(n_2217),
.A2(n_2004),
.B(n_1926),
.Y(n_2241)
);

NAND2x1p5_ASAP7_75t_L g2242 ( 
.A(n_2228),
.B(n_2208),
.Y(n_2242)
);

AOI221xp5_ASAP7_75t_L g2243 ( 
.A1(n_2204),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.C(n_210),
.Y(n_2243)
);

HB1xp67_ASAP7_75t_L g2244 ( 
.A(n_2227),
.Y(n_2244)
);

AND2x4_ASAP7_75t_L g2245 ( 
.A(n_2214),
.B(n_1926),
.Y(n_2245)
);

AOI21xp5_ASAP7_75t_L g2246 ( 
.A1(n_2212),
.A2(n_2224),
.B(n_2211),
.Y(n_2246)
);

AND2x4_ASAP7_75t_L g2247 ( 
.A(n_2215),
.B(n_2062),
.Y(n_2247)
);

NOR2x1p5_ASAP7_75t_L g2248 ( 
.A(n_2213),
.B(n_208),
.Y(n_2248)
);

NOR3xp33_ASAP7_75t_L g2249 ( 
.A(n_2219),
.B(n_211),
.C(n_212),
.Y(n_2249)
);

AND2x4_ASAP7_75t_L g2250 ( 
.A(n_2233),
.B(n_2209),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2240),
.Y(n_2251)
);

OR2x6_ASAP7_75t_L g2252 ( 
.A(n_2242),
.B(n_2225),
.Y(n_2252)
);

AOI22xp5_ASAP7_75t_L g2253 ( 
.A1(n_2247),
.A2(n_2241),
.B1(n_2235),
.B2(n_2234),
.Y(n_2253)
);

OR2x2_ASAP7_75t_L g2254 ( 
.A(n_2236),
.B(n_2210),
.Y(n_2254)
);

XNOR2x1_ASAP7_75t_L g2255 ( 
.A(n_2248),
.B(n_2207),
.Y(n_2255)
);

OR2x2_ASAP7_75t_L g2256 ( 
.A(n_2232),
.B(n_212),
.Y(n_2256)
);

INVx1_ASAP7_75t_SL g2257 ( 
.A(n_2239),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2244),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2238),
.Y(n_2259)
);

INVxp33_ASAP7_75t_L g2260 ( 
.A(n_2249),
.Y(n_2260)
);

AOI22xp33_ASAP7_75t_SL g2261 ( 
.A1(n_2230),
.A2(n_1919),
.B1(n_2036),
.B2(n_2062),
.Y(n_2261)
);

AOI22xp5_ASAP7_75t_SL g2262 ( 
.A1(n_2246),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_2262)
);

NAND3x1_ASAP7_75t_L g2263 ( 
.A(n_2243),
.B(n_213),
.C(n_214),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2237),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2245),
.B(n_216),
.Y(n_2265)
);

OAI22x1_ASAP7_75t_SL g2266 ( 
.A1(n_2231),
.A2(n_216),
.B1(n_2040),
.B2(n_2032),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_2244),
.B(n_2034),
.Y(n_2267)
);

XNOR2x2_ASAP7_75t_L g2268 ( 
.A(n_2240),
.B(n_1795),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2240),
.Y(n_2269)
);

OR2x2_ASAP7_75t_L g2270 ( 
.A(n_2242),
.B(n_1939),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2240),
.Y(n_2271)
);

BUFx6f_ASAP7_75t_L g2272 ( 
.A(n_2258),
.Y(n_2272)
);

OAI22x1_ASAP7_75t_L g2273 ( 
.A1(n_2253),
.A2(n_1875),
.B1(n_1883),
.B2(n_1935),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_2256),
.Y(n_2274)
);

NOR3xp33_ASAP7_75t_L g2275 ( 
.A(n_2251),
.B(n_2271),
.C(n_2269),
.Y(n_2275)
);

NAND4xp25_ASAP7_75t_SL g2276 ( 
.A(n_2265),
.B(n_1904),
.C(n_2017),
.D(n_2033),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2262),
.Y(n_2277)
);

AOI221xp5_ASAP7_75t_L g2278 ( 
.A1(n_2260),
.A2(n_2033),
.B1(n_2029),
.B2(n_2028),
.C(n_2044),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2250),
.Y(n_2279)
);

AOI22xp5_ASAP7_75t_L g2280 ( 
.A1(n_2264),
.A2(n_2064),
.B1(n_2029),
.B2(n_2031),
.Y(n_2280)
);

INVx3_ASAP7_75t_L g2281 ( 
.A(n_2252),
.Y(n_2281)
);

AOI21xp33_ASAP7_75t_SL g2282 ( 
.A1(n_2255),
.A2(n_382),
.B(n_384),
.Y(n_2282)
);

AOI22xp5_ASAP7_75t_L g2283 ( 
.A1(n_2257),
.A2(n_2031),
.B1(n_2028),
.B2(n_2034),
.Y(n_2283)
);

AOI31xp33_ASAP7_75t_L g2284 ( 
.A1(n_2259),
.A2(n_1935),
.A3(n_1883),
.B(n_1875),
.Y(n_2284)
);

AOI21xp5_ASAP7_75t_L g2285 ( 
.A1(n_2252),
.A2(n_1929),
.B(n_1920),
.Y(n_2285)
);

NOR2xp67_ASAP7_75t_SL g2286 ( 
.A(n_2254),
.B(n_385),
.Y(n_2286)
);

HB1xp67_ASAP7_75t_L g2287 ( 
.A(n_2263),
.Y(n_2287)
);

OAI21xp33_ASAP7_75t_L g2288 ( 
.A1(n_2270),
.A2(n_2027),
.B(n_2079),
.Y(n_2288)
);

AOI22xp5_ASAP7_75t_L g2289 ( 
.A1(n_2266),
.A2(n_2031),
.B1(n_2034),
.B2(n_1918),
.Y(n_2289)
);

XNOR2xp5_ASAP7_75t_L g2290 ( 
.A(n_2268),
.B(n_387),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2272),
.Y(n_2291)
);

AOI22x1_ASAP7_75t_L g2292 ( 
.A1(n_2287),
.A2(n_2267),
.B1(n_2261),
.B2(n_392),
.Y(n_2292)
);

AOI21xp5_ASAP7_75t_L g2293 ( 
.A1(n_2279),
.A2(n_2034),
.B(n_388),
.Y(n_2293)
);

NAND2x1p5_ASAP7_75t_L g2294 ( 
.A(n_2286),
.B(n_1918),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_2272),
.Y(n_2295)
);

AOI221xp5_ASAP7_75t_L g2296 ( 
.A1(n_2275),
.A2(n_2055),
.B1(n_2056),
.B2(n_2026),
.C(n_2060),
.Y(n_2296)
);

NAND4xp75_ASAP7_75t_L g2297 ( 
.A(n_2277),
.B(n_390),
.C(n_393),
.D(n_396),
.Y(n_2297)
);

NAND4xp25_ASAP7_75t_L g2298 ( 
.A(n_2281),
.B(n_398),
.C(n_403),
.D(n_408),
.Y(n_2298)
);

OAI221xp5_ASAP7_75t_L g2299 ( 
.A1(n_2290),
.A2(n_2274),
.B1(n_2282),
.B2(n_2289),
.C(n_2278),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_2273),
.Y(n_2300)
);

AOI221xp5_ASAP7_75t_L g2301 ( 
.A1(n_2276),
.A2(n_2055),
.B1(n_2056),
.B2(n_2026),
.C(n_2060),
.Y(n_2301)
);

AO22x2_ASAP7_75t_L g2302 ( 
.A1(n_2285),
.A2(n_1795),
.B1(n_2041),
.B2(n_2079),
.Y(n_2302)
);

OAI221xp5_ASAP7_75t_L g2303 ( 
.A1(n_2280),
.A2(n_2041),
.B1(n_2032),
.B2(n_2040),
.C(n_2027),
.Y(n_2303)
);

NAND3xp33_ASAP7_75t_SL g2304 ( 
.A(n_2288),
.B(n_409),
.C(n_411),
.Y(n_2304)
);

OR2x2_ASAP7_75t_L g2305 ( 
.A(n_2284),
.B(n_412),
.Y(n_2305)
);

AOI221xp5_ASAP7_75t_L g2306 ( 
.A1(n_2283),
.A2(n_2047),
.B1(n_2057),
.B2(n_2050),
.C(n_2058),
.Y(n_2306)
);

NOR3xp33_ASAP7_75t_L g2307 ( 
.A(n_2281),
.B(n_413),
.C(n_414),
.Y(n_2307)
);

OAI22xp5_ASAP7_75t_L g2308 ( 
.A1(n_2279),
.A2(n_2032),
.B1(n_2040),
.B2(n_2057),
.Y(n_2308)
);

NAND5xp2_ASAP7_75t_L g2309 ( 
.A(n_2291),
.B(n_415),
.C(n_416),
.D(n_417),
.E(n_420),
.Y(n_2309)
);

NAND4xp25_ASAP7_75t_L g2310 ( 
.A(n_2295),
.B(n_422),
.C(n_423),
.D(n_424),
.Y(n_2310)
);

NOR3xp33_ASAP7_75t_L g2311 ( 
.A(n_2299),
.B(n_2300),
.C(n_2305),
.Y(n_2311)
);

NAND4xp25_ASAP7_75t_SL g2312 ( 
.A(n_2293),
.B(n_1795),
.C(n_2042),
.D(n_427),
.Y(n_2312)
);

OR5x1_ASAP7_75t_L g2313 ( 
.A(n_2304),
.B(n_425),
.C(n_426),
.D(n_428),
.E(n_430),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2294),
.B(n_431),
.Y(n_2314)
);

NAND4xp75_ASAP7_75t_L g2315 ( 
.A(n_2292),
.B(n_432),
.C(n_433),
.D(n_435),
.Y(n_2315)
);

NAND3xp33_ASAP7_75t_SL g2316 ( 
.A(n_2307),
.B(n_436),
.C(n_438),
.Y(n_2316)
);

OR2x2_ASAP7_75t_L g2317 ( 
.A(n_2298),
.B(n_439),
.Y(n_2317)
);

OAI211xp5_ASAP7_75t_L g2318 ( 
.A1(n_2301),
.A2(n_440),
.B(n_441),
.C(n_442),
.Y(n_2318)
);

AOI221xp5_ASAP7_75t_L g2319 ( 
.A1(n_2303),
.A2(n_2057),
.B1(n_2047),
.B2(n_449),
.C(n_450),
.Y(n_2319)
);

AO22x2_ASAP7_75t_L g2320 ( 
.A1(n_2315),
.A2(n_2297),
.B1(n_2308),
.B2(n_2306),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2317),
.Y(n_2321)
);

HB1xp67_ASAP7_75t_L g2322 ( 
.A(n_2313),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2314),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2311),
.B(n_2296),
.Y(n_2324)
);

CKINVDCx20_ASAP7_75t_R g2325 ( 
.A(n_2316),
.Y(n_2325)
);

OAI22xp5_ASAP7_75t_SL g2326 ( 
.A1(n_2309),
.A2(n_2302),
.B1(n_1944),
.B2(n_2032),
.Y(n_2326)
);

OAI221xp5_ASAP7_75t_L g2327 ( 
.A1(n_2319),
.A2(n_2318),
.B1(n_2310),
.B2(n_2312),
.C(n_2302),
.Y(n_2327)
);

AOI22xp5_ASAP7_75t_L g2328 ( 
.A1(n_2311),
.A2(n_2032),
.B1(n_2040),
.B2(n_2057),
.Y(n_2328)
);

AOI22xp5_ASAP7_75t_L g2329 ( 
.A1(n_2311),
.A2(n_2040),
.B1(n_2047),
.B2(n_1944),
.Y(n_2329)
);

AOI22xp33_ASAP7_75t_L g2330 ( 
.A1(n_2311),
.A2(n_2058),
.B1(n_2045),
.B2(n_2050),
.Y(n_2330)
);

OAI211xp5_ASAP7_75t_L g2331 ( 
.A1(n_2311),
.A2(n_443),
.B(n_444),
.C(n_451),
.Y(n_2331)
);

NOR2x1_ASAP7_75t_L g2332 ( 
.A(n_2315),
.B(n_454),
.Y(n_2332)
);

NOR2x1_ASAP7_75t_L g2333 ( 
.A(n_2332),
.B(n_455),
.Y(n_2333)
);

XOR2xp5_ASAP7_75t_L g2334 ( 
.A(n_2325),
.B(n_456),
.Y(n_2334)
);

NAND5xp2_ASAP7_75t_L g2335 ( 
.A(n_2327),
.B(n_457),
.C(n_458),
.D(n_459),
.E(n_461),
.Y(n_2335)
);

OAI222xp33_ASAP7_75t_L g2336 ( 
.A1(n_2324),
.A2(n_2040),
.B1(n_2047),
.B2(n_2050),
.C1(n_2045),
.C2(n_2043),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_2320),
.Y(n_2337)
);

XOR2xp5_ASAP7_75t_L g2338 ( 
.A(n_2322),
.B(n_463),
.Y(n_2338)
);

INVxp67_ASAP7_75t_L g2339 ( 
.A(n_2323),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2326),
.Y(n_2340)
);

OAI22x1_ASAP7_75t_L g2341 ( 
.A1(n_2338),
.A2(n_2321),
.B1(n_2329),
.B2(n_2331),
.Y(n_2341)
);

NAND2xp33_ASAP7_75t_SL g2342 ( 
.A(n_2337),
.B(n_2330),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2333),
.Y(n_2343)
);

AOI22xp5_ASAP7_75t_L g2344 ( 
.A1(n_2342),
.A2(n_2339),
.B1(n_2340),
.B2(n_2334),
.Y(n_2344)
);

AOI21xp5_ASAP7_75t_L g2345 ( 
.A1(n_2343),
.A2(n_2335),
.B(n_2328),
.Y(n_2345)
);

AOI22x1_ASAP7_75t_L g2346 ( 
.A1(n_2345),
.A2(n_2341),
.B1(n_2336),
.B2(n_466),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_2346),
.Y(n_2347)
);

XNOR2xp5_ASAP7_75t_L g2348 ( 
.A(n_2346),
.B(n_2344),
.Y(n_2348)
);

AO21x2_ASAP7_75t_L g2349 ( 
.A1(n_2348),
.A2(n_2347),
.B(n_465),
.Y(n_2349)
);

OR2x2_ASAP7_75t_L g2350 ( 
.A(n_2347),
.B(n_464),
.Y(n_2350)
);

AOI221x1_ASAP7_75t_L g2351 ( 
.A1(n_2349),
.A2(n_467),
.B1(n_469),
.B2(n_470),
.C(n_471),
.Y(n_2351)
);

AOI211xp5_ASAP7_75t_L g2352 ( 
.A1(n_2351),
.A2(n_2350),
.B(n_474),
.C(n_477),
.Y(n_2352)
);


endmodule