module real_jpeg_20007_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_213;
wire n_202;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_0),
.A2(n_53),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_0),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_0),
.A2(n_56),
.B1(n_57),
.B2(n_61),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_0),
.A2(n_29),
.B1(n_31),
.B2(n_61),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_0),
.A2(n_39),
.B1(n_40),
.B2(n_61),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_1),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_1),
.B(n_55),
.Y(n_149)
);

AOI21xp33_ASAP7_75t_L g169 ( 
.A1(n_1),
.A2(n_16),
.B(n_29),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_1),
.A2(n_39),
.B1(n_40),
.B2(n_107),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_177),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_1),
.B(n_76),
.Y(n_190)
);

AOI21xp33_ASAP7_75t_L g207 ( 
.A1(n_1),
.A2(n_57),
.B(n_208),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_2),
.A2(n_53),
.B1(n_60),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_2),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_2),
.A2(n_56),
.B1(n_57),
.B2(n_64),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_2),
.A2(n_39),
.B1(n_40),
.B2(n_64),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_2),
.A2(n_29),
.B1(n_31),
.B2(n_64),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_3),
.A2(n_39),
.B1(n_40),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_3),
.A2(n_44),
.B1(n_56),
.B2(n_57),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_3),
.A2(n_29),
.B1(n_31),
.B2(n_44),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_4),
.A2(n_53),
.B1(n_60),
.B2(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_4),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_4),
.A2(n_56),
.B1(n_57),
.B2(n_120),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_4),
.A2(n_39),
.B1(n_40),
.B2(n_120),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_4),
.A2(n_29),
.B1(n_31),
.B2(n_120),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_5),
.A2(n_53),
.B1(n_60),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_5),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_5),
.A2(n_56),
.B1(n_57),
.B2(n_96),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_5),
.A2(n_29),
.B1(n_31),
.B2(n_96),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_5),
.A2(n_39),
.B1(n_40),
.B2(n_96),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_6),
.A2(n_39),
.B1(n_40),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_6),
.A2(n_29),
.B1(n_31),
.B2(n_46),
.Y(n_87)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_8),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_8),
.A2(n_32),
.B1(n_39),
.B2(n_40),
.Y(n_82)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_10),
.A2(n_29),
.B1(n_31),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_13),
.A2(n_56),
.B1(n_57),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_13),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_13),
.A2(n_39),
.B1(n_40),
.B2(n_69),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_13),
.A2(n_29),
.B1(n_31),
.B2(n_69),
.Y(n_152)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_14),
.A2(n_39),
.B1(n_40),
.B2(n_72),
.Y(n_74)
);

OAI32xp33_ASAP7_75t_L g202 ( 
.A1(n_14),
.A2(n_40),
.A3(n_57),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_16),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_16),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_16),
.A2(n_29),
.B1(n_31),
.B2(n_41),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_123),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_121),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_97),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_21),
.B(n_97),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_84),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_77),
.B2(n_78),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_47),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_36),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_26),
.B(n_36),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_27),
.A2(n_28),
.B(n_34),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_27),
.A2(n_87),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_27),
.A2(n_28),
.B1(n_110),
.B2(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_27),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_27),
.A2(n_111),
.B1(n_163),
.B2(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_27),
.A2(n_28),
.B1(n_165),
.B2(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_27),
.A2(n_28),
.B1(n_152),
.B2(n_195),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_28),
.B(n_107),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_29),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_31),
.B(n_181),
.Y(n_180)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_33),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_37),
.A2(n_42),
.B1(n_45),
.B2(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_37),
.A2(n_42),
.B1(n_43),
.B2(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_37),
.A2(n_42),
.B1(n_89),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_37),
.A2(n_42),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_37),
.A2(n_42),
.B1(n_173),
.B2(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_37),
.A2(n_42),
.B1(n_193),
.B2(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_37),
.A2(n_42),
.B1(n_131),
.B2(n_211),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_42),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_39),
.B(n_72),
.Y(n_203)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_40),
.A2(n_41),
.B(n_107),
.C(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_42),
.B(n_107),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_65),
.B2(n_66),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_59),
.B1(n_62),
.B2(n_63),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_50),
.A2(n_59),
.B1(n_62),
.B2(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_50),
.A2(n_62),
.B1(n_95),
.B2(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_51),
.A2(n_55),
.B1(n_106),
.B2(n_119),
.Y(n_135)
);

O2A1O1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B(n_54),
.C(n_55),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_53),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_52),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_52),
.B(n_57),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_53),
.Y(n_60)
);

HAxp5_ASAP7_75t_SL g106 ( 
.A(n_53),
.B(n_107),
.CON(n_106),
.SN(n_106)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_54),
.A2(n_56),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_72),
.B(n_73),
.C(n_74),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_72),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_56),
.B(n_107),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_71),
.B1(n_74),
.B2(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_70),
.A2(n_76),
.B1(n_146),
.B2(n_148),
.Y(n_145)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_71),
.A2(n_74),
.B1(n_92),
.B2(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_71),
.A2(n_74),
.B1(n_115),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_71),
.A2(n_74),
.B1(n_147),
.B2(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_81),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_90),
.C(n_93),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_86),
.B(n_88),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.C(n_102),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_98),
.A2(n_100),
.B1(n_101),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_98),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_102),
.A2(n_103),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_113),
.C(n_116),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_104),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_109),
.Y(n_142)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_112),
.A2(n_161),
.B1(n_162),
.B2(n_164),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_113),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_153),
.B(n_236),
.C(n_242),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_138),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_125),
.B(n_138),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_136),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_127),
.B(n_128),
.C(n_136),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_132),
.C(n_135),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_129),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_135),
.B(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.C(n_143),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_139),
.B(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.C(n_150),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_145),
.B(n_221),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_149),
.A2(n_150),
.B1(n_151),
.B2(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_149),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_235),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_230),
.B(n_234),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_216),
.B(n_229),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_197),
.B(n_215),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_185),
.B(n_196),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_174),
.B(n_184),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_166),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_166),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_170),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_179),
.B(n_183),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_178),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_187),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_194),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_192),
.C(n_194),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_199),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_205),
.B1(n_213),
.B2(n_214),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_200),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_202),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_204),
.Y(n_208)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_209),
.B1(n_210),
.B2(n_212),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_206),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_212),
.C(n_213),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_217),
.B(n_218),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_223),
.B2(n_224),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_226),
.C(n_227),
.Y(n_231)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_225),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_226),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_231),
.B(n_232),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_237),
.B(n_238),
.Y(n_242)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);


endmodule