module real_jpeg_4154_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g80 ( 
.A(n_0),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_1),
.A2(n_83),
.B1(n_86),
.B2(n_88),
.Y(n_82)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_1),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_1),
.A2(n_29),
.B1(n_88),
.B2(n_218),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_1),
.A2(n_88),
.B1(n_267),
.B2(n_269),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_1),
.A2(n_88),
.B1(n_248),
.B2(n_253),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_2),
.A2(n_158),
.B1(n_162),
.B2(n_163),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_2),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_2),
.A2(n_110),
.B1(n_163),
.B2(n_200),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_3),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_3),
.Y(n_105)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_3),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_4),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_4),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_4),
.A2(n_92),
.B1(n_248),
.B2(n_253),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_4),
.A2(n_92),
.B1(n_307),
.B2(n_309),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_5),
.A2(n_169),
.B1(n_173),
.B2(n_174),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_5),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_6),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_6),
.Y(n_205)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_8),
.A2(n_44),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_8),
.A2(n_51),
.B1(n_110),
.B2(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_8),
.A2(n_51),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_8),
.A2(n_51),
.B1(n_258),
.B2(n_262),
.Y(n_257)
);

BUFx5_ASAP7_75t_L g152 ( 
.A(n_9),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_9),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_9),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_9),
.Y(n_208)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_9),
.Y(n_280)
);

INVx8_ASAP7_75t_L g295 ( 
.A(n_9),
.Y(n_295)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_10),
.Y(n_147)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_12),
.A2(n_46),
.B1(n_121),
.B2(n_235),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_12),
.B(n_243),
.C(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_12),
.B(n_73),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_12),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_12),
.B(n_97),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_12),
.B(n_322),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_13),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_14),
.Y(n_101)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_14),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_15),
.A2(n_110),
.B1(n_113),
.B2(n_116),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_15),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_15),
.A2(n_116),
.B1(n_186),
.B2(n_188),
.Y(n_185)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_226),
.B1(n_227),
.B2(n_360),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_18),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_225),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_193),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_20),
.B(n_193),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_135),
.C(n_176),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_21),
.B(n_357),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_56),
.B2(n_134),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_22),
.B(n_57),
.C(n_95),
.Y(n_209)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_43),
.B(n_48),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_24),
.B(n_50),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_33),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_30),
.Y(n_218)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_33),
.B(n_46),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_38),
.B2(n_40),
.Y(n_33)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_36),
.Y(n_331)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_39),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_39),
.Y(n_181)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI32xp33_ASAP7_75t_L g138 ( 
.A1(n_41),
.A2(n_47),
.A3(n_139),
.B1(n_143),
.B2(n_145),
.Y(n_138)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_46),
.B(n_47),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_46),
.Y(n_47)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_46),
.A2(n_150),
.B(n_256),
.Y(n_281)
);

OAI21xp33_ASAP7_75t_SL g316 ( 
.A1(n_46),
.A2(n_317),
.B(n_320),
.Y(n_316)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_55),
.Y(n_49)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_55),
.Y(n_219)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_56),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_95),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_82),
.B1(n_89),
.B2(n_90),
.Y(n_57)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_58),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_73),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B1(n_67),
.B2(n_72),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_61),
.Y(n_336)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_62),
.Y(n_341)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_66),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_66),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

AO22x2_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_81),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_77),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_79),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_79),
.Y(n_308)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_80),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_81),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_82),
.A2(n_89),
.B(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_85),
.Y(n_319)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_89),
.B(n_180),
.Y(n_224)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_90),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_146),
.Y(n_145)
);

INVx6_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_109),
.B(n_117),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_96),
.A2(n_109),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_96),
.A2(n_197),
.B1(n_266),
.B2(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_97),
.B(n_118),
.Y(n_237)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_98),
.A2(n_117),
.B(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_102),
.B1(n_104),
.B2(n_106),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_100),
.Y(n_243)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_103),
.Y(n_188)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_103),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g244 ( 
.A(n_103),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_104),
.Y(n_162)
);

BUFx8_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_105),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g187 ( 
.A(n_105),
.Y(n_187)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_115),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_122),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_127),
.B1(n_129),
.B2(n_132),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_126),
.Y(n_241)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_126),
.Y(n_268)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_133),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_135),
.A2(n_136),
.B1(n_176),
.B2(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_148),
.B2(n_149),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_138),
.B(n_148),
.Y(n_213)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_156),
.B1(n_164),
.B2(n_167),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_150),
.A2(n_247),
.B(n_256),
.Y(n_246)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_151),
.A2(n_157),
.B1(n_185),
.B2(n_189),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_151),
.A2(n_168),
.B1(n_202),
.B2(n_207),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_151),
.B(n_257),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_151),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_161),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_161),
.Y(n_255)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_165),
.B(n_257),
.Y(n_256)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_176),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_184),
.C(n_192),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_177),
.B(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_183),
.A2(n_223),
.B(n_224),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_183),
.A2(n_224),
.B(n_316),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_184),
.B(n_192),
.Y(n_351)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_185),
.Y(n_326)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_191),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_212),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_194)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_201),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_197),
.A2(n_234),
.B(n_237),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_197),
.A2(n_237),
.B(n_306),
.Y(n_348)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_209),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_221),
.B2(n_222),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_219),
.B(n_220),
.Y(n_216)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

AOI21x1_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_354),
.B(n_359),
.Y(n_227)
);

AO21x1_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_343),
.B(n_353),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_300),
.B(n_342),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_273),
.B(n_299),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_245),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_232),
.B(n_245),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_238),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_233),
.A2(n_238),
.B1(n_239),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_233),
.Y(n_297)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_263),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_246),
.B(n_264),
.C(n_272),
.Y(n_301)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_247),
.Y(n_292)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_253),
.Y(n_277)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx8_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_255),
.Y(n_262)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_271),
.B2(n_272),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_267),
.Y(n_338)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_289),
.B(n_298),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_282),
.B(n_288),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_281),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_280),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_287),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_287),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B(n_286),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_284),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_286),
.A2(n_326),
.B(n_327),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_296),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_296),
.Y(n_298)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_301),
.B(n_302),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_324),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_314),
.B2(n_315),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_305),
.B(n_314),
.C(n_324),
.Y(n_344)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx5_ASAP7_75t_SL g310 ( 
.A(n_311),
.Y(n_310)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVxp33_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

AOI32xp33_ASAP7_75t_L g329 ( 
.A1(n_321),
.A2(n_330),
.A3(n_332),
.B1(n_334),
.B2(n_337),
.Y(n_329)
);

INVx6_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_329),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_325),
.B(n_329),
.Y(n_349)
);

INVx3_ASAP7_75t_SL g327 ( 
.A(n_328),
.Y(n_327)
);

INVx8_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

NAND2xp33_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_344),
.B(n_345),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_347),
.B1(n_350),
.B2(n_352),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_348),
.B(n_349),
.C(n_352),
.Y(n_355)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_350),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_355),
.B(n_356),
.Y(n_359)
);


endmodule