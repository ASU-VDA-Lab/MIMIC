module fake_jpeg_13267_n_265 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_225;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_207;
wire n_155;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx11_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

HAxp5_ASAP7_75t_SL g36 ( 
.A(n_17),
.B(n_0),
.CON(n_36),
.SN(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_36),
.A2(n_40),
.B(n_38),
.C(n_42),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_27),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_35),
.Y(n_39)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_0),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_41),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_42),
.A2(n_34),
.B1(n_22),
.B2(n_31),
.Y(n_68)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_46),
.B(n_30),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_20),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_47),
.B(n_58),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_30),
.B1(n_19),
.B2(n_24),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_59),
.B1(n_39),
.B2(n_35),
.Y(n_82)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_51),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_27),
.B1(n_21),
.B2(n_25),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_55),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_23),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_19),
.B1(n_24),
.B2(n_22),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_67),
.Y(n_79)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_32),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_46),
.Y(n_97)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g91 ( 
.A1(n_66),
.A2(n_41),
.B(n_37),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_25),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_35),
.Y(n_98)
);

NOR2x1_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_31),
.Y(n_75)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_73),
.B(n_79),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_75),
.A2(n_89),
.B1(n_46),
.B2(n_52),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_36),
.B(n_42),
.C(n_44),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_88),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_82),
.A2(n_94),
.B1(n_65),
.B2(n_56),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_44),
.C(n_39),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_97),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_55),
.B(n_41),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

HAxp5_ASAP7_75t_SL g103 ( 
.A(n_91),
.B(n_52),
.CON(n_103),
.SN(n_103)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_68),
.A2(n_37),
.B1(n_28),
.B2(n_20),
.Y(n_94)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_95),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_53),
.B(n_35),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_96),
.A2(n_46),
.B1(n_49),
.B2(n_69),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_101),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_54),
.B(n_32),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_100),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_54),
.B(n_29),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_53),
.B(n_29),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_62),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_102),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_103),
.A2(n_116),
.B(n_119),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_106),
.A2(n_122),
.B1(n_85),
.B2(n_78),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_76),
.A2(n_71),
.B1(n_70),
.B2(n_45),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_111),
.B1(n_112),
.B2(n_88),
.Y(n_139)
);

AND2x6_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_54),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_108),
.B(n_103),
.Y(n_154)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_75),
.A2(n_34),
.B1(n_45),
.B2(n_28),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_87),
.A2(n_45),
.B1(n_54),
.B2(n_56),
.Y(n_112)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

AOI32xp33_ASAP7_75t_L g119 ( 
.A1(n_98),
.A2(n_23),
.A3(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_88),
.A2(n_33),
.B1(n_2),
.B2(n_5),
.Y(n_122)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_127),
.Y(n_133)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_110),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_130),
.B(n_135),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_73),
.C(n_84),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_132),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_73),
.C(n_96),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_113),
.B(n_101),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_138),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_117),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_136),
.A2(n_153),
.B1(n_6),
.B2(n_8),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_92),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_137),
.B(n_149),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_102),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_139),
.A2(n_146),
.B1(n_122),
.B2(n_116),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_117),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_141),
.A2(n_145),
.B(n_1),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_118),
.A2(n_84),
.B(n_96),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_115),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_107),
.A2(n_80),
.B1(n_78),
.B2(n_77),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_80),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_151),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_85),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_85),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_104),
.B(n_77),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_152),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_106),
.A2(n_83),
.B1(n_86),
.B2(n_74),
.Y(n_153)
);

AOI322xp5_ASAP7_75t_L g166 ( 
.A1(n_154),
.A2(n_112),
.A3(n_95),
.B1(n_128),
.B2(n_127),
.C1(n_126),
.C2(n_124),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_109),
.B(n_86),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_156),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_157),
.A2(n_167),
.B1(n_169),
.B2(n_132),
.Y(n_201)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_139),
.A2(n_108),
.B1(n_125),
.B2(n_128),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_172),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_179),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_133),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_165),
.B(n_166),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_150),
.A2(n_120),
.B1(n_105),
.B2(n_74),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_138),
.A2(n_120),
.B1(n_105),
.B2(n_7),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_171),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_154),
.A2(n_33),
.B1(n_8),
.B2(n_9),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_133),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_178),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_136),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_143),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_130),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_176),
.A2(n_140),
.B(n_149),
.Y(n_183)
);

AOI21xp33_ASAP7_75t_L g219 ( 
.A1(n_183),
.A2(n_185),
.B(n_178),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_176),
.A2(n_140),
.B(n_147),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_153),
.Y(n_188)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_141),
.Y(n_191)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_180),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_192),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_137),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_196),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_197),
.A2(n_201),
.B1(n_175),
.B2(n_184),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_131),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_131),
.C(n_181),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_146),
.Y(n_200)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_200),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_168),
.B(n_181),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_134),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_212),
.C(n_214),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_194),
.A2(n_163),
.B1(n_174),
.B2(n_182),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_207),
.A2(n_215),
.B1(n_197),
.B2(n_199),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_183),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_213),
.B1(n_218),
.B2(n_189),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_151),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_201),
.A2(n_182),
.B1(n_177),
.B2(n_135),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_185),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_194),
.A2(n_177),
.B1(n_172),
.B2(n_161),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_162),
.Y(n_216)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_216),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_188),
.A2(n_159),
.B1(n_158),
.B2(n_164),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_219),
.A2(n_189),
.B1(n_187),
.B2(n_184),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_190),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_220),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_222),
.B(n_208),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_225),
.A2(n_228),
.B1(n_233),
.B2(n_207),
.Y(n_235)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_216),
.Y(n_226)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_226),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_195),
.C(n_188),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_229),
.C(n_211),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_200),
.C(n_202),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_231),
.Y(n_239)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_218),
.A2(n_187),
.B1(n_202),
.B2(n_193),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_232),
.A2(n_205),
.B1(n_211),
.B2(n_199),
.Y(n_241)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_242),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_214),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_238),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_225),
.A2(n_217),
.B1(n_215),
.B2(n_206),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_241),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_227),
.A2(n_220),
.B(n_205),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_240),
.A2(n_223),
.B(n_221),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_193),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_224),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_248),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_247),
.A2(n_249),
.B(n_222),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_232),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_242),
.A2(n_243),
.B(n_236),
.Y(n_249)
);

OAI221xp5_ASAP7_75t_L g256 ( 
.A1(n_251),
.A2(n_250),
.B1(n_156),
.B2(n_144),
.C(n_155),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_245),
.A2(n_234),
.B1(n_241),
.B2(n_186),
.Y(n_253)
);

INVxp33_ASAP7_75t_L g259 ( 
.A(n_253),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_186),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_255),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_238),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_258),
.C(n_253),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_252),
.A2(n_144),
.B(n_155),
.Y(n_258)
);

AOI322xp5_ASAP7_75t_L g262 ( 
.A1(n_260),
.A2(n_261),
.A3(n_259),
.B1(n_12),
.B2(n_15),
.C1(n_16),
.C2(n_10),
.Y(n_262)
);

AOI322xp5_ASAP7_75t_L g261 ( 
.A1(n_257),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_14),
.C2(n_15),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_262),
.B(n_12),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_263),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_16),
.Y(n_265)
);


endmodule