module real_jpeg_18915_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_6),
.B1(n_15),
.B2(n_17),
.Y(n_14)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_1),
.Y(n_76)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_1),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_2),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_3),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_3),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_3),
.B(n_51),
.Y(n_50)
);

AND2x4_ASAP7_75t_L g71 ( 
.A(n_3),
.B(n_72),
.Y(n_71)
);

NAND2x1_ASAP7_75t_L g89 ( 
.A(n_3),
.B(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_3),
.B(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_3),
.B(n_140),
.Y(n_139)
);

NAND2x1_ASAP7_75t_L g188 ( 
.A(n_3),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_4),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_4),
.B(n_229),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_4),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_4),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_4),
.B(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_5),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_5),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_5),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_5),
.B(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_5),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_5),
.B(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_9),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_9),
.Y(n_180)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_9),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_10),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_10),
.B(n_41),
.Y(n_40)
);

AND2x4_ASAP7_75t_L g55 ( 
.A(n_10),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_10),
.B(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_10),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_10),
.B(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g177 ( 
.A(n_10),
.B(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g225 ( 
.A(n_10),
.B(n_189),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_11),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g131 ( 
.A(n_12),
.Y(n_131)
);

BUFx8_ASAP7_75t_L g189 ( 
.A(n_13),
.Y(n_189)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_13),
.Y(n_247)
);

BUFx12f_ASAP7_75t_SL g15 ( 
.A(n_16),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_308),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_275),
.B(n_305),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_236),
.B(n_269),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_202),
.Y(n_21)
);

OAI21x1_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_165),
.B(n_201),
.Y(n_22)
);

AOI21x1_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_117),
.B(n_164),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_78),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_25),
.B(n_78),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_48),
.C(n_64),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_26),
.B(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_39),
.Y(n_26)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_27),
.Y(n_155)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_28),
.A2(n_40),
.B(n_47),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_34),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_29),
.A2(n_30),
.B1(n_113),
.B2(n_116),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_29),
.A2(n_30),
.B1(n_97),
.B2(n_98),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_29),
.B(n_43),
.C(n_89),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_43),
.B(n_45),
.Y(n_42)
);

NAND2x1p5_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_43),
.Y(n_45)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_33),
.Y(n_144)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_33),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_34),
.A2(n_142),
.B1(n_145),
.B2(n_146),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_34),
.Y(n_146)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_38),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_42),
.B1(n_46),
.B2(n_47),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

O2A1O1Ixp33_ASAP7_75t_R g138 ( 
.A1(n_40),
.A2(n_139),
.B(n_141),
.C(n_147),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_40),
.B(n_139),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_40),
.A2(n_46),
.B1(n_139),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_42),
.A2(n_47),
.B1(n_88),
.B2(n_89),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_43),
.A2(n_128),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_43),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_43),
.B(n_142),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_43),
.A2(n_134),
.B1(n_142),
.B2(n_145),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_43),
.A2(n_142),
.B(n_244),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_45),
.B(n_83),
.C(n_89),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_48),
.A2(n_64),
.B1(n_65),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_48),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_54),
.C(n_59),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_49),
.A2(n_50),
.B1(n_59),
.B2(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_49),
.A2(n_50),
.B1(n_177),
.B2(n_181),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_50),
.B(n_214),
.Y(n_213)
);

AO21x1_ASAP7_75t_L g250 ( 
.A1(n_50),
.A2(n_251),
.B(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_50),
.B(n_66),
.C(n_177),
.Y(n_286)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_54),
.A2(n_55),
.B1(n_96),
.B2(n_106),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_54),
.A2(n_55),
.B1(n_124),
.B2(n_126),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_55),
.A2(n_98),
.B(n_100),
.C(n_147),
.Y(n_172)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_58),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_58),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_59),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_59),
.A2(n_83),
.B1(n_91),
.B2(n_125),
.Y(n_210)
);

XNOR2x2_ASAP7_75t_L g295 ( 
.A(n_59),
.B(n_296),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_60),
.B(n_114),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_60),
.B(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_69),
.B1(n_70),
.B2(n_77),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_66),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_66),
.B(n_71),
.C(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_66),
.A2(n_77),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_71),
.A2(n_260),
.B1(n_261),
.B2(n_263),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_71),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_71),
.B(n_261),
.C(n_264),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_71),
.B(n_224),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_71),
.A2(n_187),
.B1(n_188),
.B2(n_260),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_73),
.Y(n_198)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_74),
.A2(n_110),
.B1(n_176),
.B2(n_182),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_77),
.B(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_94),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_92),
.B2(n_93),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_81),
.B(n_92),
.C(n_94),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_88),
.B1(n_89),
.B2(n_91),
.Y(n_82)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_88),
.A2(n_89),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_91),
.B(n_125),
.C(n_209),
.Y(n_257)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_107),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_95),
.B(n_108),
.C(n_112),
.Y(n_169)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_100),
.B2(n_105),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_97),
.B(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_97),
.B(n_154),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_97),
.B(n_139),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

MAJx2_ASAP7_75t_L g209 ( 
.A(n_98),
.B(n_139),
.C(n_188),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_99),
.Y(n_262)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

AO22x1_ASAP7_75t_L g296 ( 
.A1(n_100),
.A2(n_105),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_100),
.B(n_125),
.C(n_297),
.Y(n_331)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_104),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_110),
.B(n_142),
.C(n_177),
.Y(n_233)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_113),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_113),
.A2(n_116),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_113),
.B(n_225),
.C(n_228),
.Y(n_264)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_115),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_116),
.B(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_116),
.A2(n_127),
.B(n_128),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_136),
.B(n_163),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_122),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.C(n_132),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_124),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_127),
.A2(n_132),
.B1(n_133),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_151),
.B(n_162),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_148),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_148),
.Y(n_162)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_139),
.A2(n_160),
.B1(n_213),
.B2(n_218),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_139),
.B(n_215),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_142),
.A2(n_145),
.B1(n_177),
.B2(n_181),
.Y(n_176)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_158),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_157),
.B(n_161),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_155),
.B(n_156),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_160),
.B(n_214),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_167),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_183),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_170),
.C(n_183),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_173),
.B(n_175),
.C(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_174),
.B(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_176),
.Y(n_182)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_200),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_191),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_185),
.B(n_191),
.C(n_200),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_190),
.Y(n_185)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_186),
.Y(n_190)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_196),
.B(n_199),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_196),
.Y(n_199)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx4_ASAP7_75t_SL g194 ( 
.A(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_196),
.A2(n_318),
.B1(n_319),
.B2(n_320),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_196),
.Y(n_318)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_199),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_199),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_203),
.B(n_204),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_221),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_205),
.B(n_222),
.C(n_235),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_219),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_211),
.B2(n_212),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_211),
.C(n_219),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_213),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_235),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_231),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_223),
.B(n_233),
.C(n_234),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_224),
.B(n_260),
.C(n_285),
.Y(n_338)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_236),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_268),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_268),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_238),
.B(n_240),
.C(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_255),
.Y(n_239)
);

XOR2x2_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_253),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_249),
.B2(n_250),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_242),
.B(n_250),
.C(n_253),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_248),
.Y(n_243)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_255),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_267),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_265),
.B2(n_266),
.Y(n_256)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_257),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_266),
.C(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_258),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_264),
.Y(n_258)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_261),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_267),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2x1p5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_303),
.Y(n_276)
);

NOR2x1_ASAP7_75t_L g307 ( 
.A(n_277),
.B(n_303),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_278),
.B(n_281),
.C(n_312),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_292),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_291),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_289),
.B2(n_290),
.Y(n_282)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_283),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_283),
.B(n_290),
.C(n_291),
.Y(n_314)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_284),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_292),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_293),
.B(n_295),
.C(n_301),
.Y(n_333)
);

XOR2x1_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_301),
.Y(n_294)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVxp67_ASAP7_75t_SL g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_339),
.Y(n_308)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_313),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_311),
.B(n_313),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_332),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_321),
.Y(n_316)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_331),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_338),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);


endmodule