module fake_jpeg_10345_n_90 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_90);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_90;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx6_ASAP7_75t_SL g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx11_ASAP7_75t_SL g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_7),
.B(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_1),
.Y(n_26)
);

OAI21xp33_ASAP7_75t_SL g42 ( 
.A1(n_26),
.A2(n_31),
.B(n_32),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_4),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_27),
.B(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_22),
.B(n_11),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_19),
.B(n_5),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_5),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_6),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_24),
.Y(n_45)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

O2A1O1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_30),
.A2(n_20),
.B(n_15),
.C(n_14),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_23),
.B1(n_21),
.B2(n_10),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_47),
.Y(n_53)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_37),
.B(n_29),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_49),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_26),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_SL g50 ( 
.A(n_42),
.B(n_28),
.C(n_10),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_52),
.C(n_59),
.Y(n_61)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_57),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_12),
.Y(n_54)
);

FAx1_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_56),
.CI(n_41),
.CON(n_65),
.SN(n_65)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_18),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_17),
.B1(n_23),
.B2(n_21),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_9),
.Y(n_62)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_40),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_67),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_36),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_51),
.Y(n_68)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_73),
.Y(n_76)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_73),
.B(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_67),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_79),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_61),
.C(n_62),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_83),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_81),
.C(n_70),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_85),
.Y(n_86)
);

NOR2x1_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_74),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_88),
.A2(n_74),
.B(n_65),
.Y(n_89)
);

BUFx24_ASAP7_75t_SL g90 ( 
.A(n_89),
.Y(n_90)
);


endmodule