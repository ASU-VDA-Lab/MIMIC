module fake_netlist_1_5791_n_480 (n_53, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_480);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_480;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_141;
wire n_119;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_67;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_245;
wire n_70;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_68;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g67 ( .A(n_31), .Y(n_67) );
INVx1_ASAP7_75t_L g68 ( .A(n_39), .Y(n_68) );
CKINVDCx20_ASAP7_75t_R g69 ( .A(n_44), .Y(n_69) );
INVx1_ASAP7_75t_SL g70 ( .A(n_28), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_47), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_15), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_4), .Y(n_73) );
CKINVDCx20_ASAP7_75t_R g74 ( .A(n_46), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_8), .Y(n_75) );
INVxp67_ASAP7_75t_SL g76 ( .A(n_21), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_33), .Y(n_77) );
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_1), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_10), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_61), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_9), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_9), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_4), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_18), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_10), .Y(n_85) );
BUFx3_ASAP7_75t_L g86 ( .A(n_23), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_25), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_1), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_36), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_55), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_41), .Y(n_91) );
BUFx2_ASAP7_75t_L g92 ( .A(n_43), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_3), .Y(n_93) );
HB1xp67_ASAP7_75t_L g94 ( .A(n_11), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_62), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_6), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_14), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_64), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_19), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g100 ( .A(n_92), .B(n_0), .Y(n_100) );
AND2x4_ASAP7_75t_L g101 ( .A(n_92), .B(n_0), .Y(n_101) );
INVx3_ASAP7_75t_L g102 ( .A(n_83), .Y(n_102) );
BUFx12f_ASAP7_75t_L g103 ( .A(n_87), .Y(n_103) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_86), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_67), .Y(n_105) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_86), .Y(n_106) );
AND2x2_ASAP7_75t_L g107 ( .A(n_94), .B(n_2), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_67), .Y(n_108) );
NAND2xp33_ASAP7_75t_L g109 ( .A(n_91), .B(n_37), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_72), .B(n_2), .Y(n_110) );
AND2x2_ASAP7_75t_L g111 ( .A(n_83), .B(n_3), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_68), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_72), .B(n_5), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_68), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_71), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_71), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_77), .Y(n_117) );
INVx4_ASAP7_75t_L g118 ( .A(n_98), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_77), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_80), .Y(n_120) );
INVx3_ASAP7_75t_L g121 ( .A(n_80), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_84), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_84), .Y(n_123) );
BUFx2_ASAP7_75t_L g124 ( .A(n_103), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g125 ( .A(n_118), .B(n_99), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_104), .Y(n_126) );
OR2x2_ASAP7_75t_L g127 ( .A(n_100), .B(n_78), .Y(n_127) );
INVx1_ASAP7_75t_SL g128 ( .A(n_103), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_118), .B(n_95), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_115), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_115), .Y(n_131) );
OR2x2_ASAP7_75t_SL g132 ( .A(n_100), .B(n_73), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_107), .B(n_73), .Y(n_133) );
AND2x6_ASAP7_75t_L g134 ( .A(n_101), .B(n_95), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_104), .Y(n_135) );
AO22x2_ASAP7_75t_L g136 ( .A1(n_101), .A2(n_97), .B1(n_75), .B2(n_93), .Y(n_136) );
OAI21xp33_ASAP7_75t_L g137 ( .A1(n_105), .A2(n_97), .B(n_75), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_115), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_104), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_104), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_121), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_118), .B(n_88), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_116), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_116), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_116), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_104), .Y(n_146) );
AOI22xp33_ASAP7_75t_L g147 ( .A1(n_101), .A2(n_81), .B1(n_93), .B2(n_79), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_104), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_107), .B(n_81), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_121), .Y(n_150) );
INVx5_ASAP7_75t_L g151 ( .A(n_134), .Y(n_151) );
OR2x6_ASAP7_75t_L g152 ( .A(n_136), .B(n_101), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_147), .B(n_118), .Y(n_153) );
INVxp67_ASAP7_75t_L g154 ( .A(n_127), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_133), .B(n_111), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_141), .Y(n_156) );
BUFx2_ASAP7_75t_L g157 ( .A(n_136), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_133), .B(n_111), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_141), .Y(n_159) );
BUFx6f_ASAP7_75t_SL g160 ( .A(n_134), .Y(n_160) );
INVx4_ASAP7_75t_L g161 ( .A(n_134), .Y(n_161) );
BUFx4f_ASAP7_75t_L g162 ( .A(n_134), .Y(n_162) );
BUFx3_ASAP7_75t_L g163 ( .A(n_134), .Y(n_163) );
NAND2x1p5_ASAP7_75t_L g164 ( .A(n_141), .B(n_121), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_141), .Y(n_165) );
OAI21xp5_ASAP7_75t_L g166 ( .A1(n_129), .A2(n_105), .B(n_122), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_150), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_149), .B(n_110), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_150), .Y(n_169) );
HB1xp67_ASAP7_75t_L g170 ( .A(n_127), .Y(n_170) );
INVx2_ASAP7_75t_SL g171 ( .A(n_134), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_150), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_149), .B(n_103), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_142), .B(n_108), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_150), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_130), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_130), .Y(n_177) );
AND2x4_ASAP7_75t_L g178 ( .A(n_134), .B(n_110), .Y(n_178) );
BUFx12f_ASAP7_75t_L g179 ( .A(n_124), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_131), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_125), .B(n_108), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_124), .B(n_112), .Y(n_182) );
INVx5_ASAP7_75t_L g183 ( .A(n_126), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_131), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_138), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_161), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_152), .A2(n_136), .B1(n_132), .B2(n_69), .Y(n_187) );
INVx3_ASAP7_75t_L g188 ( .A(n_161), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g189 ( .A1(n_154), .A2(n_137), .B(n_113), .C(n_145), .Y(n_189) );
OR2x2_ASAP7_75t_L g190 ( .A(n_170), .B(n_128), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_180), .Y(n_191) );
NOR2xp67_ASAP7_75t_L g192 ( .A(n_161), .B(n_121), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_180), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_180), .Y(n_194) );
OR2x6_ASAP7_75t_L g195 ( .A(n_152), .B(n_136), .Y(n_195) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_179), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_168), .B(n_138), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_174), .A2(n_145), .B(n_144), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_176), .Y(n_199) );
INVx8_ASAP7_75t_L g200 ( .A(n_152), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_176), .Y(n_201) );
CKINVDCx6p67_ASAP7_75t_R g202 ( .A(n_179), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_151), .B(n_137), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_177), .Y(n_204) );
INVx6_ASAP7_75t_L g205 ( .A(n_151), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_151), .B(n_74), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_163), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_166), .A2(n_144), .B(n_143), .C(n_114), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_163), .Y(n_209) );
INVxp67_ASAP7_75t_SL g210 ( .A(n_157), .Y(n_210) );
BUFx2_ASAP7_75t_L g211 ( .A(n_152), .Y(n_211) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_157), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_173), .Y(n_213) );
INVxp67_ASAP7_75t_SL g214 ( .A(n_162), .Y(n_214) );
AOI22xp33_ASAP7_75t_L g215 ( .A1(n_168), .A2(n_143), .B1(n_122), .B2(n_114), .Y(n_215) );
CKINVDCx6p67_ASAP7_75t_R g216 ( .A(n_160), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_164), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_185), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_177), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_195), .A2(n_187), .B1(n_212), .B2(n_178), .Y(n_220) );
NAND2xp33_ASAP7_75t_SL g221 ( .A(n_211), .B(n_160), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_189), .A2(n_153), .B(n_182), .C(n_113), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_195), .A2(n_178), .B1(n_168), .B2(n_158), .Y(n_223) );
AND2x4_ASAP7_75t_L g224 ( .A(n_217), .B(n_151), .Y(n_224) );
AOI22xp33_ASAP7_75t_SL g225 ( .A1(n_200), .A2(n_160), .B1(n_155), .B2(n_158), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_195), .A2(n_178), .B1(n_162), .B2(n_185), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_195), .A2(n_155), .B1(n_158), .B2(n_162), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_202), .Y(n_228) );
AOI221xp5_ASAP7_75t_L g229 ( .A1(n_215), .A2(n_155), .B1(n_119), .B2(n_112), .C(n_96), .Y(n_229) );
BUFx2_ASAP7_75t_SL g230 ( .A(n_211), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_197), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_202), .Y(n_232) );
OR2x2_ASAP7_75t_L g233 ( .A(n_190), .B(n_132), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_195), .A2(n_89), .B1(n_171), .B2(n_184), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_201), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_210), .A2(n_184), .B1(n_151), .B2(n_171), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_201), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_197), .B(n_164), .Y(n_238) );
OAI22xp33_ASAP7_75t_L g239 ( .A1(n_200), .A2(n_164), .B1(n_156), .B2(n_181), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_199), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_SL g241 ( .A1(n_208), .A2(n_165), .B(n_172), .C(n_169), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_200), .A2(n_156), .B1(n_167), .B2(n_172), .Y(n_242) );
NAND2x1_ASAP7_75t_L g243 ( .A(n_201), .B(n_165), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_199), .A2(n_169), .B(n_167), .Y(n_244) );
NAND3xp33_ASAP7_75t_L g245 ( .A(n_222), .B(n_106), .C(n_219), .Y(n_245) );
AOI221xp5_ASAP7_75t_L g246 ( .A1(n_229), .A2(n_213), .B1(n_190), .B2(n_119), .C(n_204), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_220), .A2(n_200), .B1(n_204), .B2(n_219), .Y(n_247) );
AOI22xp33_ASAP7_75t_SL g248 ( .A1(n_230), .A2(n_200), .B1(n_196), .B2(n_217), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_231), .B(n_218), .Y(n_249) );
BUFx2_ASAP7_75t_L g250 ( .A(n_235), .Y(n_250) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_228), .Y(n_251) );
BUFx2_ASAP7_75t_L g252 ( .A(n_235), .Y(n_252) );
OAI21xp5_ASAP7_75t_L g253 ( .A1(n_244), .A2(n_198), .B(n_192), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g254 ( .A1(n_234), .A2(n_218), .B1(n_206), .B2(n_191), .Y(n_254) );
OR2x6_ASAP7_75t_L g255 ( .A(n_226), .B(n_217), .Y(n_255) );
OAI21x1_ASAP7_75t_L g256 ( .A1(n_243), .A2(n_237), .B(n_240), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_223), .A2(n_217), .B1(n_194), .B2(n_193), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_233), .A2(n_193), .B1(n_194), .B2(n_191), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_233), .A2(n_227), .B1(n_238), .B2(n_225), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_238), .A2(n_191), .B1(n_192), .B2(n_156), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_237), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_243), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_239), .B(n_159), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_221), .A2(n_216), .B1(n_203), .B2(n_188), .Y(n_264) );
INVx4_ASAP7_75t_L g265 ( .A(n_224), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_247), .A2(n_228), .B1(n_232), .B2(n_221), .Y(n_266) );
NAND3xp33_ASAP7_75t_L g267 ( .A(n_245), .B(n_109), .C(n_106), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_259), .A2(n_242), .B1(n_120), .B2(n_123), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_261), .Y(n_269) );
AOI322xp5_ASAP7_75t_L g270 ( .A1(n_246), .A2(n_79), .A3(n_82), .B1(n_85), .B2(n_102), .C1(n_232), .C2(n_120), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_261), .B(n_117), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_250), .Y(n_272) );
OA21x2_ASAP7_75t_L g273 ( .A1(n_245), .A2(n_123), .B(n_120), .Y(n_273) );
OR2x2_ASAP7_75t_L g274 ( .A(n_250), .B(n_224), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_252), .Y(n_275) );
NAND4xp25_ASAP7_75t_L g276 ( .A(n_258), .B(n_82), .C(n_102), .D(n_123), .Y(n_276) );
OR2x6_ASAP7_75t_L g277 ( .A(n_255), .B(n_224), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_251), .B(n_70), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_255), .A2(n_117), .B1(n_236), .B2(n_102), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_265), .B(n_102), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_252), .B(n_117), .Y(n_281) );
OAI211xp5_ASAP7_75t_L g282 ( .A1(n_248), .A2(n_76), .B(n_90), .C(n_241), .Y(n_282) );
AOI22xp33_ASAP7_75t_L g283 ( .A1(n_255), .A2(n_216), .B1(n_188), .B2(n_209), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g284 ( .A1(n_255), .A2(n_188), .B1(n_209), .B2(n_207), .Y(n_284) );
OAI33xp33_ASAP7_75t_L g285 ( .A1(n_249), .A2(n_148), .A3(n_140), .B1(n_146), .B2(n_8), .B3(n_11), .Y(n_285) );
AOI211xp5_ASAP7_75t_L g286 ( .A1(n_254), .A2(n_106), .B(n_148), .C(n_146), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_265), .B(n_5), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_256), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g289 ( .A1(n_268), .A2(n_257), .B1(n_265), .B2(n_254), .Y(n_289) );
AND2x2_ASAP7_75t_SL g290 ( .A(n_287), .B(n_262), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_269), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_269), .B(n_256), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_272), .B(n_262), .Y(n_293) );
INVxp67_ASAP7_75t_L g294 ( .A(n_278), .Y(n_294) );
OAI33xp33_ASAP7_75t_L g295 ( .A1(n_287), .A2(n_263), .A3(n_148), .B1(n_140), .B2(n_13), .B3(n_14), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_272), .B(n_253), .Y(n_296) );
NAND3xp33_ASAP7_75t_L g297 ( .A(n_280), .B(n_106), .C(n_260), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_275), .B(n_264), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_288), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_288), .Y(n_300) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_266), .B(n_106), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_277), .A2(n_106), .B1(n_209), .B2(n_207), .Y(n_302) );
INVxp67_ASAP7_75t_SL g303 ( .A(n_275), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_271), .B(n_6), .Y(n_304) );
NAND3xp33_ASAP7_75t_SL g305 ( .A(n_270), .B(n_7), .C(n_12), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g306 ( .A1(n_277), .A2(n_188), .B1(n_214), .B2(n_186), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_281), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_271), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_281), .B(n_7), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_273), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_274), .B(n_12), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_274), .B(n_277), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_273), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_277), .B(n_13), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g315 ( .A1(n_285), .A2(n_186), .B1(n_209), .B2(n_207), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_273), .B(n_15), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_273), .B(n_16), .Y(n_317) );
AND2x2_ASAP7_75t_SL g318 ( .A(n_279), .B(n_186), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_267), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_286), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_276), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_292), .B(n_284), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_292), .B(n_283), .Y(n_323) );
NOR2xp33_ASAP7_75t_SL g324 ( .A(n_318), .B(n_186), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_299), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_296), .B(n_139), .Y(n_326) );
INVx1_ASAP7_75t_SL g327 ( .A(n_309), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_296), .B(n_16), .Y(n_328) );
BUFx2_ASAP7_75t_L g329 ( .A(n_303), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_297), .A2(n_282), .B(n_186), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_299), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_312), .B(n_139), .Y(n_332) );
NAND2xp5_ASAP7_75t_SL g333 ( .A(n_290), .B(n_186), .Y(n_333) );
AND2x2_ASAP7_75t_SL g334 ( .A(n_290), .B(n_207), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_307), .B(n_139), .Y(n_335) );
NAND4xp25_ASAP7_75t_L g336 ( .A(n_314), .B(n_175), .C(n_159), .D(n_22), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_291), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_300), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_308), .B(n_139), .Y(n_339) );
NAND2xp5_ASAP7_75t_SL g340 ( .A(n_290), .B(n_139), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_300), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_293), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_312), .B(n_139), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_293), .B(n_135), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_308), .B(n_135), .Y(n_345) );
NAND3xp33_ASAP7_75t_L g346 ( .A(n_294), .B(n_135), .C(n_126), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_311), .B(n_135), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_316), .B(n_135), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_316), .B(n_135), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_317), .B(n_126), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_310), .B(n_126), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_310), .Y(n_352) );
AND4x1_ASAP7_75t_L g353 ( .A(n_314), .B(n_17), .C(n_20), .D(n_24), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_313), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_313), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_317), .B(n_126), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_298), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_311), .B(n_126), .Y(n_358) );
INVx3_ASAP7_75t_L g359 ( .A(n_319), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_304), .B(n_309), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_319), .Y(n_361) );
OAI22xp33_ASAP7_75t_L g362 ( .A1(n_321), .A2(n_205), .B1(n_175), .B2(n_183), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_304), .B(n_26), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_298), .B(n_27), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_321), .B(n_29), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_318), .B(n_30), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_327), .B(n_297), .Y(n_367) );
NAND4xp25_ASAP7_75t_L g368 ( .A(n_336), .B(n_305), .C(n_289), .D(n_301), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_357), .B(n_320), .Y(n_369) );
XOR2xp5_ASAP7_75t_L g370 ( .A(n_360), .B(n_306), .Y(n_370) );
NOR2x1_ASAP7_75t_L g371 ( .A(n_336), .B(n_320), .Y(n_371) );
BUFx2_ASAP7_75t_L g372 ( .A(n_329), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_342), .B(n_322), .Y(n_373) );
NOR2xp33_ASAP7_75t_SL g374 ( .A(n_324), .B(n_295), .Y(n_374) );
O2A1O1Ixp33_ASAP7_75t_L g375 ( .A1(n_365), .A2(n_306), .B(n_302), .C(n_315), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_337), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_323), .B(n_315), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_328), .B(n_32), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_342), .B(n_34), .Y(n_379) );
NAND2xp33_ASAP7_75t_SL g380 ( .A(n_363), .B(n_35), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_328), .B(n_38), .Y(n_381) );
INVxp67_ASAP7_75t_SL g382 ( .A(n_346), .Y(n_382) );
INVxp67_ASAP7_75t_L g383 ( .A(n_363), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_338), .B(n_40), .Y(n_384) );
NOR2xp67_ASAP7_75t_L g385 ( .A(n_346), .B(n_42), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_341), .B(n_45), .Y(n_386) );
NOR2xp67_ASAP7_75t_L g387 ( .A(n_366), .B(n_48), .Y(n_387) );
XOR2xp5_ASAP7_75t_SL g388 ( .A(n_366), .B(n_49), .Y(n_388) );
INVxp33_ASAP7_75t_L g389 ( .A(n_332), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_325), .B(n_50), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_353), .B(n_51), .Y(n_391) );
AND4x1_ASAP7_75t_L g392 ( .A(n_324), .B(n_52), .C(n_53), .D(n_54), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_331), .B(n_56), .Y(n_393) );
NAND2x1p5_ASAP7_75t_L g394 ( .A(n_353), .B(n_183), .Y(n_394) );
AOI21xp33_ASAP7_75t_L g395 ( .A1(n_364), .A2(n_57), .B(n_58), .Y(n_395) );
NAND2xp33_ASAP7_75t_SL g396 ( .A(n_340), .B(n_59), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_352), .B(n_60), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_332), .B(n_63), .Y(n_398) );
O2A1O1Ixp33_ASAP7_75t_L g399 ( .A1(n_362), .A2(n_65), .B(n_66), .C(n_183), .Y(n_399) );
INVxp67_ASAP7_75t_SL g400 ( .A(n_372), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_369), .B(n_355), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_373), .B(n_354), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_377), .B(n_361), .Y(n_403) );
OAI322xp33_ASAP7_75t_L g404 ( .A1(n_370), .A2(n_358), .A3(n_347), .B1(n_361), .B2(n_335), .C1(n_339), .C2(n_334), .Y(n_404) );
INVxp67_ASAP7_75t_SL g405 ( .A(n_382), .Y(n_405) );
NAND3xp33_ASAP7_75t_SL g406 ( .A(n_380), .B(n_333), .C(n_330), .Y(n_406) );
XOR2x2_ASAP7_75t_L g407 ( .A(n_388), .B(n_334), .Y(n_407) );
CKINVDCx16_ASAP7_75t_R g408 ( .A(n_371), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_367), .B(n_361), .Y(n_409) );
OAI221xp5_ASAP7_75t_L g410 ( .A1(n_368), .A2(n_359), .B1(n_364), .B2(n_348), .C(n_349), .Y(n_410) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_376), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_383), .B(n_343), .Y(n_412) );
OAI221xp5_ASAP7_75t_L g413 ( .A1(n_374), .A2(n_356), .B1(n_350), .B2(n_349), .C(n_348), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_397), .Y(n_414) );
OAI211xp5_ASAP7_75t_SL g415 ( .A1(n_381), .A2(n_334), .B(n_343), .C(n_326), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_397), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_389), .B(n_343), .Y(n_417) );
NOR2x1_ASAP7_75t_L g418 ( .A(n_385), .B(n_351), .Y(n_418) );
XNOR2xp5_ASAP7_75t_L g419 ( .A(n_392), .B(n_345), .Y(n_419) );
INVxp67_ASAP7_75t_L g420 ( .A(n_374), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_386), .Y(n_421) );
AOI211xp5_ASAP7_75t_L g422 ( .A1(n_387), .A2(n_350), .B(n_356), .C(n_345), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_378), .A2(n_351), .B1(n_344), .B2(n_205), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_390), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_393), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_391), .B(n_344), .Y(n_426) );
NAND2x1_ASAP7_75t_L g427 ( .A(n_379), .B(n_351), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_384), .Y(n_428) );
INVx2_ASAP7_75t_SL g429 ( .A(n_394), .Y(n_429) );
NOR2x1_ASAP7_75t_L g430 ( .A(n_375), .B(n_351), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_398), .Y(n_431) );
XNOR2xp5_ASAP7_75t_L g432 ( .A(n_394), .B(n_396), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_399), .Y(n_433) );
XNOR2xp5_ASAP7_75t_L g434 ( .A(n_395), .B(n_205), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_372), .B(n_183), .Y(n_435) );
NOR3xp33_ASAP7_75t_L g436 ( .A(n_368), .B(n_294), .C(n_305), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_373), .B(n_372), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_372), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_368), .A2(n_371), .B1(n_370), .B2(n_321), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_370), .B(n_294), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g441 ( .A1(n_371), .A2(n_370), .B1(n_327), .B2(n_383), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_368), .A2(n_371), .B1(n_370), .B2(n_321), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_371), .A2(n_368), .B1(n_370), .B2(n_336), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_380), .A2(n_382), .B(n_385), .Y(n_444) );
AND2x4_ASAP7_75t_L g445 ( .A(n_430), .B(n_429), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_409), .Y(n_446) );
INVx1_ASAP7_75t_SL g447 ( .A(n_437), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_440), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_443), .A2(n_439), .B1(n_442), .B2(n_420), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_442), .A2(n_439), .B1(n_420), .B2(n_408), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_444), .A2(n_407), .B(n_432), .Y(n_451) );
XNOR2xp5_ASAP7_75t_L g452 ( .A(n_407), .B(n_441), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_431), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_412), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_411), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_436), .A2(n_433), .B1(n_415), .B2(n_410), .Y(n_456) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_400), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_436), .A2(n_405), .B1(n_417), .B2(n_413), .Y(n_458) );
NOR2xp33_ASAP7_75t_R g459 ( .A(n_406), .B(n_419), .Y(n_459) );
NOR3xp33_ASAP7_75t_SL g460 ( .A(n_451), .B(n_444), .C(n_405), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_451), .A2(n_400), .B(n_435), .Y(n_461) );
AO22x2_ASAP7_75t_L g462 ( .A1(n_445), .A2(n_447), .B1(n_455), .B2(n_452), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_449), .A2(n_426), .B1(n_428), .B2(n_416), .Y(n_463) );
AO22x1_ASAP7_75t_L g464 ( .A1(n_445), .A2(n_418), .B1(n_438), .B2(n_423), .Y(n_464) );
OAI221xp5_ASAP7_75t_SL g465 ( .A1(n_456), .A2(n_422), .B1(n_403), .B2(n_434), .C(n_425), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_457), .Y(n_466) );
INVxp67_ASAP7_75t_L g467 ( .A(n_450), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_467), .Y(n_468) );
AND4x1_ASAP7_75t_L g469 ( .A(n_460), .B(n_458), .C(n_459), .D(n_448), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_466), .Y(n_470) );
OAI222xp33_ASAP7_75t_L g471 ( .A1(n_465), .A2(n_453), .B1(n_454), .B2(n_427), .C1(n_446), .C2(n_402), .Y(n_471) );
AO22x1_ASAP7_75t_L g472 ( .A1(n_469), .A2(n_462), .B1(n_464), .B2(n_461), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_470), .Y(n_473) );
NOR3xp33_ASAP7_75t_SL g474 ( .A(n_471), .B(n_404), .C(n_424), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_473), .Y(n_475) );
AO22x2_ASAP7_75t_L g476 ( .A1(n_472), .A2(n_470), .B1(n_468), .B2(n_463), .Y(n_476) );
OAI22xp33_ASAP7_75t_L g477 ( .A1(n_475), .A2(n_474), .B1(n_421), .B2(n_414), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_477), .Y(n_478) );
XNOR2xp5_ASAP7_75t_L g479 ( .A(n_478), .B(n_476), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_479), .A2(n_411), .B(n_401), .Y(n_480) );
endmodule