module fake_jpeg_28060_n_67 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_67);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_67;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;
wire n_66;

INVx1_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

BUFx5_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

BUFx5_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx2_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_18),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_15),
.B(n_17),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_0),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_14),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_15),
.B(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_23),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_16),
.C(n_19),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_22),
.Y(n_31)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_26),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_19),
.A2(n_16),
.B1(n_7),
.B2(n_13),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_7),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_29),
.A2(n_20),
.B1(n_12),
.B2(n_13),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_30),
.A2(n_35),
.B(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_32),
.B(n_27),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_23),
.B1(n_21),
.B2(n_17),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_28),
.A2(n_21),
.B1(n_23),
.B2(n_8),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_39),
.Y(n_44)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_24),
.C(n_21),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_28),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_30),
.B(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_8),
.Y(n_50)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_40),
.C(n_19),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_51),
.C(n_49),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_SL g55 ( 
.A(n_50),
.B(n_18),
.Y(n_55)
);

MAJx2_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_8),
.C(n_9),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_43),
.B1(n_44),
.B2(n_25),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_25),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_51),
.A2(n_25),
.B1(n_10),
.B2(n_6),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_54),
.B(n_56),
.Y(n_59)
);

OAI21x1_ASAP7_75t_L g58 ( 
.A1(n_55),
.A2(n_10),
.B(n_5),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_58),
.A2(n_5),
.B(n_2),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_57),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_61),
.Y(n_64)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

AOI322xp5_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_10),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_1),
.C2(n_26),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_63),
.B(n_2),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_64),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_66),
.B(n_26),
.Y(n_67)
);


endmodule