module fake_ariane_1691_n_975 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_975);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_975;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_651;
wire n_936;
wire n_347;
wire n_423;
wire n_961;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_908;
wire n_788;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_445;
wire n_379;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_885;
wire n_737;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_207;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_285;
wire n_473;
wire n_801;
wire n_202;
wire n_761;
wire n_733;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_903;
wire n_315;
wire n_871;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_331;
wire n_320;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_840;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_795;
wire n_398;
wire n_210;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_839;
wire n_821;
wire n_928;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_512;
wire n_715;
wire n_889;
wire n_935;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_658;
wire n_617;
wire n_705;
wire n_630;
wire n_616;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_747;
wire n_741;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_888;
wire n_845;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_915;
wire n_215;
wire n_252;
wire n_664;
wire n_629;
wire n_454;
wire n_966;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_213;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_931;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_963;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_882;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_174),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_18),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_29),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_126),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_16),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_20),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_5),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_124),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_167),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_10),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_3),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_136),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_42),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_123),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_141),
.Y(n_217)
);

BUFx10_ASAP7_75t_L g218 ( 
.A(n_21),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_98),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_49),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_129),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_100),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_122),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_76),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_40),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_92),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_81),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_80),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_24),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_96),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_8),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_70),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_194),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_14),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_23),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_120),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_66),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_134),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_199),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_60),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_108),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_26),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_19),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_33),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_102),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_94),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_62),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_200),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_185),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_183),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_184),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_25),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_101),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_145),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_180),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_138),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_179),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_157),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_153),
.B(n_162),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_118),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_178),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_71),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_197),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_109),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_90),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_39),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_11),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_16),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_175),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_88),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_156),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_31),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_99),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_106),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_97),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_112),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_32),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_103),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_140),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_57),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_116),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_89),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_47),
.Y(n_283)
);

OAI21x1_ASAP7_75t_L g284 ( 
.A1(n_219),
.A2(n_91),
.B(n_196),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_240),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_260),
.A2(n_223),
.B1(n_237),
.B2(n_212),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_240),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_218),
.Y(n_289)
);

OAI22x1_ASAP7_75t_R g290 ( 
.A1(n_209),
.A2(n_243),
.B1(n_231),
.B2(n_202),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_270),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_223),
.B(n_0),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_218),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_207),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_213),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_234),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_219),
.Y(n_297)
);

AND2x4_ASAP7_75t_L g298 ( 
.A(n_227),
.B(n_0),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_227),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_218),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_267),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_216),
.B(n_1),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_203),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_233),
.B(n_1),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_268),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_204),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_205),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_229),
.Y(n_308)
);

AND2x4_ASAP7_75t_L g309 ( 
.A(n_229),
.B(n_2),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_208),
.Y(n_310)
);

NAND3xp33_ASAP7_75t_L g311 ( 
.A(n_238),
.B(n_2),
.C(n_3),
.Y(n_311)
);

OAI21x1_ASAP7_75t_L g312 ( 
.A1(n_238),
.A2(n_95),
.B(n_195),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_260),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_211),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_230),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_245),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_246),
.Y(n_317)
);

CKINVDCx11_ASAP7_75t_R g318 ( 
.A(n_281),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_248),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_242),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_250),
.B(n_4),
.Y(n_321)
);

AND2x4_ASAP7_75t_L g322 ( 
.A(n_251),
.B(n_4),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_242),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_253),
.Y(n_324)
);

OA21x2_ASAP7_75t_L g325 ( 
.A1(n_261),
.A2(n_5),
.B(n_6),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_262),
.Y(n_326)
);

AND2x4_ASAP7_75t_L g327 ( 
.A(n_263),
.B(n_6),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_244),
.Y(n_328)
);

INVx5_ASAP7_75t_L g329 ( 
.A(n_259),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_266),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_244),
.Y(n_331)
);

INVx2_ASAP7_75t_SL g332 ( 
.A(n_283),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_201),
.B(n_7),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_206),
.Y(n_334)
);

INVx5_ASAP7_75t_L g335 ( 
.A(n_210),
.Y(n_335)
);

AND2x4_ASAP7_75t_L g336 ( 
.A(n_214),
.B(n_7),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_285),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_297),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_331),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_318),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_R g341 ( 
.A(n_331),
.B(n_215),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_297),
.Y(n_342)
);

AND3x2_ASAP7_75t_L g343 ( 
.A(n_304),
.B(n_8),
.C(n_9),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_318),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_313),
.Y(n_345)
);

NAND2xp33_ASAP7_75t_L g346 ( 
.A(n_292),
.B(n_217),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_295),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_320),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_328),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_298),
.B(n_309),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_285),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_334),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_285),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_285),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_288),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_288),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_323),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_293),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_297),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_289),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_R g361 ( 
.A(n_293),
.B(n_220),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_286),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_289),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_289),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_297),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_289),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_335),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_335),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_293),
.B(n_300),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_335),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_335),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_299),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_290),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_288),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_288),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_300),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_287),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_317),
.Y(n_378)
);

NOR2xp67_ASAP7_75t_L g379 ( 
.A(n_300),
.B(n_221),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_315),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_299),
.Y(n_381)
);

NOR2xp67_ASAP7_75t_L g382 ( 
.A(n_329),
.B(n_296),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_315),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_287),
.Y(n_384)
);

AND3x2_ASAP7_75t_L g385 ( 
.A(n_298),
.B(n_9),
.C(n_10),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_299),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_317),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_299),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_317),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_317),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_329),
.B(n_222),
.Y(n_391)
);

NAND2xp33_ASAP7_75t_L g392 ( 
.A(n_376),
.B(n_321),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_377),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_377),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_347),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_380),
.B(n_336),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_378),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_358),
.B(n_329),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_369),
.B(n_329),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_383),
.B(n_329),
.Y(n_400)
);

NOR3xp33_ASAP7_75t_L g401 ( 
.A(n_357),
.B(n_302),
.C(n_333),
.Y(n_401)
);

INVx2_ASAP7_75t_SL g402 ( 
.A(n_348),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_337),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_350),
.B(n_322),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_387),
.Y(n_405)
);

OR2x6_ASAP7_75t_L g406 ( 
.A(n_350),
.B(n_294),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_361),
.B(n_336),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_389),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_351),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_353),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_354),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_372),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_390),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_356),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_382),
.B(n_322),
.Y(n_415)
);

BUFx5_ASAP7_75t_L g416 ( 
.A(n_355),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_390),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_374),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_372),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_375),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_360),
.B(n_322),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_361),
.B(n_336),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_384),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_338),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_349),
.B(n_327),
.Y(n_425)
);

OR2x2_ASAP7_75t_SL g426 ( 
.A(n_373),
.B(n_301),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_372),
.Y(n_427)
);

A2O1A1Ixp33_ASAP7_75t_L g428 ( 
.A1(n_346),
.A2(n_298),
.B(n_309),
.C(n_327),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_338),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_363),
.B(n_306),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_339),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_352),
.A2(n_309),
.B1(n_327),
.B2(n_333),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_341),
.B(n_379),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_342),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_L g435 ( 
.A1(n_391),
.A2(n_332),
.B1(n_326),
.B2(n_316),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_364),
.B(n_291),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_366),
.B(n_291),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_341),
.B(n_319),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_391),
.B(n_332),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_342),
.B(n_324),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_359),
.B(n_324),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_340),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_359),
.B(n_324),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_365),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_345),
.B(n_303),
.Y(n_445)
);

NAND2xp33_ASAP7_75t_L g446 ( 
.A(n_367),
.B(n_368),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_370),
.B(n_303),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_365),
.Y(n_448)
);

NAND3xp33_ASAP7_75t_L g449 ( 
.A(n_372),
.B(n_325),
.C(n_319),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_386),
.B(n_308),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_386),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_381),
.B(n_319),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_388),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g454 ( 
.A(n_344),
.B(n_305),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_381),
.B(n_319),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_388),
.B(n_308),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_371),
.B(n_308),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_381),
.B(n_307),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_381),
.B(n_310),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_385),
.B(n_310),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_343),
.B(n_314),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_362),
.B(n_314),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_377),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_369),
.B(n_330),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_431),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_450),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_456),
.Y(n_467)
);

AO22x1_ASAP7_75t_L g468 ( 
.A1(n_402),
.A2(n_305),
.B1(n_224),
.B2(n_258),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_404),
.B(n_330),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_423),
.B(n_311),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_432),
.A2(n_401),
.B1(n_422),
.B2(n_407),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_406),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_442),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_444),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_424),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_440),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_454),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_432),
.A2(n_265),
.B1(n_226),
.B2(n_228),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_462),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_406),
.A2(n_325),
.B1(n_330),
.B2(n_269),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_445),
.B(n_330),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_425),
.B(n_225),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_406),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_441),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_L g485 ( 
.A1(n_395),
.A2(n_325),
.B1(n_271),
.B2(n_264),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_392),
.A2(n_257),
.B1(n_235),
.B2(n_282),
.Y(n_486)
);

AO22x1_ASAP7_75t_L g487 ( 
.A1(n_461),
.A2(n_275),
.B1(n_236),
.B2(n_239),
.Y(n_487)
);

BUFx8_ASAP7_75t_L g488 ( 
.A(n_393),
.Y(n_488)
);

BUFx4f_ASAP7_75t_L g489 ( 
.A(n_394),
.Y(n_489)
);

INVx5_ASAP7_75t_L g490 ( 
.A(n_412),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_447),
.B(n_232),
.Y(n_491)
);

OR2x2_ASAP7_75t_SL g492 ( 
.A(n_426),
.B(n_11),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_436),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_400),
.B(n_241),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_439),
.B(n_247),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_430),
.B(n_249),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_461),
.A2(n_278),
.B1(n_254),
.B2(n_255),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_464),
.B(n_252),
.Y(n_498)
);

NAND2x1p5_ASAP7_75t_L g499 ( 
.A(n_433),
.B(n_284),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_399),
.A2(n_312),
.B(n_284),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_398),
.B(n_421),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_428),
.B(n_256),
.Y(n_502)
);

BUFx4f_ASAP7_75t_SL g503 ( 
.A(n_438),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_460),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_412),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_415),
.B(n_272),
.Y(n_506)
);

NOR2x1_ASAP7_75t_L g507 ( 
.A(n_396),
.B(n_273),
.Y(n_507)
);

BUFx8_ASAP7_75t_L g508 ( 
.A(n_463),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_443),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_435),
.A2(n_280),
.B1(n_279),
.B2(n_277),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_448),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_437),
.B(n_12),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_419),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_457),
.A2(n_276),
.B1(n_274),
.B2(n_312),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_397),
.B(n_13),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_403),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_412),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_405),
.B(n_13),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_408),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_SL g520 ( 
.A1(n_449),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_419),
.B(n_416),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_413),
.Y(n_522)
);

AND2x6_ASAP7_75t_SL g523 ( 
.A(n_458),
.B(n_19),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_417),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_418),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_449),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_409),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_429),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_459),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_452),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_434),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_451),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_453),
.B(n_198),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_410),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_446),
.B(n_41),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_411),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_414),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_416),
.B(n_46),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_416),
.B(n_193),
.Y(n_539)
);

NOR2x1_ASAP7_75t_R g540 ( 
.A(n_416),
.B(n_48),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_416),
.B(n_427),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_420),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_427),
.B(n_53),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_427),
.B(n_192),
.Y(n_544)
);

AND3x1_ASAP7_75t_L g545 ( 
.A(n_455),
.B(n_54),
.C(n_55),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g546 ( 
.A(n_431),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_442),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_522),
.Y(n_548)
);

INVx6_ASAP7_75t_L g549 ( 
.A(n_488),
.Y(n_549)
);

O2A1O1Ixp5_ASAP7_75t_L g550 ( 
.A1(n_501),
.A2(n_506),
.B(n_496),
.C(n_500),
.Y(n_550)
);

A2O1A1Ixp33_ASAP7_75t_L g551 ( 
.A1(n_471),
.A2(n_56),
.B(n_58),
.C(n_59),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_521),
.A2(n_61),
.B(n_63),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_475),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_479),
.B(n_64),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_541),
.A2(n_65),
.B(n_67),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_473),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_517),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_470),
.B(n_68),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_498),
.A2(n_69),
.B(n_72),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_493),
.B(n_73),
.Y(n_560)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_546),
.B(n_74),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_465),
.Y(n_562)
);

INVx4_ASAP7_75t_L g563 ( 
.A(n_547),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_511),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_516),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_477),
.B(n_191),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_490),
.Y(n_567)
);

NOR3xp33_ASAP7_75t_SL g568 ( 
.A(n_519),
.B(n_75),
.C(n_77),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_476),
.A2(n_78),
.B(n_79),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_504),
.B(n_82),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_484),
.A2(n_83),
.B(n_84),
.Y(n_571)
);

NAND2x1p5_ASAP7_75t_L g572 ( 
.A(n_489),
.B(n_85),
.Y(n_572)
);

A2O1A1Ixp33_ASAP7_75t_L g573 ( 
.A1(n_478),
.A2(n_86),
.B(n_87),
.C(n_93),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_482),
.A2(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_574)
);

INVxp67_ASAP7_75t_L g575 ( 
.A(n_472),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_483),
.B(n_110),
.Y(n_576)
);

O2A1O1Ixp33_ASAP7_75t_SL g577 ( 
.A1(n_535),
.A2(n_111),
.B(n_113),
.C(n_114),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_509),
.A2(n_115),
.B(n_117),
.Y(n_578)
);

INVx4_ASAP7_75t_L g579 ( 
.A(n_490),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_491),
.A2(n_119),
.B1(n_121),
.B2(n_125),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_495),
.A2(n_127),
.B(n_128),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_492),
.B(n_130),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_503),
.B(n_131),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_489),
.B(n_132),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_534),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_525),
.B(n_133),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_480),
.A2(n_135),
.B1(n_137),
.B2(n_139),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_524),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_481),
.B(n_142),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_532),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_469),
.A2(n_143),
.B(n_144),
.Y(n_591)
);

OR2x6_ASAP7_75t_L g592 ( 
.A(n_468),
.B(n_146),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_486),
.B(n_147),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_512),
.B(n_148),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_529),
.B(n_149),
.Y(n_595)
);

NAND3xp33_ASAP7_75t_SL g596 ( 
.A(n_510),
.B(n_150),
.C(n_151),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_466),
.B(n_152),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_510),
.B(n_190),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_488),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_467),
.B(n_154),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_508),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_515),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_474),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_480),
.B(n_155),
.Y(n_604)
);

OR2x2_ASAP7_75t_L g605 ( 
.A(n_497),
.B(n_158),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_520),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_494),
.B(n_528),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_508),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_490),
.B(n_163),
.Y(n_609)
);

O2A1O1Ixp33_ASAP7_75t_L g610 ( 
.A1(n_518),
.A2(n_164),
.B(n_165),
.C(n_166),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_502),
.A2(n_168),
.B(n_169),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_507),
.B(n_170),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_556),
.Y(n_613)
);

NAND2x1p5_ASAP7_75t_L g614 ( 
.A(n_567),
.B(n_505),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_548),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_567),
.B(n_505),
.Y(n_616)
);

NAND2x1p5_ASAP7_75t_L g617 ( 
.A(n_579),
.B(n_513),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_557),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_602),
.B(n_607),
.Y(n_619)
);

OR2x6_ASAP7_75t_L g620 ( 
.A(n_549),
.B(n_536),
.Y(n_620)
);

INVx6_ASAP7_75t_L g621 ( 
.A(n_579),
.Y(n_621)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_549),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_557),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_557),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_585),
.Y(n_625)
);

OAI21xp5_ASAP7_75t_L g626 ( 
.A1(n_550),
.A2(n_514),
.B(n_499),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_563),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_588),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_575),
.Y(n_629)
);

INVx5_ASAP7_75t_L g630 ( 
.A(n_592),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_558),
.A2(n_539),
.B(n_538),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_562),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_590),
.Y(n_633)
);

OR2x6_ASAP7_75t_L g634 ( 
.A(n_599),
.B(n_530),
.Y(n_634)
);

OAI21x1_ASAP7_75t_L g635 ( 
.A1(n_589),
.A2(n_543),
.B(n_513),
.Y(n_635)
);

OAI21xp33_ASAP7_75t_SL g636 ( 
.A1(n_598),
.A2(n_485),
.B(n_544),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_553),
.Y(n_637)
);

INVx1_ASAP7_75t_SL g638 ( 
.A(n_554),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_564),
.Y(n_639)
);

OR2x6_ASAP7_75t_L g640 ( 
.A(n_601),
.B(n_563),
.Y(n_640)
);

INVx6_ASAP7_75t_L g641 ( 
.A(n_561),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_572),
.Y(n_642)
);

OAI21x1_ASAP7_75t_SL g643 ( 
.A1(n_610),
.A2(n_531),
.B(n_542),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_565),
.Y(n_644)
);

BUFx2_ASAP7_75t_SL g645 ( 
.A(n_612),
.Y(n_645)
);

AOI21x1_ASAP7_75t_L g646 ( 
.A1(n_595),
.A2(n_487),
.B(n_533),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_603),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_612),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_560),
.B(n_517),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_605),
.Y(n_650)
);

OA21x2_ASAP7_75t_L g651 ( 
.A1(n_604),
.A2(n_537),
.B(n_527),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_597),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_608),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_600),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_592),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_570),
.B(n_517),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_582),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_594),
.Y(n_658)
);

OAI21x1_ASAP7_75t_L g659 ( 
.A1(n_611),
.A2(n_545),
.B(n_526),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_576),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_566),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_586),
.B(n_540),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_583),
.B(n_523),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_574),
.Y(n_664)
);

OAI21x1_ASAP7_75t_L g665 ( 
.A1(n_559),
.A2(n_540),
.B(n_172),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_609),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_584),
.Y(n_667)
);

AO21x2_ASAP7_75t_L g668 ( 
.A1(n_593),
.A2(n_171),
.B(n_176),
.Y(n_668)
);

AO21x2_ASAP7_75t_L g669 ( 
.A1(n_596),
.A2(n_177),
.B(n_181),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_568),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_613),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_633),
.Y(n_672)
);

INVx1_ASAP7_75t_SL g673 ( 
.A(n_613),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_650),
.A2(n_587),
.B1(n_606),
.B2(n_580),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_620),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_625),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_650),
.A2(n_569),
.B1(n_578),
.B2(n_571),
.Y(n_677)
);

OAI22xp5_ASAP7_75t_L g678 ( 
.A1(n_660),
.A2(n_551),
.B1(n_573),
.B2(n_581),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g679 ( 
.A1(n_662),
.A2(n_552),
.B1(n_555),
.B2(n_591),
.Y(n_679)
);

OA21x2_ASAP7_75t_L g680 ( 
.A1(n_631),
.A2(n_577),
.B(n_187),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_633),
.Y(n_681)
);

OAI21x1_ASAP7_75t_L g682 ( 
.A1(n_635),
.A2(n_182),
.B(n_188),
.Y(n_682)
);

BUFx10_ASAP7_75t_L g683 ( 
.A(n_653),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_650),
.A2(n_189),
.B1(n_664),
.B2(n_661),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_650),
.A2(n_636),
.B1(n_638),
.B2(n_664),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_615),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_628),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_637),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_618),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_639),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_644),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_620),
.Y(n_692)
);

OAI21x1_ASAP7_75t_L g693 ( 
.A1(n_626),
.A2(n_631),
.B(n_665),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_647),
.Y(n_694)
);

BUFx2_ASAP7_75t_L g695 ( 
.A(n_634),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_632),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_618),
.Y(n_697)
);

OAI22xp33_ASAP7_75t_L g698 ( 
.A1(n_663),
.A2(n_662),
.B1(n_638),
.B2(n_657),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_647),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_629),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_619),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_619),
.Y(n_702)
);

OAI21x1_ASAP7_75t_L g703 ( 
.A1(n_626),
.A2(n_659),
.B(n_646),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_SL g704 ( 
.A1(n_645),
.A2(n_648),
.B1(n_630),
.B2(n_641),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_634),
.Y(n_705)
);

BUFx12f_ASAP7_75t_L g706 ( 
.A(n_622),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_629),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_657),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_618),
.Y(n_709)
);

AO21x2_ASAP7_75t_L g710 ( 
.A1(n_649),
.A2(n_643),
.B(n_654),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_624),
.Y(n_711)
);

HB1xp67_ASAP7_75t_L g712 ( 
.A(n_632),
.Y(n_712)
);

INVx8_ASAP7_75t_L g713 ( 
.A(n_620),
.Y(n_713)
);

CKINVDCx6p67_ASAP7_75t_R g714 ( 
.A(n_622),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_627),
.Y(n_715)
);

BUFx4f_ASAP7_75t_L g716 ( 
.A(n_648),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_618),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_624),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_623),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_623),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_652),
.Y(n_721)
);

INVx5_ASAP7_75t_L g722 ( 
.A(n_648),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_648),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_670),
.B(n_656),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_R g725 ( 
.A(n_715),
.B(n_627),
.Y(n_725)
);

NAND2xp33_ASAP7_75t_SL g726 ( 
.A(n_715),
.B(n_656),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_686),
.Y(n_727)
);

AND2x4_ASAP7_75t_SL g728 ( 
.A(n_714),
.B(n_640),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_687),
.Y(n_729)
);

OR2x6_ASAP7_75t_L g730 ( 
.A(n_713),
.B(n_655),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_712),
.B(n_634),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_713),
.Y(n_732)
);

NOR3xp33_ASAP7_75t_SL g733 ( 
.A(n_724),
.B(n_640),
.C(n_649),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_701),
.B(n_630),
.Y(n_734)
);

BUFx2_ASAP7_75t_SL g735 ( 
.A(n_671),
.Y(n_735)
);

CKINVDCx20_ASAP7_75t_R g736 ( 
.A(n_706),
.Y(n_736)
);

NAND2xp33_ASAP7_75t_R g737 ( 
.A(n_695),
.B(n_655),
.Y(n_737)
);

INVx4_ASAP7_75t_SL g738 ( 
.A(n_689),
.Y(n_738)
);

AOI211xp5_ASAP7_75t_SL g739 ( 
.A1(n_678),
.A2(n_658),
.B(n_667),
.C(n_666),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_713),
.Y(n_740)
);

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_673),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_683),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_712),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_676),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_691),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_R g746 ( 
.A(n_716),
.B(n_630),
.Y(n_746)
);

HB1xp67_ASAP7_75t_L g747 ( 
.A(n_700),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_721),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_688),
.Y(n_749)
);

NAND2xp33_ASAP7_75t_R g750 ( 
.A(n_705),
.B(n_640),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_700),
.B(n_641),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_696),
.B(n_641),
.Y(n_752)
);

INVx3_ASAP7_75t_SL g753 ( 
.A(n_683),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_702),
.B(n_630),
.Y(n_754)
);

CKINVDCx16_ASAP7_75t_R g755 ( 
.A(n_675),
.Y(n_755)
);

NAND3xp33_ASAP7_75t_L g756 ( 
.A(n_724),
.B(n_658),
.C(n_642),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_685),
.B(n_623),
.Y(n_757)
);

NAND3xp33_ASAP7_75t_SL g758 ( 
.A(n_674),
.B(n_614),
.C(n_617),
.Y(n_758)
);

BUFx2_ASAP7_75t_L g759 ( 
.A(n_696),
.Y(n_759)
);

NOR2x1_ASAP7_75t_L g760 ( 
.A(n_698),
.B(n_642),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_707),
.B(n_616),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_672),
.Y(n_762)
);

BUFx4f_ASAP7_75t_SL g763 ( 
.A(n_692),
.Y(n_763)
);

NAND2x1p5_ASAP7_75t_L g764 ( 
.A(n_722),
.B(n_623),
.Y(n_764)
);

BUFx2_ASAP7_75t_L g765 ( 
.A(n_689),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_690),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_R g767 ( 
.A(n_716),
.B(n_621),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_698),
.B(n_621),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_681),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_711),
.Y(n_770)
);

BUFx12f_ASAP7_75t_L g771 ( 
.A(n_689),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_708),
.B(n_616),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_R g773 ( 
.A(n_697),
.B(n_621),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_694),
.Y(n_774)
);

OAI21xp5_ASAP7_75t_L g775 ( 
.A1(n_674),
.A2(n_651),
.B(n_617),
.Y(n_775)
);

HB1xp67_ASAP7_75t_L g776 ( 
.A(n_717),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_R g777 ( 
.A(n_697),
.B(n_614),
.Y(n_777)
);

BUFx2_ASAP7_75t_L g778 ( 
.A(n_689),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_684),
.A2(n_651),
.B1(n_669),
.B2(n_668),
.Y(n_779)
);

CKINVDCx16_ASAP7_75t_R g780 ( 
.A(n_717),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_709),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_R g782 ( 
.A(n_709),
.B(n_669),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_743),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_747),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_748),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_759),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_727),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_751),
.B(n_699),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_780),
.B(n_710),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_729),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_731),
.B(n_774),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_781),
.Y(n_792)
);

BUFx2_ASAP7_75t_L g793 ( 
.A(n_776),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_749),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_760),
.A2(n_684),
.B1(n_704),
.B2(n_723),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_782),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_761),
.B(n_710),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_766),
.Y(n_798)
);

BUFx2_ASAP7_75t_L g799 ( 
.A(n_765),
.Y(n_799)
);

INVxp67_ASAP7_75t_L g800 ( 
.A(n_735),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_769),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_762),
.B(n_703),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_752),
.B(n_719),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_744),
.Y(n_804)
);

OR2x6_ASAP7_75t_L g805 ( 
.A(n_775),
.B(n_693),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_745),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_775),
.B(n_720),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_778),
.B(n_720),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_734),
.B(n_718),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_757),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_771),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_734),
.B(n_720),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_757),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_781),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_754),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_754),
.B(n_720),
.Y(n_816)
);

BUFx2_ASAP7_75t_L g817 ( 
.A(n_781),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_738),
.B(n_722),
.Y(n_818)
);

BUFx3_ASAP7_75t_L g819 ( 
.A(n_728),
.Y(n_819)
);

NOR2x1_ASAP7_75t_L g820 ( 
.A(n_756),
.B(n_709),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_770),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_739),
.B(n_709),
.Y(n_822)
);

OR2x2_ASAP7_75t_L g823 ( 
.A(n_756),
.B(n_680),
.Y(n_823)
);

BUFx2_ASAP7_75t_SL g824 ( 
.A(n_741),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_768),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_739),
.B(n_722),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_772),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_738),
.B(n_722),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_758),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_755),
.B(n_704),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_798),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_798),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_804),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_784),
.B(n_733),
.Y(n_834)
);

NOR3xp33_ASAP7_75t_L g835 ( 
.A(n_800),
.B(n_726),
.C(n_758),
.Y(n_835)
);

NOR2x1_ASAP7_75t_L g836 ( 
.A(n_824),
.B(n_811),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_783),
.B(n_730),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_804),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_820),
.B(n_725),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_793),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_802),
.B(n_779),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_786),
.B(n_742),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_802),
.B(n_738),
.Y(n_843)
);

OR2x2_ASAP7_75t_L g844 ( 
.A(n_793),
.B(n_730),
.Y(n_844)
);

NAND2x1p5_ASAP7_75t_L g845 ( 
.A(n_818),
.B(n_732),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_791),
.B(n_753),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_791),
.B(n_680),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_815),
.B(n_730),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_825),
.B(n_763),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_807),
.B(n_680),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_807),
.B(n_682),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_787),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_790),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_785),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_794),
.B(n_764),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_801),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_796),
.B(n_740),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_813),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_805),
.B(n_764),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_809),
.B(n_773),
.Y(n_860)
);

INVxp33_ASAP7_75t_L g861 ( 
.A(n_792),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_805),
.B(n_668),
.Y(n_862)
);

OR2x2_ASAP7_75t_L g863 ( 
.A(n_797),
.B(n_750),
.Y(n_863)
);

HB1xp67_ASAP7_75t_L g864 ( 
.A(n_799),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_799),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_813),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_803),
.B(n_777),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_806),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_841),
.B(n_805),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_854),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_854),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_841),
.B(n_805),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_847),
.B(n_808),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_847),
.B(n_808),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_843),
.B(n_803),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_843),
.B(n_789),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_858),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_864),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_866),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_840),
.B(n_812),
.Y(n_880)
);

OR2x2_ASAP7_75t_L g881 ( 
.A(n_865),
.B(n_852),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_831),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_833),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_832),
.Y(n_884)
);

BUFx2_ASAP7_75t_L g885 ( 
.A(n_857),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_834),
.A2(n_824),
.B1(n_830),
.B2(n_795),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_853),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_859),
.B(n_796),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_857),
.B(n_736),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_851),
.B(n_789),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_851),
.B(n_822),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_881),
.Y(n_892)
);

NAND4xp75_ASAP7_75t_SL g893 ( 
.A(n_889),
.B(n_862),
.C(n_849),
.D(n_836),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_885),
.Y(n_894)
);

OAI32xp33_ASAP7_75t_L g895 ( 
.A1(n_886),
.A2(n_835),
.A3(n_844),
.B1(n_823),
.B2(n_860),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_881),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_880),
.B(n_890),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_890),
.B(n_856),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_875),
.B(n_857),
.Y(n_899)
);

OR2x2_ASAP7_75t_L g900 ( 
.A(n_878),
.B(n_863),
.Y(n_900)
);

NOR2x1_ASAP7_75t_L g901 ( 
.A(n_887),
.B(n_842),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_882),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_870),
.Y(n_903)
);

OR2x2_ASAP7_75t_L g904 ( 
.A(n_878),
.B(n_848),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_884),
.Y(n_905)
);

NAND3xp33_ASAP7_75t_SL g906 ( 
.A(n_900),
.B(n_839),
.C(n_869),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_895),
.A2(n_869),
.B(n_872),
.Y(n_907)
);

OAI22xp5_ASAP7_75t_L g908 ( 
.A1(n_899),
.A2(n_872),
.B1(n_839),
.B2(n_891),
.Y(n_908)
);

NAND3xp33_ASAP7_75t_L g909 ( 
.A(n_901),
.B(n_879),
.C(n_877),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_892),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_896),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_903),
.A2(n_829),
.B1(n_862),
.B2(n_876),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_902),
.B(n_875),
.Y(n_913)
);

OAI22xp33_ASAP7_75t_SL g914 ( 
.A1(n_898),
.A2(n_821),
.B1(n_867),
.B2(n_868),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_895),
.A2(n_849),
.B(n_846),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_910),
.Y(n_916)
);

OAI31xp33_ASAP7_75t_L g917 ( 
.A1(n_914),
.A2(n_891),
.A3(n_876),
.B(n_888),
.Y(n_917)
);

AOI221x1_ASAP7_75t_L g918 ( 
.A1(n_915),
.A2(n_905),
.B1(n_821),
.B2(n_888),
.C(n_814),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_911),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_913),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_909),
.Y(n_921)
);

NOR2x1p5_ASAP7_75t_L g922 ( 
.A(n_906),
.B(n_819),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_908),
.B(n_897),
.Y(n_923)
);

OAI21xp33_ASAP7_75t_L g924 ( 
.A1(n_907),
.A2(n_904),
.B(n_874),
.Y(n_924)
);

AOI221x1_ASAP7_75t_L g925 ( 
.A1(n_921),
.A2(n_888),
.B1(n_814),
.B2(n_788),
.C(n_816),
.Y(n_925)
);

OAI322xp33_ASAP7_75t_L g926 ( 
.A1(n_923),
.A2(n_837),
.A3(n_823),
.B1(n_894),
.B2(n_850),
.C1(n_873),
.C2(n_874),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_918),
.A2(n_912),
.B(n_822),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_920),
.B(n_919),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_916),
.Y(n_929)
);

INVx5_ASAP7_75t_L g930 ( 
.A(n_928),
.Y(n_930)
);

NOR3xp33_ASAP7_75t_L g931 ( 
.A(n_929),
.B(n_924),
.C(n_923),
.Y(n_931)
);

NOR3xp33_ASAP7_75t_L g932 ( 
.A(n_928),
.B(n_916),
.C(n_811),
.Y(n_932)
);

NOR2x1_ASAP7_75t_L g933 ( 
.A(n_926),
.B(n_922),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_930),
.B(n_927),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_931),
.B(n_925),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_932),
.B(n_917),
.Y(n_936)
);

NAND3xp33_ASAP7_75t_L g937 ( 
.A(n_933),
.B(n_677),
.C(n_792),
.Y(n_937)
);

OAI211xp5_ASAP7_75t_L g938 ( 
.A1(n_935),
.A2(n_746),
.B(n_767),
.C(n_893),
.Y(n_938)
);

INVxp67_ASAP7_75t_L g939 ( 
.A(n_934),
.Y(n_939)
);

INVxp67_ASAP7_75t_L g940 ( 
.A(n_936),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_937),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_935),
.B(n_873),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_934),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_943),
.Y(n_944)
);

NAND4xp75_ASAP7_75t_L g945 ( 
.A(n_941),
.B(n_826),
.C(n_828),
.D(n_859),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_942),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_940),
.Y(n_947)
);

OR2x2_ASAP7_75t_L g948 ( 
.A(n_939),
.B(n_845),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_938),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_947),
.Y(n_950)
);

NOR2x1p5_ASAP7_75t_L g951 ( 
.A(n_944),
.B(n_946),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_949),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_945),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_948),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_951),
.Y(n_955)
);

AOI22x1_ASAP7_75t_L g956 ( 
.A1(n_952),
.A2(n_845),
.B1(n_792),
.B2(n_817),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_953),
.A2(n_954),
.B1(n_950),
.B2(n_952),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_951),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_951),
.Y(n_959)
);

CKINVDCx20_ASAP7_75t_R g960 ( 
.A(n_957),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_959),
.Y(n_961)
);

INVx4_ASAP7_75t_L g962 ( 
.A(n_955),
.Y(n_962)
);

OAI31xp33_ASAP7_75t_L g963 ( 
.A1(n_958),
.A2(n_819),
.A3(n_679),
.B(n_826),
.Y(n_963)
);

AO22x2_ASAP7_75t_L g964 ( 
.A1(n_956),
.A2(n_814),
.B1(n_855),
.B2(n_818),
.Y(n_964)
);

OAI221xp5_ASAP7_75t_SL g965 ( 
.A1(n_963),
.A2(n_677),
.B1(n_850),
.B2(n_828),
.C(n_817),
.Y(n_965)
);

AOI22xp33_ASAP7_75t_L g966 ( 
.A1(n_961),
.A2(n_855),
.B1(n_792),
.B2(n_810),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_960),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_967),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_965),
.Y(n_969)
);

NAND3xp33_ASAP7_75t_L g970 ( 
.A(n_968),
.B(n_962),
.C(n_966),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_969),
.B(n_964),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_971),
.A2(n_737),
.B1(n_792),
.B2(n_861),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_SL g973 ( 
.A1(n_970),
.A2(n_818),
.B1(n_861),
.B2(n_827),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_L g974 ( 
.A1(n_972),
.A2(n_883),
.B1(n_871),
.B2(n_810),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_974),
.A2(n_973),
.B1(n_833),
.B2(n_838),
.Y(n_975)
);


endmodule