module real_jpeg_14243_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g125 ( 
.A(n_0),
.Y(n_125)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_2),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_3),
.A2(n_67),
.B1(n_68),
.B2(n_102),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_3),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_3),
.A2(n_64),
.B(n_67),
.C(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_3),
.B(n_89),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_3),
.B(n_47),
.Y(n_174)
);

AOI21xp33_ASAP7_75t_SL g189 ( 
.A1(n_3),
.A2(n_47),
.B(n_174),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_3),
.B(n_31),
.C(n_36),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_102),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_3),
.A2(n_123),
.B1(n_124),
.B2(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_3),
.B(n_50),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_5),
.A2(n_47),
.B1(n_48),
.B2(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_5),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_5),
.A2(n_67),
.B1(n_68),
.B2(n_109),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_109),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_109),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_6),
.A2(n_67),
.B1(n_68),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_6),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_6),
.A2(n_35),
.B1(n_36),
.B2(n_72),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_72),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_6),
.A2(n_47),
.B1(n_48),
.B2(n_72),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_7),
.A2(n_67),
.B1(n_68),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_7),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_7),
.A2(n_47),
.B1(n_48),
.B2(n_74),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_74),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_74),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_8),
.A2(n_41),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_41),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_8),
.A2(n_41),
.B1(n_67),
.B2(n_68),
.Y(n_280)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_11),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_11),
.A2(n_59),
.B1(n_67),
.B2(n_68),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_59),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_11),
.A2(n_35),
.B1(n_36),
.B2(n_59),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_13),
.A2(n_67),
.B1(n_68),
.B2(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_13),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_13),
.A2(n_47),
.B1(n_48),
.B2(n_105),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_105),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_105),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_14),
.A2(n_47),
.B1(n_48),
.B2(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_14),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_111),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_14),
.A2(n_35),
.B1(n_36),
.B2(n_111),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_14),
.A2(n_67),
.B1(n_68),
.B2(n_111),
.Y(n_255)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_93),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_91),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_85),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_19),
.B(n_85),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_75),
.C(n_79),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_20),
.A2(n_75),
.B1(n_310),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_20),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_60),
.B2(n_61),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_42),
.B2(n_43),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_23),
.B(n_75),
.C(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_23),
.A2(n_24),
.B1(n_80),
.B2(n_81),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_24),
.B(n_42),
.C(n_60),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_34),
.B(n_39),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_25),
.A2(n_39),
.B(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_25),
.A2(n_167),
.B(n_169),
.Y(n_166)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_26),
.B(n_115),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_26),
.A2(n_116),
.B1(n_168),
.B2(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_26),
.A2(n_116),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_26),
.A2(n_116),
.B1(n_191),
.B2(n_201),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_26),
.A2(n_116),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_26),
.A2(n_248),
.B(n_270),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_34),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_28),
.A2(n_29),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

NAND3xp33_ASAP7_75t_SL g175 ( 
.A(n_28),
.B(n_48),
.C(n_52),
.Y(n_175)
);

INVx5_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_29),
.A2(n_53),
.B(n_173),
.C(n_175),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_29),
.B(n_198),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_34),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_34),
.A2(n_150),
.B(n_151),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_34),
.B(n_102),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_35),
.B(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_36),
.B(n_124),
.Y(n_123)
);

BUFx4f_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_40),
.B(n_116),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_54),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_44),
.A2(n_56),
.B(n_110),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_50),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_45),
.A2(n_50),
.B(n_55),
.Y(n_86)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_46),
.A2(n_56),
.B(n_84),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_47),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_48),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g130 ( 
.A1(n_47),
.A2(n_65),
.B(n_102),
.Y(n_130)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_50),
.B(n_58),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_50),
.A2(n_55),
.B1(n_83),
.B2(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_51),
.A2(n_56),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_51),
.A2(n_56),
.B1(n_108),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_51),
.A2(n_56),
.B1(n_139),
.B2(n_189),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_51),
.A2(n_54),
.B(n_277),
.Y(n_276)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_82),
.B(n_84),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_71),
.B2(n_73),
.Y(n_61)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_62),
.A2(n_73),
.B(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_62),
.A2(n_63),
.B1(n_104),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_62),
.A2(n_63),
.B1(n_144),
.B2(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_62),
.A2(n_255),
.B(n_279),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_62),
.A2(n_88),
.B(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_71),
.B(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_64),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_64),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_75),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_75),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_77),
.A2(n_89),
.B1(n_101),
.B2(n_103),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_89),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_79),
.B(n_313),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx24_ASAP7_75t_SL g323 ( 
.A(n_85),
.Y(n_323)
);

FAx1_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_87),
.CI(n_90),
.CON(n_85),
.SN(n_85)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_89),
.B(n_280),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_304),
.B(n_318),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_285),
.B(n_303),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_260),
.B(n_284),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_157),
.B(n_238),
.C(n_259),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_140),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_98),
.B(n_140),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_118),
.C(n_131),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_99),
.B(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_106),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_100),
.B(n_112),
.C(n_117),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_102),
.B(n_124),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_112),
.B1(n_113),
.B2(n_117),
.Y(n_106)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_114),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_118),
.A2(n_119),
.B1(n_131),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_128),
.B2(n_129),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_128),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_122),
.A2(n_155),
.B(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_122),
.A2(n_125),
.B1(n_203),
.B2(n_205),
.Y(n_202)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_123),
.A2(n_153),
.B(n_154),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_123),
.A2(n_124),
.B1(n_204),
.B2(n_212),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_123),
.A2(n_206),
.B(n_222),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_123),
.A2(n_124),
.B(n_267),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_135),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_125),
.A2(n_126),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_125),
.B(n_178),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_131),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_136),
.C(n_138),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_133),
.B1(n_136),
.B2(n_137),
.Y(n_165)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_134),
.B(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_138),
.B(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_147),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_141),
.B(n_148),
.C(n_156),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_143),
.B(n_145),
.C(n_146),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_156),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_149),
.B(n_152),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_150),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_151),
.B(n_169),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_236),
.B(n_237),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_179),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_160),
.B(n_163),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.C(n_170),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_166),
.A2(n_170),
.B1(n_171),
.B2(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_176),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_172),
.A2(n_176),
.B1(n_177),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_178),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_192),
.B(n_235),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_181),
.B(n_184),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.C(n_190),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_187),
.A2(n_188),
.B1(n_190),
.B2(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_229),
.B(n_234),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_218),
.B(n_228),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_207),
.B(n_217),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_202),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_202),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_199),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_213),
.B(n_216),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_215),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_220),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_224),
.C(n_227),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_222),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_226),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_233),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_233),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_258),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_258),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_242),
.C(n_250),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_250),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_246),
.B2(n_249),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_249),
.Y(n_273)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_246),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_253),
.C(n_257),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_256),
.B2(n_257),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_256),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_262),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_283),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_271),
.B1(n_281),
.B2(n_282),
.Y(n_263)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_264),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_264),
.B(n_282),
.C(n_283),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_265),
.A2(n_266),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_266),
.B(n_268),
.Y(n_296)
);

AOI21xp33_ASAP7_75t_L g311 ( 
.A1(n_266),
.A2(n_296),
.B(n_298),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_271),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_276),
.C(n_278),
.Y(n_288)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_278),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_277),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_280),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_302),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_302),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_289),
.B2(n_301),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_287),
.B(n_290),
.C(n_295),
.Y(n_316)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_289),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_295),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_293),
.B(n_294),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_291),
.B(n_293),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_307),
.C(n_311),
.Y(n_306)
);

FAx1_ASAP7_75t_SL g317 ( 
.A(n_294),
.B(n_307),
.CI(n_311),
.CON(n_317),
.SN(n_317)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_315),
.Y(n_304)
);

AOI21xp33_ASAP7_75t_L g318 ( 
.A1(n_305),
.A2(n_319),
.B(n_320),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_312),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_312),
.Y(n_320)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_317),
.Y(n_319)
);

BUFx24_ASAP7_75t_SL g322 ( 
.A(n_317),
.Y(n_322)
);


endmodule