module fake_jpeg_11106_n_437 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_437);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_437;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx5p33_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_12),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_54),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_18),
.B(n_15),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_55),
.B(n_74),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_56),
.Y(n_139)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_57),
.Y(n_132)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_58),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_59),
.Y(n_125)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_61),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

BUFx4f_ASAP7_75t_SL g63 ( 
.A(n_19),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_63),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_64),
.Y(n_140)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_13),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_66),
.B(n_69),
.Y(n_119)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_68),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_12),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_70),
.Y(n_173)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_73),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_19),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_42),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_75),
.B(n_103),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_38),
.B(n_0),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_76),
.B(n_113),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_18),
.A2(n_12),
.B(n_10),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_102),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_28),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_78),
.A2(n_22),
.B1(n_51),
.B2(n_41),
.Y(n_117)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_81),
.Y(n_150)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_82),
.Y(n_167)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_84),
.Y(n_178)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_17),
.Y(n_85)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

BUFx4f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_86),
.Y(n_180)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_87),
.Y(n_156)
);

INVx6_ASAP7_75t_SL g88 ( 
.A(n_29),
.Y(n_88)
);

INVx6_ASAP7_75t_SL g131 ( 
.A(n_88),
.Y(n_131)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

BUFx10_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_17),
.Y(n_92)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_92),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_30),
.B(n_10),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_93),
.B(n_99),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_96),
.Y(n_185)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_97),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_36),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_98),
.A2(n_76),
.B1(n_19),
.B2(n_20),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_30),
.B(n_0),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_100),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_101),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_25),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_104),
.B(n_105),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_25),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_28),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_106),
.B(n_110),
.Y(n_152)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_31),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_107),
.B(n_108),
.Y(n_168)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_35),
.Y(n_108)
);

BUFx8_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx6_ASAP7_75t_SL g136 ( 
.A(n_109),
.Y(n_136)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_39),
.Y(n_111)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_111),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_37),
.B(n_1),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_112),
.B(n_8),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_39),
.Y(n_113)
);

AND2x4_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_33),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_114),
.B(n_125),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_102),
.A2(n_48),
.B1(n_41),
.B2(n_33),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_115),
.A2(n_117),
.B1(n_123),
.B2(n_133),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_116),
.B(n_163),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_37),
.B1(n_50),
.B2(n_46),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_118),
.A2(n_145),
.B1(n_159),
.B2(n_182),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_48),
.B1(n_27),
.B2(n_35),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_103),
.A2(n_27),
.B1(n_40),
.B2(n_52),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_40),
.B1(n_51),
.B2(n_22),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_137),
.A2(n_133),
.B1(n_146),
.B2(n_181),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_99),
.A2(n_46),
.B1(n_50),
.B2(n_52),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_90),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_146),
.A2(n_177),
.B1(n_136),
.B2(n_131),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_4),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_153),
.B(n_160),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_66),
.A2(n_8),
.B1(n_69),
.B2(n_78),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_62),
.B(n_8),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_63),
.A2(n_8),
.B(n_109),
.C(n_86),
.Y(n_162)
);

AOI21xp33_ASAP7_75t_L g202 ( 
.A1(n_162),
.A2(n_169),
.B(n_184),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_64),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_73),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_164),
.B(n_166),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_84),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_94),
.B(n_95),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_172),
.B(n_174),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_101),
.B(n_55),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_55),
.B(n_74),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_175),
.B(n_116),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_88),
.A2(n_19),
.B1(n_53),
.B2(n_44),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_93),
.B(n_99),
.Y(n_184)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_186),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_188),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_121),
.A2(n_134),
.B1(n_119),
.B2(n_162),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_189),
.A2(n_191),
.B1(n_238),
.B2(n_212),
.Y(n_280)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_120),
.Y(n_190)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_190),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_121),
.A2(n_183),
.B1(n_151),
.B2(n_170),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_168),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_192),
.B(n_229),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_114),
.B(n_148),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_193),
.B(n_217),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_195),
.Y(n_255)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_132),
.Y(n_197)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_197),
.Y(n_246)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_144),
.Y(n_198)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_198),
.Y(n_258)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_147),
.Y(n_200)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_200),
.Y(n_261)
);

XNOR2x1_ASAP7_75t_SL g201 ( 
.A(n_114),
.B(n_117),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_201),
.B(n_207),
.C(n_216),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_141),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_203),
.B(n_230),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_205),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_157),
.A2(n_170),
.B1(n_180),
.B2(n_149),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_206),
.A2(n_208),
.B1(n_210),
.B2(n_212),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_152),
.A2(n_114),
.B(n_137),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_157),
.A2(n_149),
.B1(n_120),
.B2(n_130),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_209),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_130),
.A2(n_177),
.B1(n_171),
.B2(n_125),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_126),
.Y(n_211)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_211),
.Y(n_274)
);

OA22x2_ASAP7_75t_L g212 ( 
.A1(n_123),
.A2(n_122),
.B1(n_176),
.B2(n_115),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_126),
.Y(n_213)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_213),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_214),
.B(n_221),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_129),
.A2(n_143),
.B1(n_140),
.B2(n_167),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_215),
.A2(n_232),
.B1(n_187),
.B2(n_204),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_161),
.B(n_155),
.C(n_124),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_154),
.B(n_138),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_127),
.B(n_150),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_218),
.B(n_219),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_128),
.B(n_185),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_141),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_220),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_139),
.Y(n_222)
);

INVx13_ASAP7_75t_L g223 ( 
.A(n_141),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_223),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_156),
.B(n_158),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_224),
.B(n_226),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_142),
.B(n_173),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_142),
.Y(n_227)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_227),
.Y(n_285)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_173),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_228),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_167),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_135),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_135),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_231),
.B(n_220),
.Y(n_270)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_129),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_232),
.B(n_237),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_171),
.B(n_179),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_234),
.B(n_239),
.C(n_198),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_140),
.A2(n_143),
.B1(n_179),
.B2(n_139),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_235),
.A2(n_242),
.B1(n_244),
.B2(n_245),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_139),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_236),
.B(n_240),
.Y(n_281)
);

INVx4_ASAP7_75t_SL g237 ( 
.A(n_131),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_117),
.A2(n_133),
.B1(n_162),
.B2(n_177),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_114),
.B(n_134),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_168),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_134),
.A2(n_117),
.B1(n_98),
.B2(n_137),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_243),
.B(n_217),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_182),
.A2(n_19),
.B1(n_53),
.B2(n_44),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_182),
.A2(n_19),
.B1(n_53),
.B2(n_44),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_248),
.A2(n_251),
.B1(n_264),
.B2(n_269),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_189),
.A2(n_196),
.B1(n_201),
.B2(n_242),
.Y(n_251)
);

AOI32xp33_ASAP7_75t_L g254 ( 
.A1(n_193),
.A2(n_202),
.A3(n_194),
.B1(n_239),
.B2(n_221),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_254),
.B(n_190),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_221),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_260),
.B(n_276),
.C(n_234),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_263),
.B(n_265),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_241),
.B(n_199),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_196),
.A2(n_191),
.B1(n_207),
.B2(n_225),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_268),
.B(n_283),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_282),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_218),
.B(n_224),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_216),
.B(n_219),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_286),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_284),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_233),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_214),
.A2(n_212),
.B1(n_215),
.B2(n_226),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_197),
.B(n_200),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_246),
.Y(n_288)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_288),
.Y(n_324)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_246),
.Y(n_289)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_289),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_290),
.B(n_279),
.C(n_255),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_286),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_291),
.B(n_298),
.Y(n_327)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_266),
.Y(n_292)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_292),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_252),
.A2(n_212),
.B(n_234),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_294),
.A2(n_305),
.B(n_312),
.Y(n_341)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_266),
.Y(n_295)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_295),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_227),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_296),
.B(n_311),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_271),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_256),
.A2(n_186),
.B1(n_229),
.B2(n_205),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_299),
.A2(n_304),
.B1(n_315),
.B2(n_316),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_211),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_300),
.B(n_303),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_302),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_257),
.B(n_213),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_277),
.A2(n_209),
.B1(n_222),
.B2(n_228),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_256),
.A2(n_251),
.B(n_252),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_278),
.B(n_223),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_306),
.B(n_307),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_262),
.B(n_257),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_274),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_308),
.Y(n_320)
);

INVx5_ASAP7_75t_L g309 ( 
.A(n_253),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_309),
.B(n_314),
.Y(n_337)
);

AO22x1_ASAP7_75t_SL g311 ( 
.A1(n_252),
.A2(n_272),
.B1(n_276),
.B2(n_267),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_273),
.A2(n_247),
.B(n_260),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_258),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_313),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_271),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_267),
.A2(n_273),
.B1(n_249),
.B2(n_284),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_276),
.A2(n_248),
.B1(n_261),
.B2(n_258),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_271),
.B(n_275),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_317),
.B(n_318),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_261),
.B(n_285),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_319),
.A2(n_269),
.B1(n_274),
.B2(n_250),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_318),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_321),
.B(n_333),
.Y(n_355)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_317),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_323),
.B(n_330),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_312),
.A2(n_259),
.B(n_264),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_328),
.A2(n_314),
.B(n_315),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_294),
.B(n_298),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_329),
.A2(n_291),
.B(n_290),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_293),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_296),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_335),
.B(n_338),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_304),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_340),
.B(n_301),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_316),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_342),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_287),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_343),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_332),
.B(n_301),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_346),
.B(n_311),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_347),
.A2(n_341),
.B(n_328),
.Y(n_374)
);

XNOR2x2_ASAP7_75t_L g348 ( 
.A(n_332),
.B(n_287),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_SL g384 ( 
.A(n_348),
.B(n_329),
.C(n_311),
.Y(n_384)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_324),
.Y(n_349)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_349),
.Y(n_371)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_324),
.Y(n_350)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_350),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_353),
.Y(n_370)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_325),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_354),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_327),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_356),
.B(n_357),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_327),
.B(n_303),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_358),
.B(n_305),
.Y(n_375)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_325),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_359),
.B(n_362),
.Y(n_372)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_339),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_339),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_363),
.Y(n_383)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_326),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_364),
.A2(n_365),
.B1(n_336),
.B2(n_320),
.Y(n_369)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_326),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_337),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_366),
.B(n_356),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_360),
.A2(n_342),
.B1(n_334),
.B2(n_330),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_367),
.A2(n_368),
.B1(n_369),
.B2(n_352),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_360),
.A2(n_338),
.B1(n_335),
.B2(n_343),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_361),
.A2(n_297),
.B1(n_345),
.B2(n_341),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_373),
.A2(n_377),
.B1(n_352),
.B2(n_351),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_374),
.B(n_353),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_375),
.B(n_340),
.C(n_366),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_376),
.B(n_379),
.Y(n_386)
);

O2A1O1Ixp33_ASAP7_75t_L g377 ( 
.A1(n_361),
.A2(n_329),
.B(n_323),
.C(n_337),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_347),
.A2(n_329),
.B(n_351),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_382),
.B(n_358),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_384),
.B(n_346),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_385),
.B(n_387),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_388),
.B(n_389),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_381),
.B(n_331),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_390),
.A2(n_394),
.B1(n_368),
.B2(n_355),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_391),
.B(n_367),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_381),
.B(n_331),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_392),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_393),
.B(n_395),
.C(n_396),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_373),
.A2(n_333),
.B1(n_344),
.B2(n_321),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_375),
.B(n_299),
.C(n_311),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_370),
.B(n_348),
.C(n_345),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_382),
.B(n_348),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_397),
.B(n_398),
.C(n_374),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_357),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_403),
.B(n_388),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_404),
.B(n_405),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_396),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_406),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_395),
.A2(n_370),
.B1(n_302),
.B2(n_379),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_407),
.A2(n_408),
.B1(n_386),
.B2(n_393),
.Y(n_409)
);

FAx1_ASAP7_75t_SL g408 ( 
.A(n_397),
.B(n_377),
.CI(n_322),
.CON(n_408),
.SN(n_408)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_409),
.B(n_410),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_401),
.B(n_385),
.C(n_398),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_411),
.B(n_412),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_401),
.B(n_387),
.C(n_378),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_399),
.A2(n_297),
.B1(n_378),
.B2(n_369),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_414),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_406),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_415),
.A2(n_403),
.B1(n_383),
.B2(n_380),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_413),
.A2(n_399),
.B1(n_407),
.B2(n_402),
.Y(n_418)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_418),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_416),
.B(n_310),
.Y(n_419)
);

NAND3xp33_ASAP7_75t_L g428 ( 
.A(n_419),
.B(n_344),
.C(n_322),
.Y(n_428)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_420),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_411),
.B(n_400),
.C(n_364),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_422),
.B(n_420),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_417),
.A2(n_415),
.B(n_413),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_425),
.B(n_422),
.C(n_421),
.Y(n_429)
);

NOR2xp67_ASAP7_75t_SL g431 ( 
.A(n_426),
.B(n_410),
.Y(n_431)
);

AOI31xp67_ASAP7_75t_L g430 ( 
.A1(n_428),
.A2(n_423),
.A3(n_408),
.B(n_421),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_429),
.B(n_430),
.C(n_372),
.Y(n_433)
);

A2O1A1O1Ixp25_ASAP7_75t_L g432 ( 
.A1(n_431),
.A2(n_424),
.B(n_427),
.C(n_408),
.D(n_400),
.Y(n_432)
);

BUFx24_ASAP7_75t_SL g434 ( 
.A(n_432),
.Y(n_434)
);

OAI321xp33_ASAP7_75t_L g435 ( 
.A1(n_434),
.A2(n_433),
.A3(n_371),
.B1(n_380),
.B2(n_362),
.C(n_363),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_435),
.B(n_371),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_436),
.B(n_349),
.Y(n_437)
);


endmodule