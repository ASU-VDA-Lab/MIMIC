module fake_jpeg_8360_n_278 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_278);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_278;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_23),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_23),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_44),
.Y(n_56)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_42),
.Y(n_46)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_27),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_29),
.Y(n_58)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_17),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_26),
.B1(n_31),
.B2(n_34),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_67),
.B1(n_42),
.B2(n_44),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_32),
.B(n_21),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_50),
.A2(n_30),
.B(n_21),
.C(n_17),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_35),
.C(n_33),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_33),
.C(n_25),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_32),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_38),
.A2(n_26),
.B1(n_34),
.B2(n_18),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_63),
.B1(n_65),
.B2(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_24),
.Y(n_60)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_29),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_66),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_19),
.B1(n_20),
.B2(n_35),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_32),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_22),
.Y(n_69)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_74),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_42),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_75),
.B(n_80),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_65),
.B(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_78),
.B(n_84),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_62),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_83),
.Y(n_122)
);

INVx6_ASAP7_75t_SL g83 ( 
.A(n_68),
.Y(n_83)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_44),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_91),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_32),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_56),
.B(n_40),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_93),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_56),
.B(n_40),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_98),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_40),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_43),
.Y(n_121)
);

AND2x4_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_43),
.Y(n_97)
);

FAx1_ASAP7_75t_SL g111 ( 
.A(n_97),
.B(n_99),
.CI(n_30),
.CON(n_111),
.SN(n_111)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_39),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_16),
.C(n_15),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_39),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_54),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_53),
.A2(n_39),
.B1(n_30),
.B2(n_21),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_70),
.B1(n_28),
.B2(n_2),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_105),
.A2(n_80),
.B1(n_97),
.B2(n_76),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_97),
.A2(n_88),
.B1(n_94),
.B2(n_105),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_107),
.A2(n_114),
.B1(n_125),
.B2(n_130),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_129),
.B1(n_89),
.B2(n_103),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_111),
.B(n_1),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_96),
.C(n_97),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_81),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_74),
.A2(n_47),
.B1(n_53),
.B2(n_70),
.Y(n_114)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_120),
.B(n_126),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_123),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_74),
.B(n_43),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_71),
.B(n_0),
.Y(n_126)
);

NOR2x1_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_28),
.Y(n_128)
);

AO21x1_ASAP7_75t_L g149 ( 
.A1(n_128),
.A2(n_82),
.B(n_3),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_72),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_89),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_122),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_133),
.B(n_136),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_135),
.B(n_155),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_122),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_128),
.A2(n_86),
.B1(n_77),
.B2(n_95),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_149),
.B(n_106),
.Y(n_165)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_142),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_109),
.A2(n_87),
.B1(n_90),
.B2(n_100),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_141),
.A2(n_127),
.B1(n_117),
.B2(n_110),
.Y(n_181)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_101),
.B1(n_79),
.B2(n_90),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_143),
.A2(n_152),
.B1(n_127),
.B2(n_118),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_87),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_147),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_145),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_119),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_153),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_100),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_101),
.B(n_3),
.C(n_5),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_161),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_150),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_151),
.A2(n_129),
.B(n_106),
.Y(n_166)
);

AO22x2_ASAP7_75t_L g152 ( 
.A1(n_115),
.A2(n_82),
.B1(n_73),
.B2(n_79),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_156),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_131),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_5),
.Y(n_157)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_157),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_132),
.B(n_108),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_158),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_108),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_165),
.A2(n_173),
.B(n_176),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_166),
.B(n_169),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_140),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_175),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_147),
.A2(n_115),
.B(n_132),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_134),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_134),
.A2(n_124),
.B(n_110),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_SL g201 ( 
.A1(n_177),
.A2(n_149),
.B(n_137),
.C(n_154),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_152),
.A2(n_124),
.B(n_110),
.Y(n_179)
);

OAI22x1_ASAP7_75t_L g192 ( 
.A1(n_179),
.A2(n_152),
.B1(n_135),
.B2(n_148),
.Y(n_192)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_137),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_171),
.B1(n_172),
.B2(n_186),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_150),
.A2(n_111),
.B1(n_117),
.B2(n_7),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_182),
.A2(n_187),
.B1(n_5),
.B2(n_6),
.Y(n_202)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_143),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_186),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_142),
.A2(n_111),
.B1(n_6),
.B2(n_7),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_188),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_190),
.B(n_191),
.Y(n_225)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_192),
.A2(n_197),
.B(n_201),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_139),
.Y(n_194)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_187),
.A2(n_167),
.B(n_162),
.C(n_182),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_202),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_155),
.C(n_144),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_200),
.C(n_210),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_181),
.A2(n_145),
.B1(n_160),
.B2(n_161),
.Y(n_198)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

MAJx2_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_138),
.C(n_153),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_179),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_143),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_208),
.Y(n_212)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_8),
.Y(n_206)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_206),
.Y(n_216)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_164),
.Y(n_207)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_167),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_9),
.C(n_11),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_192),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_173),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_221),
.C(n_223),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_177),
.C(n_184),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_224),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_166),
.C(n_170),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_209),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_185),
.Y(n_227)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_227),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_237),
.C(n_239),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_163),
.Y(n_229)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_221),
.A2(n_189),
.B(n_197),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_231),
.A2(n_240),
.B(n_226),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_218),
.B(n_204),
.Y(n_232)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_168),
.Y(n_233)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_220),
.A2(n_198),
.B1(n_195),
.B2(n_172),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_236),
.A2(n_215),
.B1(n_222),
.B2(n_213),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_199),
.C(n_210),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_218),
.B(n_202),
.Y(n_238)
);

BUFx24_ASAP7_75t_SL g246 ( 
.A(n_238),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_189),
.C(n_165),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_201),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_211),
.C(n_217),
.Y(n_250)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_244),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_231),
.A2(n_215),
.B1(n_213),
.B2(n_220),
.Y(n_245)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_248),
.B(n_235),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_230),
.A2(n_214),
.B1(n_227),
.B2(n_226),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_249),
.A2(n_234),
.B(n_239),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_235),
.C(n_237),
.Y(n_258)
);

OAI21x1_ASAP7_75t_L g252 ( 
.A1(n_241),
.A2(n_201),
.B(n_168),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_228),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_253),
.A2(n_259),
.B(n_242),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_11),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_244),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_250),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_260),
.C(n_9),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_216),
.C(n_201),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_257),
.A2(n_251),
.B1(n_245),
.B2(n_243),
.Y(n_261)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_261),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_262),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_264),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_255),
.A2(n_247),
.B1(n_253),
.B2(n_246),
.Y(n_264)
);

BUFx24_ASAP7_75t_SL g267 ( 
.A(n_265),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_260),
.B(n_266),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_272),
.Y(n_274)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_269),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_268),
.A2(n_266),
.B(n_261),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_273),
.Y(n_275)
);

AOI321xp33_ASAP7_75t_L g276 ( 
.A1(n_274),
.A2(n_12),
.A3(n_14),
.B1(n_267),
.B2(n_270),
.C(n_271),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_276),
.B(n_275),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_12),
.Y(n_278)
);


endmodule