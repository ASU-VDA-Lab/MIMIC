module fake_jpeg_8589_n_230 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_230);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx8_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

AOI21xp33_ASAP7_75t_L g17 ( 
.A1(n_2),
.A2(n_1),
.B(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_29),
.B(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_26),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_36),
.B(n_39),
.Y(n_54)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_45),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_23),
.B(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_22),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_32),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_23),
.B1(n_33),
.B2(n_25),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_56),
.B1(n_64),
.B2(n_69),
.Y(n_82)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_47),
.Y(n_74)
);

AO21x1_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_17),
.B(n_43),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_49),
.A2(n_19),
.B1(n_28),
.B2(n_30),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_50),
.B(n_51),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_34),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_57),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_25),
.B1(n_33),
.B2(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_35),
.Y(n_72)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_24),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_63),
.A2(n_19),
.B(n_28),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_29),
.B1(n_24),
.B2(n_26),
.Y(n_64)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_42),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g102 ( 
.A(n_66),
.Y(n_102)
);

CKINVDCx12_ASAP7_75t_R g67 ( 
.A(n_42),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_67),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_27),
.Y(n_83)
);

AO22x1_ASAP7_75t_SL g69 ( 
.A1(n_37),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_20),
.Y(n_70)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_76),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

OR2x2_ASAP7_75t_SL g76 ( 
.A(n_65),
.B(n_32),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_20),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_78),
.A2(n_81),
.B(n_84),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_37),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_83),
.Y(n_103)
);

OR2x4_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_16),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_27),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_45),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_66),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_89),
.Y(n_111)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_54),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_91),
.B(n_97),
.Y(n_112)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_92),
.A2(n_58),
.B1(n_47),
.B2(n_62),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_69),
.A2(n_31),
.B1(n_27),
.B2(n_21),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_93),
.A2(n_101),
.B1(n_69),
.B2(n_58),
.Y(n_107)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_99),
.Y(n_119)
);

OR2x2_ASAP7_75t_SL g97 ( 
.A(n_61),
.B(n_19),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_64),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_0),
.Y(n_121)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_109),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_113),
.B1(n_114),
.B2(n_124),
.Y(n_134)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

AO22x1_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_56),
.B1(n_63),
.B2(n_57),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_120),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_52),
.B1(n_48),
.B2(n_59),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_82),
.A2(n_63),
.B1(n_59),
.B2(n_31),
.Y(n_114)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_117),
.B(n_121),
.Y(n_138)
);

AO22x1_ASAP7_75t_L g120 ( 
.A1(n_79),
.A2(n_30),
.B1(n_28),
.B2(n_45),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_127),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_101),
.A2(n_93),
.B1(n_97),
.B2(n_72),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_78),
.B(n_71),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_125),
.B(n_98),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_80),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_126),
.A2(n_76),
.B1(n_90),
.B2(n_75),
.Y(n_137)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_3),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_133),
.B(n_139),
.Y(n_155)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_148),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_137),
.A2(n_146),
.B1(n_106),
.B2(n_122),
.Y(n_160)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_141),
.B(n_143),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_45),
.B(n_102),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_142),
.A2(n_144),
.B(n_108),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_112),
.B(n_116),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_45),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_114),
.A2(n_92),
.B1(n_88),
.B2(n_45),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_SL g147 ( 
.A1(n_130),
.A2(n_1),
.B(n_3),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_147),
.B(n_137),
.Y(n_171)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_103),
.B(n_86),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_77),
.C(n_118),
.Y(n_165)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_10),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_153),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_116),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_132),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_159),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_148),
.A2(n_110),
.B1(n_129),
.B2(n_122),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_158),
.A2(n_161),
.B(n_166),
.Y(n_174)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_168),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_118),
.B1(n_108),
.B2(n_127),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_149),
.C(n_145),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_136),
.A2(n_146),
.B1(n_134),
.B2(n_142),
.Y(n_167)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_167),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_131),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_170),
.Y(n_183)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_154),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_138),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_154),
.Y(n_186)
);

OA21x2_ASAP7_75t_L g173 ( 
.A1(n_134),
.A2(n_4),
.B(n_5),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_153),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_182),
.C(n_188),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_178),
.A2(n_169),
.B1(n_158),
.B2(n_163),
.Y(n_190)
);

NOR3xp33_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_143),
.C(n_145),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_185),
.Y(n_191)
);

OAI21xp33_ASAP7_75t_L g180 ( 
.A1(n_166),
.A2(n_139),
.B(n_133),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_180),
.B(n_155),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_144),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_159),
.Y(n_194)
);

NOR3xp33_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_144),
.C(n_141),
.Y(n_185)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_186),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_4),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_135),
.C(n_150),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_183),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_197),
.Y(n_208)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

AO21x1_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_182),
.B(n_176),
.Y(n_210)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_194),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_157),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_195),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_177),
.A2(n_161),
.B1(n_173),
.B2(n_157),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_173),
.B1(n_170),
.B2(n_150),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_198),
.A2(n_188),
.B1(n_180),
.B2(n_189),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_200),
.C(n_178),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_5),
.Y(n_200)
);

INVxp33_ASAP7_75t_L g203 ( 
.A(n_198),
.Y(n_203)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_203),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_174),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_205),
.C(n_207),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_181),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_200),
.Y(n_216)
);

NOR2xp67_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_192),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_203),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_211),
.B(n_212),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_206),
.A2(n_192),
.B(n_199),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_209),
.C(n_206),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_216),
.Y(n_219)
);

NOR2x1_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_202),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_218),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_220),
.A2(n_208),
.B1(n_201),
.B2(n_205),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_218),
.C(n_7),
.Y(n_225)
);

NOR3xp33_ASAP7_75t_SL g222 ( 
.A(n_219),
.B(n_210),
.C(n_208),
.Y(n_222)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_222),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_R g224 ( 
.A(n_222),
.B(n_211),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_224),
.B(n_223),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_6),
.C(n_8),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_228),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_226),
.Y(n_230)
);


endmodule