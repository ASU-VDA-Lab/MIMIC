module fake_jpeg_3193_n_213 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_213);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_213;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_4),
.B(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_30),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_48),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_11),
.B(n_6),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_17),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

BUFx8_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_22),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_15),
.B(n_7),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_20),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_81),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_57),
.Y(n_85)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

BUFx10_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_86),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_64),
.B(n_55),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_89),
.A2(n_83),
.B(n_67),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_67),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_63),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_64),
.B1(n_65),
.B2(n_69),
.Y(n_91)
);

AO21x1_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_83),
.B(n_75),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_82),
.A2(n_69),
.B1(n_52),
.B2(n_62),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_92),
.A2(n_94),
.B1(n_65),
.B2(n_71),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_81),
.B(n_51),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_96),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_62),
.B1(n_60),
.B2(n_71),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_68),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_70),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_72),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_65),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_109),
.Y(n_136)
);

AND2x6_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_28),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_26),
.Y(n_123)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_97),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_108),
.B(n_110),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_111),
.B(n_114),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_87),
.Y(n_112)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_53),
.C(n_61),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_113),
.B(n_118),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_1),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_24),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_128),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_84),
.B(n_87),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_126),
.A2(n_31),
.B(n_47),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_98),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_102),
.A2(n_98),
.B1(n_88),
.B2(n_84),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_129),
.A2(n_109),
.B1(n_101),
.B2(n_59),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_88),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_137),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_1),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_134),
.B(n_138),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_2),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_105),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_139),
.B(n_106),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_140),
.B(n_145),
.Y(n_167)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_143),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_117),
.C(n_116),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_149),
.C(n_155),
.Y(n_164)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_144),
.A2(n_154),
.B1(n_135),
.B2(n_122),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_2),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_119),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_124),
.B(n_3),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_147),
.B(n_151),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_137),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_153),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_61),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

NOR3xp33_ASAP7_75t_SL g151 ( 
.A(n_135),
.B(n_59),
.C(n_61),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_136),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_29),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_157),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_25),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_12),
.Y(n_177)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_161),
.B(n_162),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_126),
.Y(n_162)
);

AO21x1_ASAP7_75t_L g169 ( 
.A1(n_163),
.A2(n_132),
.B(n_23),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_166),
.Y(n_191)
);

OAI22x1_ASAP7_75t_L g166 ( 
.A1(n_160),
.A2(n_136),
.B1(n_32),
.B2(n_34),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_174),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_136),
.B(n_50),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_170),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_142),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_172),
.A2(n_178),
.B1(n_182),
.B2(n_159),
.Y(n_187)
);

AOI221xp5_ASAP7_75t_L g174 ( 
.A1(n_149),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.C(n_12),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_146),
.A2(n_36),
.B(n_44),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_177),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_152),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_178)
);

AO21x1_ASAP7_75t_L g179 ( 
.A1(n_151),
.A2(n_38),
.B(n_42),
.Y(n_179)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_179),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_158),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_187),
.B(n_188),
.Y(n_194)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_180),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_39),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_192),
.C(n_175),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_41),
.C(n_46),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_183),
.A2(n_13),
.B1(n_16),
.B2(n_17),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_193),
.A2(n_178),
.B1(n_172),
.B2(n_177),
.Y(n_199)
);

AO22x2_ASAP7_75t_L g195 ( 
.A1(n_188),
.A2(n_181),
.B1(n_166),
.B2(n_176),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_198),
.Y(n_201)
);

XNOR2x1_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_170),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_197),
.C(n_192),
.Y(n_204)
);

BUFx24_ASAP7_75t_SL g198 ( 
.A(n_186),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_199),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_190),
.B1(n_184),
.B2(n_167),
.Y(n_200)
);

INVxp33_ASAP7_75t_L g205 ( 
.A(n_200),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_194),
.A2(n_168),
.B(n_173),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_202),
.A2(n_185),
.B1(n_195),
.B2(n_171),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_204),
.B(n_169),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_207),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_205),
.B(n_195),
.Y(n_208)
);

AOI322xp5_ASAP7_75t_L g209 ( 
.A1(n_208),
.A2(n_203),
.A3(n_201),
.B1(n_179),
.B2(n_182),
.C1(n_18),
.C2(n_16),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_209),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_211),
.A2(n_210),
.B(n_208),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_18),
.Y(n_213)
);


endmodule