module real_jpeg_30695_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_0),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_0),
.Y(n_170)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_0),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_1),
.B(n_474),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_1),
.B(n_473),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_2),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_2),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_2),
.A2(n_99),
.B1(n_221),
.B2(n_224),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_2),
.A2(n_99),
.B1(n_384),
.B2(n_385),
.Y(n_383)
);

OAI22xp33_ASAP7_75t_SL g429 ( 
.A1(n_2),
.A2(n_99),
.B1(n_430),
.B2(n_432),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_3),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_3),
.Y(n_206)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_5),
.Y(n_126)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_5),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_5),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_6),
.A2(n_152),
.B1(n_155),
.B2(n_156),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_6),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_6),
.A2(n_155),
.B1(n_242),
.B2(n_245),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_6),
.A2(n_155),
.B1(n_340),
.B2(n_344),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_7),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_7),
.Y(n_61)
);

OAI22x1_ASAP7_75t_SL g131 ( 
.A1(n_7),
.A2(n_61),
.B1(n_132),
.B2(n_135),
.Y(n_131)
);

AO22x1_ASAP7_75t_SL g235 ( 
.A1(n_7),
.A2(n_61),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

NAND2xp33_ASAP7_75t_SL g376 ( 
.A(n_7),
.B(n_377),
.Y(n_376)
);

OAI32xp33_ASAP7_75t_L g409 ( 
.A1(n_7),
.A2(n_410),
.A3(n_412),
.B1(n_414),
.B2(n_419),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_7),
.B(n_26),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_8),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_8),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_9),
.Y(n_83)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_10),
.Y(n_114)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_10),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_11),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_11),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_12),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_12),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_12),
.A2(n_74),
.B1(n_143),
.B2(n_147),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_12),
.A2(n_74),
.B1(n_172),
.B2(n_176),
.Y(n_171)
);

AO22x2_ASAP7_75t_L g253 ( 
.A1(n_12),
.A2(n_74),
.B1(n_201),
.B2(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_13),
.Y(n_474)
);

OAI31xp33_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_473),
.A3(n_475),
.B(n_492),
.Y(n_14)
);

AOI31xp33_ASAP7_75t_L g492 ( 
.A1(n_15),
.A2(n_475),
.A3(n_493),
.B(n_494),
.Y(n_492)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_358),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_326),
.Y(n_17)
);

NAND3xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_285),
.C(n_303),
.Y(n_18)
);

AOI21xp33_ASAP7_75t_L g326 ( 
.A1(n_19),
.A2(n_327),
.B(n_328),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_248),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_20),
.B(n_248),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_179),
.C(n_230),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_22),
.B(n_230),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_104),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_66),
.Y(n_23)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_24),
.Y(n_282)
);

AOI21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_39),
.B(n_56),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_26),
.B(n_229),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_26),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_26),
.B(n_220),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_26),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AO21x2_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_40),
.B(n_47),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B1(n_36),
.B2(n_38),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_29),
.Y(n_244)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_30),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_30),
.Y(n_149)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_36),
.Y(n_384)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_37),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_37),
.Y(n_139)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_39),
.Y(n_219)
);

NOR2x1_ASAP7_75t_L g257 ( 
.A(n_39),
.B(n_56),
.Y(n_257)
);

INVxp33_ASAP7_75t_L g375 ( 
.A(n_40),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_44),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_42),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_43),
.Y(n_256)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_52),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_50),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g227 ( 
.A(n_51),
.Y(n_227)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_56),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_61),
.B(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_61),
.A2(n_204),
.B(n_261),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_61),
.B(n_215),
.Y(n_318)
);

AOI32xp33_ASAP7_75t_L g369 ( 
.A1(n_61),
.A2(n_370),
.A3(n_373),
.B1(n_375),
.B2(n_376),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_61),
.B(n_415),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_R g450 ( 
.A(n_61),
.B(n_120),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_61),
.B(n_208),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVxp67_ASAP7_75t_SL g283 ( 
.A(n_66),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_95),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_77),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_68),
.B(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_72),
.Y(n_196)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_73),
.Y(n_263)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_77),
.B(n_96),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_77),
.B(n_260),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_77),
.A2(n_260),
.B(n_354),
.Y(n_353)
);

NOR2x1p5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_88),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_81),
.B1(n_84),
.B2(n_86),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_83),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_83),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_85),
.Y(n_84)
);

AO22x2_ASAP7_75t_L g88 ( 
.A1(n_86),
.A2(n_89),
.B1(n_91),
.B2(n_93),
.Y(n_88)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_88),
.B(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_88),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_88),
.Y(n_354)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_95),
.B(n_299),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

MAJx2_ASAP7_75t_L g281 ( 
.A(n_104),
.B(n_282),
.C(n_283),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_150),
.Y(n_104)
);

XOR2x2_ASAP7_75t_L g292 ( 
.A(n_105),
.B(n_150),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_140),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_106),
.B(n_397),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_131),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_107),
.B(n_142),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_107),
.Y(n_271)
);

OA21x2_ASAP7_75t_L g300 ( 
.A1(n_107),
.A2(n_131),
.B(n_141),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_107),
.B(n_383),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_120),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_112),
.B1(n_115),
.B2(n_118),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_117),
.Y(n_379)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_117),
.Y(n_387)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_124),
.B1(n_127),
.B2(n_128),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_123),
.Y(n_422)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_126),
.Y(n_236)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_130),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_130),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_130),
.Y(n_418)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_130),
.Y(n_431)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_130),
.Y(n_435)
);

NAND2xp33_ASAP7_75t_SL g336 ( 
.A(n_131),
.B(n_141),
.Y(n_336)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_140),
.A2(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_140),
.B(n_382),
.Y(n_440)
);

NAND2x1_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_141),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_141),
.B(n_383),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_143),
.B(n_420),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_146),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_149),
.Y(n_246)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_149),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_160),
.B(n_167),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_SL g207 ( 
.A1(n_151),
.A2(n_208),
.B(n_209),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_154),
.Y(n_456)
);

BUFx2_ASAP7_75t_SL g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_159),
.Y(n_166)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

AOI21x1_ASAP7_75t_L g273 ( 
.A1(n_160),
.A2(n_274),
.B(n_278),
.Y(n_273)
);

NAND2x1_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_164),
.Y(n_234)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_167),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_167),
.B(n_428),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_169),
.Y(n_446)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx4_ASAP7_75t_SL g208 ( 
.A(n_170),
.Y(n_208)
);

NAND2xp33_ASAP7_75t_SL g209 ( 
.A(n_171),
.B(n_210),
.Y(n_209)
);

AOI21xp33_ASAP7_75t_SL g231 ( 
.A1(n_171),
.A2(n_210),
.B(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_175),
.Y(n_411)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_179),
.B(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_211),
.C(n_216),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_181),
.B(n_289),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_207),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_182),
.B(n_314),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_193),
.B(n_197),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_189),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_188),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_201),
.B(n_203),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx5_ASAP7_75t_L g344 ( 
.A(n_201),
.Y(n_344)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_207),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_209),
.B(n_444),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_210),
.B(n_235),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_210),
.B(n_429),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_211),
.A2(n_217),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_211),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_212),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_213),
.B(n_299),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_214),
.B(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVxp33_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_228),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_218),
.B(n_228),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_218),
.B(n_317),
.Y(n_316)
);

NAND2xp67_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2x1p5_ASAP7_75t_L g297 ( 
.A(n_219),
.B(n_253),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_219),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_239),
.Y(n_230)
);

AOI21xp33_ASAP7_75t_L g266 ( 
.A1(n_231),
.A2(n_240),
.B(n_247),
.Y(n_266)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_232),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_235),
.Y(n_278)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_247),
.Y(n_239)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_247),
.B(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_247),
.B(n_397),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_267),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_249),
.B(n_268),
.C(n_280),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_266),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_258),
.B1(n_264),
.B2(n_265),
.Y(n_250)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_251),
.Y(n_265)
);

NOR2x1_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_257),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_252),
.Y(n_317)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_257),
.Y(n_401)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_258),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_258),
.B(n_265),
.C(n_266),
.Y(n_332)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_280),
.B1(n_281),
.B2(n_284),
.Y(n_267)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_272),
.B1(n_273),
.B2(n_279),
.Y(n_268)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_269),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_269),
.B(n_273),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_272),
.B(n_353),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_272),
.A2(n_273),
.B1(n_368),
.B2(n_369),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_272),
.A2(n_355),
.B(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_273),
.B(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_301),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_301),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_292),
.C(n_293),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_287),
.A2(n_288),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_292),
.B(n_294),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

MAJx2_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_298),
.C(n_300),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_295),
.A2(n_300),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_295),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_296),
.B(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_297),
.Y(n_346)
);

NAND3xp33_ASAP7_75t_SL g347 ( 
.A(n_297),
.B(n_335),
.C(n_348),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_300),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_304),
.B(n_471),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_323),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_306),
.B(n_323),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_312),
.C(n_315),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_307),
.B(n_389),
.Y(n_388)
);

XNOR2x1_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_311),
.B(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_313),
.B(n_315),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_318),
.C(n_319),
.Y(n_315)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_316),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_317),
.A2(n_339),
.B(n_484),
.Y(n_483)
);

XNOR2x1_ASAP7_75t_L g365 ( 
.A(n_318),
.B(n_320),
.Y(n_365)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NOR2x1_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_321),
.Y(n_454)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NOR3xp33_ASAP7_75t_L g469 ( 
.A(n_327),
.B(n_328),
.C(n_470),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_329),
.B(n_330),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_333),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_R g488 ( 
.A(n_332),
.B(n_357),
.C(n_489),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_349),
.B1(n_356),
.B2(n_357),
.Y(n_333)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_334),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_337),
.B(n_347),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_336),
.B(n_382),
.Y(n_381)
);

AOI21xp33_ASAP7_75t_R g337 ( 
.A1(n_338),
.A2(n_345),
.B(n_346),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_338),
.B(n_345),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_347),
.Y(n_485)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_349),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_349),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_351),
.B1(n_352),
.B2(n_355),
.Y(n_349)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_350),
.Y(n_355)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_353),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_469),
.B(n_472),
.Y(n_358)
);

OAI21x1_ASAP7_75t_SL g359 ( 
.A1(n_360),
.A2(n_390),
.B(n_468),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_388),
.Y(n_361)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_362),
.B(n_388),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_367),
.C(n_380),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_364),
.B(n_393),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_367),
.B(n_381),
.Y(n_393)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_381),
.Y(n_380)
);

INVx4_ASAP7_75t_SL g385 ( 
.A(n_386),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

OA21x2_ASAP7_75t_L g390 ( 
.A1(n_391),
.A2(n_404),
.B(n_467),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_394),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_392),
.B(n_394),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_398),
.C(n_402),
.Y(n_394)
);

OAI22xp33_ASAP7_75t_SL g465 ( 
.A1(n_395),
.A2(n_396),
.B1(n_399),
.B2(n_400),
.Y(n_465)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_403),
.B(n_465),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_461),
.B(n_466),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_441),
.B(n_460),
.Y(n_405)
);

NOR2xp67_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_425),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_407),
.B(n_425),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_423),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_408),
.A2(n_409),
.B1(n_423),
.B2(n_424),
.Y(n_447)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

BUFx2_ASAP7_75t_SL g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_436),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_426),
.Y(n_463)
);

AND2x4_ASAP7_75t_SL g426 ( 
.A(n_427),
.B(n_428),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_429),
.B(n_445),
.Y(n_444)
);

BUFx4f_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_437),
.A2(n_438),
.B1(n_439),
.B2(n_440),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_437),
.B(n_440),
.C(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_442),
.A2(n_448),
.B(n_459),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_447),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_443),
.B(n_447),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_444),
.B(n_454),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_446),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_449),
.A2(n_452),
.B(n_458),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_450),
.B(n_451),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_453),
.B(n_455),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_457),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_464),
.Y(n_461)
);

NOR2xp67_ASAP7_75t_L g466 ( 
.A(n_462),
.B(n_464),
.Y(n_466)
);

INVxp33_ASAP7_75t_L g493 ( 
.A(n_473),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_490),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_488),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_478),
.B(n_488),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_486),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_485),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_482),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);


endmodule