module fake_jpeg_24836_n_288 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_288);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_45;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_5),
.B(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_SL g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_9),
.B(n_0),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_28),
.B(n_32),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_15),
.B(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_28),
.A2(n_13),
.B1(n_26),
.B2(n_25),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_39),
.A2(n_44),
.B1(n_20),
.B2(n_17),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_27),
.Y(n_60)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_28),
.A2(n_13),
.B1(n_26),
.B2(n_25),
.Y(n_44)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_50),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_26),
.B1(n_25),
.B2(n_21),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_51),
.A2(n_52),
.B1(n_21),
.B2(n_20),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_17),
.B1(n_22),
.B2(n_21),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_57),
.B1(n_62),
.B2(n_69),
.Y(n_85)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_32),
.Y(n_77)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_63),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_27),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_65),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_27),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_74),
.A2(n_53),
.B1(n_17),
.B2(n_22),
.Y(n_91)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_0),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_48),
.B1(n_53),
.B2(n_41),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_91),
.B1(n_43),
.B2(n_68),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_35),
.C(n_54),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_59),
.C(n_69),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_67),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_87),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_71),
.B(n_15),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_90),
.Y(n_110)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_95),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_66),
.A2(n_53),
.B1(n_43),
.B2(n_40),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_94),
.A2(n_57),
.B1(n_68),
.B2(n_58),
.Y(n_116)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_48),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_65),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_100),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_77),
.B(n_64),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_102),
.C(n_112),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_67),
.C(n_59),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_73),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_104),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_88),
.B(n_98),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_105),
.A2(n_40),
.B1(n_46),
.B2(n_42),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_83),
.A2(n_98),
.B(n_97),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_109),
.B(n_93),
.Y(n_134)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_113),
.Y(n_125)
);

NAND2xp33_ASAP7_75t_SL g109 ( 
.A(n_88),
.B(n_86),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_85),
.A2(n_97),
.B(n_87),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_104),
.B(n_101),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_33),
.C(n_38),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_33),
.C(n_38),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_93),
.C(n_81),
.Y(n_129)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_118),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_116),
.A2(n_61),
.B1(n_40),
.B2(n_72),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_18),
.Y(n_133)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_81),
.Y(n_137)
);

NAND2xp33_ASAP7_75t_SL g123 ( 
.A(n_109),
.B(n_72),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_123),
.A2(n_76),
.B1(n_75),
.B2(n_63),
.Y(n_156)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_127),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_126),
.A2(n_100),
.B(n_117),
.Y(n_148)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_144),
.C(n_30),
.Y(n_153)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_131),
.Y(n_168)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_61),
.B1(n_58),
.B2(n_72),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_141),
.B1(n_145),
.B2(n_18),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_134),
.Y(n_162)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_138),
.B(n_142),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_108),
.A2(n_113),
.B1(n_105),
.B2(n_99),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_117),
.B1(n_42),
.B2(n_118),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_82),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_84),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_18),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_33),
.C(n_49),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

AOI22x1_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_106),
.B1(n_114),
.B2(n_112),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_SL g189 ( 
.A1(n_147),
.A2(n_165),
.B(n_135),
.C(n_14),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_148),
.A2(n_136),
.B(n_133),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_154),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_143),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_150),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_120),
.B1(n_84),
.B2(n_106),
.Y(n_151)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_159),
.C(n_164),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_129),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_125),
.A2(n_92),
.B1(n_45),
.B2(n_30),
.Y(n_157)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_131),
.B(n_22),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_158),
.B(n_137),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_45),
.C(n_20),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_130),
.A2(n_45),
.B1(n_23),
.B2(n_16),
.Y(n_161)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_170),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_23),
.C(n_16),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_169),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_126),
.A2(n_23),
.B1(n_16),
.B2(n_14),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_167),
.A2(n_138),
.B1(n_127),
.B2(n_124),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_123),
.A2(n_18),
.B1(n_16),
.B2(n_14),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_23),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_140),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_173),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_163),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_144),
.C(n_134),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_157),
.C(n_156),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_178),
.A2(n_189),
.B1(n_191),
.B2(n_0),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_155),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_2),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_152),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_181),
.A2(n_183),
.B(n_192),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_148),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_186),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_168),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_187),
.B(n_160),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_147),
.A2(n_136),
.B1(n_135),
.B2(n_14),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_147),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_12),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_164),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_182),
.B(n_149),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_194),
.B(n_208),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_161),
.Y(n_197)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_212),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_192),
.A2(n_154),
.B(n_166),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_200),
.A2(n_188),
.B(n_171),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_201),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_171),
.A2(n_151),
.B1(n_167),
.B2(n_159),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_202),
.A2(n_191),
.B1(n_178),
.B2(n_189),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_210),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_206),
.C(n_207),
.Y(n_222)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_169),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_174),
.C(n_175),
.Y(n_207)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_184),
.B(n_1),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_1),
.C(n_2),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_211),
.A2(n_185),
.B(n_173),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_1),
.Y(n_212)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_218),
.A2(n_206),
.B(n_211),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_219),
.A2(n_11),
.B1(n_4),
.B2(n_5),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_172),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_227),
.Y(n_240)
);

FAx1_ASAP7_75t_SL g225 ( 
.A(n_200),
.B(n_172),
.CI(n_179),
.CON(n_225),
.SN(n_225)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_225),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_198),
.A2(n_179),
.B(n_190),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_226),
.A2(n_202),
.B(n_195),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_190),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_11),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_212),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_224),
.B(n_208),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_229),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_204),
.C(n_199),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_242),
.C(n_243),
.Y(n_255)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_237),
.B(n_238),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_221),
.A2(n_208),
.B(n_4),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_239),
.A2(n_217),
.B1(n_230),
.B2(n_8),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_3),
.C(n_4),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_3),
.C(n_5),
.Y(n_243)
);

AO21x1_ASAP7_75t_L g244 ( 
.A1(n_223),
.A2(n_3),
.B(n_6),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_231),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_218),
.A2(n_3),
.B(n_6),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_245),
.A2(n_6),
.B(n_7),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_225),
.Y(n_247)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_247),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_246),
.A2(n_228),
.B1(n_224),
.B2(n_227),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_248),
.A2(n_233),
.B1(n_240),
.B2(n_9),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_225),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_249),
.B(n_250),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_253),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_243),
.B(n_214),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_257),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_214),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_258),
.A2(n_259),
.B(n_238),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_6),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_269),
.Y(n_273)
);

AOI211xp5_ASAP7_75t_L g261 ( 
.A1(n_256),
.A2(n_237),
.B(n_232),
.C(n_248),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_7),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_256),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_263),
.B(n_7),
.Y(n_275)
);

AOI21x1_ASAP7_75t_L g266 ( 
.A1(n_255),
.A2(n_250),
.B(n_242),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_267),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_240),
.C(n_8),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_264),
.B(n_252),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_271),
.B(n_276),
.Y(n_277)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_261),
.Y(n_272)
);

AOI21x1_ASAP7_75t_SL g278 ( 
.A1(n_272),
.A2(n_263),
.B(n_262),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_253),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_265),
.Y(n_279)
);

O2A1O1Ixp33_ASAP7_75t_SL g281 ( 
.A1(n_275),
.A2(n_8),
.B(n_10),
.C(n_11),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_278),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_279),
.B(n_280),
.Y(n_282)
);

AOI21xp33_ASAP7_75t_L g280 ( 
.A1(n_273),
.A2(n_269),
.B(n_9),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_283),
.A2(n_277),
.B(n_275),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_284),
.A2(n_282),
.B(n_281),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g286 ( 
.A(n_285),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_270),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_10),
.Y(n_288)
);


endmodule