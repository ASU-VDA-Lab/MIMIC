module fake_jpeg_25824_n_179 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_2),
.B(n_6),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_36),
.Y(n_46)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_20),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_25),
.B1(n_37),
.B2(n_32),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_4),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_5),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_40),
.B(n_36),
.Y(n_45)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_18),
.B(n_29),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_19),
.B(n_24),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_45),
.B(n_50),
.Y(n_77)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_26),
.C(n_19),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_26),
.C(n_34),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_54),
.B1(n_25),
.B2(n_15),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_19),
.Y(n_50)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_15),
.B1(n_25),
.B2(n_28),
.Y(n_54)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_34),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_39),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_68),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_59),
.A2(n_75),
.B1(n_42),
.B2(n_33),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_45),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_60),
.B(n_62),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_22),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_66),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_53),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_64),
.B(n_67),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_22),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_39),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_53),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_69),
.B(n_71),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_70),
.B(n_76),
.Y(n_83)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_42),
.A2(n_15),
.B1(n_25),
.B2(n_28),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_26),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_46),
.B(n_30),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_80),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_33),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_26),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_27),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_5),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_82),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_72),
.C(n_71),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_94),
.B1(n_82),
.B2(n_73),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_91),
.B(n_100),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_56),
.B1(n_51),
.B2(n_52),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_30),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_99),
.B(n_101),
.Y(n_107)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_100),
.B(n_96),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_27),
.Y(n_101)
);

AND2x4_ASAP7_75t_L g103 ( 
.A(n_57),
.B(n_56),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_103),
.A2(n_79),
.B1(n_82),
.B2(n_67),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_102),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_104),
.B(n_105),
.Y(n_126)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_106),
.B(n_109),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_116),
.B1(n_117),
.B2(n_51),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_83),
.B(n_77),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_113),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_83),
.B(n_64),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_114),
.Y(n_124)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_81),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_119),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_95),
.A2(n_59),
.B1(n_70),
.B2(n_69),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_87),
.C(n_103),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_63),
.Y(n_119)
);

NAND3xp33_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_84),
.C(n_103),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_24),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

NOR3xp33_ASAP7_75t_SL g147 ( 
.A(n_123),
.B(n_136),
.C(n_129),
.Y(n_147)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_133),
.C(n_110),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_118),
.A2(n_95),
.B(n_103),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_131),
.A2(n_135),
.B(n_120),
.Y(n_141)
);

AOI32xp33_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_103),
.A3(n_104),
.B1(n_116),
.B2(n_84),
.Y(n_132)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_132),
.A2(n_134),
.B(n_51),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_92),
.C(n_86),
.Y(n_133)
);

OAI31xp33_ASAP7_75t_L g134 ( 
.A1(n_106),
.A2(n_89),
.A3(n_92),
.B(n_93),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_86),
.B(n_62),
.Y(n_135)
);

BUFx12_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_139),
.Y(n_155)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_145),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_142),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_126),
.Y(n_143)
);

NOR3xp33_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_144),
.C(n_124),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_125),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_107),
.C(n_74),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_133),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_131),
.A2(n_80),
.B(n_112),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_148),
.A2(n_149),
.B1(n_135),
.B2(n_137),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_147),
.B(n_137),
.C(n_127),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_150),
.A2(n_148),
.B(n_146),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_152),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_146),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_145),
.B(n_122),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_17),
.B(n_29),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_141),
.A2(n_122),
.B1(n_132),
.B2(n_112),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g159 ( 
.A(n_158),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_161),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_142),
.C(n_139),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_139),
.C(n_138),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_164),
.C(n_154),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_165),
.A2(n_150),
.B1(n_17),
.B2(n_23),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_168),
.C(n_11),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_153),
.B1(n_155),
.B2(n_90),
.Y(n_169)
);

AOI322xp5_ASAP7_75t_L g171 ( 
.A1(n_169),
.A2(n_159),
.A3(n_160),
.B1(n_90),
.B2(n_74),
.C1(n_21),
.C2(n_5),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_18),
.B(n_23),
.C(n_12),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_170),
.A2(n_166),
.B(n_10),
.C(n_9),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_SL g175 ( 
.A1(n_171),
.A2(n_173),
.B(n_174),
.C(n_6),
.Y(n_175)
);

AOI322xp5_ASAP7_75t_L g172 ( 
.A1(n_169),
.A2(n_11),
.A3(n_14),
.B1(n_13),
.B2(n_9),
.C1(n_10),
.C2(n_74),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_172),
.A2(n_7),
.B(n_8),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_175),
.A2(n_176),
.B1(n_7),
.B2(n_21),
.Y(n_178)
);

INVxp33_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_178),
.Y(n_179)
);


endmodule