module real_jpeg_6735_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_1),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_1),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_1),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_2),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_2),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_2),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_2),
.B(n_310),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_2),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_2),
.B(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_2),
.B(n_436),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_3),
.Y(n_506)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_4),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_4),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_4),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_4),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g141 ( 
.A(n_4),
.B(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_4),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_4),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_4),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_5),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_5),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_5),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_5),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_5),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_5),
.B(n_79),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_5),
.B(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_5),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_6),
.B(n_52),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_6),
.A2(n_46),
.B(n_285),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_6),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_6),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_6),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_6),
.B(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_6),
.B(n_433),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_6),
.B(n_416),
.Y(n_443)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_8),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_8),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_8),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_8),
.B(n_202),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_8),
.B(n_244),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_8),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_8),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_8),
.B(n_353),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_9),
.Y(n_155)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_9),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_9),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_9),
.Y(n_353)
);

BUFx5_ASAP7_75t_L g416 ( 
.A(n_9),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_10),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_10),
.B(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_10),
.B(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_10),
.B(n_407),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_10),
.B(n_426),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_10),
.B(n_405),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_10),
.B(n_440),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_11),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g347 ( 
.A(n_11),
.Y(n_347)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_13),
.B(n_161),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_13),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_13),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_13),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_13),
.B(n_306),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_13),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_13),
.B(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_13),
.B(n_457),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_14),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_14),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_14),
.Y(n_281)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_15),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_16),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_16),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_16),
.Y(n_405)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_16),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_17),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_17),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_17),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_17),
.B(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g125 ( 
.A(n_17),
.B(n_126),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g154 ( 
.A(n_17),
.B(n_155),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_501),
.B(n_503),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_113),
.Y(n_19)
);

OAI21xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_73),
.B(n_112),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_21),
.B(n_73),
.Y(n_112)
);

BUFx24_ASAP7_75t_SL g509 ( 
.A(n_21),
.Y(n_509)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_62),
.CI(n_63),
.CON(n_21),
.SN(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_48),
.C(n_53),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_23),
.A2(n_24),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_42),
.B2(n_43),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_35),
.B2(n_36),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_27),
.B(n_54),
.C(n_57),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_27),
.A2(n_28),
.B1(n_54),
.B2(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_27),
.A2(n_28),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_28),
.B(n_35),
.C(n_43),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_28),
.B(n_236),
.C(n_242),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_29),
.B(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_33),
.Y(n_407)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_34),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_34),
.Y(n_277)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_34),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_35),
.A2(n_36),
.B1(n_66),
.B2(n_68),
.Y(n_65)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_36),
.B(n_187),
.C(n_188),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_36),
.B(n_233),
.Y(n_232)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_40),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_40),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_40),
.Y(n_267)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_41),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_42),
.A2(n_43),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_43),
.B(n_141),
.C(n_145),
.Y(n_170)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_47),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_48),
.A2(n_49),
.B1(n_53),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_51),
.Y(n_189)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_53),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_69),
.C(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_54),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_54),
.A2(n_106),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_54),
.A2(n_106),
.B1(n_263),
.B2(n_264),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_56),
.Y(n_135)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_56),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_56),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_57),
.A2(n_58),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_57),
.A2(n_58),
.B1(n_132),
.B2(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_58),
.B(n_130),
.C(n_132),
.Y(n_131)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_69),
.B2(n_72),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_66),
.Y(n_68)
);

MAJx2_ASAP7_75t_L g196 ( 
.A(n_66),
.B(n_197),
.C(n_201),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_66),
.A2(n_68),
.B1(n_162),
.B2(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_66),
.A2(n_68),
.B1(n_201),
.B2(n_251),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_68),
.B(n_152),
.C(n_162),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_69),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_69),
.A2(n_72),
.B1(n_77),
.B2(n_78),
.Y(n_169)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_107),
.C(n_108),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_74),
.B(n_499),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_91),
.C(n_103),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_75),
.B(n_173),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_81),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_87),
.C(n_89),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_77),
.A2(n_78),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_77),
.B(n_123),
.C(n_130),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_77),
.A2(n_78),
.B1(n_309),
.B2(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_78),
.B(n_305),
.C(n_309),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_80),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_82),
.Y(n_89)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_86),
.Y(n_248)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_86),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_87),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_91),
.B(n_103),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.C(n_101),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_92),
.A2(n_96),
.B1(n_97),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_96),
.A2(n_97),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_97),
.B(n_154),
.C(n_198),
.Y(n_197)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_100),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_101),
.B(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_106),
.B(n_263),
.C(n_268),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_107),
.B(n_108),
.Y(n_499)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AO21x1_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_496),
.B(n_500),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_253),
.B(n_493),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_210),
.Y(n_115)
);

AOI21xp33_ASAP7_75t_SL g493 ( 
.A1(n_116),
.A2(n_494),
.B(n_495),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_174),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_117),
.B(n_174),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_165),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_118),
.B(n_166),
.C(n_172),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_147),
.C(n_150),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_119),
.B(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_131),
.C(n_136),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_120),
.B(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_125),
.B1(n_129),
.B2(n_130),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_123),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_125),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_125),
.A2(n_130),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_125),
.B(n_237),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_125),
.A2(n_130),
.B1(n_236),
.B2(n_237),
.Y(n_461)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_128),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_131),
.B(n_136),
.Y(n_215)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_132),
.Y(n_185)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_134),
.Y(n_244)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

INVx6_ASAP7_75t_L g378 ( 
.A(n_135),
.Y(n_378)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_141),
.B1(n_145),
.B2(n_146),
.Y(n_138)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_141),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_141),
.B(n_224),
.Y(n_261)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_146),
.B(n_223),
.C(n_228),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_147),
.A2(n_150),
.B1(n_151),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OA22x2_ASAP7_75t_L g206 ( 
.A1(n_152),
.A2(n_153),
.B1(n_207),
.B2(n_209),
.Y(n_206)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.C(n_160),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_154),
.A2(n_160),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_154),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_154),
.A2(n_192),
.B1(n_198),
.B2(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_154),
.A2(n_192),
.B1(n_418),
.B2(n_420),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_154),
.B(n_420),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_156),
.A2(n_191),
.B1(n_194),
.B2(n_195),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_156),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_156),
.B(n_275),
.C(n_278),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_156),
.A2(n_194),
.B1(n_275),
.B2(n_342),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_160),
.Y(n_193)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_172),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.C(n_171),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_171),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.C(n_180),
.Y(n_174)
);

FAx1_ASAP7_75t_SL g252 ( 
.A(n_175),
.B(n_178),
.CI(n_180),
.CON(n_252),
.SN(n_252)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_196),
.C(n_206),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_213),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_186),
.C(n_190),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_182),
.B(n_186),
.Y(n_326)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_187),
.B(n_188),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_190),
.B(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_191),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_206),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_197),
.B(n_250),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_198),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_198),
.B(n_313),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_198),
.A2(n_221),
.B1(n_313),
.B2(n_314),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_199),
.Y(n_412)
);

INVx8_ASAP7_75t_L g434 ( 
.A(n_199),
.Y(n_434)
);

BUFx8_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g442 ( 
.A(n_200),
.Y(n_442)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_201),
.Y(n_251)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_205),
.Y(n_310)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_207),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_252),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_211),
.B(n_252),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_214),
.C(n_216),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_212),
.B(n_214),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_216),
.B(n_333),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_234),
.C(n_249),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_217),
.B(n_328),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.C(n_232),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_218),
.Y(n_298)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_222),
.B(n_232),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_261),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_234),
.B(n_249),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_243),
.C(n_245),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_235),
.B(n_295),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_236),
.A2(n_237),
.B1(n_242),
.B2(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_241),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_242),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_243),
.A2(n_245),
.B1(n_246),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_243),
.Y(n_296)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

BUFx24_ASAP7_75t_SL g508 ( 
.A(n_252),
.Y(n_508)
);

AOI221xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_391),
.B1(n_486),
.B2(n_491),
.C(n_492),
.Y(n_253)
);

NOR3xp33_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_330),
.C(n_334),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_255),
.A2(n_487),
.B(n_490),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_323),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_256),
.B(n_323),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_297),
.C(n_300),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_257),
.B(n_297),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_282),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_258),
.B(n_283),
.C(n_294),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.C(n_273),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_260),
.B(n_274),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_262),
.B(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_268),
.B(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

BUFx5_ASAP7_75t_L g419 ( 
.A(n_272),
.Y(n_419)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_275),
.Y(n_342)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_278),
.B(n_341),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_294),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_289),
.C(n_292),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_284),
.B(n_322),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_284),
.A2(n_285),
.B(n_344),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_289),
.B(n_292),
.Y(n_322)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_291),
.B(n_345),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_300),
.B(n_363),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_317),
.C(n_321),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_301),
.B(n_338),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.C(n_311),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_302),
.B(n_387),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_304),
.A2(n_311),
.B1(n_312),
.B2(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_304),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_305),
.B(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_309),
.Y(n_371)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx6_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_317),
.B(n_321),
.Y(n_338)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_329),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_327),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_327),
.C(n_329),
.Y(n_331)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_330),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_331),
.B(n_332),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_364),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_335),
.A2(n_488),
.B(n_489),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_362),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_336),
.B(n_362),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_339),
.C(n_360),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_337),
.B(n_390),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_339),
.B(n_360),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_343),
.C(n_348),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_340),
.B(n_343),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_348),
.B(n_367),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_351),
.C(n_354),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_349),
.A2(n_350),
.B1(n_474),
.B2(n_475),
.Y(n_473)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_351),
.A2(n_352),
.B1(n_354),
.B2(n_355),
.Y(n_474)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx4_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_359),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_389),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_365),
.B(n_389),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_368),
.C(n_386),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_366),
.B(n_484),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_368),
.B(n_386),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_372),
.C(n_384),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g476 ( 
.A(n_369),
.B(n_477),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_372),
.A2(n_384),
.B1(n_385),
.B2(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_372),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_376),
.C(n_379),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_373),
.A2(n_374),
.B1(n_379),
.B2(n_380),
.Y(n_466)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_376),
.B(n_466),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_378),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_377),
.B(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_378),
.Y(n_427)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx4_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx6_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_392),
.A2(n_481),
.B(n_485),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_393),
.A2(n_468),
.B(n_480),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_394),
.A2(n_452),
.B(n_467),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_395),
.A2(n_428),
.B(n_451),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_396),
.B(n_421),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_396),
.B(n_421),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_408),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_397),
.B(n_409),
.C(n_417),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_403),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_398),
.B(n_404),
.C(n_406),
.Y(n_464)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_406),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_417),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_413),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_410),
.B(n_413),
.Y(n_422)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_415),
.Y(n_413)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_418),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.C(n_424),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_422),
.B(n_448),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_423),
.A2(n_424),
.B1(n_425),
.B2(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_423),
.Y(n_449)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_445),
.B(n_450),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_430),
.A2(n_438),
.B(n_444),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_431),
.B(n_437),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_431),
.B(n_437),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_435),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_432),
.B(n_435),
.Y(n_446)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_443),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_441),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_447),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_446),
.B(n_447),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_454),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_453),
.B(n_454),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_463),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_455),
.A2(n_471),
.B1(n_472),
.B2(n_473),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_455),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_455),
.B(n_464),
.C(n_465),
.Y(n_479)
);

FAx1_ASAP7_75t_SL g455 ( 
.A(n_456),
.B(n_461),
.CI(n_462),
.CON(n_455),
.SN(n_455)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_465),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_469),
.B(n_479),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_469),
.B(n_479),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_476),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_471),
.B(n_473),
.C(n_476),
.Y(n_482)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_474),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_483),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_482),
.B(n_483),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_498),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_497),
.B(n_498),
.Y(n_500)
);

INVx6_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx5_ASAP7_75t_L g505 ( 
.A(n_502),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_506),
.Y(n_503)
);

BUFx12f_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);


endmodule