module real_jpeg_14511_n_16 (n_5, n_4, n_8, n_0, n_12, n_409, n_410, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_409;
input n_410;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_2),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_2),
.B(n_31),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_2),
.B(n_28),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_2),
.B(n_63),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_2),
.B(n_136),
.Y(n_225)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_3),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_5),
.B(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_5),
.B(n_45),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_5),
.B(n_28),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_5),
.B(n_136),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_5),
.B(n_179),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_6),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_6),
.B(n_28),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_6),
.B(n_50),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_6),
.B(n_31),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_6),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_6),
.B(n_63),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_6),
.B(n_136),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_6),
.B(n_179),
.Y(n_209)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_7),
.B(n_45),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_7),
.B(n_50),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_7),
.B(n_31),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_7),
.B(n_35),
.Y(n_174)
);

AND2x2_ASAP7_75t_SL g192 ( 
.A(n_7),
.B(n_28),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_7),
.B(n_63),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_7),
.B(n_136),
.Y(n_263)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_7),
.Y(n_301)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_10),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_10),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_10),
.B(n_35),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_10),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_10),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_11),
.B(n_45),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_11),
.B(n_50),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_11),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_11),
.B(n_35),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_11),
.B(n_28),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_11),
.B(n_136),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_12),
.Y(n_136)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_13),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_13),
.B(n_50),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_13),
.B(n_31),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_13),
.B(n_35),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_13),
.B(n_63),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_13),
.B(n_179),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_14),
.B(n_45),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_14),
.B(n_50),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_14),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_14),
.B(n_35),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_14),
.B(n_28),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_14),
.B(n_63),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_14),
.B(n_136),
.Y(n_307)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_393),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_377),
.B(n_392),
.Y(n_17)
);

OAI321xp33_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_328),
.A3(n_352),
.B1(n_375),
.B2(n_376),
.C(n_409),
.Y(n_18)
);

AOI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_250),
.A3(n_286),
.B1(n_322),
.B2(n_327),
.C(n_410),
.Y(n_19)
);

NOR3xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_183),
.C(n_245),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_144),
.B(n_182),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_109),
.B(n_143),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_78),
.B(n_108),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_53),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_25),
.B(n_53),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_37),
.C(n_47),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_26),
.A2(n_56),
.B1(n_57),
.B2(n_67),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_26),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_26),
.B(n_105),
.Y(n_104)
);

FAx1_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_30),
.CI(n_34),
.CON(n_26),
.SN(n_26)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_29),
.B(n_168),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_32),
.B(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_32),
.B(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_32),
.B(n_201),
.Y(n_200)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_SL g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_37),
.A2(n_38),
.B1(n_47),
.B2(n_106),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_43),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_39),
.B(n_43),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_42),
.Y(n_39)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_40),
.B(n_94),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_42),
.B(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_46),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_44),
.B(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_44),
.B(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_46),
.B(n_59),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_46),
.B(n_178),
.Y(n_265)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_48),
.B(n_52),
.Y(n_69)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_51),
.A2(n_52),
.B1(n_124),
.B2(n_125),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_51),
.A2(n_52),
.B1(n_172),
.B2(n_175),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_52),
.B(n_125),
.C(n_242),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_52),
.B(n_175),
.C(n_272),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_68),
.B2(n_77),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_56),
.B(n_67),
.C(n_77),
.Y(n_110)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_60),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_58),
.B(n_61),
.C(n_66),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_63),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_65),
.Y(n_66)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_69),
.B(n_71),
.C(n_72),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_73),
.A2(n_74),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_73),
.A2(n_74),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_73),
.A2(n_74),
.B1(n_119),
.B2(n_120),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_73),
.B(n_300),
.C(n_302),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_73),
.B(n_120),
.C(n_196),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_74),
.B(n_75),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_74),
.B(n_281),
.C(n_283),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_75),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_75),
.A2(n_76),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_75),
.B(n_209),
.C(n_212),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_102),
.B(n_107),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_91),
.B(n_101),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_86),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_81),
.B(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_84),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_82),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_89),
.C(n_90),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_96),
.B(n_100),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_93),
.B(n_95),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_94),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_103),
.B(n_104),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_110),
.B(n_111),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_128),
.B2(n_129),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_130),
.C(n_142),
.Y(n_145)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_121),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_122),
.C(n_123),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_117),
.C(n_120),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_119),
.A2(n_120),
.B1(n_174),
.B2(n_176),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_120),
.B(n_174),
.C(n_226),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_126),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_141),
.B2(n_142),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_140),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_137),
.C(n_139),
.Y(n_163)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_135),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_136),
.Y(n_362)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_145),
.B(n_146),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_162),
.B2(n_181),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_151),
.B2(n_161),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_149),
.B(n_161),
.C(n_181),
.Y(n_246)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_157),
.B2(n_158),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_152),
.B(n_159),
.C(n_160),
.Y(n_205)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx24_ASAP7_75t_SL g407 ( 
.A(n_153),
.Y(n_407)
);

FAx1_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_155),
.CI(n_156),
.CON(n_153),
.SN(n_153)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_154),
.B(n_155),
.C(n_156),
.Y(n_214)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

BUFx24_ASAP7_75t_SL g408 ( 
.A(n_162),
.Y(n_408)
);

FAx1_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_164),
.CI(n_170),
.CON(n_162),
.SN(n_162)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_163),
.B(n_164),
.C(n_170),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_167),
.B(n_169),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_167),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_166),
.B(n_201),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_168),
.B(n_362),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_169),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_169),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_177),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_172),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_173),
.B(n_178),
.Y(n_339)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_174),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_175),
.C(n_177),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_174),
.A2(n_176),
.B1(n_192),
.B2(n_194),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_174),
.B(n_192),
.C(n_271),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_178),
.B(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_178),
.B(n_201),
.Y(n_364)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

AOI21xp33_ASAP7_75t_L g323 ( 
.A1(n_184),
.A2(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_218),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_185),
.B(n_218),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_206),
.C(n_217),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_186),
.B(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_205),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_197),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_188),
.B(n_197),
.C(n_205),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_195),
.B2(n_196),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_191),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_192),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_193),
.C(n_196),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_192),
.A2(n_194),
.B1(n_237),
.B2(n_238),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_194),
.B(n_237),
.C(n_307),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_195),
.A2(n_196),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_204),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_202),
.C(n_204),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_206),
.A2(n_207),
.B1(n_217),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_214),
.C(n_216),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_211),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_214),
.Y(n_215)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_217),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_244),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_231),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_231),
.C(n_244),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_228),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_221),
.B(n_229),
.C(n_230),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_222),
.B(n_225),
.C(n_226),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_226),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_226),
.A2(n_227),
.B1(n_346),
.B2(n_347),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_232),
.B(n_234),
.C(n_235),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_241),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_237),
.A2(n_238),
.B1(n_263),
.B2(n_266),
.Y(n_403)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_238),
.B(n_239),
.C(n_241),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_239),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_246),
.B(n_247),
.Y(n_324)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_251),
.A2(n_323),
.B(n_326),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_252),
.B(n_253),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_285),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_255),
.B(n_256),
.C(n_285),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_277),
.B2(n_278),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_257),
.B(n_279),
.C(n_280),
.Y(n_321)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_267),
.B2(n_268),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_259),
.B(n_269),
.C(n_276),
.Y(n_292)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_261),
.B(n_263),
.C(n_265),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_263),
.Y(n_266)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_275),
.B2(n_276),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_271),
.A2(n_272),
.B1(n_368),
.B2(n_369),
.Y(n_367)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_273),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_283),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_287),
.B(n_288),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_321),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_304),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_290),
.B(n_304),
.C(n_321),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_291),
.B(n_295),
.C(n_303),
.Y(n_351)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_303),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_298),
.B2(n_302),
.Y(n_295)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_296),
.Y(n_302)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_313),
.B2(n_314),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_305),
.B(n_315),
.C(n_320),
.Y(n_331)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_309),
.B2(n_312),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_307),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_307),
.B(n_310),
.C(n_311),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_307),
.A2(n_312),
.B1(n_384),
.B2(n_385),
.Y(n_383)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_319),
.B2(n_320),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_329),
.B(n_330),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_330),
.B(n_353),
.Y(n_376)
);

FAx1_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_332),
.CI(n_351),
.CON(n_330),
.SN(n_330)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_344),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_334),
.A2(n_335),
.B1(n_336),
.B2(n_337),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_334),
.B(n_337),
.C(n_344),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_339),
.B1(n_340),
.B2(n_343),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_338),
.A2(n_339),
.B1(n_402),
.B2(n_403),
.Y(n_401)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_339),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_339),
.B(n_341),
.C(n_342),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_340),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_345),
.B(n_348),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_345),
.B(n_349),
.C(n_350),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_347),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_374),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_356),
.B1(n_372),
.B2(n_373),
.Y(n_354)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_355),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_355),
.B(n_373),
.C(n_374),
.Y(n_378)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_356),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_357),
.B(n_365),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_357),
.B(n_366),
.C(n_371),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_358),
.B(n_361),
.C(n_363),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_360),
.A2(n_361),
.B1(n_363),
.B2(n_364),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_361),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_364),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_366),
.A2(n_367),
.B1(n_370),
.B2(n_371),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_378),
.B(n_379),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_380),
.B(n_382),
.C(n_391),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_391),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_386),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_383),
.B(n_388),
.C(n_389),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_384),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_387),
.A2(n_388),
.B1(n_389),
.B2(n_390),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_388),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_390),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_405),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_396),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_395),
.B(n_396),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_404),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_398),
.A2(n_399),
.B1(n_400),
.B2(n_401),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_399),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_401),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_403),
.Y(n_402)
);


endmodule