module fake_jpeg_21461_n_336 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_42),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_22),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_32),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx5_ASAP7_75t_SL g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g85 ( 
.A(n_48),
.Y(n_85)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_50),
.Y(n_97)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_32),
.B1(n_27),
.B2(n_17),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_51),
.A2(n_32),
.B1(n_27),
.B2(n_17),
.Y(n_75)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_25),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_56),
.B(n_67),
.Y(n_84)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_41),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_69),
.B(n_72),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_70),
.Y(n_121)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_41),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_94),
.Y(n_119)
);

BUFx2_ASAP7_75t_SL g74 ( 
.A(n_63),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_74),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_75),
.A2(n_88),
.B1(n_18),
.B2(n_23),
.Y(n_116)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_52),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_79),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_46),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_82),
.A2(n_34),
.B1(n_33),
.B2(n_28),
.Y(n_123)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_55),
.A2(n_27),
.B1(n_25),
.B2(n_18),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_89),
.Y(n_125)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_59),
.A2(n_27),
.B1(n_22),
.B2(n_30),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_24),
.B1(n_34),
.B2(n_33),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_40),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_69),
.A2(n_61),
.B1(n_60),
.B2(n_57),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_99),
.A2(n_101),
.B1(n_107),
.B2(n_110),
.Y(n_136)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_94),
.A2(n_61),
.B1(n_54),
.B2(n_60),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_95),
.A2(n_57),
.B1(n_46),
.B2(n_40),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_87),
.A2(n_91),
.B1(n_78),
.B2(n_82),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_111),
.A2(n_116),
.B1(n_120),
.B2(n_85),
.Y(n_128)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_82),
.A2(n_64),
.B1(n_30),
.B2(n_22),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

AND2x2_ASAP7_75t_SL g126 ( 
.A(n_100),
.B(n_84),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_126),
.A2(n_130),
.B(n_150),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_128),
.A2(n_155),
.B1(n_102),
.B2(n_114),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_111),
.A2(n_79),
.B(n_92),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_115),
.B(n_86),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_133),
.B(n_143),
.Y(n_168)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_138),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_105),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_76),
.C(n_90),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_104),
.C(n_106),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_30),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_141),
.B(n_142),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_24),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_121),
.B(n_89),
.Y(n_143)
);

INVxp67_ASAP7_75t_SL g144 ( 
.A(n_105),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_124),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_146),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_83),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_85),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_117),
.B(n_20),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_148),
.B(n_20),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_33),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_151),
.B(n_19),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_83),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_113),
.Y(n_167)
);

BUFx8_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_101),
.A2(n_96),
.B1(n_81),
.B2(n_80),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_103),
.B1(n_107),
.B2(n_113),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_158),
.A2(n_173),
.B1(n_134),
.B2(n_154),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_160),
.B(n_175),
.Y(n_216)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_131),
.A2(n_20),
.B(n_18),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_165),
.A2(n_170),
.B(n_184),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_176),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_172),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_139),
.A2(n_103),
.B1(n_109),
.B2(n_108),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_129),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_130),
.A2(n_102),
.B1(n_114),
.B2(n_81),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_174),
.A2(n_140),
.B1(n_155),
.B2(n_132),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_109),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_129),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_131),
.A2(n_24),
.B(n_34),
.C(n_28),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_180),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_150),
.A2(n_28),
.B(n_23),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_178),
.A2(n_182),
.B(n_187),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_127),
.B(n_80),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_179),
.Y(n_198)
);

OA21x2_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_98),
.B(n_77),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_126),
.A2(n_23),
.B(n_19),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_185),
.C(n_151),
.Y(n_196)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_126),
.B(n_29),
.C(n_19),
.Y(n_184)
);

MAJx2_ASAP7_75t_L g185 ( 
.A(n_142),
.B(n_29),
.C(n_19),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_140),
.Y(n_186)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_127),
.A2(n_26),
.B(n_29),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_132),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_31),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_160),
.A2(n_136),
.B1(n_128),
.B2(n_145),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_193),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_195),
.A2(n_200),
.B1(n_206),
.B2(n_161),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_196),
.B(n_165),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_137),
.C(n_154),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_214),
.C(n_159),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_199),
.A2(n_204),
.B1(n_162),
.B2(n_157),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_174),
.A2(n_152),
.B1(n_31),
.B2(n_21),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_180),
.A2(n_31),
.B1(n_21),
.B2(n_26),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_218),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_181),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_208),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_173),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_163),
.A2(n_31),
.B1(n_26),
.B2(n_2),
.Y(n_206)
);

AOI22x1_ASAP7_75t_L g207 ( 
.A1(n_180),
.A2(n_166),
.B1(n_170),
.B2(n_158),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_211),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_156),
.Y(n_208)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_172),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_L g213 ( 
.A1(n_168),
.A2(n_14),
.B(n_12),
.Y(n_213)
);

AOI21xp33_ASAP7_75t_L g231 ( 
.A1(n_213),
.A2(n_169),
.B(n_168),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_159),
.B(n_11),
.C(n_10),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_189),
.A2(n_10),
.B1(n_1),
.B2(n_2),
.Y(n_215)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_187),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_182),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_186),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_176),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_236),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_166),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_224),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_190),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_184),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_183),
.C(n_164),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_241),
.C(n_218),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_244),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_230),
.A2(n_234),
.B1(n_239),
.B2(n_242),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_231),
.A2(n_233),
.B1(n_210),
.B2(n_192),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_194),
.B(n_188),
.Y(n_232)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_232),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_205),
.A2(n_178),
.B(n_177),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_200),
.A2(n_161),
.B1(n_162),
.B2(n_171),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_211),
.Y(n_236)
);

OA21x2_ASAP7_75t_L g240 ( 
.A1(n_201),
.A2(n_207),
.B(n_194),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_243),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_196),
.B(n_185),
.C(n_171),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_207),
.A2(n_190),
.B1(n_201),
.B2(n_193),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_191),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_205),
.B(n_157),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_191),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_209),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_221),
.B(n_214),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_254),
.Y(n_269)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_240),
.Y(n_251)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_256),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_228),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_259),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_192),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_265),
.C(n_248),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_212),
.C(n_208),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_212),
.C(n_198),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_262),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_199),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_263),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_222),
.B(n_217),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_238),
.A2(n_204),
.B1(n_206),
.B2(n_3),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_223),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_227),
.B(n_0),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_247),
.Y(n_285)
);

XNOR2x1_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_237),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_268),
.B(n_1),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_258),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_270),
.Y(n_297)
);

INVxp33_ASAP7_75t_SL g272 ( 
.A(n_251),
.Y(n_272)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_259),
.Y(n_274)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_274),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_260),
.C(n_263),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_278),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_250),
.A2(n_235),
.B1(n_226),
.B2(n_239),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_276),
.A2(n_271),
.B1(n_272),
.B2(n_270),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_255),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_246),
.A2(n_230),
.B1(n_242),
.B2(n_226),
.Y(n_281)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_281),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_282),
.A2(n_234),
.B1(n_266),
.B2(n_265),
.Y(n_288)
);

AO22x1_ASAP7_75t_L g283 ( 
.A1(n_261),
.A2(n_232),
.B1(n_240),
.B2(n_233),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_283),
.A2(n_249),
.B(n_220),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_247),
.C(n_254),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_291),
.C(n_5),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_294),
.Y(n_300)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_286),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_290),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_298),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_276),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_283),
.C(n_280),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_0),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g295 ( 
.A(n_268),
.B(n_1),
.CI(n_3),
.CON(n_295),
.SN(n_295)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_4),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_291),
.C(n_296),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_303),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_269),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_309),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_292),
.B(n_278),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_269),
.C(n_293),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_310),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_3),
.C(n_4),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_311),
.C(n_6),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_308),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_4),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_5),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_305),
.A2(n_298),
.B(n_295),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_314),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_306),
.A2(n_295),
.B(n_7),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_317),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_311),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_307),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_7),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_302),
.C(n_300),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_323),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_318),
.A2(n_309),
.B(n_301),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_312),
.A2(n_301),
.B(n_8),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_326),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_316),
.A2(n_7),
.B(n_9),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_327),
.B(n_315),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_325),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_331),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_328),
.B(n_322),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_333),
.A2(n_320),
.B1(n_317),
.B2(n_329),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_9),
.C(n_331),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_9),
.Y(n_336)
);


endmodule