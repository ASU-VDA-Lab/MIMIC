module fake_jpeg_27600_n_89 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_89);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_89;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_24),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_35),
.B(n_37),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_42),
.B(n_4),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_SL g43 ( 
.A(n_31),
.B(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_45),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_17),
.B1(n_28),
.B2(n_27),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_44),
.B(n_3),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_31),
.B(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_3),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_5),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_47),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_48),
.A2(n_38),
.B1(n_7),
.B2(n_8),
.Y(n_69)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_53),
.Y(n_60)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_40),
.B(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_5),
.Y(n_57)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_29),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_33),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_29),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_6),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_10),
.B(n_11),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_71),
.A2(n_72),
.B1(n_73),
.B2(n_66),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_62),
.B1(n_60),
.B2(n_72),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_80),
.B(n_79),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_77),
.A2(n_76),
.B1(n_78),
.B2(n_64),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_81),
.A2(n_79),
.B1(n_64),
.B2(n_71),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_83),
.C(n_81),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_84),
.A2(n_83),
.B(n_74),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_74),
.Y(n_86)
);

INVxp33_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

AOI31xp33_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_13),
.A3(n_14),
.B(n_15),
.Y(n_88)
);

AOI221xp5_ASAP7_75t_L g89 ( 
.A1(n_88),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.C(n_22),
.Y(n_89)
);


endmodule