module fake_jpeg_4339_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_24),
.B1(n_30),
.B2(n_19),
.Y(n_52)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_47),
.B(n_11),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_24),
.B1(n_30),
.B2(n_25),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_49),
.A2(n_64),
.B1(n_32),
.B2(n_23),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_52),
.A2(n_19),
.B1(n_34),
.B2(n_51),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_26),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_59),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_30),
.B1(n_24),
.B2(n_27),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_65),
.B1(n_32),
.B2(n_23),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_26),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_26),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_67),
.Y(n_96)
);

BUFx4f_ASAP7_75t_SL g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_63),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_24),
.B1(n_20),
.B2(n_25),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_37),
.A2(n_23),
.B1(n_32),
.B2(n_27),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_25),
.C(n_20),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_80),
.Y(n_102)
);

AOI32xp33_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_36),
.A3(n_44),
.B1(n_40),
.B2(n_46),
.Y(n_72)
);

FAx1_ASAP7_75t_SL g116 ( 
.A(n_72),
.B(n_78),
.CI(n_87),
.CON(n_116),
.SN(n_116)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_74),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_75),
.A2(n_76),
.B1(n_86),
.B2(n_18),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_20),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_53),
.A2(n_40),
.B1(n_27),
.B2(n_46),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_79),
.A2(n_88),
.B1(n_97),
.B2(n_18),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_48),
.Y(n_80)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_47),
.A2(n_34),
.B1(n_36),
.B2(n_28),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_17),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_50),
.A2(n_34),
.B1(n_31),
.B2(n_28),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_50),
.A2(n_18),
.B1(n_33),
.B2(n_17),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_94),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_49),
.A2(n_44),
.B1(n_31),
.B2(n_33),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_95),
.A2(n_56),
.B1(n_68),
.B2(n_60),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_51),
.A2(n_31),
.B1(n_33),
.B2(n_17),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_99),
.Y(n_118)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_107),
.Y(n_129)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_121),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_78),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_114),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_66),
.C(n_60),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_119),
.C(n_127),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_18),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_123),
.B1(n_80),
.B2(n_94),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_66),
.C(n_58),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_91),
.A2(n_68),
.B1(n_56),
.B2(n_17),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_62),
.B1(n_70),
.B2(n_66),
.Y(n_124)
);

OAI22x1_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_80),
.B1(n_97),
.B2(n_89),
.Y(n_130)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_17),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_58),
.C(n_70),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_81),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_132),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_115),
.B1(n_124),
.B2(n_100),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_126),
.B(n_81),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_131),
.B(n_134),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_109),
.B(n_96),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_105),
.B(n_84),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_104),
.B(n_0),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_139),
.Y(n_178)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_142),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_138),
.A2(n_125),
.B1(n_122),
.B2(n_117),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_77),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_105),
.B(n_71),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_140),
.B(n_101),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_113),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_141),
.Y(n_159)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_77),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_144),
.A2(n_22),
.B(n_35),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_121),
.B(n_0),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_146),
.B(n_149),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

AND2x2_ASAP7_75t_SL g148 ( 
.A(n_119),
.B(n_58),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_148),
.A2(n_158),
.B(n_33),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_111),
.B(n_0),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_118),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_150),
.Y(n_169)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_107),
.Y(n_151)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_70),
.Y(n_152)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_17),
.Y(n_153)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_154),
.B(n_108),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_17),
.Y(n_155)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_57),
.C(n_73),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_114),
.C(n_120),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_100),
.A2(n_33),
.B(n_35),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_160),
.A2(n_174),
.B1(n_151),
.B2(n_142),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_110),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_128),
.Y(n_203)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_182),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_171),
.B(n_176),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_172),
.A2(n_130),
.B1(n_143),
.B2(n_131),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_180),
.C(n_145),
.Y(n_194)
);

AO21x2_ASAP7_75t_L g174 ( 
.A1(n_130),
.A2(n_114),
.B(n_112),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_129),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_175),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_179),
.A2(n_181),
.B(n_183),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_73),
.C(n_106),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_33),
.B(n_35),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_129),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_152),
.A2(n_33),
.B(n_57),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_133),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_133),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_139),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_188),
.Y(n_219)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_189),
.A2(n_154),
.B(n_158),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_137),
.B(n_92),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_190),
.Y(n_207)
);

AO21x1_ASAP7_75t_L g191 ( 
.A1(n_135),
.A2(n_31),
.B(n_35),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_191),
.A2(n_159),
.B1(n_169),
.B2(n_166),
.Y(n_218)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_177),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_192),
.B(n_200),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_193),
.A2(n_213),
.B(n_175),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_201),
.C(n_202),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_174),
.A2(n_135),
.B1(n_138),
.B2(n_157),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_195),
.A2(n_197),
.B1(n_208),
.B2(n_216),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_218),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_174),
.A2(n_165),
.B1(n_170),
.B2(n_160),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_143),
.B1(n_132),
.B2(n_148),
.Y(n_198)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_171),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_148),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_148),
.C(n_156),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_203),
.B(n_205),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_143),
.C(n_149),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_174),
.A2(n_146),
.B1(n_136),
.B2(n_144),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_178),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_209),
.B(n_217),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_172),
.A2(n_134),
.B1(n_150),
.B2(n_141),
.Y(n_211)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_167),
.B(n_92),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_173),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_162),
.A2(n_151),
.B1(n_142),
.B2(n_147),
.Y(n_213)
);

INVxp33_ASAP7_75t_SL g215 ( 
.A(n_162),
.Y(n_215)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_215),
.Y(n_224)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_178),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_165),
.A2(n_106),
.B1(n_147),
.B2(n_35),
.Y(n_220)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_186),
.Y(n_221)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_233),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_199),
.A2(n_179),
.B(n_181),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_230),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_210),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_238),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_198),
.B(n_164),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_183),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_242),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_168),
.Y(n_235)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_235),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_214),
.B(n_159),
.Y(n_237)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_237),
.Y(n_266)
);

OA21x2_ASAP7_75t_L g238 ( 
.A1(n_204),
.A2(n_191),
.B(n_170),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_220),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_240),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_214),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_187),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_241),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_201),
.B(n_164),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_243),
.Y(n_263)
);

OAI211xp5_ASAP7_75t_L g244 ( 
.A1(n_199),
.A2(n_169),
.B(n_193),
.C(n_196),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_244),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_211),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_246),
.A2(n_35),
.B1(n_1),
.B2(n_2),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_194),
.C(n_202),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_250),
.C(n_251),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_205),
.C(n_197),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_212),
.C(n_195),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_161),
.C(n_208),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_253),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_233),
.C(n_226),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_226),
.A2(n_207),
.B1(n_182),
.B2(n_218),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_255),
.A2(n_256),
.B1(n_229),
.B2(n_222),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_227),
.A2(n_185),
.B1(n_184),
.B2(n_188),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_223),
.B(n_189),
.C(n_187),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_267),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_232),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_168),
.C(n_22),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_269),
.B(n_272),
.Y(n_294)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_259),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_277),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_247),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_264),
.A2(n_228),
.B1(n_227),
.B2(n_243),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_262),
.B(n_236),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_281),
.C(n_251),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_241),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_274),
.Y(n_297)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_263),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_275),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_221),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_256),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_248),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_258),
.A2(n_224),
.B1(n_230),
.B2(n_228),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_231),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_255),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_22),
.C(n_8),
.Y(n_298)
);

NOR2x1_ASAP7_75t_SL g289 ( 
.A(n_283),
.B(n_238),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_288),
.C(n_291),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_250),
.C(n_249),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_289),
.A2(n_12),
.B(n_6),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_268),
.C(n_284),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_254),
.C(n_252),
.Y(n_292)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_292),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_254),
.C(n_261),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_296),
.Y(n_303)
);

OAI321xp33_ASAP7_75t_L g295 ( 
.A1(n_283),
.A2(n_238),
.A3(n_239),
.B1(n_253),
.B2(n_257),
.C(n_267),
.Y(n_295)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_7),
.C(n_16),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_1),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_285),
.A2(n_275),
.B1(n_274),
.B2(n_277),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_304),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_285),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_305),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_297),
.A2(n_8),
.B1(n_16),
.B2(n_13),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_22),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_6),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_12),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_309),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_294),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_310),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_308),
.B(n_290),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_311),
.A2(n_317),
.B(n_319),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_8),
.Y(n_313)
);

XNOR2x1_ASAP7_75t_SL g324 ( 
.A(n_313),
.B(n_2),
.Y(n_324)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_314),
.Y(n_321)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_310),
.A2(n_12),
.A3(n_9),
.B1(n_10),
.B2(n_5),
.C1(n_3),
.C2(n_4),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_304),
.C(n_305),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_9),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_312),
.A2(n_301),
.B(n_303),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_320),
.A2(n_323),
.B(n_325),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_324),
.B(n_318),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_300),
.C(n_3),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_321),
.B(n_318),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_326),
.A2(n_328),
.B(n_322),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_329),
.A2(n_300),
.B1(n_327),
.B2(n_315),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_2),
.B(n_3),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_4),
.C(n_323),
.Y(n_332)
);


endmodule