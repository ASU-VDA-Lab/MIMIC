module fake_jpeg_12212_n_437 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_437);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_437;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_56),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_21),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_57),
.B(n_70),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_26),
.A2(n_10),
.B(n_16),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_58),
.B(n_112),
.C(n_52),
.Y(n_132)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_59),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_21),
.B(n_5),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_60),
.B(n_100),
.Y(n_182)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_61),
.Y(n_168)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_62),
.Y(n_131)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_65),
.Y(n_129)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_66),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_67),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_69),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_22),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_72),
.Y(n_148)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_73),
.Y(n_136)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_22),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_78),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_77),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_29),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_80),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_81),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_82),
.Y(n_185)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_83),
.Y(n_121)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_84),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_29),
.B(n_5),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_87),
.B(n_103),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_33),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_93),
.Y(n_123)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_89),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_91),
.Y(n_162)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_92),
.Y(n_167)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx6_ASAP7_75t_SL g94 ( 
.A(n_40),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_32),
.Y(n_126)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_95),
.B(n_101),
.Y(n_143)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_96),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

INVx4_ASAP7_75t_SL g98 ( 
.A(n_49),
.Y(n_98)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_98),
.Y(n_163)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_33),
.B(n_5),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_35),
.Y(n_101)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_18),
.Y(n_102)
);

BUFx10_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_35),
.B(n_10),
.Y(n_103)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_18),
.Y(n_104)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_28),
.B(n_11),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_108),
.Y(n_150)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_106),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_25),
.Y(n_107)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_54),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_54),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_109),
.B(n_110),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_27),
.Y(n_110)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_27),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_111),
.Y(n_181)
);

NOR4xp25_ASAP7_75t_SL g112 ( 
.A(n_49),
.B(n_11),
.C(n_14),
.D(n_17),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_30),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_113),
.B(n_115),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_27),
.Y(n_114)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_37),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_59),
.A2(n_43),
.B1(n_27),
.B2(n_46),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_119),
.A2(n_120),
.B1(n_122),
.B2(n_128),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_61),
.A2(n_27),
.B1(n_23),
.B2(n_46),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_94),
.A2(n_23),
.B1(n_19),
.B2(n_45),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_126),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_110),
.A2(n_32),
.B1(n_48),
.B2(n_30),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_127),
.A2(n_49),
.B1(n_163),
.B2(n_110),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_68),
.A2(n_39),
.B1(n_48),
.B2(n_41),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_132),
.B(n_187),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_69),
.A2(n_45),
.B1(n_19),
.B2(n_41),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_138),
.A2(n_146),
.B1(n_147),
.B2(n_152),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_L g145 ( 
.A1(n_64),
.A2(n_52),
.B1(n_50),
.B2(n_47),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_145),
.A2(n_149),
.B1(n_49),
.B2(n_68),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_104),
.A2(n_39),
.B1(n_31),
.B2(n_42),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_56),
.A2(n_31),
.B1(n_47),
.B2(n_42),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_L g149 ( 
.A1(n_65),
.A2(n_67),
.B1(n_86),
.B2(n_81),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_56),
.A2(n_50),
.B1(n_1),
.B2(n_2),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_77),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_153),
.A2(n_154),
.B1(n_160),
.B2(n_169),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_89),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_102),
.A2(n_3),
.B1(n_17),
.B2(n_11),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_80),
.A2(n_82),
.B1(n_85),
.B2(n_74),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_105),
.B(n_115),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_172),
.B(n_177),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_79),
.A2(n_72),
.B1(n_115),
.B2(n_75),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_175),
.A2(n_158),
.B1(n_156),
.B2(n_164),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_97),
.A2(n_114),
.B1(n_107),
.B2(n_98),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_176),
.A2(n_169),
.B1(n_119),
.B2(n_175),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_75),
.B(n_90),
.Y(n_177)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_62),
.Y(n_183)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_111),
.Y(n_186)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_186),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_90),
.B(n_96),
.Y(n_187)
);

O2A1O1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_121),
.A2(n_83),
.B(n_147),
.C(n_126),
.Y(n_188)
);

O2A1O1Ixp33_ASAP7_75t_SL g283 ( 
.A1(n_188),
.A2(n_197),
.B(n_189),
.C(n_209),
.Y(n_283)
);

OR2x4_ASAP7_75t_L g189 ( 
.A(n_125),
.B(n_83),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_189),
.B(n_244),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_140),
.B(n_162),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_190),
.B(n_200),
.Y(n_249)
);

CKINVDCx12_ASAP7_75t_R g192 ( 
.A(n_179),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_192),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_116),
.B(n_117),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_194),
.B(n_196),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_123),
.B(n_143),
.Y(n_196)
);

O2A1O1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_170),
.A2(n_146),
.B(n_122),
.C(n_165),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_198),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_181),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_199),
.B(n_229),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_167),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_124),
.Y(n_201)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_134),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_204),
.A2(n_216),
.B1(n_246),
.B2(n_237),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_136),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_206),
.B(n_207),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_141),
.B(n_173),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_150),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_208),
.B(n_214),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_138),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_209),
.B(n_215),
.Y(n_277)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_210),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_135),
.B(n_131),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_211),
.B(n_219),
.Y(n_282)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_134),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_212),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_184),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_130),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_153),
.B(n_151),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_120),
.A2(n_160),
.B1(n_139),
.B2(n_152),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_151),
.B(n_180),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_217),
.B(n_223),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_184),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_218),
.B(n_242),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_131),
.B(n_137),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_171),
.B(n_166),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_220),
.B(n_222),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_168),
.B(n_155),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_118),
.B(n_185),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_118),
.B(n_185),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_224),
.B(n_230),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_142),
.B(n_130),
.Y(n_225)
);

XNOR2x1_ASAP7_75t_L g264 ( 
.A(n_225),
.B(n_243),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_148),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_228),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_130),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_176),
.B(n_144),
.Y(n_230)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_133),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_133),
.Y(n_232)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_232),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_156),
.A2(n_158),
.B1(n_164),
.B2(n_124),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_233),
.A2(n_242),
.B1(n_215),
.B2(n_223),
.Y(n_284)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_159),
.Y(n_234)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_129),
.Y(n_235)
);

INVx11_ASAP7_75t_L g236 ( 
.A(n_159),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_129),
.B(n_154),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_238),
.B(n_204),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_163),
.A2(n_18),
.B1(n_104),
.B2(n_89),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_239),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_179),
.Y(n_240)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_240),
.Y(n_265)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_134),
.Y(n_241)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_241),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_125),
.B(n_136),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_163),
.A2(n_18),
.B1(n_104),
.B2(n_89),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_248),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_132),
.A2(n_169),
.B1(n_153),
.B2(n_58),
.Y(n_246)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_144),
.Y(n_247)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_247),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_163),
.A2(n_18),
.B1(n_104),
.B2(n_89),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_206),
.B(n_193),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_251),
.B(n_195),
.C(n_218),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_190),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_255),
.B(n_261),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_225),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_262),
.A2(n_244),
.B1(n_203),
.B2(n_212),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_283),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_208),
.B(n_226),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_270),
.B(n_240),
.Y(n_301)
);

AND2x6_ASAP7_75t_L g271 ( 
.A(n_197),
.B(n_188),
.Y(n_271)
);

A2O1A1O1Ixp25_ASAP7_75t_L g296 ( 
.A1(n_271),
.A2(n_236),
.B(n_205),
.C(n_241),
.D(n_225),
.Y(n_296)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_217),
.Y(n_272)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_207),
.Y(n_276)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_276),
.Y(n_300)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_198),
.Y(n_279)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_279),
.Y(n_318)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_243),
.Y(n_281)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_281),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_284),
.A2(n_243),
.B1(n_191),
.B2(n_232),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_251),
.B(n_246),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_287),
.B(n_304),
.C(n_268),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_288),
.B(n_289),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_284),
.A2(n_221),
.B1(n_202),
.B2(n_224),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_280),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_290),
.B(n_301),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_191),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_291),
.B(n_297),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_294),
.A2(n_303),
.B1(n_306),
.B2(n_310),
.Y(n_329)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_254),
.Y(n_295)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_295),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_296),
.A2(n_302),
.B(n_308),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_210),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_298),
.B(n_264),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_195),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_299),
.B(n_307),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_267),
.A2(n_227),
.B1(n_247),
.B2(n_213),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_262),
.A2(n_231),
.B1(n_234),
.B2(n_235),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_249),
.B(n_201),
.C(n_255),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_280),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_305),
.B(n_309),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_277),
.A2(n_272),
.B1(n_276),
.B2(n_278),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_249),
.B(n_277),
.Y(n_307)
);

OA21x2_ASAP7_75t_L g308 ( 
.A1(n_283),
.A2(n_274),
.B(n_271),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_257),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_263),
.A2(n_283),
.B1(n_259),
.B2(n_267),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_252),
.B(n_279),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_311),
.B(n_317),
.Y(n_334)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_252),
.Y(n_313)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_313),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_256),
.B(n_282),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_314),
.Y(n_326)
);

NOR2x1_ASAP7_75t_R g315 ( 
.A(n_259),
.B(n_281),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_315),
.A2(n_253),
.B(n_258),
.Y(n_341)
);

INVxp33_ASAP7_75t_L g316 ( 
.A(n_274),
.Y(n_316)
);

INVx13_ASAP7_75t_L g328 ( 
.A(n_316),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_274),
.A2(n_275),
.B1(n_285),
.B2(n_264),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_292),
.A2(n_260),
.B(n_250),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_319),
.A2(n_325),
.B(n_333),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_311),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_323),
.B(n_341),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_324),
.B(n_327),
.C(n_335),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_292),
.A2(n_260),
.B(n_269),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_287),
.B(n_253),
.Y(n_327)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_318),
.Y(n_332)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_332),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_292),
.A2(n_269),
.B(n_265),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_299),
.Y(n_336)
);

INVx13_ASAP7_75t_L g352 ( 
.A(n_336),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_297),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_338),
.B(n_342),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_293),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_318),
.Y(n_343)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_343),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_317),
.A2(n_265),
.B(n_268),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_344),
.A2(n_302),
.B(n_312),
.Y(n_364)
);

BUFx12_ASAP7_75t_L g345 ( 
.A(n_339),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_345),
.Y(n_368)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_332),
.Y(n_349)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_349),
.Y(n_369)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_343),
.Y(n_350)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_350),
.Y(n_371)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_330),
.Y(n_351)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_351),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_340),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_354),
.B(n_357),
.Y(n_376)
);

AO21x1_ASAP7_75t_L g356 ( 
.A1(n_325),
.A2(n_308),
.B(n_315),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_356),
.A2(n_358),
.B1(n_359),
.B2(n_361),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_331),
.B(n_307),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_331),
.B(n_323),
.Y(n_358)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_340),
.Y(n_359)
);

O2A1O1Ixp33_ASAP7_75t_L g360 ( 
.A1(n_320),
.A2(n_308),
.B(n_296),
.C(n_316),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_360),
.A2(n_319),
.B1(n_333),
.B2(n_334),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_320),
.A2(n_294),
.B1(n_310),
.B2(n_303),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_327),
.B(n_298),
.C(n_304),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_362),
.B(n_366),
.Y(n_380)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_330),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_363),
.B(n_337),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_364),
.A2(n_325),
.B1(n_344),
.B2(n_333),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_336),
.B(n_338),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_367),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_353),
.B(n_335),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_372),
.B(n_382),
.C(n_353),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_373),
.A2(n_374),
.B1(n_375),
.B2(n_383),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_360),
.A2(n_365),
.B1(n_334),
.B2(n_348),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_360),
.A2(n_319),
.B1(n_306),
.B2(n_321),
.Y(n_375)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_377),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_354),
.B(n_326),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_378),
.B(n_379),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_348),
.B(n_342),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_362),
.B(n_335),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_361),
.A2(n_329),
.B1(n_289),
.B2(n_321),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_365),
.A2(n_327),
.B1(n_329),
.B2(n_286),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_384),
.B(n_341),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_372),
.B(n_362),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_386),
.B(n_391),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_387),
.B(n_389),
.C(n_397),
.Y(n_407)
);

AOI32xp33_ASAP7_75t_L g388 ( 
.A1(n_368),
.A2(n_365),
.A3(n_355),
.B1(n_359),
.B2(n_356),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_388),
.B(n_398),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_382),
.B(n_353),
.C(n_324),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_376),
.B(n_337),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_393),
.B(n_357),
.Y(n_405)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_376),
.Y(n_394)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_394),
.Y(n_404)
);

O2A1O1Ixp33_ASAP7_75t_L g395 ( 
.A1(n_368),
.A2(n_366),
.B(n_364),
.C(n_356),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_395),
.A2(n_367),
.B(n_322),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_380),
.B(n_324),
.C(n_384),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_380),
.B(n_356),
.C(n_355),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_370),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_400),
.B(n_402),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_390),
.A2(n_374),
.B(n_373),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_403),
.A2(n_395),
.B(n_322),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_405),
.B(n_300),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_397),
.B(n_375),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_406),
.B(n_392),
.C(n_389),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_386),
.B(n_383),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_408),
.B(n_398),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_385),
.A2(n_329),
.B1(n_358),
.B2(n_286),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_409),
.A2(n_396),
.B1(n_369),
.B2(n_371),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_410),
.B(n_414),
.Y(n_420)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_411),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_412),
.B(n_400),
.C(n_406),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_413),
.B(n_403),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_404),
.B(n_300),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_416),
.B(n_417),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_408),
.B(n_396),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_412),
.A2(n_369),
.B1(n_371),
.B2(n_381),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_418),
.B(n_423),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_419),
.B(n_424),
.Y(n_426)
);

NOR2xp67_ASAP7_75t_SL g424 ( 
.A(n_415),
.B(n_401),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_421),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_425),
.B(n_427),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_420),
.B(n_407),
.C(n_399),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_422),
.B(n_407),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_428),
.A2(n_399),
.B(n_423),
.Y(n_431)
);

MAJx2_ASAP7_75t_L g430 ( 
.A(n_426),
.B(n_427),
.C(n_429),
.Y(n_430)
);

AOI322xp5_ASAP7_75t_L g433 ( 
.A1(n_430),
.A2(n_431),
.A3(n_352),
.B1(n_345),
.B2(n_413),
.C1(n_339),
.C2(n_328),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_433),
.B(n_434),
.Y(n_435)
);

AOI322xp5_ASAP7_75t_L g434 ( 
.A1(n_432),
.A2(n_352),
.A3(n_381),
.B1(n_345),
.B2(n_349),
.C1(n_350),
.C2(n_347),
.Y(n_434)
);

AOI321xp33_ASAP7_75t_L g436 ( 
.A1(n_435),
.A2(n_352),
.A3(n_291),
.B1(n_346),
.B2(n_347),
.C(n_363),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_436),
.B(n_351),
.Y(n_437)
);


endmodule