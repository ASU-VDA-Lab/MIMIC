module fake_ariane_960_n_1218 (n_295, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_294, n_197, n_176, n_34, n_172, n_183, n_299, n_12, n_133, n_66, n_205, n_71, n_109, n_245, n_96, n_49, n_20, n_283, n_50, n_187, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_214, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_77, n_15, n_23, n_87, n_279, n_207, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_311, n_239, n_35, n_272, n_54, n_8, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_115, n_267, n_291, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_227, n_48, n_188, n_11, n_129, n_126, n_282, n_277, n_248, n_301, n_293, n_228, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_238, n_136, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_221, n_86, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_26, n_246, n_0, n_159, n_105, n_30, n_131, n_263, n_229, n_250, n_165, n_144, n_101, n_243, n_134, n_185, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_258, n_118, n_121, n_22, n_241, n_29, n_191, n_80, n_211, n_97, n_251, n_116, n_39, n_155, n_127, n_1218);

input n_295;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_71;
input n_109;
input n_245;
input n_96;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_214;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_115;
input n_267;
input n_291;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_227;
input n_48;
input n_188;
input n_11;
input n_129;
input n_126;
input n_282;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_238;
input n_136;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_221;
input n_86;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_26;
input n_246;
input n_0;
input n_159;
input n_105;
input n_30;
input n_131;
input n_263;
input n_229;
input n_250;
input n_165;
input n_144;
input n_101;
input n_243;
input n_134;
input n_185;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_258;
input n_118;
input n_121;
input n_22;
input n_241;
input n_29;
input n_191;
input n_80;
input n_211;
input n_97;
input n_251;
input n_116;
input n_39;
input n_155;
input n_127;

output n_1218;

wire n_356;
wire n_556;
wire n_698;
wire n_1127;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_1020;
wire n_1209;
wire n_1137;
wire n_646;
wire n_1174;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_1214;
wire n_404;
wire n_943;
wire n_1118;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_479;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_836;
wire n_541;
wire n_499;
wire n_1169;
wire n_789;
wire n_788;
wire n_908;
wire n_850;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_1029;
wire n_341;
wire n_985;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_1180;
wire n_969;
wire n_1109;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_679;
wire n_643;
wire n_924;
wire n_927;
wire n_781;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_586;
wire n_443;
wire n_952;
wire n_864;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_528;
wire n_584;
wire n_424;
wire n_1154;
wire n_1166;
wire n_387;
wire n_1200;
wire n_406;
wire n_826;
wire n_1130;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_940;
wire n_466;
wire n_1016;
wire n_346;
wire n_1138;
wire n_1149;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_1196;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_1181;
wire n_379;
wire n_515;
wire n_807;
wire n_445;
wire n_765;
wire n_1131;
wire n_1187;
wire n_891;
wire n_737;
wire n_885;
wire n_441;
wire n_568;
wire n_1032;
wire n_1217;
wire n_385;
wire n_637;
wire n_917;
wire n_1208;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_1177;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_1167;
wire n_1170;
wire n_1151;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_905;
wire n_945;
wire n_702;
wire n_958;
wire n_790;
wire n_898;
wire n_857;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_1064;
wire n_633;
wire n_900;
wire n_1133;
wire n_883;
wire n_338;
wire n_1163;
wire n_995;
wire n_1093;
wire n_473;
wire n_801;
wire n_1184;
wire n_761;
wire n_733;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_779;
wire n_754;
wire n_731;
wire n_903;
wire n_315;
wire n_871;
wire n_1073;
wire n_594;
wire n_1173;
wire n_402;
wire n_1052;
wire n_1068;
wire n_829;
wire n_1198;
wire n_1062;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_1018;
wire n_597;
wire n_816;
wire n_855;
wire n_1047;
wire n_835;
wire n_808;
wire n_953;
wire n_553;
wire n_446;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_405;
wire n_557;
wire n_1201;
wire n_1107;
wire n_858;
wire n_645;
wire n_989;
wire n_1185;
wire n_320;
wire n_331;
wire n_559;
wire n_1134;
wire n_485;
wire n_401;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_1141;
wire n_350;
wire n_822;
wire n_1143;
wire n_344;
wire n_795;
wire n_381;
wire n_721;
wire n_600;
wire n_840;
wire n_481;
wire n_426;
wire n_433;
wire n_1053;
wire n_1084;
wire n_398;
wire n_1090;
wire n_529;
wire n_502;
wire n_561;
wire n_770;
wire n_821;
wire n_928;
wire n_839;
wire n_1099;
wire n_1153;
wire n_465;
wire n_486;
wire n_901;
wire n_507;
wire n_759;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_1145;
wire n_971;
wire n_369;
wire n_1192;
wire n_894;
wire n_787;
wire n_1105;
wire n_547;
wire n_1195;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_1172;
wire n_703;
wire n_478;
wire n_1207;
wire n_748;
wire n_1212;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_1160;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_997;
wire n_635;
wire n_707;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_1116;
wire n_983;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_727;
wire n_699;
wire n_1085;
wire n_467;
wire n_1152;
wire n_432;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_644;
wire n_823;
wire n_921;
wire n_620;
wire n_1197;
wire n_325;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_1165;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_455;
wire n_365;
wire n_654;
wire n_429;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_1128;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1122;
wire n_1049;
wire n_1205;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_1132;
wire n_390;
wire n_1156;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_1202;
wire n_627;
wire n_1039;
wire n_1188;
wire n_539;
wire n_1150;
wire n_728;
wire n_957;
wire n_388;
wire n_333;
wire n_612;
wire n_977;
wire n_413;
wire n_392;
wire n_376;
wire n_449;
wire n_1216;
wire n_715;
wire n_512;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_685;
wire n_911;
wire n_321;
wire n_459;
wire n_1136;
wire n_458;
wire n_361;
wire n_1190;
wire n_1144;
wire n_383;
wire n_623;
wire n_838;
wire n_1213;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_1142;
wire n_616;
wire n_617;
wire n_705;
wire n_630;
wire n_658;
wire n_1140;
wire n_570;
wire n_1055;
wire n_362;
wire n_543;
wire n_942;
wire n_709;
wire n_601;
wire n_683;
wire n_1089;
wire n_565;
wire n_1189;
wire n_628;
wire n_809;
wire n_461;
wire n_1121;
wire n_490;
wire n_743;
wire n_1194;
wire n_907;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_1159;
wire n_910;
wire n_1210;
wire n_527;
wire n_741;
wire n_772;
wire n_747;
wire n_847;
wire n_939;
wire n_1135;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1114;
wire n_676;
wire n_708;
wire n_551;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_1199;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_534;
wire n_1108;
wire n_1164;
wire n_355;
wire n_609;
wire n_851;
wire n_444;
wire n_1043;
wire n_560;
wire n_450;
wire n_890;
wire n_1193;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_1179;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_1158;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_596;
wire n_954;
wire n_912;
wire n_1168;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_1157;
wire n_555;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_982;
wire n_915;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_1182;
wire n_763;
wire n_655;
wire n_540;
wire n_544;
wire n_692;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_403;
wire n_750;
wire n_991;
wire n_834;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_812;
wire n_1126;
wire n_395;
wire n_621;
wire n_1178;
wire n_606;
wire n_951;
wire n_1026;
wire n_938;
wire n_862;
wire n_895;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_666;
wire n_1000;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_1206;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1146;
wire n_1100;
wire n_1171;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_1203;
wire n_619;
wire n_337;
wire n_697;
wire n_437;
wire n_622;
wire n_967;
wire n_998;
wire n_999;
wire n_1083;
wire n_472;
wire n_937;
wire n_746;
wire n_456;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_704;
wire n_1060;
wire n_1175;
wire n_1044;
wire n_1148;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_1211;
wire n_963;
wire n_873;
wire n_1082;
wire n_1139;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_1051;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_434;
wire n_1102;
wire n_360;
wire n_1101;
wire n_975;
wire n_1129;
wire n_563;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_1183;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_1204;
wire n_994;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_972;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_1161;
wire n_431;
wire n_1176;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1155;
wire n_1191;
wire n_1071;
wire n_712;
wire n_976;
wire n_411;
wire n_849;
wire n_909;
wire n_484;
wire n_353;
wire n_767;
wire n_736;
wire n_1025;
wire n_1215;
wire n_357;
wire n_412;
wire n_687;
wire n_964;
wire n_447;
wire n_1057;
wire n_797;
wire n_382;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_1147;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_886;
wire n_351;
wire n_471;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g314 ( 
.A(n_95),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_161),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_262),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_113),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_180),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_167),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_248),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_199),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_86),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_115),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_225),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_44),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_31),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_311),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_120),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_24),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_298),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_97),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_20),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_302),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_142),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_170),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_139),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_204),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_34),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_253),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_96),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_299),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_133),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_145),
.Y(n_343)
);

BUFx10_ASAP7_75t_L g344 ( 
.A(n_20),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_230),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_178),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_189),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_266),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_107),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_265),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_109),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_235),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_81),
.B(n_119),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_46),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_13),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_284),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_121),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_214),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_24),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_7),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_72),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_41),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_246),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_215),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_36),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_312),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_313),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_28),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_179),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_283),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_303),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_212),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_228),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_110),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_287),
.Y(n_375)
);

BUFx10_ASAP7_75t_L g376 ( 
.A(n_237),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_117),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_243),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_17),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_267),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_273),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_38),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_196),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_91),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_51),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_222),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_8),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_14),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_172),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_49),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_138),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_62),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_112),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_163),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_188),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_227),
.Y(n_396)
);

BUFx5_ASAP7_75t_L g397 ( 
.A(n_293),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_118),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_127),
.Y(n_399)
);

CKINVDCx14_ASAP7_75t_R g400 ( 
.A(n_175),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_54),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_75),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_209),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_177),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_0),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_162),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_2),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_282),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_94),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_134),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_69),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_275),
.Y(n_412)
);

INVx2_ASAP7_75t_SL g413 ( 
.A(n_59),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_80),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_153),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_21),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_198),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_11),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_156),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_68),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_305),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_229),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_285),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_234),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_90),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_61),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_122),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_251),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_200),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_45),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_186),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_193),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_147),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_71),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_148),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_50),
.Y(n_436)
);

INVx2_ASAP7_75t_SL g437 ( 
.A(n_226),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_128),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_67),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_257),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_272),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_130),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_195),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_210),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_261),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_309),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_159),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_171),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_297),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_37),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_217),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_288),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_3),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_216),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_11),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_252),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_58),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_108),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_164),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_116),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_43),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_241),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_26),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_26),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_173),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_260),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_32),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_104),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_22),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_19),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_221),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_39),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_101),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_9),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_250),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_256),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_12),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_308),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_301),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_92),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_307),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_245),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_279),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_35),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_3),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_206),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_137),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_304),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_258),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_126),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_47),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_2),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_182),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_70),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_53),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_48),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_29),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_247),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_8),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_10),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_99),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_276),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_208),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_268),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_197),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_77),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_102),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_5),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_224),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_4),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_76),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_269),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_52),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_21),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_191),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_19),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_213),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_114),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_93),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_202),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_296),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_335),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_339),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_407),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_339),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_435),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_342),
.Y(n_527)
);

INVxp67_ASAP7_75t_SL g528 ( 
.A(n_359),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_435),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_455),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_461),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_348),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_461),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_385),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_422),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_468),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_360),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_482),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_332),
.Y(n_539)
);

CKINVDCx16_ASAP7_75t_R g540 ( 
.A(n_363),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_329),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_405),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_355),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_368),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_463),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_379),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g547 ( 
.A(n_452),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_325),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_418),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_387),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_374),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_464),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_388),
.Y(n_553)
);

NOR2xp67_ASAP7_75t_L g554 ( 
.A(n_416),
.B(n_0),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_469),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_477),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_485),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_453),
.Y(n_558)
);

NOR2xp67_ASAP7_75t_L g559 ( 
.A(n_470),
.B(n_492),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_400),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_344),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_376),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_497),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_499),
.Y(n_564)
);

INVxp67_ASAP7_75t_SL g565 ( 
.A(n_508),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_376),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_500),
.Y(n_567)
);

INVx1_ASAP7_75t_SL g568 ( 
.A(n_474),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_510),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_514),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_344),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_314),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_320),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_315),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_322),
.B(n_1),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_334),
.B(n_347),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_352),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_316),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_354),
.B(n_1),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g580 ( 
.A(n_516),
.Y(n_580)
);

BUFx2_ASAP7_75t_SL g581 ( 
.A(n_384),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_465),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_521),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_317),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_319),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_321),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_358),
.B(n_4),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_364),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_323),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_365),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_366),
.Y(n_591)
);

CKINVDCx16_ASAP7_75t_R g592 ( 
.A(n_374),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_324),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_327),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_328),
.Y(n_595)
);

CKINVDCx16_ASAP7_75t_R g596 ( 
.A(n_374),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_367),
.B(n_369),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_373),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_386),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_520),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_330),
.Y(n_601)
);

INVxp67_ASAP7_75t_L g602 ( 
.A(n_391),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_392),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_394),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_331),
.Y(n_605)
);

INVxp67_ASAP7_75t_SL g606 ( 
.A(n_318),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_336),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_403),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_404),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_409),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_R g611 ( 
.A(n_337),
.B(n_30),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_338),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_340),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_343),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_345),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_414),
.B(n_5),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_417),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_346),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_349),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_419),
.B(n_6),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_421),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_350),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_351),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_423),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_430),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_436),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_439),
.Y(n_627)
);

CKINVDCx16_ASAP7_75t_R g628 ( 
.A(n_374),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_356),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_357),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_362),
.Y(n_631)
);

CKINVDCx16_ASAP7_75t_R g632 ( 
.A(n_431),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_440),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_413),
.B(n_6),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_454),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_458),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_370),
.Y(n_637)
);

CKINVDCx16_ASAP7_75t_R g638 ( 
.A(n_431),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_527),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_551),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_551),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_535),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_538),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_576),
.B(n_572),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_522),
.Y(n_645)
);

AND2x6_ASAP7_75t_L g646 ( 
.A(n_634),
.B(n_431),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_537),
.Y(n_647)
);

INVxp67_ASAP7_75t_L g648 ( 
.A(n_568),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_532),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_551),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_580),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_542),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_549),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_534),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g655 ( 
.A(n_570),
.Y(n_655)
);

CKINVDCx20_ASAP7_75t_R g656 ( 
.A(n_541),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_551),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_552),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_556),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_530),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_608),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_625),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_536),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_528),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_558),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_530),
.Y(n_666)
);

CKINVDCx16_ASAP7_75t_R g667 ( 
.A(n_540),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_573),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_574),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_547),
.B(n_578),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_584),
.B(n_460),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_565),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_562),
.B(n_333),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_585),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_577),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_588),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_590),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_616),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_591),
.B(n_467),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_589),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_598),
.B(n_475),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_603),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_545),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_594),
.Y(n_684)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_548),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_604),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_560),
.Y(n_687)
);

INVxp67_ASAP7_75t_SL g688 ( 
.A(n_524),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_609),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_595),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_617),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_592),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_605),
.B(n_607),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_612),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_596),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_621),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_613),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_614),
.Y(n_698)
);

OAI22xp5_ASAP7_75t_SL g699 ( 
.A1(n_567),
.A2(n_486),
.B1(n_487),
.B2(n_480),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_624),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_626),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_627),
.B(n_493),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_539),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_618),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_633),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_570),
.B(n_361),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_635),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_628),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_597),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_636),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_636),
.Y(n_711)
);

CKINVDCx20_ASAP7_75t_R g712 ( 
.A(n_583),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_575),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_575),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_523),
.B(n_525),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_586),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_622),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_629),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_632),
.Y(n_719)
);

HB1xp67_ASAP7_75t_L g720 ( 
.A(n_543),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_630),
.Y(n_721)
);

BUFx2_ASAP7_75t_L g722 ( 
.A(n_544),
.Y(n_722)
);

INVxp67_ASAP7_75t_L g723 ( 
.A(n_599),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_593),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_582),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_631),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_579),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_637),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_692),
.B(n_566),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_665),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_651),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_709),
.B(n_638),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_665),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_676),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_692),
.B(n_526),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_665),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_695),
.Y(n_737)
);

AND2x2_ASAP7_75t_SL g738 ( 
.A(n_667),
.B(n_529),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_695),
.B(n_546),
.Y(n_739)
);

INVx4_ASAP7_75t_L g740 ( 
.A(n_669),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_640),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_708),
.B(n_550),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_677),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_673),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_725),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_678),
.B(n_606),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_641),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_719),
.B(n_553),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_660),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_657),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_666),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_686),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_661),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_662),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_688),
.B(n_531),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_648),
.B(n_561),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_648),
.B(n_555),
.Y(n_757)
);

OR2x6_ASAP7_75t_L g758 ( 
.A(n_703),
.B(n_571),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_668),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_675),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_722),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_647),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_641),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_652),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_682),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_678),
.B(n_581),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_689),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_693),
.B(n_563),
.Y(n_768)
);

AND2x4_ASAP7_75t_L g769 ( 
.A(n_715),
.B(n_533),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_678),
.B(n_564),
.Y(n_770)
);

INVx4_ASAP7_75t_L g771 ( 
.A(n_674),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_710),
.B(n_557),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_723),
.B(n_569),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_696),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_700),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_723),
.B(n_600),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_701),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_707),
.Y(n_778)
);

INVx6_ASAP7_75t_L g779 ( 
.A(n_706),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_680),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_691),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_713),
.B(n_602),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_684),
.B(n_601),
.Y(n_783)
);

INVx1_ASAP7_75t_SL g784 ( 
.A(n_656),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_705),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_690),
.B(n_615),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_711),
.B(n_610),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_655),
.B(n_720),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_653),
.Y(n_789)
);

BUFx10_ASAP7_75t_L g790 ( 
.A(n_694),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_697),
.B(n_619),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_641),
.Y(n_792)
);

NAND3xp33_ASAP7_75t_L g793 ( 
.A(n_671),
.B(n_587),
.C(n_579),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_650),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_658),
.Y(n_795)
);

INVx5_ASAP7_75t_L g796 ( 
.A(n_646),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_664),
.B(n_623),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_659),
.Y(n_798)
);

AND2x6_ASAP7_75t_L g799 ( 
.A(n_714),
.B(n_431),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_650),
.Y(n_800)
);

NAND2x1p5_ASAP7_75t_L g801 ( 
.A(n_670),
.B(n_559),
.Y(n_801)
);

BUFx4f_ASAP7_75t_L g802 ( 
.A(n_672),
.Y(n_802)
);

NAND2xp33_ASAP7_75t_L g803 ( 
.A(n_698),
.B(n_611),
.Y(n_803)
);

AND2x6_ASAP7_75t_L g804 ( 
.A(n_727),
.B(n_496),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_650),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_644),
.B(n_587),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_646),
.Y(n_807)
);

INVx5_ASAP7_75t_L g808 ( 
.A(n_646),
.Y(n_808)
);

AND2x6_ASAP7_75t_L g809 ( 
.A(n_679),
.B(n_496),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_646),
.Y(n_810)
);

INVxp67_ASAP7_75t_L g811 ( 
.A(n_639),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_704),
.B(n_554),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_757),
.B(n_717),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_739),
.B(n_718),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_734),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_749),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_734),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_751),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_806),
.B(n_644),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_743),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_770),
.B(n_721),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_759),
.Y(n_822)
);

AO22x1_ASAP7_75t_L g823 ( 
.A1(n_797),
.A2(n_642),
.B1(n_643),
.B2(n_726),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_732),
.B(n_782),
.Y(n_824)
);

OAI22xp33_ASAP7_75t_L g825 ( 
.A1(n_793),
.A2(n_728),
.B1(n_655),
.B2(n_681),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_790),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_743),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_752),
.Y(n_828)
);

A2O1A1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_752),
.A2(n_620),
.B(n_681),
.C(n_679),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_774),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_773),
.B(n_699),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_774),
.A2(n_702),
.B(n_620),
.Y(n_832)
);

NAND2xp33_ASAP7_75t_L g833 ( 
.A(n_807),
.B(n_397),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_775),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_756),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_789),
.B(n_702),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_779),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_760),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_788),
.A2(n_735),
.B1(n_755),
.B2(n_787),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_807),
.Y(n_840)
);

OR2x6_ASAP7_75t_L g841 ( 
.A(n_745),
.B(n_712),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_737),
.B(n_716),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_765),
.Y(n_843)
);

INVx2_ASAP7_75t_SL g844 ( 
.A(n_779),
.Y(n_844)
);

NOR2x1p5_ASAP7_75t_L g845 ( 
.A(n_740),
.B(n_645),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_810),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_798),
.B(n_432),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_767),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_744),
.B(n_649),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_753),
.Y(n_850)
);

BUFx2_ASAP7_75t_L g851 ( 
.A(n_761),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_754),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_780),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_731),
.B(n_654),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_775),
.A2(n_724),
.B1(n_495),
.B2(n_502),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_746),
.B(n_457),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_777),
.B(n_371),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_777),
.B(n_372),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_778),
.Y(n_859)
);

INVx3_ASAP7_75t_L g860 ( 
.A(n_810),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_742),
.B(n_663),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_778),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_784),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_762),
.A2(n_503),
.B1(n_504),
.B2(n_498),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_764),
.A2(n_506),
.B1(n_513),
.B2(n_505),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_768),
.B(n_685),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_748),
.B(n_687),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_776),
.B(n_683),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_795),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_766),
.B(n_515),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_755),
.B(n_375),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_781),
.B(n_377),
.Y(n_872)
);

INVx8_ASAP7_75t_L g873 ( 
.A(n_758),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_771),
.B(n_378),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_802),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_781),
.B(n_380),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_811),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_729),
.B(n_381),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_785),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_785),
.B(n_382),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_787),
.B(n_383),
.Y(n_881)
);

AND2x4_ASAP7_75t_L g882 ( 
.A(n_729),
.B(n_518),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_769),
.A2(n_437),
.B1(n_473),
.B2(n_429),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_741),
.Y(n_884)
);

A2O1A1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_772),
.A2(n_353),
.B(n_517),
.C(n_490),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_730),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_733),
.Y(n_887)
);

AOI22xp5_ASAP7_75t_L g888 ( 
.A1(n_735),
.A2(n_353),
.B1(n_341),
.B2(n_326),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_772),
.B(n_733),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_747),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_800),
.A2(n_750),
.B(n_812),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_736),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_769),
.A2(n_462),
.B1(n_512),
.B2(n_511),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_736),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_853),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_841),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_813),
.B(n_738),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_831),
.A2(n_803),
.B1(n_783),
.B2(n_791),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_863),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_839),
.B(n_758),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_815),
.Y(n_901)
);

OR2x2_ASAP7_75t_L g902 ( 
.A(n_841),
.B(n_786),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_819),
.B(n_801),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_841),
.Y(n_904)
);

INVx5_ASAP7_75t_L g905 ( 
.A(n_873),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_839),
.B(n_809),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_824),
.B(n_796),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_835),
.B(n_854),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_826),
.Y(n_909)
);

BUFx2_ASAP7_75t_L g910 ( 
.A(n_851),
.Y(n_910)
);

INVxp67_ASAP7_75t_SL g911 ( 
.A(n_889),
.Y(n_911)
);

NOR3xp33_ASAP7_75t_SL g912 ( 
.A(n_877),
.B(n_814),
.C(n_825),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_R g913 ( 
.A(n_875),
.B(n_867),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_873),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_873),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_836),
.B(n_847),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_856),
.B(n_809),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_842),
.Y(n_918)
);

AOI22xp5_ASAP7_75t_L g919 ( 
.A1(n_821),
.A2(n_799),
.B1(n_804),
.B2(n_809),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_823),
.B(n_796),
.Y(n_920)
);

OR2x2_ASAP7_75t_L g921 ( 
.A(n_868),
.B(n_747),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_849),
.B(n_799),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_817),
.A2(n_808),
.B(n_796),
.C(n_390),
.Y(n_923)
);

CKINVDCx6p67_ASAP7_75t_R g924 ( 
.A(n_842),
.Y(n_924)
);

INVx3_ASAP7_75t_SL g925 ( 
.A(n_882),
.Y(n_925)
);

NOR3xp33_ASAP7_75t_SL g926 ( 
.A(n_874),
.B(n_866),
.C(n_878),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_820),
.Y(n_927)
);

INVxp67_ASAP7_75t_SL g928 ( 
.A(n_840),
.Y(n_928)
);

NOR3xp33_ASAP7_75t_SL g929 ( 
.A(n_885),
.B(n_393),
.C(n_389),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_822),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_837),
.Y(n_931)
);

INVxp67_ASAP7_75t_SL g932 ( 
.A(n_840),
.Y(n_932)
);

BUFx12f_ASAP7_75t_SL g933 ( 
.A(n_882),
.Y(n_933)
);

NAND2x1p5_ASAP7_75t_L g934 ( 
.A(n_846),
.B(n_808),
.Y(n_934)
);

OR2x4_ASAP7_75t_L g935 ( 
.A(n_869),
.B(n_763),
.Y(n_935)
);

AND2x6_ASAP7_75t_L g936 ( 
.A(n_846),
.B(n_496),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_838),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_844),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_827),
.Y(n_939)
);

BUFx12f_ASAP7_75t_SL g940 ( 
.A(n_845),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_828),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_860),
.B(n_808),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_830),
.B(n_799),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_834),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_859),
.B(n_804),
.Y(n_945)
);

INVx6_ASAP7_75t_L g946 ( 
.A(n_861),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_855),
.Y(n_947)
);

INVx4_ASAP7_75t_L g948 ( 
.A(n_860),
.Y(n_948)
);

NAND3xp33_ASAP7_75t_SL g949 ( 
.A(n_893),
.B(n_396),
.C(n_395),
.Y(n_949)
);

NAND2xp33_ASAP7_75t_SL g950 ( 
.A(n_862),
.B(n_763),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_879),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_816),
.B(n_792),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_832),
.B(n_804),
.Y(n_953)
);

INVx1_ASAP7_75t_SL g954 ( 
.A(n_910),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_947),
.B(n_855),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_911),
.B(n_903),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_908),
.B(n_832),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_898),
.B(n_829),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_901),
.B(n_871),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_927),
.B(n_939),
.Y(n_960)
);

OAI21x1_ASAP7_75t_L g961 ( 
.A1(n_953),
.A2(n_891),
.B(n_886),
.Y(n_961)
);

OAI21x1_ASAP7_75t_L g962 ( 
.A1(n_943),
.A2(n_852),
.B(n_850),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_941),
.Y(n_963)
);

AOI21x1_ASAP7_75t_SL g964 ( 
.A1(n_945),
.A2(n_858),
.B(n_857),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_944),
.B(n_893),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_897),
.B(n_881),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_951),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_916),
.A2(n_876),
.B(n_872),
.Y(n_968)
);

NAND3xp33_ASAP7_75t_L g969 ( 
.A(n_912),
.B(n_926),
.C(n_888),
.Y(n_969)
);

BUFx12f_ASAP7_75t_L g970 ( 
.A(n_914),
.Y(n_970)
);

OA21x2_ASAP7_75t_L g971 ( 
.A1(n_917),
.A2(n_870),
.B(n_880),
.Y(n_971)
);

AOI211x1_ASAP7_75t_L g972 ( 
.A1(n_949),
.A2(n_864),
.B(n_865),
.C(n_887),
.Y(n_972)
);

NOR2xp67_ASAP7_75t_SL g973 ( 
.A(n_909),
.B(n_890),
.Y(n_973)
);

AOI211x1_ASAP7_75t_L g974 ( 
.A1(n_906),
.A2(n_864),
.B(n_888),
.C(n_10),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_942),
.Y(n_975)
);

INVx5_ASAP7_75t_L g976 ( 
.A(n_914),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_930),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_923),
.A2(n_848),
.B(n_843),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_937),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_900),
.B(n_883),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_907),
.A2(n_890),
.B1(n_892),
.B2(n_894),
.Y(n_981)
);

INVx5_ASAP7_75t_L g982 ( 
.A(n_915),
.Y(n_982)
);

AOI221x1_ASAP7_75t_L g983 ( 
.A1(n_950),
.A2(n_884),
.B1(n_794),
.B2(n_805),
.C(n_792),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_925),
.B(n_818),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_952),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_899),
.B(n_794),
.Y(n_986)
);

OAI21x1_ASAP7_75t_L g987 ( 
.A1(n_934),
.A2(n_833),
.B(n_805),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_895),
.Y(n_988)
);

OAI21x1_ASAP7_75t_L g989 ( 
.A1(n_919),
.A2(n_920),
.B(n_922),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_928),
.A2(n_399),
.B(n_398),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_905),
.B(n_7),
.Y(n_991)
);

AO22x2_ASAP7_75t_L g992 ( 
.A1(n_902),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_952),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_932),
.A2(n_948),
.B(n_942),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_948),
.A2(n_402),
.B(n_401),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_929),
.A2(n_408),
.B(n_406),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_913),
.B(n_14),
.Y(n_997)
);

AOI21x1_ASAP7_75t_L g998 ( 
.A1(n_921),
.A2(n_397),
.B(n_496),
.Y(n_998)
);

OAI21x1_ASAP7_75t_L g999 ( 
.A1(n_961),
.A2(n_904),
.B(n_918),
.Y(n_999)
);

OAI21x1_ASAP7_75t_L g1000 ( 
.A1(n_962),
.A2(n_935),
.B(n_936),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_963),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_L g1002 ( 
.A1(n_964),
.A2(n_936),
.B(n_397),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_958),
.A2(n_946),
.B1(n_910),
.B2(n_896),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_967),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_968),
.A2(n_896),
.B(n_905),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_975),
.B(n_905),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_957),
.B(n_946),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_960),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_977),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_977),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_979),
.Y(n_1011)
);

OAI21x1_ASAP7_75t_L g1012 ( 
.A1(n_998),
.A2(n_936),
.B(n_397),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_979),
.Y(n_1013)
);

CKINVDCx8_ASAP7_75t_R g1014 ( 
.A(n_976),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_989),
.A2(n_397),
.B(n_940),
.Y(n_1015)
);

AOI21x1_ASAP7_75t_L g1016 ( 
.A1(n_971),
.A2(n_397),
.B(n_933),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_SL g1017 ( 
.A1(n_965),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_970),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_985),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_L g1020 ( 
.A1(n_978),
.A2(n_40),
.B(n_33),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_L g1021 ( 
.A1(n_987),
.A2(n_55),
.B(n_42),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_975),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_956),
.B(n_915),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_993),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_955),
.B(n_924),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_976),
.Y(n_1026)
);

AO21x1_ASAP7_75t_L g1027 ( 
.A1(n_981),
.A2(n_15),
.B(n_16),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_969),
.A2(n_411),
.B(n_410),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_959),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_966),
.B(n_974),
.Y(n_1030)
);

INVx5_ASAP7_75t_L g1031 ( 
.A(n_976),
.Y(n_1031)
);

AOI22xp33_ASAP7_75t_SL g1032 ( 
.A1(n_992),
.A2(n_895),
.B1(n_938),
.B2(n_931),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_986),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_992),
.A2(n_938),
.B1(n_931),
.B2(n_23),
.Y(n_1034)
);

NAND2x1_ASAP7_75t_L g1035 ( 
.A(n_994),
.B(n_56),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_971),
.A2(n_60),
.B(n_57),
.Y(n_1036)
);

AOI22xp33_ASAP7_75t_L g1037 ( 
.A1(n_980),
.A2(n_519),
.B1(n_509),
.B2(n_507),
.Y(n_1037)
);

AOI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_1034),
.A2(n_991),
.B1(n_954),
.B2(n_997),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_1030),
.A2(n_972),
.B1(n_991),
.B2(n_996),
.Y(n_1039)
);

AND2x4_ASAP7_75t_SL g1040 ( 
.A(n_1006),
.B(n_984),
.Y(n_1040)
);

OAI221xp5_ASAP7_75t_L g1041 ( 
.A1(n_1034),
.A2(n_973),
.B1(n_988),
.B2(n_990),
.C(n_995),
.Y(n_1041)
);

BUFx10_ASAP7_75t_L g1042 ( 
.A(n_1025),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_1018),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1001),
.Y(n_1044)
);

OAI22xp33_ASAP7_75t_L g1045 ( 
.A1(n_1003),
.A2(n_982),
.B1(n_983),
.B2(n_501),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1010),
.Y(n_1046)
);

OAI211xp5_ASAP7_75t_L g1047 ( 
.A1(n_1028),
.A2(n_982),
.B(n_494),
.C(n_491),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_1007),
.B(n_982),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_SL g1049 ( 
.A1(n_1003),
.A2(n_489),
.B1(n_488),
.B2(n_484),
.Y(n_1049)
);

NOR2xp67_ASAP7_75t_L g1050 ( 
.A(n_1005),
.B(n_63),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_1004),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_1007),
.B(n_18),
.Y(n_1052)
);

INVx4_ASAP7_75t_L g1053 ( 
.A(n_1031),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_1028),
.A2(n_415),
.B(n_412),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_1030),
.A2(n_483),
.B1(n_481),
.B2(n_479),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_1031),
.B(n_420),
.Y(n_1056)
);

CKINVDCx16_ASAP7_75t_R g1057 ( 
.A(n_1006),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1013),
.Y(n_1058)
);

INVx1_ASAP7_75t_SL g1059 ( 
.A(n_1031),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_1029),
.B(n_18),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_1015),
.A2(n_65),
.B(n_64),
.Y(n_1061)
);

AOI21xp33_ASAP7_75t_SL g1062 ( 
.A1(n_1032),
.A2(n_22),
.B(n_23),
.Y(n_1062)
);

CKINVDCx8_ASAP7_75t_R g1063 ( 
.A(n_1014),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_1026),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_1037),
.A2(n_478),
.B1(n_476),
.B2(n_472),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_1026),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1008),
.B(n_25),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1023),
.B(n_25),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_1009),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_1011),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_1022),
.Y(n_1071)
);

NAND2xp33_ASAP7_75t_R g1072 ( 
.A(n_1023),
.B(n_471),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1019),
.Y(n_1073)
);

OR2x6_ASAP7_75t_L g1074 ( 
.A(n_1005),
.B(n_66),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_1035),
.A2(n_466),
.B(n_459),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_1027),
.A2(n_456),
.B1(n_451),
.B2(n_450),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_1038),
.A2(n_1017),
.B1(n_1033),
.B2(n_1022),
.Y(n_1077)
);

AOI221xp5_ASAP7_75t_L g1078 ( 
.A1(n_1062),
.A2(n_1024),
.B1(n_424),
.B2(n_443),
.C(n_444),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_1046),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_1076),
.A2(n_999),
.B1(n_1000),
.B2(n_1020),
.Y(n_1080)
);

AOI222xp33_ASAP7_75t_L g1081 ( 
.A1(n_1054),
.A2(n_1052),
.B1(n_1039),
.B2(n_1060),
.C1(n_1067),
.C2(n_1068),
.Y(n_1081)
);

OAI221xp5_ASAP7_75t_L g1082 ( 
.A1(n_1049),
.A2(n_1016),
.B1(n_425),
.B2(n_442),
.C(n_445),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_1051),
.A2(n_1036),
.B1(n_1021),
.B2(n_1002),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_1048),
.B(n_1066),
.Y(n_1084)
);

OR2x2_ASAP7_75t_L g1085 ( 
.A(n_1044),
.B(n_27),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_1069),
.A2(n_1012),
.B1(n_449),
.B2(n_448),
.Y(n_1086)
);

AOI221xp5_ASAP7_75t_L g1087 ( 
.A1(n_1062),
.A2(n_447),
.B1(n_446),
.B2(n_441),
.C(n_438),
.Y(n_1087)
);

OAI211xp5_ASAP7_75t_SL g1088 ( 
.A1(n_1041),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_1088)
);

AO31x2_ASAP7_75t_L g1089 ( 
.A1(n_1070),
.A2(n_73),
.A3(n_74),
.B(n_78),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_1057),
.B(n_426),
.Y(n_1090)
);

AOI221xp5_ASAP7_75t_L g1091 ( 
.A1(n_1055),
.A2(n_434),
.B1(n_433),
.B2(n_428),
.C(n_427),
.Y(n_1091)
);

OAI221xp5_ASAP7_75t_L g1092 ( 
.A1(n_1047),
.A2(n_79),
.B1(n_82),
.B2(n_83),
.C(n_84),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_1045),
.A2(n_1064),
.B1(n_1074),
.B2(n_1063),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_1074),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1071),
.A2(n_1043),
.B1(n_1056),
.B2(n_1059),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1073),
.B(n_89),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_SL g1097 ( 
.A1(n_1040),
.A2(n_98),
.B1(n_100),
.B2(n_103),
.Y(n_1097)
);

AOI221xp5_ASAP7_75t_L g1098 ( 
.A1(n_1065),
.A2(n_105),
.B1(n_106),
.B2(n_111),
.C(n_123),
.Y(n_1098)
);

OAI221xp5_ASAP7_75t_L g1099 ( 
.A1(n_1072),
.A2(n_124),
.B1(n_125),
.B2(n_129),
.C(n_131),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1058),
.Y(n_1100)
);

AO22x2_ASAP7_75t_L g1101 ( 
.A1(n_1071),
.A2(n_132),
.B1(n_135),
.B2(n_136),
.Y(n_1101)
);

INVx11_ASAP7_75t_L g1102 ( 
.A(n_1042),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1042),
.B(n_1053),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_1053),
.B(n_140),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1050),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1050),
.A2(n_141),
.B(n_143),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_1061),
.A2(n_144),
.B(n_146),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1075),
.A2(n_149),
.B(n_150),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_SL g1109 ( 
.A1(n_1039),
.A2(n_151),
.B1(n_152),
.B2(n_154),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1044),
.B(n_155),
.Y(n_1110)
);

OAI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1038),
.A2(n_157),
.B1(n_158),
.B2(n_160),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_SL g1112 ( 
.A1(n_1039),
.A2(n_165),
.B1(n_166),
.B2(n_168),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_1102),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1079),
.Y(n_1114)
);

OR2x2_ASAP7_75t_L g1115 ( 
.A(n_1100),
.B(n_169),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1084),
.B(n_310),
.Y(n_1116)
);

HB1xp67_ASAP7_75t_L g1117 ( 
.A(n_1105),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1103),
.B(n_174),
.Y(n_1118)
);

AND2x4_ASAP7_75t_SL g1119 ( 
.A(n_1104),
.B(n_176),
.Y(n_1119)
);

HB1xp67_ASAP7_75t_L g1120 ( 
.A(n_1096),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1090),
.B(n_181),
.Y(n_1121)
);

INVx4_ASAP7_75t_L g1122 ( 
.A(n_1101),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1089),
.Y(n_1123)
);

AND2x4_ASAP7_75t_L g1124 ( 
.A(n_1085),
.B(n_183),
.Y(n_1124)
);

OR2x2_ASAP7_75t_L g1125 ( 
.A(n_1095),
.B(n_184),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1089),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1089),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1110),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1077),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1101),
.Y(n_1130)
);

NOR2x1_ASAP7_75t_SL g1131 ( 
.A(n_1093),
.B(n_185),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1094),
.A2(n_1088),
.B(n_1081),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_1099),
.B(n_187),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1107),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1080),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1092),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1111),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1114),
.B(n_1112),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1117),
.B(n_1109),
.Y(n_1139)
);

INVx1_ASAP7_75t_SL g1140 ( 
.A(n_1121),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_1113),
.Y(n_1141)
);

AOI221xp5_ASAP7_75t_L g1142 ( 
.A1(n_1132),
.A2(n_1078),
.B1(n_1087),
.B2(n_1098),
.C(n_1091),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_1122),
.B(n_1097),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_1117),
.B(n_1083),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_1119),
.Y(n_1145)
);

OAI31xp33_ASAP7_75t_L g1146 ( 
.A1(n_1136),
.A2(n_1082),
.A3(n_1106),
.B(n_1108),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1120),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1120),
.B(n_1086),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1128),
.B(n_190),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1147),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_1144),
.B(n_1130),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1148),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1139),
.B(n_1135),
.Y(n_1153)
);

AND2x4_ASAP7_75t_L g1154 ( 
.A(n_1145),
.B(n_1122),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1139),
.B(n_1129),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1138),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1140),
.Y(n_1157)
);

BUFx2_ASAP7_75t_SL g1158 ( 
.A(n_1141),
.Y(n_1158)
);

OR2x2_ASAP7_75t_L g1159 ( 
.A(n_1145),
.B(n_1116),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1152),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1154),
.B(n_1143),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1154),
.B(n_1143),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1153),
.B(n_1134),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1150),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1155),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1151),
.B(n_1118),
.Y(n_1166)
);

OAI221xp5_ASAP7_75t_L g1167 ( 
.A1(n_1163),
.A2(n_1156),
.B1(n_1146),
.B2(n_1136),
.C(n_1133),
.Y(n_1167)
);

INVx3_ASAP7_75t_SL g1168 ( 
.A(n_1166),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1165),
.B(n_1157),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1160),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1163),
.Y(n_1171)
);

OR2x2_ASAP7_75t_L g1172 ( 
.A(n_1161),
.B(n_1159),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1162),
.B(n_1151),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1166),
.B(n_1158),
.Y(n_1174)
);

NOR3xp33_ASAP7_75t_L g1175 ( 
.A(n_1164),
.B(n_1142),
.C(n_1137),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1164),
.Y(n_1176)
);

NOR3xp33_ASAP7_75t_L g1177 ( 
.A(n_1167),
.B(n_1142),
.C(n_1133),
.Y(n_1177)
);

OR2x2_ASAP7_75t_L g1178 ( 
.A(n_1169),
.B(n_1172),
.Y(n_1178)
);

OAI32xp33_ASAP7_75t_L g1179 ( 
.A1(n_1175),
.A2(n_1125),
.A3(n_1115),
.B1(n_1131),
.B2(n_1149),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1168),
.A2(n_1119),
.B1(n_1124),
.B2(n_1126),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1169),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1173),
.Y(n_1182)
);

HB1xp67_ASAP7_75t_L g1183 ( 
.A(n_1182),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1178),
.B(n_1174),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1181),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1177),
.B(n_1170),
.Y(n_1186)
);

AOI31xp33_ASAP7_75t_L g1187 ( 
.A1(n_1180),
.A2(n_1171),
.A3(n_1124),
.B(n_1176),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1179),
.B(n_1127),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1186),
.B(n_1127),
.Y(n_1189)
);

XNOR2xp5_ASAP7_75t_L g1190 ( 
.A(n_1184),
.B(n_1126),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1183),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1185),
.B(n_1123),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1191),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1192),
.Y(n_1194)
);

AOI221xp5_ASAP7_75t_L g1195 ( 
.A1(n_1189),
.A2(n_1187),
.B1(n_1188),
.B2(n_1123),
.C(n_203),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1193),
.A2(n_1187),
.B(n_1190),
.Y(n_1196)
);

NOR4xp25_ASAP7_75t_L g1197 ( 
.A(n_1194),
.B(n_192),
.C(n_194),
.D(n_201),
.Y(n_1197)
);

O2A1O1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1195),
.A2(n_205),
.B(n_207),
.C(n_211),
.Y(n_1198)
);

NOR2x1_ASAP7_75t_L g1199 ( 
.A(n_1196),
.B(n_218),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1198),
.A2(n_219),
.B(n_220),
.C(n_223),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_1199),
.Y(n_1201)
);

OAI21xp33_ASAP7_75t_L g1202 ( 
.A1(n_1201),
.A2(n_1197),
.B(n_1200),
.Y(n_1202)
);

NAND3xp33_ASAP7_75t_L g1203 ( 
.A(n_1201),
.B(n_306),
.C(n_232),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1202),
.Y(n_1204)
);

NAND4xp25_ASAP7_75t_L g1205 ( 
.A(n_1203),
.B(n_231),
.C(n_233),
.D(n_236),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1204),
.B(n_238),
.Y(n_1206)
);

INVx4_ASAP7_75t_L g1207 ( 
.A(n_1205),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1204),
.A2(n_300),
.B(n_240),
.Y(n_1208)
);

HB1xp67_ASAP7_75t_L g1209 ( 
.A(n_1208),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1209),
.Y(n_1210)
);

AOI31xp33_ASAP7_75t_L g1211 ( 
.A1(n_1210),
.A2(n_1206),
.A3(n_1207),
.B(n_244),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1210),
.A2(n_239),
.B1(n_242),
.B2(n_249),
.Y(n_1212)
);

AOI222xp33_ASAP7_75t_L g1213 ( 
.A1(n_1212),
.A2(n_254),
.B1(n_255),
.B2(n_259),
.C1(n_263),
.C2(n_264),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1211),
.A2(n_270),
.B1(n_271),
.B2(n_274),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1214),
.A2(n_1213),
.B1(n_278),
.B2(n_280),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_SL g1216 ( 
.A1(n_1214),
.A2(n_277),
.B1(n_281),
.B2(n_286),
.Y(n_1216)
);

AOI221xp5_ASAP7_75t_L g1217 ( 
.A1(n_1215),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.C(n_292),
.Y(n_1217)
);

AOI211xp5_ASAP7_75t_L g1218 ( 
.A1(n_1217),
.A2(n_1216),
.B(n_294),
.C(n_295),
.Y(n_1218)
);


endmodule