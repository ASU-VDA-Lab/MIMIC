module fake_jpeg_16931_n_336 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_7),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_43),
.B(n_45),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_7),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_23),
.B(n_8),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_50),
.B(n_52),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_23),
.B(n_13),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_18),
.B(n_2),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_55),
.B(n_58),
.Y(n_108)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_19),
.B(n_2),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_25),
.B(n_9),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_59),
.B(n_61),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_28),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_28),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_64),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_30),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_63),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g79 ( 
.A(n_66),
.B(n_44),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

CKINVDCx12_ASAP7_75t_R g70 ( 
.A(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_70),
.B(n_90),
.Y(n_118)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_38),
.A2(n_30),
.B1(n_21),
.B2(n_48),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_74),
.A2(n_83),
.B1(n_99),
.B2(n_116),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_57),
.A2(n_30),
.B1(n_36),
.B2(n_25),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_76),
.A2(n_97),
.B1(n_20),
.B2(n_27),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_61),
.B(n_37),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_77),
.B(n_85),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_79),
.B(n_87),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_63),
.A2(n_34),
.B1(n_18),
.B2(n_35),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_34),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_34),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_36),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_58),
.B(n_26),
.Y(n_91)
);

XNOR2x1_ASAP7_75t_L g134 ( 
.A(n_91),
.B(n_22),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_93),
.B(n_4),
.Y(n_164)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

AO22x1_ASAP7_75t_SL g97 ( 
.A1(n_63),
.A2(n_22),
.B1(n_27),
.B2(n_5),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_17),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_98),
.B(n_113),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_53),
.A2(n_17),
.B1(n_31),
.B2(n_35),
.Y(n_99)
);

CKINVDCx9p33_ASAP7_75t_R g101 ( 
.A(n_67),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_101),
.Y(n_153)
);

CKINVDCx12_ASAP7_75t_R g103 ( 
.A(n_49),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_107),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_39),
.B(n_26),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_47),
.B(n_14),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_32),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_31),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_41),
.A2(n_15),
.B1(n_32),
.B2(n_14),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_56),
.B1(n_51),
.B2(n_12),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_120),
.A2(n_150),
.B1(n_163),
.B2(n_151),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_123),
.B(n_133),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_82),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_124),
.B(n_143),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_126),
.A2(n_143),
.B1(n_124),
.B2(n_150),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_27),
.Y(n_127)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_88),
.B(n_22),
.Y(n_128)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_44),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_129),
.B(n_151),
.Y(n_178)
);

NOR2xp67_ASAP7_75t_L g133 ( 
.A(n_91),
.B(n_20),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_145),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_137),
.B(n_141),
.Y(n_194)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_138),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_75),
.B(n_10),
.Y(n_139)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_139),
.Y(n_190)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_140),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_73),
.Y(n_141)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_142),
.B(n_144),
.Y(n_197)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_80),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_106),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_146),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_68),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_147),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_73),
.B(n_10),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_71),
.B(n_12),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_74),
.A2(n_44),
.B1(n_4),
.B2(n_5),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_93),
.B(n_3),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_89),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_152),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_155),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_83),
.B(n_3),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_158),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_97),
.B(n_3),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_157),
.A2(n_111),
.B1(n_99),
.B2(n_76),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_115),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_72),
.Y(n_159)
);

OA22x2_ASAP7_75t_L g173 ( 
.A1(n_159),
.A2(n_86),
.B1(n_72),
.B2(n_109),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_116),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_161),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_89),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_L g163 ( 
.A1(n_102),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_163)
);

O2A1O1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_92),
.B(n_6),
.C(n_4),
.Y(n_177)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_135),
.A2(n_69),
.B1(n_102),
.B2(n_86),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_168),
.A2(n_176),
.B1(n_184),
.B2(n_159),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_170),
.A2(n_182),
.B(n_198),
.Y(n_220)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_160),
.A2(n_92),
.B1(n_68),
.B2(n_111),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_177),
.A2(n_146),
.B1(n_138),
.B2(n_152),
.Y(n_222)
);

OA22x2_ASAP7_75t_L g180 ( 
.A1(n_134),
.A2(n_78),
.B1(n_84),
.B2(n_96),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_195),
.B1(n_200),
.B2(n_159),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_6),
.B(n_84),
.Y(n_182)
);

BUFx8_ASAP7_75t_L g183 ( 
.A(n_119),
.Y(n_183)
);

INVx13_ASAP7_75t_L g235 ( 
.A(n_183),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_129),
.B(n_96),
.C(n_71),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_189),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_78),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_130),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_120),
.B(n_154),
.C(n_122),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_122),
.C(n_144),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_203),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_157),
.A2(n_126),
.B1(n_162),
.B2(n_163),
.Y(n_198)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_132),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_147),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_157),
.A2(n_140),
.B1(n_145),
.B2(n_136),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_125),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_202),
.B(n_153),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_158),
.B(n_125),
.C(n_131),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_204),
.A2(n_205),
.B1(n_231),
.B2(n_176),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_187),
.A2(n_131),
.B1(n_161),
.B2(n_136),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_206),
.A2(n_173),
.B1(n_201),
.B2(n_199),
.Y(n_256)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_209),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_183),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_212),
.B(n_228),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_121),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_214),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_118),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_183),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_215),
.B(n_217),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_142),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_177),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_218),
.B(n_221),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_172),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_222),
.A2(n_182),
.B(n_170),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_178),
.B(n_119),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_229),
.C(n_234),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_224),
.B(n_225),
.Y(n_249)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_227),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_166),
.B(n_130),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_178),
.B(n_186),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_171),
.B(n_141),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_233),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_185),
.A2(n_184),
.B1(n_188),
.B2(n_168),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_203),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_232),
.B(n_236),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_190),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_189),
.B(n_185),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_173),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_238),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_209),
.B(n_191),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_241),
.B(n_246),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_245),
.A2(n_251),
.B1(n_256),
.B2(n_262),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_225),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_174),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_247),
.B(n_253),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_231),
.A2(n_198),
.B1(n_180),
.B2(n_174),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_180),
.Y(n_253)
);

AOI221xp5_ASAP7_75t_L g254 ( 
.A1(n_220),
.A2(n_180),
.B1(n_179),
.B2(n_165),
.C(n_169),
.Y(n_254)
);

OAI322xp33_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_221),
.A3(n_232),
.B1(n_218),
.B2(n_219),
.C1(n_216),
.C2(n_222),
.Y(n_268)
);

MAJx2_ASAP7_75t_L g255 ( 
.A(n_220),
.B(n_165),
.C(n_169),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_255),
.B(n_204),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_208),
.B(n_192),
.Y(n_258)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_258),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_215),
.B(n_167),
.Y(n_259)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_226),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_262),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_236),
.A2(n_173),
.B(n_175),
.Y(n_262)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_264),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_246),
.Y(n_287)
);

NAND3xp33_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_257),
.C(n_242),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_216),
.C(n_219),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_286),
.C(n_255),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_271),
.A2(n_274),
.B1(n_277),
.B2(n_279),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_249),
.B(n_205),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_275),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_245),
.A2(n_207),
.B1(n_227),
.B2(n_175),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_242),
.B(n_210),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_239),
.A2(n_207),
.B1(n_235),
.B2(n_210),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_239),
.B(n_253),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_278),
.A2(n_263),
.B(n_240),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_240),
.A2(n_241),
.B1(n_251),
.B2(n_238),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_248),
.Y(n_281)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_244),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_284),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_252),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_249),
.B(n_237),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_263),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_247),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_291),
.Y(n_307)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_288),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_266),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_299),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_255),
.C(n_243),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_302),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_266),
.B(n_237),
.Y(n_297)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_297),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_298),
.Y(n_311)
);

NAND3xp33_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_250),
.C(n_243),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_276),
.A2(n_256),
.B1(n_250),
.B2(n_244),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_300),
.A2(n_274),
.B1(n_271),
.B2(n_277),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_264),
.Y(n_301)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_301),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_273),
.C(n_282),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_284),
.Y(n_305)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_305),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_295),
.A2(n_278),
.B1(n_276),
.B2(n_300),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_312),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_295),
.A2(n_278),
.B1(n_279),
.B2(n_265),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_296),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_303),
.A2(n_292),
.B(n_289),
.Y(n_315)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_315),
.Y(n_325)
);

INVx11_ASAP7_75t_L g317 ( 
.A(n_309),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_313),
.Y(n_326)
);

AOI31xp67_ASAP7_75t_L g318 ( 
.A1(n_308),
.A2(n_290),
.A3(n_287),
.B(n_282),
.Y(n_318)
);

O2A1O1Ixp33_ASAP7_75t_SL g328 ( 
.A1(n_318),
.A2(n_323),
.B(n_273),
.C(n_310),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_314),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_306),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_320),
.B(n_322),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_270),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_306),
.A2(n_293),
.B1(n_291),
.B2(n_302),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_324),
.A2(n_328),
.B(n_323),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_326),
.B(n_321),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_324),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_330),
.B(n_331),
.C(n_327),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_325),
.A2(n_318),
.B1(n_311),
.B2(n_316),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_333),
.C(n_319),
.Y(n_334)
);

OAI321xp33_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_307),
.A3(n_310),
.B1(n_312),
.B2(n_317),
.C(n_329),
.Y(n_335)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_335),
.Y(n_336)
);


endmodule