module fake_jpeg_23788_n_43 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_37;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx8_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

BUFx5_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_1),
.B(n_2),
.Y(n_9)
);

BUFx8_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_9),
.B(n_4),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_17),
.A2(n_18),
.B(n_19),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g18 ( 
.A1(n_7),
.A2(n_4),
.B1(n_5),
.B2(n_14),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_L g19 ( 
.A1(n_7),
.A2(n_14),
.B1(n_11),
.B2(n_8),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_13),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_23),
.Y(n_33)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx24_ASAP7_75t_SL g30 ( 
.A(n_24),
.Y(n_30)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_10),
.B(n_9),
.C(n_13),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_27),
.B(n_25),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_30),
.C(n_26),
.Y(n_38)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_35),
.B(n_36),
.Y(n_37)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_10),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_29),
.Y(n_39)
);

AOI31xp67_ASAP7_75t_SL g41 ( 
.A1(n_39),
.A2(n_40),
.A3(n_18),
.B(n_24),
.Y(n_41)
);

AOI21xp33_ASAP7_75t_L g42 ( 
.A1(n_41),
.A2(n_32),
.B(n_28),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_19),
.C(n_22),
.Y(n_43)
);


endmodule