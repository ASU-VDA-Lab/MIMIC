module fake_jpeg_19296_n_157 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_157);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_157;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_6),
.B(n_18),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_9),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_2),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_4),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_12),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_48),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_25),
.C(n_43),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_66),
.Y(n_88)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_46),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_75),
.B(n_54),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_87),
.Y(n_94)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_88),
.Y(n_105)
);

AOI21xp33_ASAP7_75t_SL g91 ( 
.A1(n_78),
.A2(n_74),
.B(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_92),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_68),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_104),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_90),
.A2(n_55),
.B1(n_61),
.B2(n_72),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_100),
.B(n_62),
.C(n_60),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_84),
.A2(n_47),
.B1(n_54),
.B2(n_68),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_74),
.B1(n_59),
.B2(n_63),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_102),
.A2(n_71),
.B1(n_70),
.B2(n_69),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVxp33_ASAP7_75t_SL g106 ( 
.A(n_97),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_57),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_109),
.A2(n_119),
.B(n_53),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_59),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_113),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_102),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_120),
.B1(n_121),
.B2(n_58),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_67),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_117),
.Y(n_130)
);

INVxp33_ASAP7_75t_SL g116 ( 
.A(n_99),
.Y(n_116)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_98),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_65),
.B1(n_52),
.B2(n_4),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_57),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g125 ( 
.A1(n_118),
.A2(n_56),
.B1(n_28),
.B2(n_44),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_125),
.A2(n_127),
.B1(n_110),
.B2(n_3),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_110),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_128),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_24),
.B1(n_42),
.B2(n_41),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_108),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_131),
.B(n_133),
.Y(n_136)
);

OAI32xp33_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_20),
.A3(n_37),
.B1(n_34),
.B2(n_32),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_107),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_134),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

INVxp33_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_129),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_141),
.A2(n_130),
.B1(n_127),
.B2(n_132),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_125),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_146),
.B(n_145),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_136),
.B(n_138),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_135),
.B(n_144),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_132),
.C(n_142),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_140),
.Y(n_152)
);

NOR3xp33_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_140),
.C(n_135),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_124),
.C(n_5),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_21),
.B(n_38),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_155),
.A2(n_19),
.B(n_30),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_10),
.Y(n_157)
);


endmodule