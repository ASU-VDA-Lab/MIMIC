module fake_netlist_6_383_n_1681 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1681);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1681;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_110),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_54),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_43),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_2),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_124),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_155),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_102),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_67),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_45),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_35),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_88),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_120),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_145),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_144),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_39),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_56),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_147),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_85),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_83),
.Y(n_183)
);

BUFx10_ASAP7_75t_L g184 ( 
.A(n_105),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_89),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_133),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_68),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_9),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_1),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_72),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_139),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_17),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_5),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_96),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_29),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_43),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_61),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_5),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_2),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_127),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_162),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_100),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_135),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_81),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_87),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_103),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_4),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_156),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_9),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_79),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_76),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_134),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_39),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_160),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_42),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_95),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_16),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_0),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_116),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_77),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_70),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_18),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_157),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_20),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_37),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_10),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_18),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_53),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_66),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_29),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_11),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_117),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_42),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_49),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_65),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_31),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_71),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_136),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_163),
.Y(n_239)
);

BUFx8_ASAP7_75t_SL g240 ( 
.A(n_108),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_32),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_114),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_109),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_24),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_40),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_122),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_58),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_101),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_21),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_28),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_24),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_33),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_16),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_28),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_90),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_130),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_17),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_63),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_4),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_69),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_115),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_3),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_44),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_149),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_158),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_148),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_154),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_86),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_33),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_11),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_91),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_6),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_137),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_132),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_57),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_153),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_47),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_22),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_52),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_112),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_152),
.Y(n_281)
);

BUFx2_ASAP7_75t_SL g282 ( 
.A(n_12),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_20),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_26),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_23),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_118),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_14),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_1),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_150),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_30),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_37),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_30),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_12),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_106),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_97),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_13),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_99),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_21),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_146),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_142),
.Y(n_300)
);

BUFx2_ASAP7_75t_SL g301 ( 
.A(n_31),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_51),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_113),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_138),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_27),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_6),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_80),
.Y(n_307)
);

BUFx10_ASAP7_75t_L g308 ( 
.A(n_129),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_123),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_82),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_125),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_107),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_73),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_119),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_46),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_151),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_44),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_131),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_111),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_13),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_121),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_159),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_32),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_47),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_64),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_60),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_23),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_74),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_169),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_263),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_263),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_L g332 ( 
.A(n_195),
.B(n_0),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_240),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_189),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_195),
.B(n_3),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_263),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_263),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_263),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_197),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_298),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_177),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_200),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_302),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_201),
.Y(n_344)
);

NOR2xp67_ASAP7_75t_L g345 ( 
.A(n_257),
.B(n_7),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_202),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_298),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_307),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_203),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_298),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_298),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_204),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_214),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_298),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_205),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_206),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_216),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_208),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_199),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_210),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_211),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_221),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_199),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_228),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_217),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_189),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_217),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_253),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_253),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_192),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_166),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_229),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_237),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_238),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_242),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_167),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_246),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_194),
.Y(n_378)
);

INVxp33_ASAP7_75t_SL g379 ( 
.A(n_192),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_258),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_261),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_173),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_264),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_174),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_265),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_266),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_218),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_233),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_254),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_259),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_R g391 ( 
.A(n_267),
.B(n_50),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_272),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_268),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_215),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_278),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_283),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_290),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_293),
.Y(n_398)
);

NOR2xp67_ASAP7_75t_L g399 ( 
.A(n_257),
.B(n_7),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_271),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_273),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_305),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_281),
.Y(n_403)
);

INVxp33_ASAP7_75t_SL g404 ( 
.A(n_193),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_247),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_289),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_315),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_317),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_248),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_219),
.B(n_8),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_330),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_330),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_329),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_331),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_410),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_334),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_337),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_337),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_340),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_339),
.B(n_342),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_344),
.B(n_280),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_331),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_336),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_340),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_360),
.Y(n_425)
);

INVx5_ASAP7_75t_L g426 ( 
.A(n_347),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_336),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_338),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_346),
.B(n_279),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_338),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_350),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_361),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_350),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_394),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_351),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_351),
.Y(n_436)
);

NOR2xp67_ASAP7_75t_L g437 ( 
.A(n_349),
.B(n_190),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_352),
.B(n_219),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_378),
.A2(n_405),
.B1(n_409),
.B2(n_353),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_354),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_364),
.Y(n_441)
);

NAND2xp33_ASAP7_75t_L g442 ( 
.A(n_335),
.B(n_193),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_380),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_347),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_381),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_341),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_354),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_376),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_385),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_376),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_359),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_343),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_371),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_371),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_355),
.B(n_279),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_366),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_359),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_363),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_363),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_365),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_365),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_370),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_382),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_382),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_384),
.Y(n_465)
);

AND2x6_ASAP7_75t_L g466 ( 
.A(n_335),
.B(n_303),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_356),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_357),
.B(n_184),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_332),
.B(n_300),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_348),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_367),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_367),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_368),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_386),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_358),
.Y(n_475)
);

INVx4_ASAP7_75t_L g476 ( 
.A(n_362),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_368),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_372),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_384),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_369),
.Y(n_480)
);

OAI21x1_ASAP7_75t_L g481 ( 
.A1(n_369),
.A2(n_239),
.B(n_223),
.Y(n_481)
);

NOR2xp67_ASAP7_75t_L g482 ( 
.A(n_373),
.B(n_300),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_387),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_387),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_412),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_482),
.B(n_374),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_429),
.B(n_375),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_415),
.B(n_484),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_455),
.B(n_377),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_440),
.Y(n_490)
);

BUFx4f_ASAP7_75t_L g491 ( 
.A(n_466),
.Y(n_491)
);

INVx4_ASAP7_75t_L g492 ( 
.A(n_411),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_414),
.Y(n_493)
);

INVx5_ASAP7_75t_L g494 ( 
.A(n_466),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_438),
.B(n_383),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_469),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_484),
.B(n_388),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_411),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_411),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_417),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_414),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_434),
.Y(n_502)
);

BUFx4f_ASAP7_75t_L g503 ( 
.A(n_466),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_469),
.A2(n_399),
.B1(n_345),
.B2(n_332),
.Y(n_504)
);

NAND2xp33_ASAP7_75t_L g505 ( 
.A(n_466),
.B(n_303),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_484),
.B(n_408),
.Y(n_506)
);

NAND2xp33_ASAP7_75t_SL g507 ( 
.A(n_469),
.B(n_277),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_417),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g509 ( 
.A1(n_469),
.A2(n_345),
.B1(n_399),
.B2(n_277),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_481),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_425),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_453),
.B(n_388),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_462),
.B(n_393),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_425),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_422),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_442),
.A2(n_379),
.B1(n_404),
.B2(n_323),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_419),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_421),
.B(n_400),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_419),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_447),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_420),
.B(n_401),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_437),
.B(n_403),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_447),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_466),
.A2(n_324),
.B1(n_282),
.B2(n_301),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_416),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_416),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_411),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_481),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_422),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_453),
.B(n_408),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_454),
.Y(n_531)
);

AND2x6_ASAP7_75t_L g532 ( 
.A(n_454),
.B(n_223),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_466),
.B(n_406),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_476),
.B(n_462),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_476),
.B(n_333),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_418),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_423),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_418),
.Y(n_538)
);

INVx6_ASAP7_75t_L g539 ( 
.A(n_418),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_466),
.B(n_212),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_423),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_418),
.Y(n_542)
);

OR2x6_ASAP7_75t_L g543 ( 
.A(n_467),
.B(n_179),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_463),
.B(n_407),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_427),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_418),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_463),
.Y(n_547)
);

INVx4_ASAP7_75t_SL g548 ( 
.A(n_424),
.Y(n_548)
);

AND2x6_ASAP7_75t_L g549 ( 
.A(n_464),
.B(n_239),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_476),
.B(n_456),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_427),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_439),
.B(n_391),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_432),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_424),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_468),
.A2(n_226),
.B1(n_292),
.B2(n_291),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_475),
.A2(n_309),
.B1(n_328),
.B2(n_187),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_428),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_464),
.B(n_389),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_428),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_430),
.B(n_235),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_424),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_465),
.B(n_243),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_430),
.B(n_260),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_431),
.B(n_294),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_431),
.B(n_256),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_444),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_444),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_465),
.B(n_479),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_444),
.Y(n_569)
);

AND2x6_ASAP7_75t_L g570 ( 
.A(n_479),
.B(n_256),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_433),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_433),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_444),
.Y(n_573)
);

CKINVDCx6p67_ASAP7_75t_R g574 ( 
.A(n_478),
.Y(n_574)
);

AND2x6_ASAP7_75t_L g575 ( 
.A(n_435),
.B(n_275),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_444),
.Y(n_576)
);

INVxp67_ASAP7_75t_SL g577 ( 
.A(n_435),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_432),
.B(n_184),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_436),
.B(n_451),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_436),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_451),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_426),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_451),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_451),
.B(n_275),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_451),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_483),
.A2(n_318),
.B1(n_303),
.B2(n_398),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_457),
.B(n_389),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_448),
.A2(n_318),
.B1(n_303),
.B2(n_407),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_446),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_413),
.B(n_188),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_460),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_460),
.B(n_170),
.Y(n_592)
);

BUFx10_ASAP7_75t_L g593 ( 
.A(n_441),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_460),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_460),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_441),
.A2(n_181),
.B1(n_297),
.B2(n_187),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_460),
.B(n_175),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_471),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_448),
.B(n_164),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_461),
.B(n_164),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_471),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_461),
.A2(n_303),
.B1(n_398),
.B2(n_397),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_471),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_471),
.Y(n_604)
);

BUFx10_ASAP7_75t_L g605 ( 
.A(n_443),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_461),
.B(n_390),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_472),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_472),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_477),
.A2(n_402),
.B1(n_397),
.B2(n_396),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_457),
.B(n_402),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_477),
.A2(n_396),
.B1(n_395),
.B2(n_392),
.Y(n_611)
);

INVx1_ASAP7_75t_SL g612 ( 
.A(n_443),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_472),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_472),
.Y(n_614)
);

BUFx8_ASAP7_75t_SL g615 ( 
.A(n_452),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_477),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_458),
.B(n_459),
.Y(n_617)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_426),
.Y(n_618)
);

OR2x6_ASAP7_75t_L g619 ( 
.A(n_458),
.B(n_390),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_445),
.B(n_184),
.Y(n_620)
);

INVxp67_ASAP7_75t_SL g621 ( 
.A(n_473),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_480),
.B(n_180),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_450),
.A2(n_395),
.B1(n_392),
.B2(n_286),
.Y(n_623)
);

INVxp67_ASAP7_75t_SL g624 ( 
.A(n_480),
.Y(n_624)
);

INVx5_ASAP7_75t_L g625 ( 
.A(n_426),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_450),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_513),
.B(n_262),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_502),
.B(n_445),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_568),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_485),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_496),
.B(n_191),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_491),
.B(n_220),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_491),
.B(n_234),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_488),
.B(n_255),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_491),
.B(n_274),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_488),
.A2(n_276),
.B(n_295),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_525),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_487),
.B(n_299),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_513),
.B(n_270),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_568),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_489),
.B(n_313),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_504),
.B(n_325),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_495),
.B(n_165),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_510),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_525),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_503),
.B(n_168),
.Y(n_646)
);

OAI21xp5_ASAP7_75t_L g647 ( 
.A1(n_503),
.A2(n_186),
.B(n_168),
.Y(n_647)
);

INVx2_ASAP7_75t_SL g648 ( 
.A(n_526),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_577),
.B(n_171),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_621),
.B(n_171),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_530),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_510),
.A2(n_224),
.B1(n_227),
.B2(n_250),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_624),
.B(n_172),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_600),
.B(n_172),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_606),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_SL g656 ( 
.A1(n_514),
.A2(n_269),
.B1(n_470),
.B2(n_449),
.Y(n_656)
);

NAND2xp33_ASAP7_75t_L g657 ( 
.A(n_533),
.B(n_176),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_530),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_485),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_526),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_521),
.B(n_176),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_580),
.B(n_178),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_528),
.A2(n_306),
.B1(n_320),
.B2(n_327),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_518),
.B(n_178),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_552),
.B(n_181),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_550),
.B(n_182),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_580),
.B(n_182),
.Y(n_667)
);

NOR2xp67_ASAP7_75t_L g668 ( 
.A(n_556),
.B(n_449),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_590),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_534),
.B(n_183),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_503),
.B(n_183),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_540),
.A2(n_311),
.B1(n_328),
.B2(n_326),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_494),
.B(n_185),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_531),
.B(n_185),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_494),
.B(n_186),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_615),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_547),
.B(n_297),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_494),
.B(n_304),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_490),
.B(n_493),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_544),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_494),
.B(n_304),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_590),
.Y(n_682)
);

OR2x6_ASAP7_75t_L g683 ( 
.A(n_589),
.B(n_474),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_490),
.B(n_309),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_493),
.B(n_310),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_501),
.B(n_310),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_L g687 ( 
.A1(n_516),
.A2(n_311),
.B1(n_312),
.B2(n_314),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_501),
.B(n_515),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_544),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_522),
.B(n_312),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_615),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_515),
.B(n_314),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_562),
.B(n_474),
.Y(n_693)
);

NOR2xp67_ASAP7_75t_L g694 ( 
.A(n_596),
.B(n_316),
.Y(n_694)
);

INVx4_ASAP7_75t_L g695 ( 
.A(n_494),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_616),
.B(n_316),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_529),
.B(n_319),
.Y(n_697)
);

OAI221xp5_ASAP7_75t_L g698 ( 
.A1(n_509),
.A2(n_251),
.B1(n_198),
.B2(n_207),
.C(n_209),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_528),
.A2(n_306),
.B1(n_327),
.B2(n_320),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_626),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_543),
.A2(n_326),
.B1(n_322),
.B2(n_321),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_512),
.B(n_213),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_529),
.B(n_322),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_616),
.B(n_321),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_500),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_524),
.A2(n_319),
.B1(n_245),
.B2(n_244),
.Y(n_706)
);

OAI221xp5_ASAP7_75t_L g707 ( 
.A1(n_609),
.A2(n_249),
.B1(n_222),
.B2(n_296),
.C(n_288),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_587),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_564),
.B(n_196),
.Y(n_709)
);

NAND2xp33_ASAP7_75t_L g710 ( 
.A(n_532),
.B(n_241),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_508),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_543),
.B(n_225),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_537),
.B(n_426),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_512),
.B(n_558),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_587),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_610),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_497),
.A2(n_252),
.B1(n_231),
.B2(n_287),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_512),
.B(n_230),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_508),
.Y(n_719)
);

OR2x6_ASAP7_75t_L g720 ( 
.A(n_589),
.B(n_308),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_541),
.B(n_285),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_610),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_606),
.Y(n_723)
);

AND2x6_ASAP7_75t_SL g724 ( 
.A(n_543),
.B(n_284),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_545),
.B(n_236),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_543),
.B(n_8),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_560),
.B(n_308),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_619),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_619),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_517),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_563),
.B(n_308),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_517),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_519),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_545),
.B(n_551),
.Y(n_734)
);

INVx5_ASAP7_75t_L g735 ( 
.A(n_575),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_551),
.B(n_232),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_557),
.B(n_232),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_581),
.B(n_232),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_586),
.A2(n_59),
.B1(n_143),
.B2(n_141),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_606),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_581),
.B(n_48),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_583),
.B(n_55),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_557),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_559),
.B(n_161),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_559),
.B(n_140),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_555),
.B(n_10),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_571),
.B(n_128),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_571),
.B(n_126),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_519),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_619),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_514),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_497),
.A2(n_14),
.B1(n_15),
.B2(n_19),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_506),
.A2(n_15),
.B1(n_19),
.B2(n_22),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_617),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_602),
.A2(n_62),
.B1(n_94),
.B2(n_93),
.Y(n_755)
);

OR2x6_ASAP7_75t_L g756 ( 
.A(n_535),
.B(n_25),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_558),
.B(n_25),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_572),
.B(n_98),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_520),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_572),
.B(n_92),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_523),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_486),
.B(n_26),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_617),
.B(n_506),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_578),
.B(n_27),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_599),
.B(n_84),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_511),
.B(n_34),
.Y(n_766)
);

O2A1O1Ixp33_ASAP7_75t_L g767 ( 
.A1(n_565),
.A2(n_34),
.B(n_35),
.C(n_36),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_583),
.B(n_78),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_507),
.A2(n_620),
.B1(n_619),
.B2(n_549),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_585),
.B(n_594),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_579),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_585),
.B(n_75),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_527),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_612),
.B(n_36),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_507),
.B(n_38),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_538),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_591),
.B(n_38),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_538),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_532),
.A2(n_40),
.B1(n_41),
.B2(n_45),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_627),
.B(n_553),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_627),
.B(n_605),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_763),
.A2(n_505),
.B(n_492),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_695),
.A2(n_505),
.B(n_492),
.Y(n_783)
);

OR2x6_ASAP7_75t_L g784 ( 
.A(n_683),
.B(n_574),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_639),
.B(n_553),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_639),
.B(n_605),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_634),
.A2(n_576),
.B(n_566),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_771),
.B(n_595),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_770),
.A2(n_576),
.B(n_566),
.Y(n_789)
);

AO21x1_ASAP7_75t_L g790 ( 
.A1(n_765),
.A2(n_584),
.B(n_597),
.Y(n_790)
);

A2O1A1Ixp33_ASAP7_75t_L g791 ( 
.A1(n_665),
.A2(n_622),
.B(n_592),
.C(n_603),
.Y(n_791)
);

AOI21x1_ASAP7_75t_L g792 ( 
.A1(n_713),
.A2(n_613),
.B(n_598),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_754),
.A2(n_527),
.B(n_546),
.Y(n_793)
);

OAI21xp5_ASAP7_75t_L g794 ( 
.A1(n_632),
.A2(n_613),
.B(n_598),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_754),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_629),
.B(n_601),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_640),
.B(n_601),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_723),
.Y(n_798)
);

OAI321xp33_ASAP7_75t_L g799 ( 
.A1(n_746),
.A2(n_623),
.A3(n_611),
.B1(n_588),
.B2(n_614),
.C(n_591),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_750),
.B(n_593),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_645),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_693),
.B(n_593),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_643),
.B(n_569),
.Y(n_803)
);

INVx1_ASAP7_75t_SL g804 ( 
.A(n_628),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_643),
.B(n_569),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_638),
.B(n_569),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_740),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_655),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_750),
.B(n_605),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_641),
.B(n_554),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_735),
.A2(n_546),
.B(n_561),
.Y(n_811)
);

AOI21xp33_ASAP7_75t_L g812 ( 
.A1(n_665),
.A2(n_607),
.B(n_614),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_666),
.B(n_554),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_632),
.A2(n_608),
.B(n_607),
.Y(n_814)
);

A2O1A1Ixp33_ASAP7_75t_L g815 ( 
.A1(n_727),
.A2(n_604),
.B(n_608),
.C(n_542),
.Y(n_815)
);

BUFx4f_ASAP7_75t_L g816 ( 
.A(n_750),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_752),
.A2(n_574),
.B1(n_573),
.B2(n_542),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_L g818 ( 
.A1(n_633),
.A2(n_635),
.B(n_636),
.Y(n_818)
);

A2O1A1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_727),
.A2(n_604),
.B(n_573),
.C(n_561),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_669),
.B(n_593),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_666),
.B(n_536),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_700),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_709),
.B(n_536),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_709),
.B(n_661),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_679),
.A2(n_734),
.B(n_688),
.Y(n_825)
);

CKINVDCx10_ASAP7_75t_R g826 ( 
.A(n_683),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_633),
.A2(n_498),
.B(n_499),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_635),
.A2(n_498),
.B(n_499),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_644),
.Y(n_829)
);

AOI21x1_ASAP7_75t_L g830 ( 
.A1(n_673),
.A2(n_539),
.B(n_548),
.Y(n_830)
);

AO21x1_ASAP7_75t_L g831 ( 
.A1(n_746),
.A2(n_570),
.B(n_549),
.Y(n_831)
);

NAND3xp33_ASAP7_75t_SL g832 ( 
.A(n_652),
.B(n_532),
.C(n_570),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_743),
.B(n_570),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_644),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_752),
.A2(n_536),
.B1(n_567),
.B2(n_539),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_651),
.B(n_570),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_773),
.A2(n_567),
.B(n_582),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_682),
.B(n_637),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_658),
.B(n_680),
.Y(n_839)
);

INVx1_ASAP7_75t_SL g840 ( 
.A(n_648),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_689),
.B(n_570),
.Y(n_841)
);

INVx4_ASAP7_75t_L g842 ( 
.A(n_644),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_660),
.B(n_567),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_753),
.A2(n_539),
.B1(n_532),
.B2(n_549),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_708),
.B(n_549),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_714),
.A2(n_549),
.B1(n_570),
.B2(n_532),
.Y(n_846)
);

O2A1O1Ixp5_ASAP7_75t_L g847 ( 
.A1(n_631),
.A2(n_671),
.B(n_646),
.C(n_654),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_773),
.A2(n_582),
.B(n_618),
.Y(n_848)
);

CKINVDCx10_ASAP7_75t_R g849 ( 
.A(n_683),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_773),
.A2(n_582),
.B(n_618),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_630),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_646),
.A2(n_618),
.B(n_625),
.Y(n_852)
);

OR2x2_ASAP7_75t_L g853 ( 
.A(n_652),
.B(n_41),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_715),
.B(n_549),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_664),
.B(n_539),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_671),
.A2(n_625),
.B(n_548),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_716),
.A2(n_575),
.B(n_625),
.Y(n_857)
);

OAI321xp33_ASAP7_75t_L g858 ( 
.A1(n_753),
.A2(n_46),
.A3(n_548),
.B1(n_575),
.B2(n_625),
.C(n_764),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_631),
.A2(n_575),
.B(n_657),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_722),
.A2(n_575),
.B(n_647),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_664),
.A2(n_575),
.B1(n_731),
.B2(n_690),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_659),
.Y(n_862)
);

INVx1_ASAP7_75t_SL g863 ( 
.A(n_751),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_644),
.B(n_757),
.Y(n_864)
);

NOR2xp67_ASAP7_75t_L g865 ( 
.A(n_731),
.B(n_670),
.Y(n_865)
);

CKINVDCx16_ASAP7_75t_R g866 ( 
.A(n_656),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_776),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_690),
.A2(n_769),
.B1(n_670),
.B2(n_762),
.Y(n_868)
);

AOI21x1_ASAP7_75t_L g869 ( 
.A1(n_673),
.A2(n_678),
.B(n_675),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_779),
.A2(n_699),
.B1(n_663),
.B2(n_717),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_650),
.A2(n_653),
.B(n_778),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_642),
.B(n_649),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_712),
.B(n_701),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_772),
.A2(n_745),
.B(n_758),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_744),
.A2(n_748),
.B(n_760),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_721),
.B(n_725),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_747),
.A2(n_662),
.B(n_667),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_676),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_762),
.B(n_764),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_759),
.A2(n_761),
.B(n_681),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_779),
.A2(n_663),
.B1(n_699),
.B2(n_717),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_696),
.A2(n_704),
.B(n_681),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_775),
.A2(n_756),
.B1(n_698),
.B2(n_726),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_SL g884 ( 
.A(n_691),
.B(n_668),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_675),
.A2(n_678),
.B(n_705),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_685),
.B(n_703),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_696),
.A2(n_704),
.B1(n_718),
.B2(n_702),
.Y(n_887)
);

AO32x2_ASAP7_75t_L g888 ( 
.A1(n_755),
.A2(n_739),
.A3(n_687),
.B1(n_706),
.B2(n_777),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_686),
.B(n_692),
.Y(n_889)
);

BUFx2_ASAP7_75t_L g890 ( 
.A(n_766),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_712),
.A2(n_672),
.B1(n_697),
.B2(n_684),
.Y(n_891)
);

A2O1A1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_775),
.A2(n_737),
.B(n_736),
.C(n_694),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_711),
.A2(n_732),
.B(n_730),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_719),
.A2(n_733),
.B(n_749),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_777),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_774),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_674),
.A2(n_677),
.B(n_729),
.C(n_728),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_756),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_741),
.A2(n_742),
.B(n_768),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_710),
.A2(n_738),
.B1(n_756),
.B2(n_707),
.Y(n_900)
);

A2O1A1Ixp33_ASAP7_75t_L g901 ( 
.A1(n_738),
.A2(n_767),
.B(n_724),
.C(n_720),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_720),
.A2(n_503),
.B(n_491),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_720),
.B(n_488),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_763),
.A2(n_503),
.B(n_491),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_637),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_655),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_627),
.B(n_502),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_643),
.B(n_488),
.Y(n_908)
);

A2O1A1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_665),
.A2(n_643),
.B(n_731),
.C(n_727),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_754),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_643),
.B(n_488),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_750),
.B(n_502),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_754),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_628),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_750),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_763),
.B(n_488),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_763),
.A2(n_503),
.B(n_491),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_750),
.B(n_502),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_754),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_627),
.B(n_502),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_752),
.A2(n_753),
.B1(n_779),
.B2(n_504),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_627),
.B(n_502),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_763),
.A2(n_503),
.B(n_491),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_665),
.A2(n_643),
.B(n_731),
.C(n_727),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_750),
.B(n_502),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_763),
.A2(n_503),
.B(n_491),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_763),
.B(n_488),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_754),
.Y(n_928)
);

AND2x6_ASAP7_75t_SL g929 ( 
.A(n_683),
.B(n_628),
.Y(n_929)
);

NOR2xp67_ASAP7_75t_L g930 ( 
.A(n_682),
.B(n_476),
.Y(n_930)
);

AO21x1_ASAP7_75t_L g931 ( 
.A1(n_765),
.A2(n_641),
.B(n_638),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_763),
.A2(n_503),
.B(n_491),
.Y(n_932)
);

AND2x2_ASAP7_75t_SL g933 ( 
.A(n_652),
.B(n_413),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_763),
.A2(n_503),
.B(n_491),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_754),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_754),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_754),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_655),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_763),
.B(n_488),
.Y(n_939)
);

BUFx2_ASAP7_75t_L g940 ( 
.A(n_637),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_643),
.B(n_488),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_763),
.B(n_488),
.Y(n_942)
);

O2A1O1Ixp5_ASAP7_75t_L g943 ( 
.A1(n_638),
.A2(n_641),
.B(n_633),
.C(n_635),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_915),
.B(n_800),
.Y(n_944)
);

OAI21xp33_ASAP7_75t_L g945 ( 
.A1(n_870),
.A2(n_881),
.B(n_921),
.Y(n_945)
);

OAI21x1_ASAP7_75t_L g946 ( 
.A1(n_880),
.A2(n_830),
.B(n_828),
.Y(n_946)
);

NAND2x1p5_ASAP7_75t_L g947 ( 
.A(n_816),
.B(n_915),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_916),
.A2(n_939),
.B(n_927),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_824),
.B(n_908),
.Y(n_949)
);

OAI21x1_ASAP7_75t_L g950 ( 
.A1(n_827),
.A2(n_789),
.B(n_792),
.Y(n_950)
);

AOI21xp33_ASAP7_75t_L g951 ( 
.A1(n_870),
.A2(n_881),
.B(n_921),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_909),
.A2(n_924),
.B(n_916),
.Y(n_952)
);

AO21x2_ASAP7_75t_L g953 ( 
.A1(n_790),
.A2(n_818),
.B(n_812),
.Y(n_953)
);

OA21x2_ASAP7_75t_L g954 ( 
.A1(n_819),
.A2(n_815),
.B(n_847),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_927),
.A2(n_942),
.B(n_939),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_915),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_822),
.Y(n_957)
);

OAI21xp33_ASAP7_75t_L g958 ( 
.A1(n_873),
.A2(n_922),
.B(n_879),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_940),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_942),
.A2(n_825),
.B(n_874),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_868),
.A2(n_865),
.B(n_861),
.C(n_876),
.Y(n_961)
);

NAND2x1p5_ASAP7_75t_L g962 ( 
.A(n_816),
.B(n_842),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_907),
.B(n_920),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_878),
.Y(n_964)
);

AOI21x1_ASAP7_75t_L g965 ( 
.A1(n_813),
.A2(n_821),
.B(n_823),
.Y(n_965)
);

OA21x2_ASAP7_75t_L g966 ( 
.A1(n_794),
.A2(n_812),
.B(n_943),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_875),
.A2(n_917),
.B(n_904),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_781),
.B(n_804),
.Y(n_968)
);

BUFx10_ASAP7_75t_L g969 ( 
.A(n_802),
.Y(n_969)
);

AND3x2_ASAP7_75t_L g970 ( 
.A(n_786),
.B(n_785),
.C(n_780),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_914),
.Y(n_971)
);

AOI21x1_ASAP7_75t_SL g972 ( 
.A1(n_864),
.A2(n_872),
.B(n_886),
.Y(n_972)
);

INVxp33_ASAP7_75t_SL g973 ( 
.A(n_884),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_911),
.B(n_941),
.Y(n_974)
);

OAI21x1_ASAP7_75t_L g975 ( 
.A1(n_793),
.A2(n_787),
.B(n_934),
.Y(n_975)
);

BUFx4_ASAP7_75t_SL g976 ( 
.A(n_784),
.Y(n_976)
);

NOR2x1_ASAP7_75t_L g977 ( 
.A(n_930),
.B(n_842),
.Y(n_977)
);

CKINVDCx11_ASAP7_75t_R g978 ( 
.A(n_929),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_905),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_923),
.A2(n_932),
.B(n_926),
.Y(n_980)
);

INVx1_ASAP7_75t_SL g981 ( 
.A(n_863),
.Y(n_981)
);

CKINVDCx14_ASAP7_75t_R g982 ( 
.A(n_784),
.Y(n_982)
);

OAI21x1_ASAP7_75t_L g983 ( 
.A1(n_885),
.A2(n_814),
.B(n_899),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_891),
.B(n_795),
.Y(n_984)
);

NAND2x1_ASAP7_75t_L g985 ( 
.A(n_834),
.B(n_829),
.Y(n_985)
);

OAI22x1_ASAP7_75t_L g986 ( 
.A1(n_853),
.A2(n_900),
.B1(n_887),
.B2(n_890),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_877),
.A2(n_871),
.B(n_805),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_882),
.A2(n_892),
.B(n_883),
.C(n_858),
.Y(n_988)
);

NAND2x2_ASAP7_75t_L g989 ( 
.A(n_898),
.B(n_801),
.Y(n_989)
);

INVx6_ASAP7_75t_L g990 ( 
.A(n_784),
.Y(n_990)
);

NOR3xp33_ASAP7_75t_L g991 ( 
.A(n_883),
.B(n_901),
.C(n_903),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_809),
.B(n_798),
.Y(n_992)
);

OAI21x1_ASAP7_75t_L g993 ( 
.A1(n_811),
.A2(n_837),
.B(n_893),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_860),
.A2(n_782),
.B(n_791),
.Y(n_994)
);

OAI21x1_ASAP7_75t_L g995 ( 
.A1(n_894),
.A2(n_869),
.B(n_859),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_896),
.B(n_820),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_835),
.A2(n_841),
.B(n_836),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_840),
.Y(n_998)
);

INVx4_ASAP7_75t_L g999 ( 
.A(n_834),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_834),
.Y(n_1000)
);

OAI21x1_ASAP7_75t_L g1001 ( 
.A1(n_852),
.A2(n_856),
.B(n_857),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_803),
.A2(n_855),
.B(n_864),
.Y(n_1002)
);

INVx4_ASAP7_75t_L g1003 ( 
.A(n_829),
.Y(n_1003)
);

OAI21x1_ASAP7_75t_L g1004 ( 
.A1(n_783),
.A2(n_850),
.B(n_848),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_933),
.B(n_838),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_928),
.B(n_935),
.Y(n_1006)
);

OAI21x1_ASAP7_75t_L g1007 ( 
.A1(n_835),
.A2(n_788),
.B(n_796),
.Y(n_1007)
);

AO31x2_ASAP7_75t_L g1008 ( 
.A1(n_931),
.A2(n_831),
.A3(n_844),
.B(n_897),
.Y(n_1008)
);

AOI211x1_ASAP7_75t_L g1009 ( 
.A1(n_839),
.A2(n_936),
.B(n_913),
.C(n_919),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_806),
.A2(n_810),
.B(n_788),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_910),
.B(n_937),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_839),
.B(n_889),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_836),
.A2(n_841),
.B(n_807),
.C(n_845),
.Y(n_1013)
);

AO31x2_ASAP7_75t_L g1014 ( 
.A1(n_844),
.A2(n_817),
.A3(n_833),
.B(n_854),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_796),
.A2(n_797),
.B(n_833),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_895),
.A2(n_797),
.B1(n_846),
.B2(n_938),
.Y(n_1016)
);

OAI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_845),
.A2(n_854),
.B(n_817),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_895),
.B(n_843),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_895),
.B(n_938),
.Y(n_1019)
);

OAI22x1_ASAP7_75t_L g1020 ( 
.A1(n_912),
.A2(n_925),
.B1(n_918),
.B2(n_866),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_808),
.A2(n_906),
.B(n_832),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_808),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_906),
.A2(n_799),
.B(n_862),
.C(n_851),
.Y(n_1023)
);

AND2x4_ASAP7_75t_SL g1024 ( 
.A(n_867),
.B(n_826),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_867),
.B(n_888),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_888),
.B(n_849),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_SL g1027 ( 
.A1(n_888),
.A2(n_933),
.B1(n_921),
.B2(n_873),
.Y(n_1027)
);

O2A1O1Ixp5_ASAP7_75t_L g1028 ( 
.A1(n_909),
.A2(n_924),
.B(n_879),
.C(n_931),
.Y(n_1028)
);

OAI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_909),
.A2(n_924),
.B(n_916),
.Y(n_1029)
);

OR2x2_ASAP7_75t_L g1030 ( 
.A(n_907),
.B(n_502),
.Y(n_1030)
);

INVx5_ASAP7_75t_L g1031 ( 
.A(n_834),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_922),
.B(n_502),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_824),
.B(n_908),
.Y(n_1033)
);

AO31x2_ASAP7_75t_L g1034 ( 
.A1(n_790),
.A2(n_931),
.A3(n_815),
.B(n_819),
.Y(n_1034)
);

AND2x2_ASAP7_75t_SL g1035 ( 
.A(n_933),
.B(n_786),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_916),
.B(n_927),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_907),
.B(n_920),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_842),
.Y(n_1038)
);

OAI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_909),
.A2(n_924),
.B(n_916),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_916),
.A2(n_503),
.B(n_491),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_880),
.A2(n_830),
.B(n_828),
.Y(n_1041)
);

AND2x6_ASAP7_75t_L g1042 ( 
.A(n_834),
.B(n_915),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_915),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_916),
.A2(n_503),
.B(n_491),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_916),
.A2(n_503),
.B(n_491),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_916),
.A2(n_503),
.B(n_491),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_909),
.A2(n_924),
.B(n_916),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_907),
.B(n_920),
.Y(n_1048)
);

OR2x2_ASAP7_75t_L g1049 ( 
.A(n_907),
.B(n_502),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_922),
.B(n_502),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_915),
.B(n_714),
.Y(n_1051)
);

OA22x2_ASAP7_75t_L g1052 ( 
.A1(n_870),
.A2(n_881),
.B1(n_921),
.B2(n_502),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_907),
.B(n_502),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_SL g1054 ( 
.A1(n_921),
.A2(n_831),
.B(n_902),
.Y(n_1054)
);

INVx1_ASAP7_75t_SL g1055 ( 
.A(n_940),
.Y(n_1055)
);

O2A1O1Ixp5_ASAP7_75t_L g1056 ( 
.A1(n_909),
.A2(n_924),
.B(n_879),
.C(n_931),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_SL g1057 ( 
.A1(n_921),
.A2(n_831),
.B(n_902),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_915),
.B(n_714),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_915),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_916),
.B(n_927),
.Y(n_1060)
);

INVx2_ASAP7_75t_SL g1061 ( 
.A(n_940),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_921),
.A2(n_870),
.B1(n_881),
.B2(n_909),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_824),
.B(n_908),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_824),
.B(n_908),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_SL g1065 ( 
.A1(n_933),
.A2(n_921),
.B1(n_873),
.B2(n_881),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_824),
.B(n_908),
.Y(n_1066)
);

OAI22x1_ASAP7_75t_L g1067 ( 
.A1(n_780),
.A2(n_785),
.B1(n_873),
.B2(n_922),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_822),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_822),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_824),
.B(n_908),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_822),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_865),
.B(n_502),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_957),
.Y(n_1073)
);

OAI21xp33_ASAP7_75t_L g1074 ( 
.A1(n_1032),
.A2(n_1050),
.B(n_958),
.Y(n_1074)
);

INVx2_ASAP7_75t_SL g1075 ( 
.A(n_998),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_1030),
.B(n_1049),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_964),
.Y(n_1077)
);

INVx3_ASAP7_75t_SL g1078 ( 
.A(n_1024),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_1055),
.Y(n_1079)
);

AOI221x1_ASAP7_75t_L g1080 ( 
.A1(n_1062),
.A2(n_1067),
.B1(n_951),
.B2(n_945),
.C(n_988),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_958),
.A2(n_945),
.B(n_1065),
.C(n_951),
.Y(n_1081)
);

A2O1A1Ixp33_ASAP7_75t_SL g1082 ( 
.A1(n_952),
.A2(n_1039),
.B(n_1047),
.C(n_1029),
.Y(n_1082)
);

OAI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_1062),
.A2(n_1056),
.B(n_1028),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_1037),
.B(n_1048),
.Y(n_1084)
);

INVx5_ASAP7_75t_SL g1085 ( 
.A(n_956),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_1051),
.B(n_1058),
.Y(n_1086)
);

OR2x6_ASAP7_75t_L g1087 ( 
.A(n_990),
.B(n_947),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_1027),
.A2(n_1064),
.B1(n_1063),
.B2(n_1070),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_1066),
.A2(n_1052),
.B1(n_1035),
.B2(n_1036),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_979),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_960),
.A2(n_987),
.B(n_967),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_973),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_959),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1036),
.B(n_1060),
.Y(n_1094)
);

AND2x6_ASAP7_75t_L g1095 ( 
.A(n_1038),
.B(n_1051),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_1061),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_956),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_1055),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1060),
.B(n_974),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_974),
.B(n_1012),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_SL g1101 ( 
.A1(n_1054),
.A2(n_1057),
.B(n_984),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_1058),
.B(n_944),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_944),
.B(n_992),
.Y(n_1103)
);

CKINVDCx6p67_ASAP7_75t_R g1104 ( 
.A(n_981),
.Y(n_1104)
);

O2A1O1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_961),
.A2(n_952),
.B(n_1029),
.C(n_1039),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_968),
.B(n_963),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_1043),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1068),
.Y(n_1108)
);

BUFx12f_ASAP7_75t_L g1109 ( 
.A(n_978),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_SL g1110 ( 
.A(n_969),
.Y(n_1110)
);

AOI222xp33_ASAP7_75t_L g1111 ( 
.A1(n_1026),
.A2(n_1005),
.B1(n_1047),
.B2(n_986),
.C1(n_1071),
.C2(n_1069),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_990),
.Y(n_1112)
);

CKINVDCx11_ASAP7_75t_R g1113 ( 
.A(n_981),
.Y(n_1113)
);

OR2x6_ASAP7_75t_L g1114 ( 
.A(n_962),
.B(n_1043),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_976),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_991),
.A2(n_1053),
.B1(n_970),
.B2(n_1072),
.Y(n_1116)
);

OR2x6_ASAP7_75t_L g1117 ( 
.A(n_1043),
.B(n_1059),
.Y(n_1117)
);

OAI21xp33_ASAP7_75t_L g1118 ( 
.A1(n_971),
.A2(n_996),
.B(n_1020),
.Y(n_1118)
);

AOI222xp33_ASAP7_75t_L g1119 ( 
.A1(n_971),
.A2(n_992),
.B1(n_1011),
.B2(n_1017),
.C1(n_1025),
.C2(n_1006),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_948),
.B(n_955),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_L g1121 ( 
.A1(n_989),
.A2(n_1019),
.B1(n_1018),
.B2(n_1016),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_994),
.A2(n_1002),
.B(n_1010),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1009),
.B(n_1017),
.Y(n_1123)
);

HB1xp67_ASAP7_75t_L g1124 ( 
.A(n_1059),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_1059),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_1042),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1009),
.Y(n_1127)
);

AOI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_1016),
.A2(n_1022),
.B1(n_982),
.B2(n_997),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1007),
.B(n_1014),
.Y(n_1129)
);

INVxp67_ASAP7_75t_SL g1130 ( 
.A(n_1038),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_1022),
.B(n_1000),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_1021),
.A2(n_994),
.B(n_1013),
.C(n_997),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1014),
.B(n_1023),
.Y(n_1133)
);

NAND2x1p5_ASAP7_75t_L g1134 ( 
.A(n_1031),
.B(n_999),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_1000),
.B(n_999),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1015),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1014),
.Y(n_1137)
);

INVx6_ASAP7_75t_SL g1138 ( 
.A(n_1031),
.Y(n_1138)
);

OA21x2_ASAP7_75t_L g1139 ( 
.A1(n_983),
.A2(n_995),
.B(n_980),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1042),
.Y(n_1140)
);

INVx6_ASAP7_75t_SL g1141 ( 
.A(n_972),
.Y(n_1141)
);

INVx5_ASAP7_75t_L g1142 ( 
.A(n_1042),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1040),
.A2(n_1044),
.B1(n_1046),
.B2(n_1045),
.Y(n_1143)
);

INVx4_ASAP7_75t_L g1144 ( 
.A(n_954),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_953),
.A2(n_966),
.B(n_975),
.Y(n_1145)
);

NAND2x1p5_ASAP7_75t_L g1146 ( 
.A(n_977),
.B(n_985),
.Y(n_1146)
);

INVx2_ASAP7_75t_SL g1147 ( 
.A(n_1008),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1008),
.B(n_953),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1008),
.B(n_965),
.Y(n_1149)
);

BUFx2_ASAP7_75t_L g1150 ( 
.A(n_1034),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1034),
.B(n_950),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_993),
.Y(n_1152)
);

INVx5_ASAP7_75t_L g1153 ( 
.A(n_1001),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_946),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1041),
.A2(n_1004),
.B(n_924),
.C(n_909),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_1051),
.B(n_1058),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_958),
.A2(n_909),
.B(n_924),
.C(n_868),
.Y(n_1157)
);

AOI221xp5_ASAP7_75t_L g1158 ( 
.A1(n_951),
.A2(n_1062),
.B1(n_870),
.B2(n_881),
.C(n_945),
.Y(n_1158)
);

A2O1A1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_958),
.A2(n_909),
.B(n_924),
.C(n_868),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_949),
.B(n_1033),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1037),
.B(n_1048),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1037),
.B(n_1048),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_960),
.A2(n_987),
.B(n_967),
.Y(n_1163)
);

INVx2_ASAP7_75t_SL g1164 ( 
.A(n_998),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1065),
.A2(n_921),
.B1(n_870),
.B2(n_881),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_1055),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1065),
.A2(n_870),
.B1(n_881),
.B2(n_873),
.Y(n_1167)
);

INVx2_ASAP7_75t_SL g1168 ( 
.A(n_998),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1037),
.B(n_1048),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_957),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_957),
.Y(n_1171)
);

HB1xp67_ASAP7_75t_L g1172 ( 
.A(n_1055),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1032),
.B(n_1050),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_964),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_957),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1037),
.B(n_1048),
.Y(n_1176)
);

CKINVDCx20_ASAP7_75t_R g1177 ( 
.A(n_964),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_956),
.Y(n_1178)
);

O2A1O1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1062),
.A2(n_924),
.B(n_909),
.C(n_879),
.Y(n_1179)
);

INVx1_ASAP7_75t_SL g1180 ( 
.A(n_1055),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_998),
.Y(n_1181)
);

OAI21xp33_ASAP7_75t_L g1182 ( 
.A1(n_1032),
.A2(n_922),
.B(n_639),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_949),
.B(n_1033),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_1003),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_957),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_957),
.Y(n_1186)
);

BUFx12f_ASAP7_75t_L g1187 ( 
.A(n_964),
.Y(n_1187)
);

BUFx3_ASAP7_75t_L g1188 ( 
.A(n_998),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_1051),
.B(n_1058),
.Y(n_1189)
);

INVx4_ASAP7_75t_SL g1190 ( 
.A(n_1042),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_957),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_960),
.A2(n_987),
.B(n_967),
.Y(n_1192)
);

OR2x2_ASAP7_75t_L g1193 ( 
.A(n_963),
.B(n_1030),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_956),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_998),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_957),
.Y(n_1196)
);

HB1xp67_ASAP7_75t_L g1197 ( 
.A(n_1055),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_949),
.B(n_1033),
.Y(n_1198)
);

NAND2xp33_ASAP7_75t_SL g1199 ( 
.A(n_1067),
.B(n_921),
.Y(n_1199)
);

BUFx12f_ASAP7_75t_L g1200 ( 
.A(n_964),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_1098),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_SL g1202 ( 
.A1(n_1165),
.A2(n_1088),
.B1(n_1089),
.B2(n_1083),
.Y(n_1202)
);

BUFx2_ASAP7_75t_R g1203 ( 
.A(n_1077),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1079),
.Y(n_1204)
);

BUFx2_ASAP7_75t_L g1205 ( 
.A(n_1181),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1182),
.A2(n_1159),
.B(n_1157),
.Y(n_1206)
);

AO21x1_ASAP7_75t_SL g1207 ( 
.A1(n_1167),
.A2(n_1083),
.B(n_1123),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_1177),
.Y(n_1208)
);

INVx6_ASAP7_75t_L g1209 ( 
.A(n_1142),
.Y(n_1209)
);

OA21x2_ASAP7_75t_L g1210 ( 
.A1(n_1145),
.A2(n_1122),
.B(n_1091),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1188),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1175),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1099),
.B(n_1094),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1099),
.B(n_1094),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1165),
.A2(n_1199),
.B1(n_1158),
.B2(n_1111),
.Y(n_1215)
);

CKINVDCx14_ASAP7_75t_R g1216 ( 
.A(n_1113),
.Y(n_1216)
);

AO22x1_ASAP7_75t_L g1217 ( 
.A1(n_1092),
.A2(n_1160),
.B1(n_1198),
.B2(n_1183),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1195),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1183),
.B(n_1084),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1103),
.B(n_1102),
.Y(n_1220)
);

INVx1_ASAP7_75t_SL g1221 ( 
.A(n_1180),
.Y(n_1221)
);

HB1xp67_ASAP7_75t_L g1222 ( 
.A(n_1166),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_1142),
.Y(n_1223)
);

BUFx2_ASAP7_75t_SL g1224 ( 
.A(n_1075),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1095),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1100),
.B(n_1081),
.Y(n_1226)
);

OAI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1116),
.A2(n_1173),
.B1(n_1080),
.B2(n_1193),
.Y(n_1227)
);

INVxp67_ASAP7_75t_L g1228 ( 
.A(n_1172),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1108),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1158),
.A2(n_1111),
.B1(n_1074),
.B2(n_1088),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1170),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1171),
.Y(n_1232)
);

OR2x2_ASAP7_75t_L g1233 ( 
.A(n_1089),
.B(n_1082),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1185),
.Y(n_1234)
);

INVx2_ASAP7_75t_SL g1235 ( 
.A(n_1090),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1161),
.A2(n_1162),
.B1(n_1169),
.B2(n_1176),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1100),
.B(n_1128),
.Y(n_1237)
);

OR2x6_ASAP7_75t_L g1238 ( 
.A(n_1105),
.B(n_1179),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1186),
.Y(n_1239)
);

INVx5_ASAP7_75t_L g1240 ( 
.A(n_1095),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1118),
.A2(n_1106),
.B1(n_1076),
.B2(n_1121),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1197),
.Y(n_1242)
);

OAI22x1_ASAP7_75t_L g1243 ( 
.A1(n_1150),
.A2(n_1147),
.B1(n_1144),
.B2(n_1127),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1101),
.A2(n_1103),
.B1(n_1119),
.B2(n_1156),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1180),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1148),
.B(n_1119),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1191),
.B(n_1196),
.Y(n_1247)
);

CKINVDCx20_ASAP7_75t_R g1248 ( 
.A(n_1174),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1086),
.A2(n_1189),
.B1(n_1168),
.B2(n_1164),
.Y(n_1249)
);

INVx6_ASAP7_75t_L g1250 ( 
.A(n_1190),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1093),
.Y(n_1251)
);

OA21x2_ASAP7_75t_L g1252 ( 
.A1(n_1120),
.A2(n_1132),
.B(n_1129),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1130),
.Y(n_1253)
);

OR2x2_ASAP7_75t_L g1254 ( 
.A(n_1123),
.B(n_1133),
.Y(n_1254)
);

OA21x2_ASAP7_75t_L g1255 ( 
.A1(n_1120),
.A2(n_1129),
.B(n_1133),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1096),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1124),
.Y(n_1257)
);

AO21x2_ASAP7_75t_L g1258 ( 
.A1(n_1143),
.A2(n_1155),
.B(n_1136),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1130),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1179),
.B(n_1149),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1131),
.Y(n_1261)
);

CKINVDCx6p67_ASAP7_75t_R g1262 ( 
.A(n_1078),
.Y(n_1262)
);

INVx3_ASAP7_75t_L g1263 ( 
.A(n_1095),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1137),
.B(n_1105),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1144),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1151),
.B(n_1135),
.Y(n_1266)
);

BUFx12f_ASAP7_75t_L g1267 ( 
.A(n_1115),
.Y(n_1267)
);

CKINVDCx11_ASAP7_75t_R g1268 ( 
.A(n_1109),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1112),
.Y(n_1269)
);

AOI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1104),
.A2(n_1110),
.B1(n_1087),
.B2(n_1187),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1140),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1152),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1117),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1087),
.B(n_1114),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1114),
.B(n_1184),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1117),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1117),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1154),
.A2(n_1139),
.B(n_1146),
.Y(n_1278)
);

CKINVDCx16_ASAP7_75t_R g1279 ( 
.A(n_1200),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1139),
.A2(n_1146),
.B(n_1184),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1141),
.A2(n_1110),
.B1(n_1114),
.B2(n_1125),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1153),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1190),
.B(n_1194),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_SL g1284 ( 
.A1(n_1126),
.A2(n_1085),
.B1(n_1153),
.B2(n_1134),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1097),
.B(n_1194),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_1141),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1138),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1097),
.B(n_1107),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_SL g1289 ( 
.A1(n_1085),
.A2(n_1153),
.B1(n_1134),
.B2(n_1107),
.Y(n_1289)
);

CKINVDCx11_ASAP7_75t_R g1290 ( 
.A(n_1178),
.Y(n_1290)
);

OAI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1194),
.A2(n_1067),
.B1(n_921),
.B2(n_881),
.Y(n_1291)
);

BUFx8_ASAP7_75t_L g1292 ( 
.A(n_1110),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1120),
.A2(n_1192),
.B(n_1163),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1167),
.B(n_1065),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1098),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1098),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1182),
.A2(n_924),
.B(n_909),
.Y(n_1297)
);

CKINVDCx11_ASAP7_75t_R g1298 ( 
.A(n_1109),
.Y(n_1298)
);

OA21x2_ASAP7_75t_L g1299 ( 
.A1(n_1145),
.A2(n_1122),
.B(n_1091),
.Y(n_1299)
);

INVx1_ASAP7_75t_SL g1300 ( 
.A(n_1113),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1073),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1073),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1079),
.Y(n_1303)
);

AND2x4_ASAP7_75t_L g1304 ( 
.A(n_1103),
.B(n_1102),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1265),
.B(n_1282),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1245),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1213),
.B(n_1214),
.Y(n_1307)
);

INVxp67_ASAP7_75t_L g1308 ( 
.A(n_1204),
.Y(n_1308)
);

OR2x6_ASAP7_75t_L g1309 ( 
.A(n_1293),
.B(n_1238),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1260),
.B(n_1246),
.Y(n_1310)
);

INVx3_ASAP7_75t_L g1311 ( 
.A(n_1280),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1255),
.B(n_1238),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1255),
.B(n_1238),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1272),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1252),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1213),
.B(n_1214),
.Y(n_1316)
);

INVx2_ASAP7_75t_SL g1317 ( 
.A(n_1247),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1260),
.B(n_1246),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1266),
.B(n_1264),
.Y(n_1319)
);

BUFx2_ASAP7_75t_L g1320 ( 
.A(n_1272),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1264),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1266),
.B(n_1238),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1243),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1226),
.B(n_1202),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1226),
.B(n_1254),
.Y(n_1325)
);

INVxp67_ASAP7_75t_L g1326 ( 
.A(n_1222),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1243),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1208),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1219),
.B(n_1205),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_1242),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1253),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1254),
.B(n_1207),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1297),
.A2(n_1206),
.B(n_1230),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1233),
.B(n_1258),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_1303),
.Y(n_1335)
);

OA21x2_ASAP7_75t_L g1336 ( 
.A1(n_1233),
.A2(n_1278),
.B(n_1215),
.Y(n_1336)
);

INVx2_ASAP7_75t_SL g1337 ( 
.A(n_1247),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1210),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1299),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1237),
.B(n_1294),
.Y(n_1340)
);

CKINVDCx6p67_ASAP7_75t_R g1341 ( 
.A(n_1248),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1237),
.B(n_1294),
.Y(n_1342)
);

BUFx12f_ASAP7_75t_L g1343 ( 
.A(n_1268),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_1221),
.Y(n_1344)
);

INVx4_ASAP7_75t_L g1345 ( 
.A(n_1240),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1229),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1227),
.B(n_1241),
.Y(n_1347)
);

AO21x2_ASAP7_75t_L g1348 ( 
.A1(n_1291),
.A2(n_1259),
.B(n_1271),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_1201),
.Y(n_1349)
);

INVx3_ASAP7_75t_L g1350 ( 
.A(n_1240),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1231),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1261),
.Y(n_1352)
);

AOI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1217),
.A2(n_1253),
.B(n_1277),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1240),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1232),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1234),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1239),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1228),
.B(n_1236),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1212),
.Y(n_1359)
);

AND2x4_ASAP7_75t_L g1360 ( 
.A(n_1225),
.B(n_1263),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1208),
.Y(n_1361)
);

AO21x2_ASAP7_75t_L g1362 ( 
.A1(n_1273),
.A2(n_1276),
.B(n_1301),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1302),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1244),
.A2(n_1304),
.B1(n_1220),
.B2(n_1249),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1257),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1274),
.B(n_1275),
.Y(n_1366)
);

INVx2_ASAP7_75t_SL g1367 ( 
.A(n_1274),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1312),
.B(n_1288),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1312),
.B(n_1288),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1331),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1310),
.B(n_1296),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1311),
.B(n_1263),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1313),
.B(n_1285),
.Y(n_1373)
);

INVxp67_ASAP7_75t_L g1374 ( 
.A(n_1362),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1313),
.B(n_1285),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1315),
.B(n_1275),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1310),
.B(n_1289),
.Y(n_1377)
);

NOR2x1p5_ASAP7_75t_L g1378 ( 
.A(n_1347),
.B(n_1225),
.Y(n_1378)
);

NAND3xp33_ASAP7_75t_SL g1379 ( 
.A(n_1333),
.B(n_1281),
.C(n_1270),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1362),
.Y(n_1380)
);

OR2x2_ASAP7_75t_L g1381 ( 
.A(n_1334),
.B(n_1201),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1362),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1328),
.Y(n_1383)
);

NAND3xp33_ASAP7_75t_L g1384 ( 
.A(n_1324),
.B(n_1292),
.C(n_1218),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1318),
.B(n_1284),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1314),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1321),
.B(n_1295),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1325),
.B(n_1321),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1325),
.B(n_1295),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1323),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1309),
.B(n_1304),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_SL g1392 ( 
.A1(n_1324),
.A2(n_1216),
.B1(n_1292),
.B2(n_1209),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1309),
.B(n_1304),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1309),
.B(n_1319),
.Y(n_1394)
);

BUFx2_ASAP7_75t_L g1395 ( 
.A(n_1323),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1309),
.B(n_1220),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1327),
.B(n_1235),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1309),
.B(n_1305),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1319),
.B(n_1336),
.Y(n_1399)
);

OA21x2_ASAP7_75t_L g1400 ( 
.A1(n_1374),
.A2(n_1339),
.B(n_1338),
.Y(n_1400)
);

INVxp67_ASAP7_75t_SL g1401 ( 
.A(n_1386),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1379),
.A2(n_1345),
.B(n_1348),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_SL g1403 ( 
.A(n_1392),
.B(n_1329),
.Y(n_1403)
);

NAND3xp33_ASAP7_75t_L g1404 ( 
.A(n_1384),
.B(n_1358),
.C(n_1352),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1371),
.B(n_1330),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_SL g1406 ( 
.A(n_1392),
.B(n_1349),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_SL g1407 ( 
.A(n_1384),
.B(n_1360),
.Y(n_1407)
);

AOI221xp5_ASAP7_75t_L g1408 ( 
.A1(n_1379),
.A2(n_1308),
.B1(n_1326),
.B2(n_1365),
.C(n_1335),
.Y(n_1408)
);

NAND4xp25_ASAP7_75t_L g1409 ( 
.A(n_1397),
.B(n_1340),
.C(n_1342),
.D(n_1365),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1388),
.B(n_1306),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1385),
.A2(n_1342),
.B1(n_1340),
.B2(n_1364),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1368),
.B(n_1322),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1388),
.B(n_1307),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1368),
.B(n_1322),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1385),
.A2(n_1344),
.B1(n_1316),
.B2(n_1216),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1387),
.B(n_1332),
.Y(n_1416)
);

OAI221xp5_ASAP7_75t_SL g1417 ( 
.A1(n_1377),
.A2(n_1332),
.B1(n_1327),
.B2(n_1300),
.C(n_1341),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1368),
.B(n_1366),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1369),
.B(n_1366),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1369),
.B(n_1314),
.Y(n_1420)
);

AOI221x1_ASAP7_75t_SL g1421 ( 
.A1(n_1377),
.A2(n_1357),
.B1(n_1356),
.B2(n_1346),
.C(n_1351),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1378),
.A2(n_1317),
.B1(n_1337),
.B2(n_1341),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1373),
.B(n_1320),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1373),
.B(n_1375),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1375),
.B(n_1320),
.Y(n_1425)
);

AOI211xp5_ASAP7_75t_SL g1426 ( 
.A1(n_1381),
.A2(n_1350),
.B(n_1354),
.C(n_1360),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1375),
.B(n_1367),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1389),
.B(n_1346),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1381),
.B(n_1351),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1386),
.B(n_1355),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_SL g1431 ( 
.A(n_1391),
.B(n_1360),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1397),
.B(n_1376),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1397),
.B(n_1355),
.Y(n_1433)
);

NAND3xp33_ASAP7_75t_L g1434 ( 
.A(n_1374),
.B(n_1363),
.C(n_1359),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1399),
.B(n_1336),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1399),
.B(n_1317),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1378),
.A2(n_1337),
.B1(n_1250),
.B2(n_1353),
.Y(n_1437)
);

OAI211xp5_ASAP7_75t_L g1438 ( 
.A1(n_1390),
.A2(n_1353),
.B(n_1357),
.C(n_1286),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1424),
.B(n_1394),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1432),
.B(n_1390),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1424),
.B(n_1394),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1401),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1433),
.Y(n_1443)
);

NAND3xp33_ASAP7_75t_L g1444 ( 
.A(n_1408),
.B(n_1382),
.C(n_1380),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1430),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1436),
.B(n_1398),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1434),
.Y(n_1447)
);

INVx4_ASAP7_75t_L g1448 ( 
.A(n_1400),
.Y(n_1448)
);

INVx2_ASAP7_75t_SL g1449 ( 
.A(n_1412),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1434),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1420),
.B(n_1395),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1412),
.B(n_1398),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1429),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1414),
.B(n_1398),
.Y(n_1454)
);

INVx2_ASAP7_75t_SL g1455 ( 
.A(n_1414),
.Y(n_1455)
);

NOR2xp33_ASAP7_75t_L g1456 ( 
.A(n_1405),
.B(n_1361),
.Y(n_1456)
);

AOI21xp33_ASAP7_75t_SL g1457 ( 
.A1(n_1415),
.A2(n_1279),
.B(n_1383),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1428),
.Y(n_1458)
);

INVxp67_ASAP7_75t_SL g1459 ( 
.A(n_1416),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1423),
.B(n_1395),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1400),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1431),
.B(n_1398),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1400),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1425),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1406),
.A2(n_1396),
.B1(n_1391),
.B2(n_1393),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1418),
.B(n_1419),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1435),
.B(n_1370),
.Y(n_1467)
);

AND2x4_ASAP7_75t_L g1468 ( 
.A(n_1418),
.B(n_1398),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1421),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1421),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1419),
.B(n_1435),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1426),
.B(n_1391),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1447),
.B(n_1450),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1472),
.B(n_1426),
.Y(n_1474)
);

INVx3_ASAP7_75t_L g1475 ( 
.A(n_1448),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1442),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1472),
.B(n_1413),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1442),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1447),
.B(n_1402),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1450),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1467),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1462),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1462),
.B(n_1372),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1468),
.B(n_1407),
.Y(n_1484)
);

INVxp33_ASAP7_75t_L g1485 ( 
.A(n_1456),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1461),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1467),
.Y(n_1487)
);

NAND4xp25_ASAP7_75t_L g1488 ( 
.A(n_1444),
.B(n_1404),
.C(n_1417),
.D(n_1415),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1462),
.B(n_1468),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1448),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1468),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1448),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1469),
.B(n_1410),
.Y(n_1493)
);

AOI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1469),
.A2(n_1404),
.B1(n_1403),
.B2(n_1411),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1443),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1471),
.B(n_1452),
.Y(n_1496)
);

INVxp67_ASAP7_75t_L g1497 ( 
.A(n_1470),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1443),
.Y(n_1498)
);

INVxp67_ASAP7_75t_SL g1499 ( 
.A(n_1463),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1471),
.B(n_1427),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1445),
.Y(n_1501)
);

INVxp67_ASAP7_75t_L g1502 ( 
.A(n_1470),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1445),
.Y(n_1503)
);

INVxp67_ASAP7_75t_L g1504 ( 
.A(n_1453),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1440),
.Y(n_1505)
);

INVx1_ASAP7_75t_SL g1506 ( 
.A(n_1493),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1476),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1489),
.B(n_1452),
.Y(n_1508)
);

INVx2_ASAP7_75t_SL g1509 ( 
.A(n_1482),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1494),
.B(n_1459),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1504),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1474),
.B(n_1454),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1473),
.B(n_1451),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1476),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1486),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1474),
.B(n_1454),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1489),
.B(n_1439),
.Y(n_1517)
);

NOR2x1p5_ASAP7_75t_SL g1518 ( 
.A(n_1490),
.B(n_1463),
.Y(n_1518)
);

XOR2x2_ASAP7_75t_L g1519 ( 
.A(n_1494),
.B(n_1411),
.Y(n_1519)
);

INVxp67_ASAP7_75t_L g1520 ( 
.A(n_1493),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1473),
.B(n_1451),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1477),
.B(n_1453),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1478),
.Y(n_1523)
);

NOR2xp67_ASAP7_75t_L g1524 ( 
.A(n_1489),
.B(n_1343),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1477),
.B(n_1458),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1504),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1489),
.B(n_1439),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1479),
.B(n_1497),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_SL g1529 ( 
.A(n_1479),
.B(n_1457),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1505),
.B(n_1460),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1491),
.B(n_1441),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1491),
.B(n_1441),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1482),
.B(n_1446),
.Y(n_1533)
);

AOI32xp33_ASAP7_75t_L g1534 ( 
.A1(n_1484),
.A2(n_1465),
.A3(n_1422),
.B1(n_1437),
.B2(n_1455),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1478),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1501),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1484),
.B(n_1446),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1501),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1496),
.B(n_1449),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1503),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1503),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_1483),
.B(n_1455),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1495),
.Y(n_1543)
);

NAND2x1_ASAP7_75t_L g1544 ( 
.A(n_1483),
.B(n_1475),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1497),
.B(n_1458),
.Y(n_1545)
);

INVxp67_ASAP7_75t_L g1546 ( 
.A(n_1480),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1485),
.B(n_1343),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1536),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1538),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1519),
.A2(n_1488),
.B1(n_1480),
.B2(n_1505),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1512),
.B(n_1502),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1519),
.A2(n_1488),
.B1(n_1409),
.B2(n_1393),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1512),
.B(n_1502),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1516),
.B(n_1483),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1506),
.B(n_1481),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_1547),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1511),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1540),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1529),
.B(n_1268),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1541),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1516),
.B(n_1483),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1528),
.B(n_1481),
.Y(n_1562)
);

AOI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1529),
.A2(n_1498),
.B(n_1495),
.Y(n_1563)
);

AOI222xp33_ASAP7_75t_L g1564 ( 
.A1(n_1510),
.A2(n_1487),
.B1(n_1499),
.B2(n_1498),
.C1(n_1438),
.C2(n_1437),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1509),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_1520),
.B(n_1298),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1524),
.B(n_1298),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1513),
.Y(n_1568)
);

NAND3xp33_ASAP7_75t_L g1569 ( 
.A(n_1526),
.B(n_1492),
.C(n_1490),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1513),
.B(n_1487),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1537),
.B(n_1500),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1543),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1537),
.B(n_1500),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1521),
.B(n_1466),
.Y(n_1574)
);

INVx1_ASAP7_75t_SL g1575 ( 
.A(n_1521),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_L g1576 ( 
.A1(n_1527),
.A2(n_1409),
.B1(n_1396),
.B2(n_1393),
.Y(n_1576)
);

AO21x2_ASAP7_75t_L g1577 ( 
.A1(n_1515),
.A2(n_1499),
.B(n_1492),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1507),
.Y(n_1578)
);

CKINVDCx16_ASAP7_75t_R g1579 ( 
.A(n_1509),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1545),
.B(n_1464),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1514),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_1530),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1515),
.Y(n_1583)
);

AOI322xp5_ASAP7_75t_L g1584 ( 
.A1(n_1550),
.A2(n_1552),
.A3(n_1559),
.B1(n_1557),
.B2(n_1553),
.C1(n_1551),
.C2(n_1582),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_1556),
.B(n_1267),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1551),
.B(n_1517),
.Y(n_1586)
);

AOI21xp33_ASAP7_75t_SL g1587 ( 
.A1(n_1564),
.A2(n_1534),
.B(n_1546),
.Y(n_1587)
);

AOI22xp5_ASAP7_75t_SL g1588 ( 
.A1(n_1567),
.A2(n_1248),
.B1(n_1527),
.B2(n_1508),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1548),
.Y(n_1589)
);

INVxp67_ASAP7_75t_SL g1590 ( 
.A(n_1553),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1568),
.B(n_1531),
.Y(n_1591)
);

AOI22xp33_ASAP7_75t_SL g1592 ( 
.A1(n_1579),
.A2(n_1527),
.B1(n_1531),
.B2(n_1532),
.Y(n_1592)
);

INVxp67_ASAP7_75t_L g1593 ( 
.A(n_1566),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1575),
.B(n_1565),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1548),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1565),
.B(n_1532),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1549),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1549),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1554),
.B(n_1517),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1555),
.Y(n_1600)
);

AOI21xp33_ASAP7_75t_L g1601 ( 
.A1(n_1569),
.A2(n_1544),
.B(n_1535),
.Y(n_1601)
);

INVxp67_ASAP7_75t_L g1602 ( 
.A(n_1555),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1563),
.B(n_1533),
.Y(n_1603)
);

INVxp33_ASAP7_75t_L g1604 ( 
.A(n_1562),
.Y(n_1604)
);

OAI321xp33_ASAP7_75t_L g1605 ( 
.A1(n_1562),
.A2(n_1530),
.A3(n_1522),
.B1(n_1523),
.B2(n_1525),
.C(n_1422),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1580),
.B(n_1267),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1571),
.B(n_1573),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1571),
.B(n_1533),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_R g1609 ( 
.A(n_1578),
.B(n_1292),
.Y(n_1609)
);

OAI221xp5_ASAP7_75t_L g1610 ( 
.A1(n_1576),
.A2(n_1492),
.B1(n_1490),
.B2(n_1475),
.C(n_1539),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1600),
.B(n_1570),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1599),
.B(n_1586),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1590),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1589),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1595),
.Y(n_1615)
);

INVx1_ASAP7_75t_SL g1616 ( 
.A(n_1609),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1608),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1593),
.B(n_1574),
.Y(n_1618)
);

NAND2x1p5_ASAP7_75t_L g1619 ( 
.A(n_1585),
.B(n_1211),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1592),
.B(n_1554),
.Y(n_1620)
);

INVx3_ASAP7_75t_L g1621 ( 
.A(n_1597),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1584),
.B(n_1573),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1607),
.Y(n_1623)
);

NAND2xp33_ASAP7_75t_L g1624 ( 
.A(n_1609),
.B(n_1583),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1587),
.A2(n_1574),
.B1(n_1508),
.B2(n_1561),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1591),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1598),
.Y(n_1627)
);

INVx2_ASAP7_75t_SL g1628 ( 
.A(n_1596),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1594),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_SL g1630 ( 
.A(n_1585),
.B(n_1203),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1612),
.Y(n_1631)
);

INVxp33_ASAP7_75t_L g1632 ( 
.A(n_1618),
.Y(n_1632)
);

OAI221xp5_ASAP7_75t_L g1633 ( 
.A1(n_1622),
.A2(n_1588),
.B1(n_1603),
.B2(n_1601),
.C(n_1602),
.Y(n_1633)
);

AOI211x1_ASAP7_75t_L g1634 ( 
.A1(n_1620),
.A2(n_1610),
.B(n_1581),
.C(n_1560),
.Y(n_1634)
);

NOR3xp33_ASAP7_75t_L g1635 ( 
.A(n_1616),
.B(n_1605),
.C(n_1606),
.Y(n_1635)
);

OAI211xp5_ASAP7_75t_SL g1636 ( 
.A1(n_1624),
.A2(n_1606),
.B(n_1558),
.C(n_1560),
.Y(n_1636)
);

NOR3xp33_ASAP7_75t_SL g1637 ( 
.A(n_1613),
.B(n_1572),
.C(n_1558),
.Y(n_1637)
);

AOI222xp33_ASAP7_75t_L g1638 ( 
.A1(n_1629),
.A2(n_1604),
.B1(n_1518),
.B2(n_1572),
.C1(n_1583),
.C2(n_1561),
.Y(n_1638)
);

OAI21xp33_ASAP7_75t_L g1639 ( 
.A1(n_1620),
.A2(n_1612),
.B(n_1625),
.Y(n_1639)
);

AOI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1624),
.A2(n_1604),
.B(n_1577),
.Y(n_1640)
);

AOI221xp5_ASAP7_75t_L g1641 ( 
.A1(n_1628),
.A2(n_1577),
.B1(n_1570),
.B2(n_1475),
.C(n_1486),
.Y(n_1641)
);

NOR3xp33_ASAP7_75t_L g1642 ( 
.A(n_1633),
.B(n_1639),
.C(n_1636),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1631),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1632),
.B(n_1623),
.Y(n_1644)
);

NOR3xp33_ASAP7_75t_L g1645 ( 
.A(n_1635),
.B(n_1626),
.C(n_1623),
.Y(n_1645)
);

NOR3xp33_ASAP7_75t_L g1646 ( 
.A(n_1640),
.B(n_1626),
.C(n_1617),
.Y(n_1646)
);

NOR2x1_ASAP7_75t_SL g1647 ( 
.A(n_1637),
.B(n_1611),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1634),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1638),
.Y(n_1649)
);

OAI211xp5_ASAP7_75t_SL g1650 ( 
.A1(n_1641),
.A2(n_1614),
.B(n_1627),
.C(n_1617),
.Y(n_1650)
);

OAI211xp5_ASAP7_75t_SL g1651 ( 
.A1(n_1642),
.A2(n_1649),
.B(n_1648),
.C(n_1645),
.Y(n_1651)
);

AOI211xp5_ASAP7_75t_L g1652 ( 
.A1(n_1650),
.A2(n_1611),
.B(n_1628),
.C(n_1615),
.Y(n_1652)
);

NOR3xp33_ASAP7_75t_L g1653 ( 
.A(n_1644),
.B(n_1621),
.C(n_1615),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1643),
.Y(n_1654)
);

NOR3x1_ASAP7_75t_L g1655 ( 
.A(n_1647),
.B(n_1619),
.C(n_1630),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1655),
.B(n_1621),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1653),
.Y(n_1657)
);

NOR2x1_ASAP7_75t_L g1658 ( 
.A(n_1651),
.B(n_1621),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1652),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1654),
.B(n_1646),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1652),
.A2(n_1619),
.B1(n_1508),
.B2(n_1542),
.Y(n_1661)
);

OAI211xp5_ASAP7_75t_L g1662 ( 
.A1(n_1659),
.A2(n_1650),
.B(n_1287),
.C(n_1256),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1656),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1658),
.B(n_1577),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1660),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1657),
.B(n_1619),
.Y(n_1666)
);

OAI21xp33_ASAP7_75t_L g1667 ( 
.A1(n_1663),
.A2(n_1661),
.B(n_1518),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1664),
.Y(n_1668)
);

NAND2xp33_ASAP7_75t_SL g1669 ( 
.A(n_1666),
.B(n_1287),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1668),
.Y(n_1670)
);

OAI221xp5_ASAP7_75t_L g1671 ( 
.A1(n_1670),
.A2(n_1667),
.B1(n_1662),
.B2(n_1669),
.C(n_1665),
.Y(n_1671)
);

NAND4xp75_ASAP7_75t_L g1672 ( 
.A(n_1671),
.B(n_1662),
.C(n_1664),
.D(n_1262),
.Y(n_1672)
);

OAI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1671),
.A2(n_1256),
.B(n_1251),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_SL g1674 ( 
.A(n_1673),
.B(n_1251),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1672),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1675),
.B(n_1211),
.Y(n_1676)
);

AOI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1674),
.A2(n_1235),
.B(n_1269),
.Y(n_1677)
);

NAND3xp33_ASAP7_75t_L g1678 ( 
.A(n_1676),
.B(n_1269),
.C(n_1290),
.Y(n_1678)
);

AOI22xp5_ASAP7_75t_SL g1679 ( 
.A1(n_1678),
.A2(n_1677),
.B1(n_1262),
.B2(n_1224),
.Y(n_1679)
);

OAI221xp5_ASAP7_75t_R g1680 ( 
.A1(n_1679),
.A2(n_1475),
.B1(n_1486),
.B2(n_1290),
.C(n_1542),
.Y(n_1680)
);

AOI211xp5_ASAP7_75t_L g1681 ( 
.A1(n_1680),
.A2(n_1286),
.B(n_1283),
.C(n_1223),
.Y(n_1681)
);


endmodule