module fake_jpeg_23085_n_191 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_191);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_191;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx2_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_9),
.B(n_7),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_33),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_36),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_38),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_26),
.B(n_1),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_20),
.Y(n_48)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_30),
.B1(n_21),
.B2(n_24),
.Y(n_54)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_42),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_45),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_1),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_21),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_25),
.B(n_1),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_49),
.Y(n_77)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_52),
.Y(n_82)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_30),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_67),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_54),
.A2(n_4),
.B(n_5),
.Y(n_89)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_58),
.Y(n_99)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_61),
.Y(n_80)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_25),
.Y(n_64)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_33),
.A2(n_23),
.B1(n_31),
.B2(n_30),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_69),
.B1(n_18),
.B2(n_22),
.Y(n_78)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

OR2x4_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_19),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_33),
.B(n_26),
.Y(n_68)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_40),
.A2(n_29),
.B1(n_22),
.B2(n_17),
.Y(n_69)
);

CKINVDCx12_ASAP7_75t_R g71 ( 
.A(n_36),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_2),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_74),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_29),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_73),
.B(n_51),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_28),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_28),
.C(n_20),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_85),
.C(n_86),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_78),
.A2(n_93),
.B1(n_69),
.B2(n_47),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_18),
.B1(n_27),
.B2(n_15),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_83),
.A2(n_89),
.B1(n_90),
.B2(n_98),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_27),
.C(n_19),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_19),
.C(n_5),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_19),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_95),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_4),
.C(n_6),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_95),
.C(n_85),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_65),
.A2(n_8),
.B1(n_14),
.B2(n_11),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_10),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_49),
.A2(n_13),
.B1(n_14),
.B2(n_50),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_100),
.B(n_56),
.Y(n_118)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_107),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_79),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_111),
.C(n_121),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_99),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_106),
.B(n_117),
.Y(n_133)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_87),
.A2(n_49),
.B(n_70),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_72),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_112),
.B(n_114),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_76),
.B1(n_77),
.B2(n_93),
.Y(n_123)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_59),
.Y(n_116)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_118),
.B(n_122),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_69),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_120),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_63),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_132),
.B1(n_134),
.B2(n_136),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_77),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_130),
.C(n_137),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_93),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_75),
.B(n_117),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_86),
.C(n_70),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_114),
.A2(n_89),
.B1(n_93),
.B2(n_96),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_81),
.B1(n_62),
.B2(n_52),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_110),
.A2(n_92),
.B1(n_91),
.B2(n_55),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_94),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_138),
.A2(n_102),
.B1(n_109),
.B2(n_121),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_139),
.B(n_141),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_123),
.B(n_111),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_147),
.Y(n_158)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_143),
.B(n_144),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_109),
.C(n_104),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_107),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_152),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

INVx3_ASAP7_75t_SL g159 ( 
.A(n_149),
.Y(n_159)
);

FAx1_ASAP7_75t_SL g161 ( 
.A(n_150),
.B(n_153),
.CI(n_154),
.CON(n_161),
.SN(n_161)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_134),
.A2(n_46),
.B1(n_63),
.B2(n_13),
.Y(n_151)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_151),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_46),
.C(n_108),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_46),
.C(n_130),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_140),
.C(n_126),
.Y(n_154)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_149),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_163),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_146),
.Y(n_163)
);

OAI31xp33_ASAP7_75t_SL g165 ( 
.A1(n_142),
.A2(n_127),
.A3(n_129),
.B(n_132),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_129),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_147),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_145),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_167),
.A2(n_173),
.B(n_174),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_135),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_169),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_145),
.C(n_153),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_139),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_170),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_171),
.A2(n_175),
.B1(n_165),
.B2(n_163),
.Y(n_176)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_128),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_176),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_172),
.A2(n_171),
.B(n_156),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_180),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_169),
.A2(n_156),
.B(n_161),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_161),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_184),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_162),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_178),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_183),
.Y(n_190)
);

AOI322xp5_ASAP7_75t_L g188 ( 
.A1(n_182),
.A2(n_181),
.A3(n_177),
.B1(n_180),
.B2(n_161),
.C1(n_158),
.C2(n_162),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_188),
.A2(n_183),
.B(n_187),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_189),
.B(n_190),
.Y(n_191)
);


endmodule