module fake_jpeg_16951_n_143 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_143);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx2_ASAP7_75t_SL g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_42),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_30),
.A2(n_22),
.B1(n_18),
.B2(n_19),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_13),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_14),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_24),
.B1(n_18),
.B2(n_19),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_22),
.B1(n_13),
.B2(n_23),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_27),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_53),
.B(n_59),
.Y(n_68)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NOR2x1_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_24),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_57),
.Y(n_69)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_46),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_58),
.Y(n_78)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_15),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_60),
.B(n_64),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_48),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_61),
.B(n_48),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_20),
.B1(n_26),
.B2(n_25),
.Y(n_77)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_48),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_51),
.B(n_15),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_75),
.B(n_10),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_32),
.B1(n_31),
.B2(n_29),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_40),
.B1(n_37),
.B2(n_52),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_81),
.B1(n_37),
.B2(n_25),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_SL g79 ( 
.A1(n_55),
.A2(n_25),
.B(n_16),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_79),
.A2(n_65),
.B1(n_20),
.B2(n_57),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_55),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_94),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_85),
.B(n_89),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_53),
.B(n_59),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_48),
.B(n_28),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_63),
.B(n_52),
.C(n_28),
.Y(n_88)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_73),
.B(n_78),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_66),
.B1(n_56),
.B2(n_40),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_90),
.B(n_91),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_95),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_82),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_0),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_96),
.B(n_86),
.Y(n_104)
);

OAI321xp33_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_80),
.A3(n_71),
.B1(n_81),
.B2(n_67),
.C(n_82),
.Y(n_100)
);

NAND3xp33_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_104),
.C(n_96),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_71),
.Y(n_103)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_104),
.C(n_83),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_116),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_107),
.A2(n_84),
.B1(n_90),
.B2(n_88),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_113),
.B1(n_97),
.B2(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_105),
.B(n_94),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_112),
.B(n_114),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_99),
.A2(n_96),
.B1(n_74),
.B2(n_67),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_99),
.B(n_9),
.Y(n_114)
);

A2O1A1O1Ixp25_ASAP7_75t_L g116 ( 
.A1(n_97),
.A2(n_14),
.B(n_16),
.C(n_4),
.D(n_5),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_106),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_124),
.C(n_118),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_121),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_101),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_120),
.A2(n_117),
.B(n_113),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_128),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_129),
.B(n_130),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_123),
.A2(n_116),
.B(n_11),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_14),
.Y(n_129)
);

INVxp33_ASAP7_75t_SL g131 ( 
.A(n_121),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_131),
.Y(n_134)
);

AOI31xp67_ASAP7_75t_L g135 ( 
.A1(n_131),
.A2(n_122),
.A3(n_125),
.B(n_3),
.Y(n_135)
);

OAI221xp5_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_7),
.B1(n_11),
.B2(n_12),
.C(n_4),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_133),
.A2(n_122),
.B(n_7),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_136),
.A2(n_132),
.B(n_14),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_138),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_134),
.A2(n_12),
.B(n_3),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_139),
.Y(n_143)
);


endmodule