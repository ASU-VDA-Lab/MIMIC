module fake_jpeg_3299_n_611 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_611);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_611;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_539;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_7),
.B(n_17),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_SL g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_8),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_14),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_L g60 ( 
.A1(n_31),
.A2(n_9),
.B(n_17),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_60),
.B(n_118),
.C(n_39),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_61),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_62),
.Y(n_155)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_64),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_31),
.B(n_9),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_65),
.B(n_19),
.Y(n_136)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_67),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_35),
.B(n_9),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_68),
.B(n_101),
.Y(n_132)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_69),
.Y(n_184)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_72),
.Y(n_190)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_73),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_74),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_75),
.Y(n_181)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_77),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_80),
.Y(n_161)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g156 ( 
.A(n_82),
.Y(n_156)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_85),
.Y(n_178)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_87),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_88),
.Y(n_177)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_89),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_52),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_93),
.A2(n_33),
.B1(n_38),
.B2(n_37),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_95),
.Y(n_149)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_97),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_99),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_100),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_23),
.B(n_8),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_102),
.Y(n_167)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_103),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_104),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_105),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_106),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_107),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_108),
.Y(n_170)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_109),
.Y(n_192)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_23),
.Y(n_110)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_20),
.B(n_11),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_122),
.Y(n_123)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_40),
.Y(n_112)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_23),
.Y(n_113)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_115),
.Y(n_180)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_42),
.Y(n_116)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_116),
.Y(n_183)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_47),
.Y(n_117)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_117),
.Y(n_189)
);

AOI21xp33_ASAP7_75t_L g118 ( 
.A1(n_54),
.A2(n_41),
.B(n_19),
.Y(n_118)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_120),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_121),
.Y(n_148)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_19),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_65),
.B(n_20),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_133),
.B(n_168),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_136),
.A2(n_1),
.B(n_2),
.Y(n_262)
);

AOI21xp33_ASAP7_75t_SL g236 ( 
.A1(n_137),
.A2(n_51),
.B(n_26),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_68),
.A2(n_36),
.B1(n_22),
.B2(n_55),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_138),
.A2(n_172),
.B1(n_179),
.B2(n_32),
.Y(n_204)
);

HAxp5_ASAP7_75t_SL g142 ( 
.A(n_101),
.B(n_48),
.CON(n_142),
.SN(n_142)
);

NAND2xp33_ASAP7_75t_SL g261 ( 
.A(n_142),
.B(n_153),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_67),
.A2(n_36),
.B1(n_40),
.B2(n_39),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_150),
.A2(n_151),
.B1(n_201),
.B2(n_32),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_98),
.A2(n_36),
.B1(n_40),
.B2(n_39),
.Y(n_151)
);

AO22x2_ASAP7_75t_L g153 ( 
.A1(n_63),
.A2(n_48),
.B1(n_41),
.B2(n_42),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_89),
.B(n_28),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_158),
.B(n_159),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_73),
.B(n_28),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_164),
.A2(n_32),
.B1(n_29),
.B2(n_33),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_113),
.B(n_30),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_114),
.B(n_41),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_188),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_61),
.A2(n_26),
.B1(n_55),
.B2(n_53),
.Y(n_172)
);

AND2x2_ASAP7_75t_SL g174 ( 
.A(n_62),
.B(n_42),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_174),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_64),
.A2(n_33),
.B1(n_29),
.B2(n_38),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_115),
.B(n_59),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_186),
.B(n_187),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_120),
.Y(n_187)
);

NAND3xp33_ASAP7_75t_L g188 ( 
.A(n_121),
.B(n_59),
.C(n_53),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_72),
.B(n_21),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_197),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_74),
.B(n_22),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_78),
.A2(n_58),
.B1(n_38),
.B2(n_37),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_202),
.A2(n_212),
.B1(n_221),
.B2(n_232),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_204),
.B(n_246),
.Y(n_280)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_205),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_206),
.Y(n_287)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_127),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_207),
.Y(n_317)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_145),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_208),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_140),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_209),
.Y(n_285)
);

BUFx12_ASAP7_75t_L g210 ( 
.A(n_140),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_210),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_L g212 ( 
.A1(n_201),
.A2(n_108),
.B1(n_107),
.B2(n_106),
.Y(n_212)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_194),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_214),
.Y(n_307)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_149),
.Y(n_216)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_216),
.Y(n_305)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_198),
.Y(n_217)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_217),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_135),
.Y(n_218)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_218),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_136),
.A2(n_105),
.B1(n_104),
.B2(n_102),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g328 ( 
.A1(n_219),
.A2(n_270),
.B1(n_1),
.B2(n_3),
.Y(n_328)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_154),
.Y(n_220)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_220),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_123),
.A2(n_24),
.B1(n_30),
.B2(n_21),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_162),
.Y(n_222)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_222),
.Y(n_319)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_166),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_223),
.Y(n_284)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_191),
.Y(n_224)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_224),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_132),
.B(n_51),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_225),
.B(n_240),
.Y(n_311)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_191),
.Y(n_226)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_226),
.Y(n_288)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_145),
.Y(n_227)
);

INVx8_ASAP7_75t_L g289 ( 
.A(n_227),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_228),
.Y(n_301)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_181),
.Y(n_230)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_230),
.Y(n_292)
);

INVx8_ASAP7_75t_L g231 ( 
.A(n_155),
.Y(n_231)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_231),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_148),
.A2(n_58),
.B1(n_37),
.B2(n_34),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_153),
.A2(n_58),
.B1(n_34),
.B2(n_29),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_233),
.A2(n_234),
.B1(n_238),
.B2(n_243),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_188),
.A2(n_171),
.B1(n_156),
.B2(n_170),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_125),
.Y(n_235)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_235),
.Y(n_297)
);

AOI21xp33_ASAP7_75t_L g298 ( 
.A1(n_236),
.A2(n_273),
.B(n_146),
.Y(n_298)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_152),
.Y(n_237)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_237),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_153),
.A2(n_34),
.B1(n_24),
.B2(n_88),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_176),
.Y(n_239)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_239),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_157),
.B(n_94),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_142),
.A2(n_90),
.B1(n_87),
.B2(n_42),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_241),
.B(n_262),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_124),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_242),
.B(n_256),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_179),
.A2(n_42),
.B1(n_48),
.B2(n_12),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_126),
.Y(n_244)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_244),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_135),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_245),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_161),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_155),
.Y(n_247)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_247),
.Y(n_320)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_128),
.Y(n_248)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_248),
.Y(n_331)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_134),
.Y(n_249)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_249),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_131),
.B(n_42),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_250),
.B(n_266),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_192),
.B(n_11),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_251),
.B(n_267),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_175),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_252),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_180),
.A2(n_48),
.B(n_2),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_253),
.A2(n_1),
.B(n_3),
.Y(n_313)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_161),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_254),
.B(n_257),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_175),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_255),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_169),
.B(n_11),
.Y(n_256)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_165),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_199),
.A2(n_11),
.B1(n_16),
.B2(n_15),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_258),
.A2(n_196),
.B1(n_193),
.B2(n_163),
.Y(n_318)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_190),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_259),
.Y(n_306)
);

INVx11_ASAP7_75t_L g260 ( 
.A(n_151),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_260),
.Y(n_312)
);

BUFx4f_ASAP7_75t_SL g263 ( 
.A(n_178),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_263),
.B(n_265),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_160),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_264),
.Y(n_329)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_183),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_139),
.B(n_7),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_143),
.Y(n_267)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_129),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_268),
.B(n_269),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_160),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_150),
.A2(n_12),
.B1(n_15),
.B2(n_5),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_144),
.B(n_5),
.C(n_6),
.Y(n_272)
);

AND2x2_ASAP7_75t_SL g324 ( 
.A(n_272),
.B(n_274),
.Y(n_324)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_147),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_174),
.B(n_5),
.C(n_6),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_182),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_275),
.B(n_278),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_215),
.B(n_182),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_211),
.B(n_163),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_279),
.B(n_316),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_238),
.A2(n_156),
.B1(n_184),
.B2(n_141),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_282),
.A2(n_286),
.B1(n_304),
.B2(n_325),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_229),
.A2(n_184),
.B1(n_141),
.B2(n_177),
.Y(n_286)
);

NOR3xp33_ASAP7_75t_SL g347 ( 
.A(n_298),
.B(n_228),
.C(n_242),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_229),
.A2(n_177),
.B1(n_173),
.B2(n_193),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_313),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_271),
.B(n_196),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_318),
.B(n_246),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_203),
.B(n_173),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_323),
.B(n_327),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_206),
.A2(n_200),
.B1(n_190),
.B2(n_167),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_274),
.B(n_200),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_328),
.A2(n_280),
.B1(n_278),
.B2(n_279),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_261),
.B(n_3),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_330),
.B(n_332),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_272),
.B(n_5),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_233),
.A2(n_129),
.B1(n_130),
.B2(n_167),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_333),
.A2(n_263),
.B1(n_231),
.B2(n_208),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_330),
.A2(n_253),
.B(n_232),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_336),
.A2(n_340),
.B(n_355),
.Y(n_387)
);

AO22x2_ASAP7_75t_L g339 ( 
.A1(n_293),
.A2(n_260),
.B1(n_212),
.B2(n_241),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_339),
.B(n_349),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_313),
.A2(n_213),
.B(n_258),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_287),
.A2(n_217),
.B1(n_257),
.B2(n_214),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g400 ( 
.A1(n_341),
.A2(n_343),
.B1(n_359),
.B2(n_376),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_280),
.A2(n_130),
.B1(n_227),
.B2(n_259),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_342),
.A2(n_348),
.B1(n_351),
.B2(n_371),
.Y(n_397)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_277),
.Y(n_345)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_345),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_347),
.B(n_307),
.Y(n_409)
);

BUFx5_ASAP7_75t_L g350 ( 
.A(n_308),
.Y(n_350)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_350),
.Y(n_394)
);

OAI22xp33_ASAP7_75t_L g351 ( 
.A1(n_312),
.A2(n_287),
.B1(n_280),
.B2(n_325),
.Y(n_351)
);

INVx6_ASAP7_75t_L g352 ( 
.A(n_289),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g395 ( 
.A(n_352),
.Y(n_395)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_315),
.Y(n_353)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_353),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_276),
.A2(n_209),
.B(n_254),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_315),
.Y(n_356)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_356),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_314),
.Y(n_357)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_357),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_320),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_358),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_291),
.A2(n_268),
.B1(n_255),
.B2(n_252),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_276),
.A2(n_287),
.B(n_312),
.Y(n_360)
);

O2A1O1Ixp33_ASAP7_75t_L g419 ( 
.A1(n_360),
.A2(n_364),
.B(n_365),
.C(n_381),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_304),
.B(n_224),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g404 ( 
.A(n_361),
.Y(n_404)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_315),
.Y(n_362)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_362),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_282),
.A2(n_247),
.B1(n_264),
.B2(n_245),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_363),
.A2(n_370),
.B1(n_378),
.B2(n_382),
.Y(n_406)
);

OAI22x1_ASAP7_75t_L g364 ( 
.A1(n_323),
.A2(n_230),
.B1(n_218),
.B2(n_226),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_316),
.A2(n_263),
.B(n_210),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_303),
.Y(n_367)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_367),
.Y(n_410)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_303),
.Y(n_368)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_368),
.Y(n_416)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_277),
.Y(n_369)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_369),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_333),
.A2(n_210),
.B1(n_12),
.B2(n_13),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_327),
.A2(n_18),
.B1(n_6),
.B2(n_13),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_309),
.Y(n_372)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_372),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_311),
.B(n_6),
.Y(n_373)
);

CKINVDCx14_ASAP7_75t_R g389 ( 
.A(n_373),
.Y(n_389)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_309),
.Y(n_374)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_374),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_326),
.B(n_13),
.C(n_324),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_375),
.B(n_377),
.C(n_310),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_295),
.A2(n_321),
.B1(n_311),
.B2(n_275),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_326),
.B(n_324),
.C(n_332),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_286),
.A2(n_306),
.B1(n_324),
.B2(n_281),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_317),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_379),
.B(n_380),
.Y(n_392)
);

INVx5_ASAP7_75t_L g380 ( 
.A(n_289),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_299),
.A2(n_314),
.B(n_292),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_306),
.A2(n_281),
.B1(n_300),
.B2(n_296),
.Y(n_382)
);

BUFx5_ASAP7_75t_L g383 ( 
.A(n_308),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_383),
.Y(n_405)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_297),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_384),
.B(n_283),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_344),
.B(n_300),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_386),
.B(n_403),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_379),
.B(n_292),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_388),
.B(n_413),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_360),
.A2(n_314),
.B(n_329),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_391),
.A2(n_393),
.B(n_424),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_336),
.A2(n_329),
.B(n_301),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_377),
.B(n_335),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_396),
.B(n_398),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_375),
.B(n_335),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_354),
.B(n_310),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_399),
.B(n_421),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_351),
.A2(n_296),
.B1(n_320),
.B2(n_302),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_402),
.A2(n_423),
.B1(n_374),
.B2(n_367),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_354),
.B(n_307),
.Y(n_403)
);

OAI21x1_ASAP7_75t_L g433 ( 
.A1(n_409),
.A2(n_338),
.B(n_365),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_352),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_412),
.B(n_414),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_346),
.B(n_297),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_380),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_415),
.B(n_420),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_371),
.B(n_307),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_378),
.A2(n_302),
.B1(n_331),
.B2(n_319),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_355),
.A2(n_301),
.B(n_283),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_425),
.A2(n_338),
.B1(n_337),
.B2(n_340),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_426),
.A2(n_431),
.B1(n_446),
.B2(n_449),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_415),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_427),
.B(n_433),
.Y(n_477)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_410),
.Y(n_428)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_428),
.Y(n_462)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_410),
.Y(n_429)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_429),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_389),
.B(n_398),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_430),
.B(n_440),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_SL g431 ( 
.A1(n_404),
.A2(n_343),
.B1(n_342),
.B2(n_361),
.Y(n_431)
);

A2O1A1O1Ixp25_ASAP7_75t_L g432 ( 
.A1(n_387),
.A2(n_366),
.B(n_362),
.C(n_356),
.D(n_353),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_432),
.A2(n_424),
.B(n_419),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_409),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_434),
.B(n_444),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_425),
.A2(n_337),
.B1(n_339),
.B2(n_343),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_435),
.A2(n_404),
.B1(n_401),
.B2(n_420),
.Y(n_484)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_416),
.Y(n_436)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_436),
.Y(n_472)
);

OA22x2_ASAP7_75t_L g437 ( 
.A1(n_402),
.A2(n_348),
.B1(n_363),
.B2(n_370),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_437),
.B(n_445),
.Y(n_479)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_416),
.Y(n_438)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_438),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_386),
.B(n_334),
.Y(n_440)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_418),
.Y(n_442)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_442),
.Y(n_475)
);

MAJx2_ASAP7_75t_L g443 ( 
.A(n_396),
.B(n_347),
.C(n_357),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_443),
.B(n_421),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_392),
.Y(n_444)
);

OA22x2_ASAP7_75t_L g445 ( 
.A1(n_397),
.A2(n_339),
.B1(n_382),
.B2(n_364),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_425),
.A2(n_339),
.B1(n_381),
.B2(n_361),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_403),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_448),
.B(n_422),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_400),
.A2(n_339),
.B1(n_372),
.B2(n_368),
.Y(n_451)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_451),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_408),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_453),
.B(n_456),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_397),
.A2(n_384),
.B1(n_358),
.B2(n_369),
.Y(n_454)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_454),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_419),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_399),
.B(n_345),
.Y(n_457)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_457),
.Y(n_488)
);

AO22x2_ASAP7_75t_L g458 ( 
.A1(n_406),
.A2(n_319),
.B1(n_288),
.B2(n_331),
.Y(n_458)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_458),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_406),
.A2(n_302),
.B1(n_288),
.B2(n_284),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_459),
.A2(n_423),
.B1(n_385),
.B2(n_407),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_385),
.B(n_285),
.Y(n_461)
);

CKINVDCx14_ASAP7_75t_R g476 ( 
.A(n_461),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_463),
.A2(n_484),
.B1(n_461),
.B2(n_453),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_464),
.B(n_426),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_439),
.B(n_407),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_466),
.B(n_481),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_460),
.B(n_455),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_467),
.B(n_473),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_470),
.A2(n_452),
.B1(n_429),
.B2(n_436),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_460),
.B(n_387),
.Y(n_473)
);

XNOR2x1_ASAP7_75t_SL g480 ( 
.A(n_441),
.B(n_390),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_480),
.B(n_445),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_450),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_455),
.B(n_390),
.C(n_401),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_482),
.B(n_485),
.C(n_490),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_456),
.A2(n_393),
.B(n_391),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_483),
.A2(n_434),
.B(n_447),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_443),
.B(n_422),
.C(n_418),
.Y(n_485)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_489),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_457),
.B(n_414),
.C(n_334),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_441),
.B(n_412),
.C(n_417),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_491),
.B(n_450),
.Y(n_496)
);

FAx1_ASAP7_75t_SL g493 ( 
.A(n_432),
.B(n_405),
.CI(n_417),
.CON(n_493),
.SN(n_493)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_493),
.B(n_458),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_494),
.B(n_510),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_495),
.B(n_496),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_487),
.A2(n_446),
.B(n_447),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_498),
.B(n_515),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_467),
.B(n_435),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_499),
.B(n_502),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_478),
.A2(n_452),
.B1(n_444),
.B2(n_459),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_500),
.A2(n_509),
.B1(n_511),
.B2(n_517),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_501),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_482),
.B(n_458),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_471),
.Y(n_503)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_503),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_504),
.A2(n_479),
.B1(n_492),
.B2(n_487),
.Y(n_539)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_469),
.Y(n_505)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_505),
.Y(n_528)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_471),
.Y(n_506)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_506),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_478),
.A2(n_445),
.B1(n_458),
.B2(n_442),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_468),
.A2(n_445),
.B1(n_458),
.B2(n_438),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_462),
.Y(n_513)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_513),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_SL g514 ( 
.A(n_473),
.B(n_428),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_514),
.B(n_516),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_485),
.B(n_437),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_476),
.A2(n_395),
.B1(n_437),
.B2(n_408),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_466),
.B(n_411),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_518),
.B(n_519),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_486),
.A2(n_395),
.B1(n_437),
.B2(n_405),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_479),
.A2(n_395),
.B1(n_411),
.B2(n_394),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_520),
.B(n_470),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_508),
.B(n_491),
.C(n_490),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_521),
.B(n_523),
.Y(n_562)
);

NOR3xp33_ASAP7_75t_SL g522 ( 
.A(n_512),
.B(n_497),
.C(n_477),
.Y(n_522)
);

OAI221xp5_ASAP7_75t_L g559 ( 
.A1(n_522),
.A2(n_525),
.B1(n_472),
.B2(n_475),
.C(n_394),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_508),
.B(n_464),
.C(n_488),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_496),
.B(n_465),
.Y(n_524)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_524),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_516),
.B(n_465),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_507),
.B(n_514),
.C(n_499),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_529),
.B(n_530),
.C(n_535),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_507),
.B(n_488),
.C(n_463),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_494),
.B(n_480),
.C(n_481),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_539),
.B(n_510),
.Y(n_545)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_540),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_502),
.B(n_483),
.C(n_484),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_542),
.B(n_520),
.C(n_509),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_545),
.B(n_561),
.Y(n_567)
);

FAx1_ASAP7_75t_SL g546 ( 
.A(n_535),
.B(n_523),
.CI(n_530),
.CON(n_546),
.SN(n_546)
);

AOI22xp33_ASAP7_75t_SL g570 ( 
.A1(n_546),
.A2(n_529),
.B1(n_543),
.B2(n_541),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_521),
.B(n_500),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_547),
.B(n_558),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_538),
.A2(n_486),
.B1(n_498),
.B2(n_479),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_548),
.A2(n_560),
.B1(n_528),
.B2(n_290),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_542),
.B(n_495),
.Y(n_549)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_549),
.Y(n_564)
);

AOI21x1_ASAP7_75t_L g551 ( 
.A1(n_526),
.A2(n_493),
.B(n_474),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_551),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_552),
.B(n_556),
.Y(n_575)
);

A2O1A1Ixp33_ASAP7_75t_L g553 ( 
.A1(n_539),
.A2(n_492),
.B(n_493),
.C(n_469),
.Y(n_553)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_553),
.Y(n_565)
);

INVxp33_ASAP7_75t_SL g554 ( 
.A(n_533),
.Y(n_554)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_554),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_SL g556 ( 
.A1(n_522),
.A2(n_513),
.B(n_511),
.Y(n_556)
);

FAx1_ASAP7_75t_L g557 ( 
.A(n_531),
.B(n_474),
.CI(n_462),
.CON(n_557),
.SN(n_557)
);

OAI21xp5_ASAP7_75t_SL g568 ( 
.A1(n_557),
.A2(n_537),
.B(n_536),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_531),
.B(n_475),
.Y(n_558)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_559),
.Y(n_573)
);

OAI221xp5_ASAP7_75t_L g560 ( 
.A1(n_527),
.A2(n_472),
.B1(n_284),
.B2(n_322),
.C(n_305),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_532),
.B(n_305),
.Y(n_561)
);

CKINVDCx16_ASAP7_75t_R g566 ( 
.A(n_557),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_566),
.B(n_569),
.Y(n_583)
);

INVxp67_ASAP7_75t_L g586 ( 
.A(n_568),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_SL g569 ( 
.A(n_544),
.B(n_534),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_570),
.A2(n_574),
.B(n_383),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_572),
.B(n_550),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_547),
.B(n_532),
.C(n_541),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_SL g577 ( 
.A1(n_557),
.A2(n_543),
.B(n_350),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_SL g579 ( 
.A1(n_577),
.A2(n_549),
.B(n_553),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_573),
.B(n_555),
.Y(n_578)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_578),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_579),
.B(n_580),
.Y(n_591)
);

XOR2xp5_ASAP7_75t_L g580 ( 
.A(n_567),
.B(n_552),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_574),
.B(n_562),
.Y(n_581)
);

NOR2x1_ASAP7_75t_SL g592 ( 
.A(n_581),
.B(n_571),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_573),
.A2(n_554),
.B1(n_545),
.B2(n_558),
.Y(n_582)
);

OAI21x1_ASAP7_75t_L g593 ( 
.A1(n_582),
.A2(n_587),
.B(n_589),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_SL g584 ( 
.A1(n_565),
.A2(n_546),
.B1(n_550),
.B2(n_561),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_584),
.A2(n_588),
.B(n_577),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_564),
.B(n_576),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_585),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_564),
.B(n_285),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_SL g590 ( 
.A1(n_587),
.A2(n_575),
.B(n_563),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_L g600 ( 
.A1(n_590),
.A2(n_584),
.B(n_586),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_592),
.Y(n_601)
);

AOI21x1_ASAP7_75t_L g598 ( 
.A1(n_595),
.A2(n_583),
.B(n_571),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_581),
.A2(n_563),
.B(n_565),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_596),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_L g604 ( 
.A1(n_598),
.A2(n_597),
.B1(n_586),
.B2(n_591),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_594),
.B(n_582),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_599),
.B(n_568),
.Y(n_605)
);

AOI21x1_ASAP7_75t_L g603 ( 
.A1(n_600),
.A2(n_593),
.B(n_591),
.Y(n_603)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_603),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_604),
.B(n_605),
.C(n_602),
.Y(n_606)
);

AOI21xp33_ASAP7_75t_L g608 ( 
.A1(n_606),
.A2(n_601),
.B(n_580),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_608),
.B(n_607),
.C(n_567),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_609),
.B(n_322),
.C(n_294),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g611 ( 
.A(n_610),
.B(n_294),
.Y(n_611)
);


endmodule