module fake_jpeg_26418_n_308 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_308);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_44),
.B(n_48),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_42),
.A2(n_31),
.B1(n_18),
.B2(n_22),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_45),
.A2(n_34),
.B1(n_33),
.B2(n_32),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_46),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_38),
.C(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_22),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_53),
.B(n_18),
.Y(n_77)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_23),
.C(n_26),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_37),
.Y(n_74)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_65),
.Y(n_69)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_66),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_34),
.B1(n_41),
.B2(n_38),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_67),
.A2(n_71),
.B1(n_89),
.B2(n_64),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_41),
.B1(n_34),
.B2(n_31),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_16),
.B1(n_21),
.B2(n_20),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_74),
.A2(n_77),
.B(n_32),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_37),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_36),
.Y(n_111)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_81),
.A2(n_87),
.B1(n_73),
.B2(n_32),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_51),
.B(n_37),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_84),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_33),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_50),
.B(n_39),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_37),
.Y(n_96)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_50),
.A2(n_27),
.B1(n_21),
.B2(n_20),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_59),
.A2(n_41),
.B1(n_28),
.B2(n_26),
.Y(n_89)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_93),
.B(n_98),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_111),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_27),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_97),
.B(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_43),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_106),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_71),
.A2(n_64),
.B1(n_55),
.B2(n_43),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_112),
.B1(n_73),
.B2(n_80),
.Y(n_126)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_103),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_79),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_104),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_101),
.B1(n_102),
.B2(n_109),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_39),
.C(n_47),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_70),
.A2(n_0),
.B(n_1),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_110),
.Y(n_124)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_115),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_54),
.C(n_40),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_73),
.A2(n_61),
.B1(n_41),
.B2(n_56),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_33),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_85),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_30),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_68),
.B(n_30),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_24),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_91),
.B1(n_69),
.B2(n_56),
.Y(n_146)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_126),
.A2(n_130),
.B1(n_78),
.B2(n_112),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_136),
.Y(n_158)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_128),
.A2(n_40),
.B1(n_23),
.B2(n_26),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_135),
.B(n_97),
.Y(n_160)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_144),
.Y(n_165)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_105),
.A2(n_85),
.B1(n_88),
.B2(n_80),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_140),
.A2(n_142),
.B1(n_61),
.B2(n_79),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_100),
.A2(n_82),
.B1(n_90),
.B2(n_88),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_24),
.B1(n_75),
.B2(n_40),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_92),
.A2(n_85),
.B1(n_82),
.B2(n_90),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_93),
.B(n_91),
.Y(n_145)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_146),
.A2(n_104),
.B(n_115),
.Y(n_154)
);

AOI32xp33_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_111),
.A3(n_106),
.B1(n_110),
.B2(n_113),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_147),
.A2(n_149),
.B(n_150),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_143),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_148),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_129),
.A2(n_111),
.B(n_107),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_129),
.A2(n_117),
.B(n_106),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_110),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_163),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_133),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_153),
.B(n_168),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_154),
.A2(n_166),
.B1(n_172),
.B2(n_176),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_116),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_160),
.Y(n_191)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_98),
.B(n_114),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_157),
.A2(n_134),
.B1(n_123),
.B2(n_24),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_142),
.A2(n_108),
.B(n_1),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_159),
.A2(n_175),
.B(n_0),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_78),
.C(n_75),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_170),
.B1(n_139),
.B2(n_143),
.Y(n_179)
);

OAI22x1_ASAP7_75t_SL g166 ( 
.A1(n_140),
.A2(n_79),
.B1(n_75),
.B2(n_28),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_141),
.Y(n_168)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_121),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_120),
.Y(n_190)
);

XOR2x2_ASAP7_75t_L g173 ( 
.A(n_124),
.B(n_25),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_120),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_136),
.A2(n_138),
.B1(n_144),
.B2(n_130),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_174),
.A2(n_145),
.B1(n_128),
.B2(n_125),
.Y(n_182)
);

AND2x4_ASAP7_75t_L g175 ( 
.A(n_127),
.B(n_25),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_179),
.A2(n_193),
.B1(n_17),
.B2(n_19),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_131),
.B1(n_132),
.B2(n_134),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_180),
.A2(n_197),
.B1(n_198),
.B2(n_201),
.Y(n_213)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_186),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_182),
.A2(n_167),
.B1(n_156),
.B2(n_152),
.Y(n_205)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_184),
.A2(n_171),
.B1(n_152),
.B2(n_165),
.Y(n_206)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_158),
.Y(n_208)
);

INVxp33_ASAP7_75t_SL g189 ( 
.A(n_173),
.Y(n_189)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_189),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_190),
.Y(n_207)
);

AOI322xp5_ASAP7_75t_L g192 ( 
.A1(n_175),
.A2(n_149),
.A3(n_150),
.B1(n_151),
.B2(n_154),
.C1(n_155),
.C2(n_174),
.Y(n_192)
);

BUFx24_ASAP7_75t_SL g222 ( 
.A(n_192),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_162),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_194),
.Y(n_218)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_202),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_196),
.A2(n_199),
.B(n_172),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_169),
.A2(n_137),
.B1(n_121),
.B2(n_28),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_169),
.A2(n_28),
.B1(n_26),
.B2(n_23),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_175),
.A2(n_0),
.B(n_1),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_162),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_200),
.B(n_19),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_175),
.A2(n_19),
.B1(n_17),
.B2(n_25),
.Y(n_201)
);

AO22x1_ASAP7_75t_SL g202 ( 
.A1(n_159),
.A2(n_19),
.B1(n_17),
.B2(n_4),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_203),
.A2(n_212),
.B(n_217),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_205),
.A2(n_219),
.B1(n_220),
.B2(n_211),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_206),
.A2(n_216),
.B1(n_180),
.B2(n_179),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_210),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_158),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_196),
.A2(n_160),
.B(n_19),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_214),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_215),
.A2(n_178),
.B1(n_181),
.B2(n_194),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_184),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_187),
.A2(n_15),
.B(n_14),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_182),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_183),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_177),
.B(n_15),
.C(n_14),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_188),
.C(n_193),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_199),
.A2(n_2),
.B(n_3),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_224),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_187),
.A2(n_2),
.B(n_5),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_185),
.A2(n_5),
.B(n_6),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_225),
.Y(n_230)
);

INVxp33_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_226),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_195),
.Y(n_227)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_227),
.Y(n_251)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_228),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_231),
.B(n_237),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_218),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_232),
.Y(n_247)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_235),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_236),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_220),
.A2(n_197),
.B1(n_198),
.B2(n_186),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_204),
.B(n_201),
.Y(n_238)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_238),
.B(n_213),
.CI(n_219),
.CON(n_258),
.SN(n_258)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_204),
.A2(n_202),
.B1(n_6),
.B2(n_7),
.Y(n_242)
);

INVx3_ASAP7_75t_SL g252 ( 
.A(n_242),
.Y(n_252)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_205),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_208),
.C(n_210),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_213),
.A2(n_202),
.B1(n_191),
.B2(n_5),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_246),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_211),
.A2(n_191),
.B1(n_8),
.B2(n_11),
.Y(n_246)
);

MAJx2_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_245),
.C(n_246),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_234),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_254),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_224),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_207),
.C(n_221),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_230),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_258),
.A2(n_245),
.B1(n_241),
.B2(n_229),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_227),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_259),
.Y(n_272)
);

NAND2x1_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_203),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_228),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_231),
.C(n_222),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_265),
.Y(n_279)
);

NOR2xp67_ASAP7_75t_SL g263 ( 
.A(n_260),
.B(n_217),
.Y(n_263)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_250),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_237),
.C(n_238),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_250),
.B(n_239),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_225),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_243),
.C(n_244),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_271),
.Y(n_284)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_252),
.A2(n_230),
.B1(n_229),
.B2(n_207),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_269),
.A2(n_257),
.B1(n_261),
.B2(n_258),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_247),
.C(n_254),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_273),
.A2(n_252),
.B1(n_248),
.B2(n_251),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_274),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_275),
.A2(n_274),
.B(n_269),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_285),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_280),
.A2(n_10),
.B1(n_12),
.B2(n_15),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_257),
.C(n_258),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_270),
.C(n_272),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_272),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_283),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_279),
.B(n_281),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_289),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_288),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_284),
.A2(n_212),
.B(n_223),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_291),
.A2(n_282),
.B1(n_278),
.B2(n_277),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_12),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_293),
.B(n_277),
.Y(n_298)
);

INVx11_ASAP7_75t_L g294 ( 
.A(n_290),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_296),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_299),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_292),
.B(n_275),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_293),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_295),
.Y(n_303)
);

OAI311xp33_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_295),
.A3(n_301),
.B1(n_294),
.C1(n_296),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_300),
.C(n_10),
.Y(n_305)
);

OAI21x1_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_10),
.B(n_8),
.Y(n_306)
);

BUFx24_ASAP7_75t_SL g307 ( 
.A(n_306),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_8),
.Y(n_308)
);


endmodule