module fake_jpeg_11536_n_146 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_146);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_28),
.B(n_14),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_11),
.Y(n_55)
);

INVx11_ASAP7_75t_SL g56 ( 
.A(n_34),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_3),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_17),
.B(n_7),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_62),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_66),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_67),
.B(n_69),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_1),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_47),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_61),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_77),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_46),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_57),
.B1(n_60),
.B2(n_50),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_78),
.A2(n_54),
.B1(n_48),
.B2(n_68),
.Y(n_92)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_45),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_76),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_45),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_82),
.B(n_1),
.Y(n_98)
);

HAxp5_ASAP7_75t_SL g84 ( 
.A(n_66),
.B(n_56),
.CON(n_84),
.SN(n_84)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_55),
.C(n_52),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_78),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_99),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_88),
.A2(n_95),
.B(n_2),
.Y(n_102)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_91),
.B(n_98),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_92),
.A2(n_8),
.B1(n_9),
.B2(n_12),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_46),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_97),
.Y(n_117)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_74),
.A2(n_56),
.B1(n_54),
.B2(n_3),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_23),
.C(n_39),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

AND2x6_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_21),
.Y(n_100)
);

NOR2x1_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_27),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_13),
.B(n_18),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_109),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_89),
.B(n_5),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_103),
.B(n_114),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_7),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_105),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_111),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_101),
.A2(n_8),
.B1(n_9),
.B2(n_83),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_118),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_113),
.A2(n_31),
.B(n_33),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_85),
.B(n_86),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_100),
.B(n_20),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_24),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_36),
.C(n_37),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_115),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_123),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_25),
.C(n_30),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_124),
.C(n_128),
.Y(n_133)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_125),
.Y(n_136)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_105),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_134),
.C(n_122),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_107),
.C(n_112),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_135),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_138),
.C(n_139),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_129),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_123),
.B(n_127),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_131),
.B(n_133),
.Y(n_142)
);

AOI322xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_116),
.A3(n_106),
.B1(n_130),
.B2(n_109),
.C1(n_42),
.C2(n_38),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_110),
.B(n_130),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_106),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_110),
.Y(n_146)
);


endmodule