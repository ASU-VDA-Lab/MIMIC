module fake_jpeg_12978_n_124 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_124);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_124;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx2_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_2),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g71 ( 
.A(n_51),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_52),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_19),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_56),
.Y(n_60)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_55),
.Y(n_70)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_58),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_0),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_37),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_62),
.B(n_6),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_56),
.A2(n_46),
.B1(n_44),
.B2(n_35),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_63),
.A2(n_67),
.B1(n_40),
.B2(n_42),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_51),
.A2(n_46),
.B1(n_44),
.B2(n_33),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_72),
.Y(n_75)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_74),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_41),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_79),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_64),
.A2(n_45),
.B1(n_36),
.B2(n_42),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_80),
.B1(n_75),
.B2(n_86),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_63),
.A2(n_71),
.B1(n_64),
.B2(n_65),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_1),
.B(n_3),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_6),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_83),
.Y(n_97)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_1),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_85),
.Y(n_98)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_4),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_87),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_4),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_7),
.Y(n_100)
);

AO21x2_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_22),
.B(n_28),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_96),
.Y(n_112)
);

AND2x6_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_31),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_94),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

AND2x6_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_21),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_102),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_82),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_103),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_7),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_87),
.B(n_13),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_104),
.A2(n_18),
.B(n_23),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_16),
.C(n_17),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_110),
.B(n_104),
.C(n_97),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_101),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_112),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_113),
.B(n_115),
.Y(n_117)
);

OA21x2_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_90),
.B(n_98),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_116),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_117),
.B(n_114),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_118),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_109),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_111),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_111),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_108),
.Y(n_124)
);


endmodule