module real_aes_6370_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g107 ( .A(n_0), .Y(n_107) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_1), .A2(n_130), .B(n_134), .C(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g183 ( .A(n_2), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_3), .A2(n_125), .B(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_4), .B(n_147), .Y(n_466) );
AOI21xp33_ASAP7_75t_L g151 ( .A1(n_5), .A2(n_125), .B(n_152), .Y(n_151) );
AND2x6_ASAP7_75t_L g130 ( .A(n_6), .B(n_131), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_7), .A2(n_233), .B(n_234), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_8), .B(n_40), .Y(n_108) );
INVx1_ASAP7_75t_L g522 ( .A(n_9), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_10), .B(n_156), .Y(n_501) );
INVx1_ASAP7_75t_L g158 ( .A(n_11), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_12), .B(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g123 ( .A(n_13), .Y(n_123) );
INVx1_ASAP7_75t_L g239 ( .A(n_14), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_15), .A2(n_142), .B(n_240), .C(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_16), .B(n_147), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_17), .B(n_139), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_18), .B(n_125), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_19), .B(n_550), .Y(n_549) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_20), .A2(n_166), .B(n_225), .C(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_21), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_22), .B(n_156), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_23), .A2(n_237), .B(n_238), .C(n_240), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_24), .B(n_156), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g446 ( .A(n_25), .Y(n_446) );
INVx1_ASAP7_75t_L g472 ( .A(n_26), .Y(n_472) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_27), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_28), .Y(n_497) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_29), .A2(n_43), .B1(n_101), .B2(n_714), .C1(n_715), .C2(n_719), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_30), .B(n_156), .Y(n_185) );
INVx1_ASAP7_75t_L g547 ( .A(n_31), .Y(n_547) );
INVx1_ASAP7_75t_L g172 ( .A(n_32), .Y(n_172) );
INVx2_ASAP7_75t_L g128 ( .A(n_33), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_34), .Y(n_503) );
A2O1A1Ixp33_ASAP7_75t_L g463 ( .A1(n_35), .A2(n_143), .B(n_225), .C(n_464), .Y(n_463) );
INVxp67_ASAP7_75t_L g548 ( .A(n_36), .Y(n_548) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_37), .A2(n_130), .B(n_134), .C(n_197), .Y(n_196) );
CKINVDCx14_ASAP7_75t_R g462 ( .A(n_38), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_39), .A2(n_134), .B(n_471), .C(n_476), .Y(n_470) );
INVx1_ASAP7_75t_L g170 ( .A(n_41), .Y(n_170) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_42), .A2(n_99), .B1(n_722), .B2(n_731), .C1(n_738), .C2(n_744), .Y(n_98) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_42), .A2(n_436), .B1(n_437), .B2(n_733), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_42), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_43), .Y(n_714) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_44), .A2(n_155), .B(n_201), .C(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_45), .B(n_156), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_46), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_47), .Y(n_544) );
INVx1_ASAP7_75t_L g487 ( .A(n_48), .Y(n_487) );
CKINVDCx16_ASAP7_75t_R g173 ( .A(n_49), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_50), .B(n_125), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g165 ( .A1(n_51), .A2(n_134), .B1(n_166), .B2(n_168), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_52), .Y(n_205) );
CKINVDCx16_ASAP7_75t_R g180 ( .A(n_53), .Y(n_180) );
A2O1A1Ixp33_ASAP7_75t_L g154 ( .A1(n_54), .A2(n_143), .B(n_155), .C(n_157), .Y(n_154) );
CKINVDCx14_ASAP7_75t_R g519 ( .A(n_55), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_56), .Y(n_215) );
INVx1_ASAP7_75t_L g153 ( .A(n_57), .Y(n_153) );
INVx1_ASAP7_75t_L g131 ( .A(n_58), .Y(n_131) );
INVx1_ASAP7_75t_L g122 ( .A(n_59), .Y(n_122) );
INVx1_ASAP7_75t_SL g465 ( .A(n_60), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_61), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_62), .B(n_147), .Y(n_491) );
INVx1_ASAP7_75t_L g449 ( .A(n_63), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_SL g138 ( .A1(n_64), .A2(n_139), .B(n_140), .C(n_143), .Y(n_138) );
INVxp67_ASAP7_75t_L g141 ( .A(n_65), .Y(n_141) );
INVx1_ASAP7_75t_L g726 ( .A(n_66), .Y(n_726) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_67), .A2(n_125), .B(n_518), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_68), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_69), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_70), .A2(n_125), .B(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g208 ( .A(n_71), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_72), .B(n_736), .Y(n_737) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_73), .A2(n_233), .B(n_543), .Y(n_542) );
CKINVDCx16_ASAP7_75t_R g469 ( .A(n_74), .Y(n_469) );
INVx1_ASAP7_75t_L g507 ( .A(n_75), .Y(n_507) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_76), .A2(n_130), .B(n_134), .C(n_210), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_77), .A2(n_125), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g510 ( .A(n_78), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_79), .B(n_184), .Y(n_198) );
INVx2_ASAP7_75t_L g120 ( .A(n_80), .Y(n_120) );
INVx1_ASAP7_75t_L g500 ( .A(n_81), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_82), .B(n_139), .Y(n_199) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_83), .A2(n_130), .B(n_134), .C(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g105 ( .A(n_84), .Y(n_105) );
OR2x2_ASAP7_75t_L g435 ( .A(n_84), .B(n_106), .Y(n_435) );
OR2x2_ASAP7_75t_L g730 ( .A(n_84), .B(n_718), .Y(n_730) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_85), .A2(n_134), .B(n_448), .C(n_452), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_86), .B(n_160), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_87), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_88), .A2(n_130), .B(n_134), .C(n_222), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_89), .Y(n_229) );
INVx1_ASAP7_75t_L g137 ( .A(n_90), .Y(n_137) );
CKINVDCx16_ASAP7_75t_R g235 ( .A(n_91), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_92), .B(n_184), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_93), .B(n_118), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_94), .B(n_118), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g124 ( .A1(n_95), .A2(n_125), .B(n_132), .Y(n_124) );
INVx2_ASAP7_75t_L g490 ( .A(n_96), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_97), .B(n_726), .Y(n_725) );
INVxp67_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AOI22xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_109), .B1(n_434), .B2(n_436), .Y(n_102) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_103), .A2(n_434), .B1(n_437), .B2(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
OR2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
NOR2x2_ASAP7_75t_L g717 ( .A(n_105), .B(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_106), .Y(n_718) );
AND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
INVx2_ASAP7_75t_L g721 ( .A(n_109), .Y(n_721) );
INVx3_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND4x1_ASAP7_75t_L g110 ( .A(n_111), .B(n_352), .C(n_399), .D(n_419), .Y(n_110) );
NOR3xp33_ASAP7_75t_SL g111 ( .A(n_112), .B(n_282), .C(n_307), .Y(n_111) );
OAI211xp5_ASAP7_75t_SL g112 ( .A1(n_113), .A2(n_190), .B(n_242), .C(n_272), .Y(n_112) );
INVxp67_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_161), .Y(n_114) );
INVx3_ASAP7_75t_SL g324 ( .A(n_115), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_115), .B(n_255), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_115), .B(n_177), .Y(n_405) );
AND2x2_ASAP7_75t_L g428 ( .A(n_115), .B(n_294), .Y(n_428) );
AND2x4_ASAP7_75t_L g115 ( .A(n_116), .B(n_149), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AND2x2_ASAP7_75t_L g246 ( .A(n_117), .B(n_150), .Y(n_246) );
INVx3_ASAP7_75t_L g259 ( .A(n_117), .Y(n_259) );
AND2x2_ASAP7_75t_L g264 ( .A(n_117), .B(n_149), .Y(n_264) );
OR2x2_ASAP7_75t_L g315 ( .A(n_117), .B(n_256), .Y(n_315) );
BUFx2_ASAP7_75t_L g335 ( .A(n_117), .Y(n_335) );
AND2x2_ASAP7_75t_L g345 ( .A(n_117), .B(n_256), .Y(n_345) );
AND2x2_ASAP7_75t_L g351 ( .A(n_117), .B(n_162), .Y(n_351) );
OA21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_124), .B(n_146), .Y(n_117) );
INVx4_ASAP7_75t_L g148 ( .A(n_118), .Y(n_148) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_118), .Y(n_459) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g163 ( .A(n_119), .Y(n_163) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
AND2x2_ASAP7_75t_SL g160 ( .A(n_120), .B(n_121), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
BUFx2_ASAP7_75t_L g233 ( .A(n_125), .Y(n_233) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_130), .Y(n_125) );
NAND2x1p5_ASAP7_75t_L g174 ( .A(n_126), .B(n_130), .Y(n_174) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_129), .Y(n_126) );
INVx1_ASAP7_75t_L g475 ( .A(n_127), .Y(n_475) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g135 ( .A(n_128), .Y(n_135) );
INVx1_ASAP7_75t_L g167 ( .A(n_128), .Y(n_167) );
INVx1_ASAP7_75t_L g136 ( .A(n_129), .Y(n_136) );
INVx1_ASAP7_75t_L g139 ( .A(n_129), .Y(n_139) );
INVx3_ASAP7_75t_L g142 ( .A(n_129), .Y(n_142) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_129), .Y(n_156) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_129), .Y(n_169) );
INVx4_ASAP7_75t_SL g145 ( .A(n_130), .Y(n_145) );
BUFx3_ASAP7_75t_L g476 ( .A(n_130), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_137), .B(n_138), .C(n_145), .Y(n_132) );
O2A1O1Ixp33_ASAP7_75t_L g152 ( .A1(n_133), .A2(n_145), .B(n_153), .C(n_154), .Y(n_152) );
O2A1O1Ixp33_ASAP7_75t_L g234 ( .A1(n_133), .A2(n_145), .B(n_235), .C(n_236), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_133), .A2(n_145), .B(n_462), .C(n_463), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_SL g486 ( .A1(n_133), .A2(n_145), .B(n_487), .C(n_488), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_SL g506 ( .A1(n_133), .A2(n_145), .B(n_507), .C(n_508), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_SL g518 ( .A1(n_133), .A2(n_145), .B(n_519), .C(n_520), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_SL g543 ( .A1(n_133), .A2(n_145), .B(n_544), .C(n_545), .Y(n_543) );
INVx5_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x6_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_135), .Y(n_144) );
BUFx3_ASAP7_75t_L g202 ( .A(n_135), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_142), .B(n_158), .Y(n_157) );
INVx5_ASAP7_75t_L g184 ( .A(n_142), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_142), .B(n_522), .Y(n_521) );
INVx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_144), .Y(n_226) );
OAI22xp33_ASAP7_75t_L g164 ( .A1(n_145), .A2(n_165), .B1(n_173), .B2(n_174), .Y(n_164) );
INVx1_ASAP7_75t_L g452 ( .A(n_145), .Y(n_452) );
OA21x2_ASAP7_75t_L g150 ( .A1(n_147), .A2(n_151), .B(n_159), .Y(n_150) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NOR2xp33_ASAP7_75t_SL g204 ( .A(n_148), .B(n_205), .Y(n_204) );
AO21x2_ASAP7_75t_L g444 ( .A1(n_148), .A2(n_445), .B(n_453), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_148), .B(n_478), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_148), .B(n_503), .Y(n_502) );
INVx1_ASAP7_75t_SL g149 ( .A(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_150), .B(n_256), .Y(n_270) );
INVx2_ASAP7_75t_L g280 ( .A(n_150), .Y(n_280) );
AND2x2_ASAP7_75t_L g293 ( .A(n_150), .B(n_259), .Y(n_293) );
OR2x2_ASAP7_75t_L g304 ( .A(n_150), .B(n_256), .Y(n_304) );
AND2x2_ASAP7_75t_SL g350 ( .A(n_150), .B(n_351), .Y(n_350) );
BUFx2_ASAP7_75t_L g362 ( .A(n_150), .Y(n_362) );
AND2x2_ASAP7_75t_L g408 ( .A(n_150), .B(n_162), .Y(n_408) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx4_ASAP7_75t_L g225 ( .A(n_156), .Y(n_225) );
INVx1_ASAP7_75t_L g189 ( .A(n_160), .Y(n_189) );
INVx2_ASAP7_75t_L g219 ( .A(n_160), .Y(n_219) );
OA21x2_ASAP7_75t_L g231 ( .A1(n_160), .A2(n_232), .B(n_241), .Y(n_231) );
O2A1O1Ixp33_ASAP7_75t_L g468 ( .A1(n_160), .A2(n_174), .B(n_469), .C(n_470), .Y(n_468) );
OA21x2_ASAP7_75t_L g516 ( .A1(n_160), .A2(n_517), .B(n_523), .Y(n_516) );
INVx3_ASAP7_75t_SL g281 ( .A(n_161), .Y(n_281) );
OR2x2_ASAP7_75t_L g334 ( .A(n_161), .B(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_177), .Y(n_161) );
INVx3_ASAP7_75t_L g256 ( .A(n_162), .Y(n_256) );
AND2x2_ASAP7_75t_L g323 ( .A(n_162), .B(n_178), .Y(n_323) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_162), .Y(n_391) );
AOI33xp33_ASAP7_75t_L g395 ( .A1(n_162), .A2(n_324), .A3(n_331), .B1(n_340), .B2(n_396), .B3(n_397), .Y(n_395) );
AO21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .B(n_175), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_163), .B(n_176), .Y(n_175) );
AO21x2_ASAP7_75t_L g178 ( .A1(n_163), .A2(n_179), .B(n_187), .Y(n_178) );
INVx2_ASAP7_75t_L g203 ( .A(n_163), .Y(n_203) );
INVx2_ASAP7_75t_L g186 ( .A(n_166), .Y(n_186) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
OAI22xp5_ASAP7_75t_SL g168 ( .A1(n_169), .A2(n_170), .B1(n_171), .B2(n_172), .Y(n_168) );
INVx2_ASAP7_75t_L g171 ( .A(n_169), .Y(n_171) );
INVx4_ASAP7_75t_L g237 ( .A(n_169), .Y(n_237) );
INVx2_ASAP7_75t_L g450 ( .A(n_171), .Y(n_450) );
OAI21xp5_ASAP7_75t_L g179 ( .A1(n_174), .A2(n_180), .B(n_181), .Y(n_179) );
OAI21xp5_ASAP7_75t_L g207 ( .A1(n_174), .A2(n_208), .B(n_209), .Y(n_207) );
OAI21xp5_ASAP7_75t_L g445 ( .A1(n_174), .A2(n_446), .B(n_447), .Y(n_445) );
OAI21xp5_ASAP7_75t_L g496 ( .A1(n_174), .A2(n_497), .B(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g244 ( .A(n_177), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_177), .B(n_259), .Y(n_258) );
NOR3xp33_ASAP7_75t_L g318 ( .A(n_177), .B(n_319), .C(n_321), .Y(n_318) );
AND2x2_ASAP7_75t_L g344 ( .A(n_177), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_177), .B(n_351), .Y(n_354) );
AND2x2_ASAP7_75t_L g407 ( .A(n_177), .B(n_408), .Y(n_407) );
INVx3_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx3_ASAP7_75t_L g263 ( .A(n_178), .Y(n_263) );
OR2x2_ASAP7_75t_L g357 ( .A(n_178), .B(n_256), .Y(n_357) );
O2A1O1Ixp33_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_185), .C(n_186), .Y(n_182) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_184), .A2(n_472), .B(n_473), .C(n_474), .Y(n_471) );
OAI22xp33_ASAP7_75t_L g546 ( .A1(n_184), .A2(n_237), .B1(n_547), .B2(n_548), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_189), .B(n_215), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_189), .B(n_229), .Y(n_228) );
AO21x2_ASAP7_75t_L g495 ( .A1(n_189), .A2(n_496), .B(n_502), .Y(n_495) );
OR2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_216), .Y(n_190) );
AOI32xp33_ASAP7_75t_L g308 ( .A1(n_191), .A2(n_309), .A3(n_311), .B1(n_313), .B2(n_316), .Y(n_308) );
NOR2xp67_ASAP7_75t_L g381 ( .A(n_191), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g411 ( .A(n_191), .Y(n_411) );
INVx4_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g343 ( .A(n_192), .B(n_327), .Y(n_343) );
AND2x2_ASAP7_75t_L g363 ( .A(n_192), .B(n_289), .Y(n_363) );
AND2x2_ASAP7_75t_L g431 ( .A(n_192), .B(n_349), .Y(n_431) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_206), .Y(n_192) );
INVx3_ASAP7_75t_L g252 ( .A(n_193), .Y(n_252) );
AND2x2_ASAP7_75t_L g266 ( .A(n_193), .B(n_250), .Y(n_266) );
OR2x2_ASAP7_75t_L g271 ( .A(n_193), .B(n_249), .Y(n_271) );
INVx1_ASAP7_75t_L g278 ( .A(n_193), .Y(n_278) );
AND2x2_ASAP7_75t_L g286 ( .A(n_193), .B(n_260), .Y(n_286) );
AND2x2_ASAP7_75t_L g288 ( .A(n_193), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_193), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g341 ( .A(n_193), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_193), .B(n_426), .Y(n_425) );
OR2x6_ASAP7_75t_L g193 ( .A(n_194), .B(n_204), .Y(n_193) );
AOI21xp5_ASAP7_75t_SL g194 ( .A1(n_195), .A2(n_196), .B(n_203), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_200), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_200), .A2(n_211), .B(n_212), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_L g448 ( .A1(n_200), .A2(n_449), .B(n_450), .C(n_451), .Y(n_448) );
O2A1O1Ixp5_ASAP7_75t_L g499 ( .A1(n_200), .A2(n_450), .B(n_500), .C(n_501), .Y(n_499) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g240 ( .A(n_202), .Y(n_240) );
INVx1_ASAP7_75t_L g213 ( .A(n_203), .Y(n_213) );
INVx2_ASAP7_75t_L g250 ( .A(n_206), .Y(n_250) );
AND2x2_ASAP7_75t_L g296 ( .A(n_206), .B(n_217), .Y(n_296) );
AND2x2_ASAP7_75t_L g306 ( .A(n_206), .B(n_231), .Y(n_306) );
AO21x2_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_213), .B(n_214), .Y(n_206) );
INVx1_ASAP7_75t_L g541 ( .A(n_213), .Y(n_541) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_213), .A2(n_558), .B(n_559), .Y(n_557) );
INVx2_ASAP7_75t_L g426 ( .A(n_216), .Y(n_426) );
OR2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_230), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_217), .B(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g267 ( .A(n_217), .Y(n_267) );
AND2x2_ASAP7_75t_L g311 ( .A(n_217), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g327 ( .A(n_217), .B(n_290), .Y(n_327) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g275 ( .A(n_218), .Y(n_275) );
AND2x2_ASAP7_75t_L g289 ( .A(n_218), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g340 ( .A(n_218), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_218), .B(n_250), .Y(n_372) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_228), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_219), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g550 ( .A(n_219), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_221), .B(n_227), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_226), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_225), .B(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g251 ( .A(n_230), .B(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g312 ( .A(n_230), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_230), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g349 ( .A(n_230), .Y(n_349) );
INVx1_ASAP7_75t_L g382 ( .A(n_230), .Y(n_382) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g260 ( .A(n_231), .B(n_250), .Y(n_260) );
INVx1_ASAP7_75t_L g290 ( .A(n_231), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_237), .B(n_239), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_237), .B(n_490), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_237), .B(n_510), .Y(n_509) );
AOI221xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_247), .B1(n_253), .B2(n_260), .C(n_261), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_244), .B(n_264), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_244), .B(n_327), .Y(n_404) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_246), .B(n_294), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_246), .B(n_255), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_246), .B(n_269), .Y(n_398) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_251), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g320 ( .A(n_250), .Y(n_320) );
AND2x2_ASAP7_75t_L g295 ( .A(n_251), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g373 ( .A(n_251), .Y(n_373) );
AND2x2_ASAP7_75t_L g305 ( .A(n_252), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_252), .B(n_275), .Y(n_321) );
AND2x2_ASAP7_75t_L g385 ( .A(n_252), .B(n_311), .Y(n_385) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_257), .Y(n_254) );
BUFx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g294 ( .A(n_256), .B(n_263), .Y(n_294) );
AND2x2_ASAP7_75t_L g390 ( .A(n_257), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_259), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_260), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_260), .B(n_267), .Y(n_355) );
AND2x2_ASAP7_75t_L g375 ( .A(n_260), .B(n_275), .Y(n_375) );
AND2x2_ASAP7_75t_L g396 ( .A(n_260), .B(n_340), .Y(n_396) );
OAI32xp33_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_265), .A3(n_267), .B1(n_268), .B2(n_271), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx1_ASAP7_75t_SL g269 ( .A(n_263), .Y(n_269) );
NAND2x1_ASAP7_75t_L g310 ( .A(n_263), .B(n_293), .Y(n_310) );
OR2x2_ASAP7_75t_L g314 ( .A(n_263), .B(n_315), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_263), .B(n_362), .Y(n_415) );
INVx1_ASAP7_75t_L g283 ( .A(n_264), .Y(n_283) );
OAI221xp5_ASAP7_75t_SL g401 ( .A1(n_265), .A2(n_356), .B1(n_402), .B2(n_405), .C(n_406), .Y(n_401) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g273 ( .A(n_266), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g316 ( .A(n_266), .B(n_289), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_266), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g394 ( .A(n_266), .B(n_327), .Y(n_394) );
INVxp67_ASAP7_75t_L g330 ( .A(n_267), .Y(n_330) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
AND2x2_ASAP7_75t_L g400 ( .A(n_269), .B(n_387), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_269), .B(n_350), .Y(n_423) );
INVx1_ASAP7_75t_L g298 ( .A(n_271), .Y(n_298) );
NAND2xp5_ASAP7_75t_SL g379 ( .A(n_271), .B(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g416 ( .A(n_271), .B(n_417), .Y(n_416) );
OAI21xp5_ASAP7_75t_SL g272 ( .A1(n_273), .A2(n_276), .B(n_279), .Y(n_272) );
AND2x2_ASAP7_75t_L g285 ( .A(n_274), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g369 ( .A(n_278), .B(n_289), .Y(n_369) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
AND2x2_ASAP7_75t_L g387 ( .A(n_280), .B(n_345), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_280), .B(n_344), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_281), .B(n_293), .Y(n_367) );
OAI211xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_284), .B(n_287), .C(n_297), .Y(n_282) );
AOI221xp5_ASAP7_75t_L g317 ( .A1(n_283), .A2(n_318), .B1(n_322), .B2(n_325), .C(n_328), .Y(n_317) );
AOI31xp33_ASAP7_75t_L g412 ( .A1(n_283), .A2(n_413), .A3(n_414), .B(n_416), .Y(n_412) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_291), .B1(n_293), .B2(n_295), .Y(n_287) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx1_ASAP7_75t_L g413 ( .A(n_293), .Y(n_413) );
INVx1_ASAP7_75t_L g376 ( .A(n_294), .Y(n_376) );
O2A1O1Ixp33_ASAP7_75t_L g419 ( .A1(n_296), .A2(n_420), .B(n_422), .C(n_424), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B1(n_301), .B2(n_305), .Y(n_297) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_302), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OAI221xp5_ASAP7_75t_SL g392 ( .A1(n_304), .A2(n_338), .B1(n_357), .B2(n_393), .C(n_395), .Y(n_392) );
INVx1_ASAP7_75t_L g388 ( .A(n_305), .Y(n_388) );
INVx1_ASAP7_75t_L g342 ( .A(n_306), .Y(n_342) );
NAND3xp33_ASAP7_75t_SL g307 ( .A(n_308), .B(n_317), .C(n_332), .Y(n_307) );
OAI21xp33_ASAP7_75t_L g358 ( .A1(n_309), .A2(n_359), .B(n_363), .Y(n_358) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_311), .B(n_411), .Y(n_410) );
INVxp67_ASAP7_75t_L g418 ( .A(n_312), .Y(n_418) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g356 ( .A(n_319), .B(n_339), .Y(n_356) );
INVx1_ASAP7_75t_L g331 ( .A(n_320), .Y(n_331) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g329 ( .A(n_323), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_323), .B(n_361), .Y(n_360) );
NOR4xp25_ASAP7_75t_L g328 ( .A(n_324), .B(n_329), .C(n_330), .D(n_331), .Y(n_328) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AOI222xp33_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_337), .B1(n_343), .B2(n_344), .C1(n_346), .C2(n_350), .Y(n_332) );
NAND2xp5_ASAP7_75t_SL g333 ( .A(n_334), .B(n_336), .Y(n_333) );
INVx1_ASAP7_75t_L g430 ( .A(n_334), .Y(n_430) );
INVx1_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_342), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_346), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OAI21xp5_ASAP7_75t_SL g406 ( .A1(n_351), .A2(n_407), .B(n_409), .Y(n_406) );
NOR4xp25_ASAP7_75t_L g352 ( .A(n_353), .B(n_364), .C(n_377), .D(n_392), .Y(n_352) );
OAI221xp5_ASAP7_75t_SL g353 ( .A1(n_354), .A2(n_355), .B1(n_356), .B2(n_357), .C(n_358), .Y(n_353) );
INVx1_ASAP7_75t_L g433 ( .A(n_354), .Y(n_433) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_361), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
OAI222xp33_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_368), .B1(n_370), .B2(n_371), .C1(n_374), .C2(n_376), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AOI211xp5_ASAP7_75t_L g399 ( .A1(n_369), .A2(n_400), .B(n_401), .C(n_412), .Y(n_399) );
OR2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
INVx1_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
OAI222xp33_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_383), .B1(n_384), .B2(n_386), .C1(n_388), .C2(n_389), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVxp67_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_394), .A2(n_397), .B1(n_430), .B2(n_431), .Y(n_429) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OAI211xp5_ASAP7_75t_SL g424 ( .A1(n_425), .A2(n_427), .B(n_429), .C(n_432), .Y(n_424) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx3_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_SL g437 ( .A(n_438), .B(n_669), .Y(n_437) );
NOR4xp25_ASAP7_75t_L g438 ( .A(n_439), .B(n_606), .C(n_640), .D(n_656), .Y(n_438) );
NAND4xp25_ASAP7_75t_SL g439 ( .A(n_440), .B(n_536), .C(n_570), .D(n_586), .Y(n_439) );
AOI222xp33_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_479), .B1(n_512), .B2(n_524), .C1(n_529), .C2(n_535), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AOI31xp33_ASAP7_75t_L g702 ( .A1(n_442), .A2(n_703), .A3(n_704), .B(n_706), .Y(n_702) );
OR2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_455), .Y(n_442) );
AND2x2_ASAP7_75t_L g677 ( .A(n_443), .B(n_457), .Y(n_677) );
BUFx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_SL g528 ( .A(n_444), .Y(n_528) );
AND2x2_ASAP7_75t_L g535 ( .A(n_444), .B(n_467), .Y(n_535) );
AND2x2_ASAP7_75t_L g591 ( .A(n_444), .B(n_458), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_455), .B(n_621), .Y(n_620) );
INVx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_456), .B(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_456), .B(n_539), .Y(n_581) );
AND2x2_ASAP7_75t_L g674 ( .A(n_456), .B(n_614), .Y(n_674) );
OAI321xp33_ASAP7_75t_L g708 ( .A1(n_456), .A2(n_528), .A3(n_681), .B1(n_709), .B2(n_711), .C(n_712), .Y(n_708) );
NAND4xp25_ASAP7_75t_L g712 ( .A(n_456), .B(n_515), .C(n_621), .D(n_713), .Y(n_712) );
AND2x4_ASAP7_75t_L g456 ( .A(n_457), .B(n_467), .Y(n_456) );
AND2x2_ASAP7_75t_L g576 ( .A(n_457), .B(n_526), .Y(n_576) );
AND2x2_ASAP7_75t_L g595 ( .A(n_457), .B(n_528), .Y(n_595) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g527 ( .A(n_458), .B(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g551 ( .A(n_458), .B(n_467), .Y(n_551) );
AND2x2_ASAP7_75t_L g637 ( .A(n_458), .B(n_526), .Y(n_637) );
OA21x2_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_460), .B(n_466), .Y(n_458) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_459), .A2(n_485), .B(n_491), .Y(n_484) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_459), .A2(n_505), .B(n_511), .Y(n_504) );
INVx3_ASAP7_75t_SL g526 ( .A(n_467), .Y(n_526) );
AND2x2_ASAP7_75t_L g569 ( .A(n_467), .B(n_556), .Y(n_569) );
OR2x2_ASAP7_75t_L g602 ( .A(n_467), .B(n_528), .Y(n_602) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_467), .Y(n_609) );
AND2x2_ASAP7_75t_L g638 ( .A(n_467), .B(n_527), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_467), .B(n_611), .Y(n_653) );
AND2x2_ASAP7_75t_L g685 ( .A(n_467), .B(n_677), .Y(n_685) );
AND2x2_ASAP7_75t_L g694 ( .A(n_467), .B(n_540), .Y(n_694) );
OR2x6_ASAP7_75t_L g467 ( .A(n_468), .B(n_477), .Y(n_467) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_475), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_492), .Y(n_480) );
INVx1_ASAP7_75t_SL g662 ( .A(n_481), .Y(n_662) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g531 ( .A(n_482), .B(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g514 ( .A(n_483), .B(n_494), .Y(n_514) );
AND2x2_ASAP7_75t_L g598 ( .A(n_483), .B(n_516), .Y(n_598) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g568 ( .A(n_484), .B(n_504), .Y(n_568) );
OR2x2_ASAP7_75t_L g579 ( .A(n_484), .B(n_516), .Y(n_579) );
AND2x2_ASAP7_75t_L g605 ( .A(n_484), .B(n_516), .Y(n_605) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_484), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_492), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_492), .B(n_662), .Y(n_661) );
INVx2_ASAP7_75t_SL g492 ( .A(n_493), .Y(n_492) );
OR2x2_ASAP7_75t_L g578 ( .A(n_493), .B(n_579), .Y(n_578) );
AOI322xp5_ASAP7_75t_L g664 ( .A1(n_493), .A2(n_568), .A3(n_574), .B1(n_605), .B2(n_655), .C1(n_665), .C2(n_667), .Y(n_664) );
OR2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_504), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_494), .B(n_515), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_494), .B(n_516), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_494), .B(n_532), .Y(n_585) );
AND2x2_ASAP7_75t_L g639 ( .A(n_494), .B(n_605), .Y(n_639) );
INVx1_ASAP7_75t_L g643 ( .A(n_494), .Y(n_643) );
AND2x2_ASAP7_75t_L g655 ( .A(n_494), .B(n_504), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_494), .B(n_531), .Y(n_687) );
INVx4_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g552 ( .A(n_495), .B(n_504), .Y(n_552) );
BUFx3_ASAP7_75t_L g566 ( .A(n_495), .Y(n_566) );
AND3x2_ASAP7_75t_L g648 ( .A(n_495), .B(n_628), .C(n_649), .Y(n_648) );
NAND3xp33_ASAP7_75t_L g513 ( .A(n_504), .B(n_514), .C(n_515), .Y(n_513) );
INVx1_ASAP7_75t_SL g532 ( .A(n_504), .Y(n_532) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_504), .Y(n_633) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g627 ( .A(n_514), .B(n_628), .Y(n_627) );
INVxp67_ASAP7_75t_L g634 ( .A(n_514), .Y(n_634) );
AND2x2_ASAP7_75t_L g672 ( .A(n_515), .B(n_650), .Y(n_672) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx3_ASAP7_75t_L g553 ( .A(n_516), .Y(n_553) );
AND2x2_ASAP7_75t_L g628 ( .A(n_516), .B(n_532), .Y(n_628) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
OR2x2_ASAP7_75t_L g572 ( .A(n_526), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g691 ( .A(n_526), .B(n_591), .Y(n_691) );
AND2x2_ASAP7_75t_L g705 ( .A(n_526), .B(n_528), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_527), .B(n_540), .Y(n_646) );
AND2x2_ASAP7_75t_L g693 ( .A(n_527), .B(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g556 ( .A(n_528), .B(n_557), .Y(n_556) );
OR2x2_ASAP7_75t_L g573 ( .A(n_528), .B(n_540), .Y(n_573) );
INVx1_ASAP7_75t_L g583 ( .A(n_528), .Y(n_583) );
AND2x2_ASAP7_75t_L g614 ( .A(n_528), .B(n_540), .Y(n_614) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OAI221xp5_ASAP7_75t_L g656 ( .A1(n_530), .A2(n_657), .B1(n_661), .B2(n_663), .C(n_664), .Y(n_656) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_531), .B(n_533), .Y(n_530) );
AND2x2_ASAP7_75t_L g560 ( .A(n_531), .B(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_534), .B(n_567), .Y(n_710) );
AOI322xp5_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_552), .A3(n_553), .B1(n_554), .B2(n_560), .C1(n_562), .C2(n_569), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_551), .Y(n_538) );
NAND2x1p5_ASAP7_75t_L g590 ( .A(n_539), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_539), .B(n_601), .Y(n_600) );
O2A1O1Ixp33_ASAP7_75t_L g624 ( .A1(n_539), .A2(n_551), .B(n_625), .C(n_626), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_539), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_539), .B(n_595), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_539), .B(n_677), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_539), .B(n_705), .Y(n_704) );
BUFx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_540), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_540), .B(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g666 ( .A(n_540), .B(n_553), .Y(n_666) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B(n_549), .Y(n_540) );
INVx1_ASAP7_75t_L g558 ( .A(n_542), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_549), .Y(n_559) );
INVx1_ASAP7_75t_L g641 ( .A(n_551), .Y(n_641) );
OAI31xp33_ASAP7_75t_L g651 ( .A1(n_551), .A2(n_576), .A3(n_652), .B(n_654), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_551), .B(n_557), .Y(n_703) );
INVx1_ASAP7_75t_SL g564 ( .A(n_552), .Y(n_564) );
AND2x2_ASAP7_75t_L g597 ( .A(n_552), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g678 ( .A(n_552), .B(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g563 ( .A(n_553), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g588 ( .A(n_553), .Y(n_588) );
AND2x2_ASAP7_75t_L g615 ( .A(n_553), .B(n_568), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_553), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g707 ( .A(n_553), .B(n_655), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_555), .B(n_625), .Y(n_698) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g594 ( .A(n_557), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_SL g612 ( .A(n_557), .Y(n_612) );
NAND2xp33_ASAP7_75t_SL g562 ( .A(n_563), .B(n_565), .Y(n_562) );
OAI211xp5_ASAP7_75t_SL g606 ( .A1(n_564), .A2(n_607), .B(n_613), .C(n_629), .Y(n_606) );
OR2x2_ASAP7_75t_L g681 ( .A(n_564), .B(n_662), .Y(n_681) );
OR2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
CKINVDCx16_ASAP7_75t_R g618 ( .A(n_566), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_566), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g587 ( .A(n_568), .B(n_588), .Y(n_587) );
O2A1O1Ixp33_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_574), .B(n_577), .C(n_580), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_SL g621 ( .A(n_573), .Y(n_621) );
INVx1_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_576), .B(n_614), .Y(n_619) );
INVx1_ASAP7_75t_L g625 ( .A(n_576), .Y(n_625) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g584 ( .A(n_579), .B(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g617 ( .A(n_579), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g679 ( .A(n_579), .Y(n_679) );
AOI21xp33_ASAP7_75t_SL g580 ( .A1(n_581), .A2(n_582), .B(n_584), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_582), .A2(n_593), .B(n_596), .Y(n_592) );
AOI211xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_589), .B(n_592), .C(n_599), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_587), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_590), .B(n_681), .Y(n_680) );
INVx2_ASAP7_75t_SL g603 ( .A(n_591), .Y(n_603) );
OAI21xp5_ASAP7_75t_L g658 ( .A1(n_593), .A2(n_659), .B(n_660), .Y(n_658) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_598), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_SL g623 ( .A(n_598), .Y(n_623) );
AOI21xp33_ASAP7_75t_SL g599 ( .A1(n_600), .A2(n_603), .B(n_604), .Y(n_599) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g654 ( .A(n_605), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_611), .B(n_637), .Y(n_663) );
AND2x2_ASAP7_75t_L g676 ( .A(n_611), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g690 ( .A(n_611), .B(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g700 ( .A(n_611), .B(n_638), .Y(n_700) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AOI211xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_615), .B(n_616), .C(n_624), .Y(n_613) );
INVx1_ASAP7_75t_L g660 ( .A(n_614), .Y(n_660) );
OAI22xp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_619), .B1(n_620), .B2(n_622), .Y(n_616) );
OR2x2_ASAP7_75t_L g622 ( .A(n_618), .B(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_618), .B(n_679), .Y(n_701) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g695 ( .A(n_628), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_635), .B1(n_638), .B2(n_639), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .Y(n_631) );
INVx1_ASAP7_75t_L g713 ( .A(n_633), .Y(n_713) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g659 ( .A(n_637), .Y(n_659) );
OAI211xp5_ASAP7_75t_SL g640 ( .A1(n_641), .A2(n_642), .B(n_644), .C(n_651), .Y(n_640) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
INVx2_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
INVxp67_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVxp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_659), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NOR5xp2_ASAP7_75t_L g669 ( .A(n_670), .B(n_688), .C(n_696), .D(n_702), .E(n_708), .Y(n_669) );
OAI211xp5_ASAP7_75t_SL g670 ( .A1(n_671), .A2(n_673), .B(n_675), .C(n_682), .Y(n_670) );
INVxp67_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_678), .B(n_680), .Y(n_675) );
OAI21xp33_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_685), .B(n_686), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_685), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AOI21xp33_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_692), .B(n_695), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_SL g711 ( .A(n_691), .Y(n_711) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AOI21xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_699), .B(n_701), .Y(n_696) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
NAND2xp33_ASAP7_75t_L g723 ( .A(n_724), .B(n_728), .Y(n_723) );
NOR2xp33_ASAP7_75t_SL g724 ( .A(n_725), .B(n_727), .Y(n_724) );
INVx1_ASAP7_75t_SL g743 ( .A(n_725), .Y(n_743) );
INVx1_ASAP7_75t_L g742 ( .A(n_727), .Y(n_742) );
OA21x2_ASAP7_75t_L g745 ( .A1(n_727), .A2(n_743), .B(n_746), .Y(n_745) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g736 ( .A(n_730), .Y(n_736) );
BUFx2_ASAP7_75t_L g746 ( .A(n_730), .Y(n_746) );
OAI21xp5_ASAP7_75t_SL g731 ( .A1(n_732), .A2(n_734), .B(n_737), .Y(n_731) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
CKINVDCx6p67_ASAP7_75t_R g739 ( .A(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_743), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_745), .Y(n_744) );
endmodule