module fake_jpeg_13811_n_639 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_639);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_639;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_378;
wire n_133;
wire n_419;
wire n_132;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_8),
.B(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_14),
.B(n_15),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_0),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_60),
.Y(n_142)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_54),
.B(n_18),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_63),
.B(n_64),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_30),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_67),
.B(n_22),
.Y(n_195)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_68),
.Y(n_155)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_69),
.Y(n_160)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVxp67_ASAP7_75t_SL g206 ( 
.A(n_71),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_72),
.Y(n_146)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_73),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_74),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_75),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g182 ( 
.A(n_76),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_21),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_77),
.B(n_86),
.Y(n_153)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_78),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_80),
.Y(n_188)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_81),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_83),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_85),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_21),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_21),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_87),
.B(n_93),
.Y(n_154)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_89),
.Y(n_176)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_90),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_91),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_44),
.B(n_16),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_94),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_95),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_44),
.B(n_16),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_96),
.B(n_121),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_21),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_97),
.B(n_99),
.Y(n_170)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_98),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_21),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_100),
.Y(n_174)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_101),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_57),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_102),
.B(n_103),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_33),
.B(n_16),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_32),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_104),
.Y(n_211)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_105),
.Y(n_190)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

INVx11_ASAP7_75t_L g158 ( 
.A(n_106),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_28),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_107),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_33),
.B(n_14),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_119),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_57),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_109),
.B(n_115),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

INVx3_ASAP7_75t_SL g152 ( 
.A(n_110),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_111),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_39),
.Y(n_112)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

BUFx8_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_113),
.Y(n_173)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_32),
.Y(n_114)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_114),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_57),
.Y(n_115)
);

BUFx10_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g213 ( 
.A(n_116),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

INVx3_ASAP7_75t_SL g215 ( 
.A(n_117),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_39),
.Y(n_118)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_43),
.B(n_0),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_43),
.Y(n_120)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_120),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_42),
.B(n_27),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_42),
.B(n_13),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_122),
.B(n_13),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_22),
.Y(n_123)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_34),
.Y(n_124)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_124),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_50),
.Y(n_125)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_125),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_39),
.Y(n_126)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_50),
.Y(n_127)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_127),
.Y(n_172)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_22),
.Y(n_128)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_128),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_106),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_129),
.B(n_139),
.Y(n_246)
);

INVx4_ASAP7_75t_SL g130 ( 
.A(n_116),
.Y(n_130)
);

INVx4_ASAP7_75t_SL g280 ( 
.A(n_130),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_67),
.A2(n_49),
.B1(n_37),
.B2(n_55),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_133),
.A2(n_159),
.B1(n_74),
.B2(n_126),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_36),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_137),
.B(n_151),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_116),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_104),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_143),
.B(n_163),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_60),
.A2(n_49),
.B1(n_55),
.B2(n_37),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_148),
.A2(n_26),
.B1(n_22),
.B2(n_117),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_36),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_68),
.A2(n_49),
.B1(n_37),
.B2(n_55),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_88),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_169),
.Y(n_288)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_127),
.Y(n_180)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_125),
.Y(n_183)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_183),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_95),
.B(n_24),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_197),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_95),
.B(n_24),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_186),
.B(n_189),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_107),
.B(n_25),
.Y(n_189)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_90),
.Y(n_194)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_194),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_198),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_107),
.B(n_25),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_94),
.B(n_58),
.Y(n_198)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_98),
.Y(n_201)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_201),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_71),
.Y(n_202)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_202),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_79),
.B(n_23),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_203),
.B(n_207),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_128),
.B(n_23),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_59),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_101),
.B(n_59),
.Y(n_207)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_80),
.Y(n_209)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_209),
.Y(n_256)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_73),
.Y(n_210)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_210),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_66),
.B(n_45),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_51),
.Y(n_227)
);

NOR2x1_ASAP7_75t_R g216 ( 
.A(n_212),
.B(n_69),
.Y(n_216)
);

XNOR2x1_ASAP7_75t_SL g307 ( 
.A(n_216),
.B(n_287),
.Y(n_307)
);

CKINVDCx12_ASAP7_75t_R g217 ( 
.A(n_173),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_217),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_218),
.A2(n_251),
.B1(n_286),
.B2(n_289),
.Y(n_327)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_208),
.Y(n_219)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_219),
.Y(n_311)
);

OAI22x1_ASAP7_75t_L g308 ( 
.A1(n_220),
.A2(n_213),
.B1(n_215),
.B2(n_152),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_211),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_223),
.B(n_272),
.Y(n_300)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_135),
.Y(n_225)
);

INVx3_ASAP7_75t_SL g333 ( 
.A(n_225),
.Y(n_333)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_135),
.Y(n_226)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_226),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_227),
.B(n_253),
.Y(n_294)
);

BUFx12f_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_229),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_230),
.B(n_232),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_153),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_170),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_233),
.B(n_238),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_200),
.Y(n_234)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_234),
.Y(n_312)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_171),
.Y(n_235)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_235),
.Y(n_298)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_142),
.Y(n_237)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_237),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_134),
.B(n_38),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_146),
.Y(n_240)
);

INVx8_ASAP7_75t_L g304 ( 
.A(n_240),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_198),
.A2(n_85),
.B1(n_81),
.B2(n_105),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_241),
.A2(n_264),
.B1(n_291),
.B2(n_206),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_242),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_175),
.B(n_45),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_244),
.B(n_247),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_136),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_245),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_154),
.B(n_47),
.Y(n_247)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_182),
.Y(n_248)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_248),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_146),
.Y(n_249)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_249),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_159),
.A2(n_123),
.B1(n_62),
.B2(n_72),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_181),
.B(n_27),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_150),
.B(n_38),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_254),
.B(n_257),
.Y(n_309)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_208),
.Y(n_255)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_255),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_179),
.B(n_58),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_131),
.B(n_51),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_258),
.B(n_261),
.Y(n_325)
);

BUFx2_ASAP7_75t_R g259 ( 
.A(n_173),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_259),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_144),
.B(n_47),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_145),
.B(n_35),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_262),
.B(n_265),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_187),
.Y(n_263)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_263),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_147),
.A2(n_110),
.B1(n_92),
.B2(n_75),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_162),
.B(n_34),
.Y(n_265)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_187),
.Y(n_266)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_266),
.Y(n_334)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_165),
.Y(n_268)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_268),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_168),
.B(n_56),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_269),
.B(n_270),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_174),
.B(n_204),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_193),
.B(n_56),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_271),
.B(n_276),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_195),
.B(n_118),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_211),
.Y(n_273)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_273),
.Y(n_292)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_169),
.Y(n_274)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_274),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_136),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_275),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_172),
.B(n_35),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_141),
.B(n_13),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_277),
.B(n_166),
.Y(n_335)
);

BUFx5_ASAP7_75t_L g278 ( 
.A(n_158),
.Y(n_278)
);

BUFx4f_ASAP7_75t_SL g338 ( 
.A(n_278),
.Y(n_338)
);

CKINVDCx12_ASAP7_75t_R g279 ( 
.A(n_130),
.Y(n_279)
);

BUFx8_ASAP7_75t_L g318 ( 
.A(n_279),
.Y(n_318)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_156),
.Y(n_281)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_281),
.Y(n_299)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_149),
.Y(n_282)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_282),
.Y(n_303)
);

INVx5_ASAP7_75t_L g283 ( 
.A(n_182),
.Y(n_283)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_149),
.Y(n_284)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_284),
.Y(n_313)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_156),
.Y(n_285)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_285),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_133),
.A2(n_112),
.B1(n_26),
.B2(n_111),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_141),
.B(n_113),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_188),
.A2(n_26),
.B1(n_91),
.B2(n_89),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_188),
.Y(n_290)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_290),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_152),
.A2(n_26),
.B1(n_84),
.B2(n_76),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_221),
.B(n_140),
.C(n_160),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_295),
.B(n_310),
.Y(n_355)
);

OAI21xp33_ASAP7_75t_L g296 ( 
.A1(n_221),
.A2(n_206),
.B(n_158),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_296),
.A2(n_341),
.B(n_336),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_286),
.A2(n_251),
.B1(n_216),
.B2(n_264),
.Y(n_302)
);

OA22x2_ASAP7_75t_L g384 ( 
.A1(n_302),
.A2(n_210),
.B1(n_177),
.B2(n_313),
.Y(n_384)
);

OAI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_276),
.A2(n_192),
.B1(n_155),
.B2(n_178),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_305),
.A2(n_320),
.B1(n_342),
.B2(n_349),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_308),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_228),
.B(n_252),
.C(n_272),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_288),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_321),
.B(n_231),
.Y(n_351)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_246),
.Y(n_323)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_323),
.Y(n_357)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_256),
.Y(n_326)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_326),
.Y(n_383)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_236),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_328),
.Y(n_353)
);

NAND3xp33_ASAP7_75t_L g369 ( 
.A(n_335),
.B(n_259),
.C(n_280),
.Y(n_369)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_237),
.Y(n_337)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_337),
.Y(n_362)
);

OAI22xp33_ASAP7_75t_L g342 ( 
.A1(n_220),
.A2(n_157),
.B1(n_164),
.B2(n_190),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_268),
.Y(n_343)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_343),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_267),
.A2(n_178),
.B(n_155),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_345),
.A2(n_223),
.B(n_275),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_224),
.B(n_196),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_348),
.B(n_245),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_241),
.A2(n_215),
.B1(n_157),
.B2(n_192),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_351),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_329),
.B(n_222),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_354),
.B(n_359),
.Y(n_407)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_344),
.Y(n_356)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_356),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_332),
.B(n_250),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_310),
.B(n_243),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_360),
.Y(n_403)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_344),
.Y(n_361)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_361),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_340),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_363),
.B(n_365),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_327),
.A2(n_308),
.B1(n_300),
.B2(n_342),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_SL g412 ( 
.A1(n_364),
.A2(n_381),
.B1(n_394),
.B2(n_333),
.Y(n_412)
);

AOI32xp33_ASAP7_75t_L g365 ( 
.A1(n_345),
.A2(n_166),
.A3(n_202),
.B1(n_229),
.B2(n_182),
.Y(n_365)
);

INVx13_ASAP7_75t_L g366 ( 
.A(n_318),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_366),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_295),
.B(n_239),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_367),
.B(n_368),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_347),
.B(n_239),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_369),
.B(n_370),
.Y(n_433)
);

NAND3xp33_ASAP7_75t_L g370 ( 
.A(n_322),
.B(n_280),
.C(n_287),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_316),
.B(n_235),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_371),
.B(n_376),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_372),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_325),
.B(n_260),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_373),
.B(n_380),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_327),
.A2(n_307),
.B1(n_296),
.B2(n_300),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_374),
.A2(n_213),
.B1(n_167),
.B2(n_161),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_300),
.Y(n_375)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_375),
.Y(n_414)
);

FAx1_ASAP7_75t_SL g376 ( 
.A(n_307),
.B(n_283),
.CI(n_248),
.CON(n_376),
.SN(n_376)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_377),
.B(n_385),
.Y(n_410)
);

INVx13_ASAP7_75t_L g378 ( 
.A(n_318),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_378),
.Y(n_398)
);

OAI22x1_ASAP7_75t_SL g379 ( 
.A1(n_333),
.A2(n_138),
.B1(n_184),
.B2(n_176),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_379),
.A2(n_358),
.B1(n_375),
.B2(n_138),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_330),
.B(n_255),
.Y(n_380)
);

INVx3_ASAP7_75t_SL g381 ( 
.A(n_304),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_301),
.Y(n_382)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_382),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_384),
.A2(n_379),
.B1(n_352),
.B2(n_177),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_309),
.B(n_285),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_318),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_387),
.B(n_392),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_297),
.A2(n_219),
.B(n_234),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_388),
.A2(n_391),
.B(n_336),
.Y(n_418)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_350),
.Y(n_389)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_389),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_304),
.Y(n_390)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_390),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_294),
.B(n_281),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_292),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_393),
.Y(n_400)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_311),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_303),
.B(n_284),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_395),
.B(n_396),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_317),
.B(n_282),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_391),
.A2(n_306),
.B(n_341),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_397),
.A2(n_402),
.B(n_418),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_372),
.A2(n_374),
.B(n_358),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_355),
.B(n_315),
.C(n_299),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_404),
.B(n_406),
.C(n_380),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_355),
.B(n_314),
.C(n_350),
.Y(n_406)
);

NOR2xp67_ASAP7_75t_SL g409 ( 
.A(n_376),
.B(n_338),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_409),
.A2(n_413),
.B(n_419),
.Y(n_459)
);

XNOR2x1_ASAP7_75t_L g411 ( 
.A(n_367),
.B(n_338),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_411),
.B(n_429),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_412),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_384),
.A2(n_319),
.B1(n_334),
.B2(n_301),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_415),
.A2(n_423),
.B1(n_362),
.B2(n_389),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_376),
.A2(n_312),
.B(n_339),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_422),
.A2(n_378),
.B(n_366),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_384),
.A2(n_334),
.B1(n_346),
.B2(n_331),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_424),
.A2(n_176),
.B1(n_184),
.B2(n_166),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_396),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_428),
.B(n_373),
.Y(n_437)
);

XOR2x2_ASAP7_75t_L g429 ( 
.A(n_368),
.B(n_338),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_352),
.A2(n_290),
.B1(n_226),
.B2(n_266),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_432),
.A2(n_434),
.B1(n_381),
.B2(n_388),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_384),
.A2(n_331),
.B1(n_240),
.B2(n_249),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_436),
.B(n_461),
.C(n_467),
.Y(n_489)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_437),
.Y(n_498)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_438),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_425),
.B(n_395),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_439),
.B(n_445),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_434),
.A2(n_353),
.B1(n_382),
.B2(n_390),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_441),
.A2(n_463),
.B1(n_468),
.B2(n_423),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_430),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_442),
.B(n_451),
.Y(n_473)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_430),
.Y(n_444)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_444),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_400),
.B(n_353),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_400),
.B(n_357),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_446),
.B(n_447),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_407),
.B(n_383),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_428),
.B(n_386),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_448),
.B(n_449),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_421),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_435),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_450),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_407),
.B(n_356),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_421),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_452),
.B(n_453),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_398),
.B(n_386),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_454),
.B(n_455),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_398),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_420),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_456),
.B(n_457),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_410),
.B(n_362),
.Y(n_457)
);

CKINVDCx12_ASAP7_75t_R g458 ( 
.A(n_420),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_458),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_419),
.A2(n_346),
.B1(n_361),
.B2(n_225),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_460),
.B(n_462),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_404),
.B(n_324),
.C(n_312),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_410),
.B(n_394),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_408),
.B(n_324),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_464),
.B(n_465),
.Y(n_502)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_435),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_466),
.A2(n_416),
.B(n_414),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_406),
.B(n_339),
.C(n_317),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_426),
.A2(n_263),
.B1(n_311),
.B2(n_298),
.Y(n_468)
);

OAI21xp33_ASAP7_75t_SL g470 ( 
.A1(n_402),
.A2(n_191),
.B(n_298),
.Y(n_470)
);

OAI21xp33_ASAP7_75t_L g493 ( 
.A1(n_470),
.A2(n_414),
.B(n_413),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_445),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_471),
.B(n_480),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_449),
.B(n_427),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_474),
.B(n_491),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_443),
.A2(n_409),
.B(n_422),
.Y(n_476)
);

NAND2xp33_ASAP7_75t_SL g525 ( 
.A(n_476),
.B(n_484),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_436),
.B(n_408),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_478),
.B(n_490),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_479),
.A2(n_493),
.B1(n_424),
.B2(n_459),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_446),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_453),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_482),
.B(n_485),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_443),
.A2(n_397),
.B(n_418),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_483),
.B(n_488),
.Y(n_527)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_451),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_459),
.A2(n_405),
.B(n_416),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_440),
.B(n_411),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_452),
.B(n_405),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_447),
.B(n_403),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_492),
.B(n_494),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_448),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_467),
.B(n_429),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_499),
.B(n_468),
.Y(n_529)
);

CKINVDCx16_ASAP7_75t_R g503 ( 
.A(n_462),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_503),
.B(n_458),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_489),
.B(n_461),
.C(n_440),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_505),
.B(n_515),
.C(n_524),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_478),
.B(n_429),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_506),
.B(n_507),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_489),
.B(n_444),
.Y(n_507)
);

OA21x2_ASAP7_75t_L g508 ( 
.A1(n_500),
.A2(n_438),
.B(n_415),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_508),
.B(n_486),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_500),
.A2(n_442),
.B1(n_469),
.B2(n_441),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_510),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_475),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_511),
.B(n_521),
.Y(n_541)
);

BUFx10_ASAP7_75t_L g512 ( 
.A(n_477),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_512),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_499),
.B(n_490),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_513),
.B(n_481),
.Y(n_534)
);

NOR2x1_ASAP7_75t_L g514 ( 
.A(n_475),
.B(n_425),
.Y(n_514)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_514),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_501),
.B(n_488),
.C(n_483),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_495),
.Y(n_516)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_516),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_498),
.A2(n_433),
.B1(n_437),
.B2(n_457),
.Y(n_517)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_517),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_496),
.A2(n_460),
.B1(n_454),
.B2(n_432),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_519),
.A2(n_523),
.B1(n_533),
.B2(n_471),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_520),
.A2(n_482),
.B1(n_481),
.B2(n_495),
.Y(n_545)
);

NOR3xp33_ASAP7_75t_SL g521 ( 
.A(n_498),
.B(n_433),
.C(n_439),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_496),
.A2(n_455),
.B1(n_450),
.B2(n_465),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_501),
.B(n_464),
.C(n_466),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_473),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_526),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_SL g538 ( 
.A(n_529),
.B(n_486),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_484),
.B(n_417),
.C(n_401),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_530),
.B(n_529),
.C(n_524),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_480),
.A2(n_463),
.B1(n_456),
.B2(n_431),
.Y(n_531)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_531),
.Y(n_552)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_532),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_479),
.A2(n_431),
.B1(n_417),
.B2(n_401),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_534),
.B(n_538),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_537),
.A2(n_543),
.B1(n_545),
.B2(n_508),
.Y(n_568)
);

BUFx12f_ASAP7_75t_SL g539 ( 
.A(n_521),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_539),
.B(n_527),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_SL g563 ( 
.A1(n_540),
.A2(n_516),
.B1(n_518),
.B2(n_508),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_542),
.B(n_553),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_519),
.A2(n_494),
.B1(n_503),
.B2(n_476),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_505),
.B(n_477),
.C(n_502),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_549),
.B(n_550),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_507),
.B(n_504),
.C(n_513),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_504),
.B(n_502),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_506),
.B(n_399),
.C(n_487),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_554),
.B(n_555),
.C(n_512),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_515),
.B(n_399),
.C(n_487),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_522),
.B(n_523),
.Y(n_556)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_556),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_560),
.B(n_574),
.Y(n_592)
);

CKINVDCx14_ASAP7_75t_R g561 ( 
.A(n_541),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_561),
.B(n_562),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_558),
.A2(n_509),
.B1(n_528),
.B2(n_533),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_563),
.A2(n_568),
.B1(n_556),
.B2(n_555),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g566 ( 
.A(n_557),
.Y(n_566)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_566),
.Y(n_583)
);

INVx13_ASAP7_75t_L g567 ( 
.A(n_546),
.Y(n_567)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_567),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_569),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_536),
.B(n_530),
.C(n_525),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_570),
.B(n_573),
.Y(n_591)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_548),
.Y(n_572)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_572),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_549),
.B(n_497),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_536),
.B(n_512),
.C(n_487),
.Y(n_574)
);

NOR3xp33_ASAP7_75t_SL g575 ( 
.A(n_539),
.B(n_497),
.C(n_514),
.Y(n_575)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_575),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_SL g576 ( 
.A1(n_551),
.A2(n_472),
.B1(n_293),
.B2(n_242),
.Y(n_576)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_576),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_534),
.B(n_472),
.Y(n_577)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_577),
.B(n_542),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_SL g578 ( 
.A1(n_535),
.A2(n_552),
.B1(n_544),
.B2(n_540),
.Y(n_578)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_578),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_L g579 ( 
.A1(n_543),
.A2(n_293),
.B(n_132),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_579),
.B(n_537),
.Y(n_580)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_580),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_SL g609 ( 
.A(n_581),
.B(n_596),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_SL g601 ( 
.A1(n_582),
.A2(n_594),
.B1(n_580),
.B2(n_595),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_574),
.B(n_554),
.Y(n_585)
);

OAI21x1_ASAP7_75t_L g600 ( 
.A1(n_585),
.A2(n_564),
.B(n_560),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_SL g586 ( 
.A1(n_578),
.A2(n_538),
.B1(n_553),
.B2(n_547),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_586),
.A2(n_570),
.B1(n_565),
.B2(n_571),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_568),
.A2(n_550),
.B1(n_547),
.B2(n_199),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_593),
.B(n_567),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_L g596 ( 
.A(n_571),
.B(n_229),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_582),
.A2(n_559),
.B1(n_576),
.B2(n_566),
.Y(n_597)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_597),
.Y(n_615)
);

XOR2xp5_ASAP7_75t_L g612 ( 
.A(n_598),
.B(n_601),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_590),
.A2(n_579),
.B(n_575),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_599),
.A2(n_600),
.B(n_608),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_SL g602 ( 
.A(n_588),
.B(n_564),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_SL g620 ( 
.A(n_602),
.B(n_596),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_591),
.B(n_577),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_603),
.B(n_604),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_592),
.B(n_278),
.C(n_132),
.Y(n_605)
);

NOR2xp67_ASAP7_75t_SL g613 ( 
.A(n_605),
.B(n_585),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_587),
.B(n_214),
.Y(n_606)
);

CKINVDCx16_ASAP7_75t_R g614 ( 
.A(n_606),
.Y(n_614)
);

OAI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_584),
.A2(n_113),
.B(n_111),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_581),
.B(n_0),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_610),
.B(n_583),
.Y(n_616)
);

AOI21x1_ASAP7_75t_L g628 ( 
.A1(n_613),
.A2(n_1),
.B(n_2),
.Y(n_628)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_616),
.B(n_618),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g618 ( 
.A(n_605),
.B(n_592),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_609),
.B(n_586),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_619),
.A2(n_621),
.B(n_607),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_SL g626 ( 
.A1(n_620),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_SL g621 ( 
.A(n_599),
.B(n_589),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_622),
.B(n_626),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_611),
.A2(n_601),
.B(n_597),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_L g632 ( 
.A1(n_624),
.A2(n_625),
.B(n_627),
.Y(n_632)
);

AOI21xp33_ASAP7_75t_L g625 ( 
.A1(n_617),
.A2(n_609),
.B(n_2),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_612),
.A2(n_11),
.B(n_2),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_628),
.B(n_1),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_630),
.B(n_631),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_623),
.B(n_614),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_629),
.B(n_612),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_634),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_635),
.A2(n_615),
.B1(n_633),
.B2(n_632),
.Y(n_636)
);

OAI21xp5_ASAP7_75t_SL g637 ( 
.A1(n_636),
.A2(n_616),
.B(n_7),
.Y(n_637)
);

AOI322xp5_ASAP7_75t_L g638 ( 
.A1(n_637),
.A2(n_4),
.A3(n_7),
.B1(n_8),
.B2(n_10),
.C1(n_400),
.C2(n_567),
.Y(n_638)
);

XOR2xp5_ASAP7_75t_L g639 ( 
.A(n_638),
.B(n_8),
.Y(n_639)
);


endmodule