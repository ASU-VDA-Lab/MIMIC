module fake_jpeg_5208_n_280 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_280);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_280;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_11),
.B(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_38),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_20),
.B(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_40),
.B(n_33),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_0),
.C(n_1),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_0),
.Y(n_50)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_51),
.Y(n_60)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_31),
.B1(n_18),
.B2(n_27),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_44),
.A2(n_22),
.B1(n_33),
.B2(n_30),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_45),
.B(n_53),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_31),
.B1(n_21),
.B2(n_27),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_49),
.B1(n_37),
.B2(n_35),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_34),
.A2(n_27),
.B1(n_31),
.B2(n_24),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_39),
.B(n_20),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_30),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_55),
.Y(n_59)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_38),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_54),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_61),
.B(n_63),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_62),
.B(n_65),
.Y(n_109)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_79),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_43),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_66),
.A2(n_69),
.B1(n_91),
.B2(n_48),
.Y(n_112)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_68),
.B(n_71),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_55),
.A2(n_35),
.B1(n_36),
.B2(n_40),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_54),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_70),
.Y(n_95)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_38),
.B1(n_36),
.B2(n_28),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_72),
.A2(n_74),
.B1(n_85),
.B2(n_48),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_50),
.A2(n_38),
.B1(n_16),
.B2(n_28),
.Y(n_74)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_29),
.Y(n_76)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_77),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_78),
.Y(n_93)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_52),
.B(n_17),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_83),
.Y(n_96)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_46),
.A2(n_21),
.B1(n_17),
.B2(n_30),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_86),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_46),
.A2(n_33),
.B1(n_19),
.B2(n_22),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_42),
.Y(n_88)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_40),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_23),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_44),
.A2(n_19),
.B1(n_22),
.B2(n_23),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_59),
.A2(n_51),
.B(n_49),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_91),
.C(n_81),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_112),
.B1(n_115),
.B2(n_64),
.Y(n_121)
);

FAx1_ASAP7_75t_SL g149 ( 
.A(n_102),
.B(n_116),
.CI(n_16),
.CON(n_149),
.SN(n_149)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_51),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_97),
.Y(n_142)
);

FAx1_ASAP7_75t_SL g110 ( 
.A(n_69),
.B(n_38),
.CI(n_29),
.CON(n_110),
.SN(n_110)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_110),
.B(n_68),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_59),
.A2(n_48),
.B1(n_46),
.B2(n_19),
.Y(n_115)
);

AOI32xp33_ASAP7_75t_L g116 ( 
.A1(n_62),
.A2(n_48),
.A3(n_46),
.B1(n_29),
.B2(n_28),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_67),
.A2(n_26),
.B(n_23),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_79),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_113),
.B1(n_116),
.B2(n_120),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_105),
.A2(n_82),
.B1(n_70),
.B2(n_89),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_122),
.Y(n_168)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_126),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_97),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_84),
.Y(n_125)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_106),
.A2(n_67),
.B1(n_66),
.B2(n_72),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_127),
.A2(n_131),
.B1(n_145),
.B2(n_147),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_77),
.Y(n_128)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_96),
.B(n_65),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_143),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_90),
.Y(n_130)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_93),
.A2(n_74),
.B1(n_81),
.B2(n_71),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_111),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_132),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_133),
.A2(n_141),
.B(n_16),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_60),
.C(n_80),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_107),
.C(n_32),
.Y(n_177)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_136),
.Y(n_175)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_88),
.Y(n_137)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_137),
.Y(n_176)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_93),
.B1(n_97),
.B2(n_98),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_139),
.A2(n_133),
.B1(n_149),
.B2(n_134),
.Y(n_173)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_102),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_88),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_105),
.A2(n_63),
.B1(n_86),
.B2(n_92),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_32),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_148),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_94),
.A2(n_73),
.B1(n_28),
.B2(n_16),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_114),
.B(n_10),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_32),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_150),
.A2(n_165),
.B1(n_169),
.B2(n_173),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_156),
.Y(n_184)
);

AND2x6_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_95),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_0),
.Y(n_191)
);

AND2x6_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_95),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_163),
.Y(n_195)
);

OR2x2_ASAP7_75t_SL g161 ( 
.A(n_124),
.B(n_96),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_161),
.A2(n_178),
.B(n_32),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_127),
.A2(n_110),
.B1(n_99),
.B2(n_103),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_162),
.A2(n_149),
.B1(n_131),
.B2(n_135),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_110),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_121),
.A2(n_99),
.B1(n_101),
.B2(n_108),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_139),
.A2(n_108),
.B1(n_107),
.B2(n_119),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_170),
.B(n_1),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_147),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_144),
.C(n_32),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_179),
.B(n_180),
.Y(n_209)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_175),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_181),
.B(n_191),
.Y(n_207)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_185),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_156),
.A2(n_140),
.B1(n_136),
.B2(n_132),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_183),
.A2(n_200),
.B1(n_157),
.B2(n_163),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_32),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_194),
.C(n_197),
.Y(n_214)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_189),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_10),
.Y(n_188)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_190),
.A2(n_193),
.B(n_167),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_25),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_168),
.A2(n_25),
.B1(n_2),
.B2(n_3),
.Y(n_196)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_25),
.C(n_2),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_25),
.C(n_2),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_202),
.C(n_160),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_25),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_171),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_159),
.A2(n_170),
.B1(n_157),
.B2(n_168),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_151),
.B(n_25),
.Y(n_201)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_201),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_1),
.C(n_5),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_183),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_208),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_211),
.A2(n_219),
.B1(n_192),
.B2(n_195),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_217),
.Y(n_222)
);

OA21x2_ASAP7_75t_L g215 ( 
.A1(n_191),
.A2(n_171),
.B(n_161),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_215),
.A2(n_221),
.B(n_198),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_196),
.Y(n_217)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_218),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_192),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_155),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_195),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_190),
.A2(n_164),
.B(n_154),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_194),
.C(n_201),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_225),
.C(n_234),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_220),
.C(n_206),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_226),
.A2(n_233),
.B1(n_204),
.B2(n_217),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_235),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_228),
.A2(n_232),
.B1(n_204),
.B2(n_215),
.Y(n_246)
);

XNOR2x1_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_184),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_231),
.B(n_207),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_212),
.A2(n_181),
.B1(n_197),
.B2(n_202),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_212),
.A2(n_154),
.B1(n_172),
.B2(n_7),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_5),
.C(n_6),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_6),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_7),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_216),
.C(n_209),
.Y(n_249)
);

MAJx2_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_237),
.C(n_215),
.Y(n_257)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_245),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_203),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_242),
.A2(n_218),
.B(n_205),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_205),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_246),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_244),
.Y(n_256)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_222),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_235),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_247),
.B(n_248),
.Y(n_251)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_234),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_249),
.A2(n_228),
.B(n_225),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_249),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_243),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_257),
.C(n_240),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_254),
.A2(n_255),
.B1(n_258),
.B2(n_232),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_238),
.A2(n_223),
.B1(n_231),
.B2(n_229),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_241),
.A2(n_229),
.B(n_230),
.Y(n_258)
);

BUFx24_ASAP7_75t_SL g260 ( 
.A(n_252),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_260),
.B(n_264),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_262),
.C(n_263),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_203),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_256),
.A2(n_241),
.B1(n_224),
.B2(n_213),
.Y(n_265)
);

AOI322xp5_ASAP7_75t_L g270 ( 
.A1(n_265),
.A2(n_255),
.A3(n_9),
.B1(n_11),
.B2(n_12),
.C1(n_7),
.C2(n_14),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_240),
.C(n_9),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_257),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g267 ( 
.A(n_266),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_267),
.A2(n_269),
.B(n_13),
.Y(n_272)
);

NOR2xp67_ASAP7_75t_SL g274 ( 
.A(n_270),
.B(n_14),
.Y(n_274)
);

NOR3xp33_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_273),
.C(n_274),
.Y(n_276)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_271),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_272),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_268),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_277),
.Y(n_278)
);

AO21x1_ASAP7_75t_L g279 ( 
.A1(n_278),
.A2(n_276),
.B(n_15),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_15),
.Y(n_280)
);


endmodule