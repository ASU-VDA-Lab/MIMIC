module fake_jpeg_19688_n_73 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_73);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_73;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_71;
wire n_52;
wire n_68;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_9),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_2),
.Y(n_11)
);

INVx6_ASAP7_75t_SL g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_26),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_1),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_25),
.Y(n_30)
);

BUFx2_ASAP7_75t_SL g23 ( 
.A(n_19),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_23),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_1),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_4),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_10),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_22),
.A2(n_11),
.B(n_19),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_28),
.A2(n_19),
.B(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_21),
.A2(n_13),
.B(n_17),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_13),
.C(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_18),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_36),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_20),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_29),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_24),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_32),
.B1(n_31),
.B2(n_35),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_44),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_31),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_24),
.C(n_14),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_12),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_41),
.B1(n_43),
.B2(n_42),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_12),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_58),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_47),
.C(n_39),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_38),
.B1(n_3),
.B2(n_6),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_59),
.B(n_56),
.Y(n_62)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_62),
.B(n_64),
.Y(n_66)
);

AO221x1_ASAP7_75t_L g64 ( 
.A1(n_60),
.A2(n_51),
.B1(n_53),
.B2(n_3),
.C(n_49),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_61),
.A2(n_48),
.B(n_62),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_67),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_58),
.C(n_50),
.Y(n_67)
);

FAx1_ASAP7_75t_SL g69 ( 
.A(n_66),
.B(n_52),
.CI(n_63),
.CON(n_69),
.SN(n_69)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_4),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_71),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_7),
.B(n_68),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_68),
.C(n_7),
.Y(n_73)
);


endmodule