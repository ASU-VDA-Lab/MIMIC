module fake_jpeg_5824_n_216 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_216);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

AND2x6_ASAP7_75t_L g25 ( 
.A(n_3),
.B(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_11),
.B(n_9),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_35),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_36),
.B(n_48),
.Y(n_79)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_7),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_38),
.B(n_51),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_18),
.Y(n_39)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_43),
.Y(n_57)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_45),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_25),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_47),
.Y(n_73)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_26),
.B(n_0),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_30),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_32),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_52),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_16),
.B(n_7),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_0),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_19),
.B(n_8),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_54),
.B(n_33),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_17),
.A2(n_1),
.B(n_2),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_21),
.C(n_20),
.Y(n_81)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_28),
.Y(n_63)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_30),
.B1(n_17),
.B2(n_34),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_59),
.A2(n_62),
.B1(n_66),
.B2(n_55),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_29),
.B1(n_31),
.B2(n_16),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_63),
.B(n_78),
.Y(n_109)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_67),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_29),
.B1(n_27),
.B2(n_24),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_68),
.A2(n_75),
.B1(n_82),
.B2(n_15),
.Y(n_108)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_71),
.Y(n_101)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_35),
.B(n_24),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_83),
.Y(n_118)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_36),
.B(n_28),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_89),
.B(n_54),
.Y(n_100)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_21),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_84),
.B(n_91),
.Y(n_115)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_45),
.A2(n_29),
.B1(n_27),
.B2(n_20),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_90),
.B(n_8),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_56),
.B(n_52),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_88),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_73),
.A2(n_49),
.B1(n_44),
.B2(n_40),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_94),
.A2(n_102),
.B1(n_64),
.B2(n_61),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_50),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_99),
.Y(n_123)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_103),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_15),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_100),
.B(n_70),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_44),
.B1(n_43),
.B2(n_30),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_57),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_110),
.Y(n_121)
);

AND2x6_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_15),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_116),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_60),
.B(n_15),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_80),
.Y(n_124)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g110 ( 
.A(n_72),
.Y(n_110)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

OAI22x1_ASAP7_75t_L g112 ( 
.A1(n_59),
.A2(n_62),
.B1(n_66),
.B2(n_69),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_116),
.C(n_118),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_117),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_59),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_129),
.B1(n_100),
.B2(n_111),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_127),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_75),
.B(n_68),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_126),
.A2(n_134),
.B(n_114),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_80),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_74),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_128),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_137),
.B1(n_97),
.B2(n_93),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_88),
.Y(n_131)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_115),
.Y(n_132)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_76),
.C(n_86),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_86),
.C(n_96),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_102),
.A2(n_82),
.B(n_61),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_138),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_98),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_83),
.Y(n_139)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_2),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_127),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_141),
.A2(n_112),
.B1(n_94),
.B2(n_92),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_150),
.B1(n_153),
.B2(n_158),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_135),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_147),
.Y(n_171)
);

NAND4xp25_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_156),
.C(n_130),
.D(n_131),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_109),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_123),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_141),
.A2(n_97),
.B1(n_109),
.B2(n_105),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_160),
.C(n_133),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_119),
.A2(n_93),
.B1(n_5),
.B2(n_7),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_155),
.A2(n_128),
.B1(n_157),
.B2(n_132),
.Y(n_168)
);

NOR4xp25_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_4),
.C(n_5),
.D(n_8),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_121),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_159),
.B(n_121),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_114),
.C(n_104),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_166),
.C(n_142),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_146),
.A2(n_126),
.B1(n_119),
.B2(n_137),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_163),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_143),
.Y(n_164)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_165),
.A2(n_168),
.B(n_151),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_141),
.Y(n_167)
);

AOI321xp33_ASAP7_75t_L g189 ( 
.A1(n_167),
.A2(n_173),
.A3(n_151),
.B1(n_152),
.B2(n_147),
.C(n_125),
.Y(n_189)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_140),
.Y(n_173)
);

O2A1O1Ixp33_ASAP7_75t_SL g175 ( 
.A1(n_144),
.A2(n_159),
.B(n_129),
.C(n_122),
.Y(n_175)
);

AO22x1_ASAP7_75t_SL g176 ( 
.A1(n_158),
.A2(n_122),
.B1(n_134),
.B2(n_129),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_142),
.A2(n_122),
.B1(n_139),
.B2(n_123),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_174),
.Y(n_178)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_154),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_181),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_180),
.A2(n_152),
.B1(n_176),
.B2(n_171),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_150),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_182),
.B(n_183),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_160),
.C(n_125),
.Y(n_183)
);

NOR3xp33_ASAP7_75t_SL g186 ( 
.A(n_176),
.B(n_165),
.C(n_156),
.Y(n_186)
);

AOI322xp5_ASAP7_75t_L g192 ( 
.A1(n_186),
.A2(n_167),
.A3(n_177),
.B1(n_163),
.B2(n_176),
.C1(n_171),
.C2(n_170),
.Y(n_192)
);

AOI321xp33_ASAP7_75t_L g195 ( 
.A1(n_189),
.A2(n_173),
.A3(n_168),
.B1(n_175),
.B2(n_155),
.C(n_120),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_193),
.B1(n_188),
.B2(n_189),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_195),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_178),
.A2(n_172),
.B1(n_175),
.B2(n_167),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_187),
.A2(n_120),
.B1(n_145),
.B2(n_169),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_196),
.A2(n_184),
.B1(n_183),
.B2(n_136),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_196),
.B(n_185),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_199),
.A2(n_203),
.B(n_195),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_200),
.A2(n_182),
.B1(n_181),
.B2(n_190),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_202),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_197),
.A2(n_184),
.B(n_186),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_145),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_204),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_148),
.C(n_104),
.Y(n_211)
);

MAJx2_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_190),
.C(n_194),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_206),
.A2(n_207),
.B(n_11),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_198),
.A2(n_179),
.B(n_194),
.Y(n_207)
);

AOI322xp5_ASAP7_75t_L g209 ( 
.A1(n_208),
.A2(n_202),
.A3(n_200),
.B1(n_148),
.B2(n_114),
.C1(n_14),
.C2(n_9),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_211),
.Y(n_213)
);

AOI31xp33_ASAP7_75t_L g214 ( 
.A1(n_212),
.A2(n_210),
.A3(n_12),
.B(n_13),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_12),
.C(n_13),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_213),
.Y(n_216)
);


endmodule