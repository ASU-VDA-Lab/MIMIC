module real_aes_5888_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_93;
wire n_182;
wire n_449;
wire n_417;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_87;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
HB1xp67_ASAP7_75t_L g195 ( .A(n_0), .Y(n_195) );
INVx1_ASAP7_75t_L g411 ( .A(n_0), .Y(n_411) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_1), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g158 ( .A1(n_2), .A2(n_68), .B1(n_159), .B2(n_162), .Y(n_158) );
AOI22xp33_ASAP7_75t_L g143 ( .A1(n_3), .A2(n_22), .B1(n_144), .B2(n_146), .Y(n_143) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_4), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_5), .B(n_277), .Y(n_361) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_5), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g362 ( .A(n_6), .B(n_363), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_7), .A2(n_35), .B1(n_276), .B2(n_328), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g87 ( .A1(n_8), .A2(n_20), .B1(n_88), .B2(n_113), .Y(n_87) );
AOI22xp5_ASAP7_75t_L g239 ( .A1(n_9), .A2(n_37), .B1(n_240), .B2(n_244), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_10), .A2(n_51), .B1(n_254), .B2(n_376), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_11), .B(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g406 ( .A(n_12), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g151 ( .A1(n_13), .A2(n_76), .B1(n_152), .B2(n_156), .Y(n_151) );
AOI22xp33_ASAP7_75t_L g131 ( .A1(n_14), .A2(n_57), .B1(n_132), .B2(n_136), .Y(n_131) );
INVx1_ASAP7_75t_L g110 ( .A(n_15), .Y(n_110) );
INVxp67_ASAP7_75t_L g180 ( .A(n_15), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_15), .B(n_60), .Y(n_186) );
INVx1_ASAP7_75t_L g409 ( .A(n_16), .Y(n_409) );
OA21x2_ASAP7_75t_L g262 ( .A1(n_17), .A2(n_55), .B(n_263), .Y(n_262) );
OA21x2_ASAP7_75t_L g270 ( .A1(n_17), .A2(n_55), .B(n_263), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g106 ( .A(n_18), .B(n_94), .Y(n_106) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_19), .A2(n_53), .B1(n_254), .B2(n_376), .Y(n_375) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_21), .Y(n_206) );
INVx1_ASAP7_75t_L g403 ( .A(n_23), .Y(n_403) );
BUFx3_ASAP7_75t_L g216 ( .A(n_24), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_25), .Y(n_203) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_26), .Y(n_94) );
AO22x1_ASAP7_75t_L g356 ( .A1(n_27), .A2(n_63), .B1(n_289), .B2(n_357), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_28), .Y(n_280) );
AND2x2_ASAP7_75t_L g299 ( .A(n_29), .B(n_244), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_30), .B(n_289), .Y(n_288) );
AOI22x1_ASAP7_75t_L g251 ( .A1(n_31), .A2(n_75), .B1(n_252), .B2(n_254), .Y(n_251) );
INVx1_ASAP7_75t_L g95 ( .A(n_32), .Y(n_95) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_32), .B(n_59), .Y(n_177) );
AOI22xp33_ASAP7_75t_L g170 ( .A1(n_33), .A2(n_42), .B1(n_171), .B2(n_181), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_34), .B(n_260), .Y(n_331) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_36), .B(n_307), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g122 ( .A1(n_38), .A2(n_67), .B1(n_123), .B2(n_128), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_39), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_40), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g263 ( .A(n_41), .Y(n_263) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_43), .Y(n_227) );
AND2x4_ASAP7_75t_L g265 ( .A(n_43), .B(n_225), .Y(n_265) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_44), .Y(n_250) );
INVx2_ASAP7_75t_L g378 ( .A(n_45), .Y(n_378) );
INVxp33_ASAP7_75t_SL g196 ( .A(n_46), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_46), .A2(n_61), .B1(n_252), .B2(n_276), .Y(n_324) );
CKINVDCx14_ASAP7_75t_R g365 ( .A(n_47), .Y(n_365) );
AND2x2_ASAP7_75t_L g304 ( .A(n_48), .B(n_289), .Y(n_304) );
OA22x2_ASAP7_75t_L g100 ( .A1(n_49), .A2(n_60), .B1(n_94), .B2(n_98), .Y(n_100) );
INVx1_ASAP7_75t_L g119 ( .A(n_49), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_50), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_52), .B(n_337), .Y(n_336) );
NAND2x1p5_ASAP7_75t_L g308 ( .A(n_54), .B(n_295), .Y(n_308) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_56), .Y(n_81) );
CKINVDCx14_ASAP7_75t_R g267 ( .A(n_58), .Y(n_267) );
INVx1_ASAP7_75t_L g112 ( .A(n_59), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_59), .B(n_117), .Y(n_189) );
HB1xp67_ASAP7_75t_L g219 ( .A(n_59), .Y(n_219) );
OAI21xp33_ASAP7_75t_L g120 ( .A1(n_60), .A2(n_64), .B(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_62), .B(n_277), .Y(n_342) );
INVx1_ASAP7_75t_L g97 ( .A(n_64), .Y(n_97) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_64), .B(n_74), .Y(n_187) );
INVx1_ASAP7_75t_L g243 ( .A(n_65), .Y(n_243) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_65), .Y(n_247) );
BUFx5_ASAP7_75t_L g256 ( .A(n_65), .Y(n_256) );
INVx2_ASAP7_75t_L g413 ( .A(n_66), .Y(n_413) );
NAND2xp33_ASAP7_75t_L g301 ( .A(n_69), .B(n_253), .Y(n_301) );
INVx2_ASAP7_75t_SL g225 ( .A(n_70), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_71), .B(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_72), .B(n_307), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_73), .A2(n_82), .B1(n_83), .B2(n_655), .Y(n_654) );
CKINVDCx5p33_ASAP7_75t_R g655 ( .A(n_73), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_74), .B(n_105), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_77), .B(n_293), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_211), .B1(n_228), .B2(n_642), .C(n_648), .Y(n_78) );
XNOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_191), .Y(n_79) );
AOI22xp33_ASAP7_75t_SL g80 ( .A1(n_81), .A2(n_82), .B1(n_83), .B2(n_190), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_81), .Y(n_190) );
AOI22xp33_ASAP7_75t_SL g649 ( .A1(n_82), .A2(n_83), .B1(n_650), .B2(n_651), .Y(n_649) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_83), .Y(n_82) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
NAND2xp5_ASAP7_75t_L g84 ( .A(n_85), .B(n_149), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
NAND4xp25_ASAP7_75t_SL g86 ( .A(n_87), .B(n_122), .C(n_131), .D(n_143), .Y(n_86) );
BUFx6f_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
AND2x4_ASAP7_75t_L g89 ( .A(n_90), .B(n_101), .Y(n_89) );
AND2x4_ASAP7_75t_L g133 ( .A(n_90), .B(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g140 ( .A(n_90), .B(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g145 ( .A(n_90), .B(n_126), .Y(n_145) );
AND2x4_ASAP7_75t_L g90 ( .A(n_91), .B(n_99), .Y(n_90) );
AND2x2_ASAP7_75t_L g155 ( .A(n_91), .B(n_100), .Y(n_155) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
AND2x2_ASAP7_75t_L g125 ( .A(n_92), .B(n_100), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g92 ( .A(n_93), .B(n_96), .Y(n_92) );
NAND2xp33_ASAP7_75t_L g93 ( .A(n_94), .B(n_95), .Y(n_93) );
INVx2_ASAP7_75t_L g98 ( .A(n_94), .Y(n_98) );
INVx3_ASAP7_75t_L g105 ( .A(n_94), .Y(n_105) );
NAND2xp33_ASAP7_75t_L g111 ( .A(n_94), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g121 ( .A(n_94), .Y(n_121) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_94), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_95), .B(n_119), .Y(n_118) );
INVxp67_ASAP7_75t_L g220 ( .A(n_95), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g96 ( .A(n_97), .B(n_98), .Y(n_96) );
OAI21xp5_ASAP7_75t_L g179 ( .A1(n_97), .A2(n_121), .B(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
AND2x2_ASAP7_75t_L g178 ( .A(n_100), .B(n_179), .Y(n_178) );
AND2x4_ASAP7_75t_L g114 ( .A(n_101), .B(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx2_ASAP7_75t_L g130 ( .A(n_102), .Y(n_130) );
OR2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_107), .Y(n_102) );
AND2x4_ASAP7_75t_L g126 ( .A(n_103), .B(n_127), .Y(n_126) );
AND2x4_ASAP7_75t_L g134 ( .A(n_103), .B(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g142 ( .A(n_103), .Y(n_142) );
AND2x2_ASAP7_75t_L g174 ( .A(n_103), .B(n_175), .Y(n_174) );
AND2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_105), .B(n_110), .Y(n_109) );
INVxp67_ASAP7_75t_L g117 ( .A(n_105), .Y(n_117) );
NAND3xp33_ASAP7_75t_L g188 ( .A(n_106), .B(n_116), .C(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g127 ( .A(n_107), .Y(n_127) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g135 ( .A(n_108), .Y(n_135) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
BUFx12f_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x4_ASAP7_75t_L g148 ( .A(n_115), .B(n_126), .Y(n_148) );
AND2x4_ASAP7_75t_L g157 ( .A(n_115), .B(n_141), .Y(n_157) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_120), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_119), .Y(n_221) );
BUFx8_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
AND2x4_ASAP7_75t_L g129 ( .A(n_125), .B(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g164 ( .A(n_125), .B(n_134), .Y(n_164) );
AND2x2_ASAP7_75t_L g169 ( .A(n_125), .B(n_141), .Y(n_169) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x4_ASAP7_75t_L g161 ( .A(n_134), .B(n_155), .Y(n_161) );
AND2x4_ASAP7_75t_L g141 ( .A(n_135), .B(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x4_ASAP7_75t_L g154 ( .A(n_141), .B(n_155), .Y(n_154) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx4_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx8_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NAND4xp25_ASAP7_75t_L g150 ( .A(n_151), .B(n_158), .C(n_165), .D(n_170), .Y(n_150) );
INVx2_ASAP7_75t_SL g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
BUFx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx4_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx5_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AND2x4_ASAP7_75t_L g173 ( .A(n_174), .B(n_178), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
INVx1_ASAP7_75t_L g184 ( .A(n_176), .Y(n_184) );
HB1xp67_ASAP7_75t_L g217 ( .A(n_177), .Y(n_217) );
INVx2_ASAP7_75t_SL g181 ( .A(n_182), .Y(n_181) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AO21x2_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_188), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_186), .B(n_187), .Y(n_185) );
OAI22xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B1(n_205), .B2(n_210), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_199), .B1(n_200), .B2(n_204), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_194), .Y(n_204) );
OAI22xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B1(n_197), .B2(n_198), .Y(n_194) );
INVx1_ASAP7_75t_L g197 ( .A(n_195), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_196), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_200), .Y(n_199) );
XNOR2xp5_ASAP7_75t_L g200 ( .A(n_201), .B(n_202), .Y(n_200) );
HB1xp67_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g210 ( .A(n_205), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B1(n_208), .B2(n_209), .Y(n_205) );
INVx1_ASAP7_75t_L g208 ( .A(n_206), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_207), .Y(n_209) );
BUFx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_214), .B(n_222), .Y(n_213) );
INVxp67_ASAP7_75t_SL g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g653 ( .A(n_215), .B(n_222), .Y(n_653) );
AOI211xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_218), .C(n_221), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_223), .B(n_226), .Y(n_222) );
OR2x2_ASAP7_75t_L g657 ( .A(n_223), .B(n_227), .Y(n_657) );
INVx1_ASAP7_75t_L g660 ( .A(n_223), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_223), .B(n_226), .Y(n_661) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_231), .B(n_531), .Y(n_230) );
NOR3xp33_ASAP7_75t_L g231 ( .A(n_232), .B(n_455), .C(n_501), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_421), .Y(n_232) );
AOI21xp33_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_332), .B(n_366), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_271), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_235), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_236), .B(n_429), .Y(n_617) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x4_ASAP7_75t_L g388 ( .A(n_237), .B(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g497 ( .A(n_237), .B(n_297), .Y(n_497) );
AND2x2_ASAP7_75t_L g593 ( .A(n_237), .B(n_297), .Y(n_593) );
AO31x2_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_259), .A3(n_264), .B(n_266), .Y(n_237) );
AO31x2_ASAP7_75t_L g434 ( .A1(n_238), .A2(n_259), .A3(n_264), .B(n_266), .Y(n_434) );
OAI22x1_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_248), .B1(n_251), .B2(n_257), .Y(n_238) );
INVx3_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g359 ( .A(n_243), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_244), .B(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g253 ( .A(n_246), .Y(n_253) );
INVx1_ASAP7_75t_L g307 ( .A(n_246), .Y(n_307) );
INVx6_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g283 ( .A(n_247), .Y(n_283) );
INVx2_ASAP7_75t_L g287 ( .A(n_247), .Y(n_287) );
INVx3_ASAP7_75t_L g330 ( .A(n_247), .Y(n_330) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_249), .B(n_322), .Y(n_326) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_250), .Y(n_258) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_250), .Y(n_291) );
INVxp67_ASAP7_75t_L g302 ( .A(n_250), .Y(n_302) );
INVx4_ASAP7_75t_L g373 ( .A(n_250), .Y(n_373) );
INVx3_ASAP7_75t_L g382 ( .A(n_250), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_250), .B(n_403), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_250), .B(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g277 ( .A(n_256), .Y(n_277) );
INVx2_ASAP7_75t_L g289 ( .A(n_256), .Y(n_289) );
INVx2_ASAP7_75t_L g347 ( .A(n_256), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_257), .B(n_279), .Y(n_278) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_257), .Y(n_645) );
INVx4_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g275 ( .A1(n_258), .A2(n_276), .B1(n_278), .B2(n_281), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_258), .B(n_322), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_258), .A2(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_262), .B(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g374 ( .A(n_262), .Y(n_374) );
OAI21x1_ASAP7_75t_L g274 ( .A1(n_264), .A2(n_275), .B(n_284), .Y(n_274) );
AND2x2_ASAP7_75t_L g643 ( .A(n_264), .B(n_644), .Y(n_643) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx3_ASAP7_75t_L g315 ( .A(n_265), .Y(n_315) );
INVx3_ASAP7_75t_L g323 ( .A(n_265), .Y(n_323) );
INVx1_ASAP7_75t_L g353 ( .A(n_265), .Y(n_353) );
NOR2xp67_ASAP7_75t_SL g266 ( .A(n_267), .B(n_268), .Y(n_266) );
OR2x2_ASAP7_75t_L g364 ( .A(n_268), .B(n_365), .Y(n_364) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OA21x2_ASAP7_75t_L g273 ( .A1(n_269), .A2(n_274), .B(n_292), .Y(n_273) );
OA21x2_ASAP7_75t_L g393 ( .A1(n_269), .A2(n_274), .B(n_292), .Y(n_393) );
BUFx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx4_ASAP7_75t_L g296 ( .A(n_270), .Y(n_296) );
INVx2_ASAP7_75t_L g338 ( .A(n_270), .Y(n_338) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_317), .Y(n_271) );
INVx2_ASAP7_75t_L g494 ( .A(n_272), .Y(n_494) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_297), .Y(n_272) );
NAND2x1_ASAP7_75t_L g467 ( .A(n_273), .B(n_433), .Y(n_467) );
AND2x2_ASAP7_75t_L g508 ( .A(n_273), .B(n_319), .Y(n_508) );
AND2x2_ASAP7_75t_L g513 ( .A(n_273), .B(n_420), .Y(n_513) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_288), .B(n_290), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_286), .B(n_405), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_286), .A2(n_289), .B1(n_408), .B2(n_410), .Y(n_407) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g647 ( .A(n_287), .Y(n_647) );
INVxp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_SL g310 ( .A(n_291), .Y(n_310) );
INVx1_ASAP7_75t_L g348 ( .A(n_291), .Y(n_348) );
INVx1_ASAP7_75t_L g355 ( .A(n_291), .Y(n_355) );
OR2x2_ASAP7_75t_L g352 ( .A(n_293), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g377 ( .A(n_294), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx3_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g313 ( .A(n_296), .Y(n_313) );
AND2x4_ASAP7_75t_L g484 ( .A(n_297), .B(n_429), .Y(n_484) );
AO21x2_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_303), .B(n_311), .Y(n_297) );
AO21x2_ASAP7_75t_L g390 ( .A1(n_298), .A2(n_303), .B(n_311), .Y(n_390) );
OAI21x1_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_300), .B(n_302), .Y(n_298) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OAI21x1_ASAP7_75t_SL g303 ( .A1(n_304), .A2(n_305), .B(n_309), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_308), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g316 ( .A(n_308), .Y(n_316) );
AOI21x1_ASAP7_75t_L g360 ( .A1(n_310), .A2(n_361), .B(n_362), .Y(n_360) );
AOI21xp33_ASAP7_75t_SL g311 ( .A1(n_312), .A2(n_314), .B(n_316), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND3xp33_ASAP7_75t_SL g372 ( .A(n_314), .B(n_373), .C(n_374), .Y(n_372) );
NAND3xp33_ASAP7_75t_L g380 ( .A(n_314), .B(n_374), .C(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NOR2x1_ASAP7_75t_L g349 ( .A(n_315), .B(n_337), .Y(n_349) );
INVx1_ASAP7_75t_L g589 ( .A(n_317), .Y(n_589) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g458 ( .A(n_318), .Y(n_458) );
OR2x2_ASAP7_75t_L g553 ( .A(n_318), .B(n_467), .Y(n_553) );
AND2x2_ASAP7_75t_L g561 ( .A(n_318), .B(n_432), .Y(n_561) );
INVx2_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_325), .Y(n_319) );
NAND2x1p5_ASAP7_75t_L g420 ( .A(n_320), .B(n_325), .Y(n_420) );
OR2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_324), .Y(n_320) );
OA21x2_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_327), .B(n_331), .Y(n_325) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g376 ( .A(n_329), .Y(n_376) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g345 ( .A(n_330), .Y(n_345) );
INVx1_ASAP7_75t_L g363 ( .A(n_330), .Y(n_363) );
AOI32xp33_ASAP7_75t_L g557 ( .A1(n_332), .A2(n_554), .A3(n_558), .B1(n_560), .B2(n_561), .Y(n_557) );
AOI221x1_ASAP7_75t_L g575 ( .A1(n_332), .A2(n_576), .B1(n_579), .B2(n_581), .C(n_582), .Y(n_575) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g443 ( .A(n_333), .B(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g586 ( .A(n_334), .B(n_474), .Y(n_586) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_350), .Y(n_334) );
INVx3_ASAP7_75t_L g386 ( .A(n_335), .Y(n_386) );
INVx2_ASAP7_75t_L g473 ( .A(n_335), .Y(n_473) );
AND2x2_ASAP7_75t_L g488 ( .A(n_335), .B(n_351), .Y(n_488) );
AND2x4_ASAP7_75t_L g335 ( .A(n_336), .B(n_339), .Y(n_335) );
INVx3_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_338), .B(n_413), .Y(n_412) );
OAI21x1_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_343), .B(n_349), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_346), .B(n_348), .Y(n_343) );
INVx1_ASAP7_75t_L g414 ( .A(n_350), .Y(n_414) );
INVx1_ASAP7_75t_L g441 ( .A(n_350), .Y(n_441) );
AND2x2_ASAP7_75t_L g549 ( .A(n_350), .B(n_397), .Y(n_549) );
INVx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g385 ( .A(n_351), .B(n_386), .Y(n_385) );
OAI21x1_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_354), .B(n_364), .Y(n_351) );
OAI21xp5_ASAP7_75t_L g454 ( .A1(n_352), .A2(n_354), .B(n_364), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_353), .B(n_399), .Y(n_398) );
AOI21x1_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_356), .B(n_360), .Y(n_354) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OAI22xp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_387), .B1(n_394), .B2(n_415), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_367), .A2(n_477), .B1(n_580), .B2(n_611), .Y(n_610) );
OR2x2_ASAP7_75t_SL g367 ( .A(n_368), .B(n_384), .Y(n_367) );
OR2x2_ASAP7_75t_L g461 ( .A(n_368), .B(n_439), .Y(n_461) );
INVx2_ASAP7_75t_L g559 ( .A(n_368), .Y(n_559) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g631 ( .A(n_369), .B(n_452), .Y(n_631) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NOR2x1_ASAP7_75t_L g425 ( .A(n_370), .B(n_426), .Y(n_425) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_370), .Y(n_451) );
AND2x2_ASAP7_75t_L g463 ( .A(n_370), .B(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g475 ( .A(n_370), .Y(n_475) );
AND2x2_ASAP7_75t_L g500 ( .A(n_370), .B(n_397), .Y(n_500) );
INVx1_ASAP7_75t_L g520 ( .A(n_370), .Y(n_520) );
INVx1_ASAP7_75t_L g547 ( .A(n_370), .Y(n_547) );
AND2x2_ASAP7_75t_L g623 ( .A(n_370), .B(n_386), .Y(n_623) );
OR2x6_ASAP7_75t_L g370 ( .A(n_371), .B(n_379), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_375), .B(n_377), .Y(n_371) );
NOR2xp33_ASAP7_75t_SL g408 ( .A(n_373), .B(n_409), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_373), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g399 ( .A(n_374), .Y(n_399) );
NOR2xp67_ASAP7_75t_L g379 ( .A(n_380), .B(n_383), .Y(n_379) );
INVx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g580 ( .A(n_384), .B(n_547), .Y(n_580) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x4_ASAP7_75t_L g424 ( .A(n_385), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g462 ( .A(n_385), .B(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g440 ( .A(n_386), .Y(n_440) );
OAI22xp33_ASAP7_75t_L g442 ( .A1(n_387), .A2(n_443), .B1(n_445), .B2(n_449), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_391), .Y(n_387) );
AND2x4_ASAP7_75t_L g571 ( .A(n_388), .B(n_508), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_388), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g448 ( .A(n_389), .Y(n_448) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g417 ( .A(n_390), .Y(n_417) );
INVxp67_ASAP7_75t_L g459 ( .A(n_390), .Y(n_459) );
AND2x2_ASAP7_75t_L g510 ( .A(n_390), .B(n_433), .Y(n_510) );
AND3x2_ASAP7_75t_L g457 ( .A(n_391), .B(n_458), .C(n_459), .Y(n_457) );
OR2x2_ASAP7_75t_L g496 ( .A(n_391), .B(n_497), .Y(n_496) );
OR2x2_ASAP7_75t_L g577 ( .A(n_391), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_392), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g437 ( .A(n_392), .B(n_420), .Y(n_437) );
AND2x2_ASAP7_75t_L g640 ( .A(n_392), .B(n_434), .Y(n_640) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g429 ( .A(n_393), .Y(n_429) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_393), .Y(n_447) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_414), .Y(n_395) );
NOR2xp67_ASAP7_75t_SL g438 ( .A(n_396), .B(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g481 ( .A(n_396), .Y(n_481) );
AND2x2_ASAP7_75t_L g568 ( .A(n_396), .B(n_472), .Y(n_568) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g426 ( .A(n_397), .Y(n_426) );
OR2x2_ASAP7_75t_L g453 ( .A(n_397), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g464 ( .A(n_397), .Y(n_464) );
INVxp67_ASAP7_75t_L g517 ( .A(n_397), .Y(n_517) );
AO21x2_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_400), .B(n_412), .Y(n_397) );
NAND3xp33_ASAP7_75t_SL g400 ( .A(n_401), .B(n_404), .C(n_407), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_414), .B(n_463), .Y(n_587) );
OR2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_418), .Y(n_415) );
INVx1_ASAP7_75t_L g469 ( .A(n_416), .Y(n_469) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_417), .B(n_420), .Y(n_578) );
INVxp67_ASAP7_75t_L g566 ( .A(n_418), .Y(n_566) );
AND2x2_ASAP7_75t_L g538 ( .A(n_419), .B(n_433), .Y(n_538) );
AND2x2_ASAP7_75t_L g584 ( .A(n_419), .B(n_484), .Y(n_584) );
INVx1_ASAP7_75t_L g621 ( .A(n_419), .Y(n_621) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g487 ( .A(n_420), .Y(n_487) );
INVx1_ASAP7_75t_L g597 ( .A(n_420), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_422), .B(n_442), .Y(n_421) );
OAI21xp5_ASAP7_75t_SL g422 ( .A1(n_423), .A2(n_427), .B(n_435), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g444 ( .A(n_425), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_430), .Y(n_427) );
INVxp67_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g492 ( .A(n_430), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g436 ( .A(n_431), .B(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g483 ( .A(n_431), .B(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g541 ( .A(n_432), .Y(n_541) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g527 ( .A(n_433), .Y(n_527) );
INVx3_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NAND2x1p5_ASAP7_75t_L g435 ( .A(n_436), .B(n_438), .Y(n_435) );
INVx1_ASAP7_75t_L g628 ( .A(n_436), .Y(n_628) );
INVx1_ASAP7_75t_L g542 ( .A(n_437), .Y(n_542) );
OR2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
INVx1_ASAP7_75t_L g598 ( .A(n_440), .Y(n_598) );
INVxp67_ASAP7_75t_SL g607 ( .A(n_441), .Y(n_607) );
INVx1_ASAP7_75t_L g560 ( .A(n_443), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g602 ( .A1(n_443), .A2(n_587), .B(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g609 ( .A(n_444), .B(n_472), .Y(n_609) );
INVxp33_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
INVx1_ASAP7_75t_L g639 ( .A(n_448), .Y(n_639) );
INVx2_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g503 ( .A(n_450), .Y(n_503) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_451), .Y(n_536) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g523 ( .A(n_453), .Y(n_523) );
OR2x2_ASAP7_75t_L g534 ( .A(n_453), .B(n_473), .Y(n_534) );
BUFx2_ASAP7_75t_L g519 ( .A(n_454), .Y(n_519) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_479), .C(n_489), .Y(n_455) );
AOI222xp33_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_460), .B1(n_462), .B2(n_465), .C1(n_470), .C2(n_476), .Y(n_456) );
NAND2x1_ASAP7_75t_L g603 ( .A(n_458), .B(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_458), .B(n_510), .Y(n_611) );
AND2x2_ASAP7_75t_L g619 ( .A(n_458), .B(n_593), .Y(n_619) );
INVx1_ASAP7_75t_L g478 ( .A(n_459), .Y(n_478) );
AND2x2_ASAP7_75t_L g512 ( .A(n_459), .B(n_513), .Y(n_512) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_459), .Y(n_633) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_462), .B(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g474 ( .A(n_464), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_466), .B(n_468), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_L g477 ( .A(n_467), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_474), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_473), .B(n_517), .Y(n_516) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_473), .Y(n_522) );
AND2x2_ASAP7_75t_L g546 ( .A(n_473), .B(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND3xp33_ASAP7_75t_L g479 ( .A(n_480), .B(n_482), .C(n_485), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_480), .A2(n_592), .B1(n_594), .B2(n_599), .Y(n_591) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
O2A1O1Ixp5_ASAP7_75t_L g605 ( .A1(n_483), .A2(n_606), .B(n_608), .C(n_610), .Y(n_605) );
AND2x4_ASAP7_75t_SL g526 ( .A(n_484), .B(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_488), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g555 ( .A(n_487), .Y(n_555) );
INVx1_ASAP7_75t_L g601 ( .A(n_487), .Y(n_601) );
AND2x2_ASAP7_75t_L g499 ( .A(n_488), .B(n_500), .Y(n_499) );
OAI21xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_495), .B(n_498), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g556 ( .A(n_497), .Y(n_556) );
INVx2_ASAP7_75t_L g604 ( .A(n_497), .Y(n_604) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g606 ( .A(n_500), .B(n_607), .Y(n_606) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_500), .Y(n_627) );
OAI211xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_504), .B(n_514), .C(n_528), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_511), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_509), .Y(n_506) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx3_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_510), .B(n_621), .Y(n_620) );
INVx2_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
O2A1O1Ixp5_ASAP7_75t_L g563 ( .A1(n_512), .A2(n_564), .B(n_567), .C(n_569), .Y(n_563) );
INVx1_ASAP7_75t_L g530 ( .A(n_513), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_513), .B(n_636), .Y(n_635) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_521), .B(n_524), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_515), .A2(n_544), .B1(n_550), .B2(n_554), .Y(n_543) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_518), .Y(n_515) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_517), .Y(n_574) );
AND2x2_ASAP7_75t_L g567 ( .A(n_518), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_518), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_523), .Y(n_521) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g636 ( .A(n_527), .Y(n_636) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NOR3xp33_ASAP7_75t_L g531 ( .A(n_532), .B(n_562), .C(n_612), .Y(n_531) );
OAI211xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_537), .B(n_543), .C(n_557), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_534), .Y(n_637) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AOI21x1_ASAP7_75t_L g569 ( .A1(n_540), .A2(n_570), .B(n_572), .Y(n_569) );
OR2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NAND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_548), .Y(n_545) );
BUFx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x4_ASAP7_75t_L g622 ( .A(n_549), .B(n_623), .Y(n_622) );
INVxp67_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_559), .A2(n_591), .B(n_602), .Y(n_590) );
NAND4xp25_ASAP7_75t_L g562 ( .A(n_563), .B(n_575), .C(n_590), .D(n_605), .Y(n_562) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g581 ( .A(n_578), .Y(n_581) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OAI22x1_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_585), .B1(n_587), .B2(n_588), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g600 ( .A(n_593), .B(n_601), .Y(n_600) );
INVx2_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g630 ( .A(n_595), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g641 ( .A(n_606), .Y(n_641) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_629), .Y(n_612) );
AOI21xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_622), .B(n_624), .Y(n_613) );
NAND3xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_618), .C(n_620), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g625 ( .A(n_623), .Y(n_625) );
AOI21xp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_626), .B(n_628), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AOI21xp33_ASAP7_75t_SL g629 ( .A1(n_630), .A2(n_632), .B(n_634), .Y(n_629) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_637), .B1(n_638), .B2(n_641), .Y(n_634) );
NAND2x1p5_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
BUFx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OA21x2_ASAP7_75t_L g659 ( .A1(n_644), .A2(n_660), .B(n_661), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OAI222xp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_651), .B1(n_652), .B2(n_654), .C1(n_656), .C2(n_658), .Y(n_648) );
CKINVDCx16_ASAP7_75t_R g651 ( .A(n_650), .Y(n_651) );
INVx1_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
BUFx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
endmodule