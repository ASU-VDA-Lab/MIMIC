module real_jpeg_26667_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_314, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_314;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_0),
.A2(n_35),
.B1(n_36),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_0),
.A2(n_46),
.B1(n_53),
.B2(n_54),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_46),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_0),
.A2(n_46),
.B1(n_60),
.B2(n_62),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_1),
.Y(n_90)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_1),
.Y(n_93)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_1),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_2),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_99),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_2),
.A2(n_53),
.B1(n_54),
.B2(n_99),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_2),
.A2(n_60),
.B1(n_62),
.B2(n_99),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_3),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_SL g161 ( 
.A1(n_3),
.A2(n_32),
.B(n_36),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_160),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_3),
.B(n_34),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_3),
.A2(n_53),
.B(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_3),
.B(n_53),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_3),
.B(n_57),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_3),
.A2(n_88),
.B1(n_250),
.B2(n_254),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_3),
.A2(n_35),
.B(n_266),
.Y(n_265)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_5),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_156),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_5),
.A2(n_53),
.B1(n_54),
.B2(n_156),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_5),
.A2(n_60),
.B1(n_62),
.B2(n_156),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_6),
.A2(n_35),
.B1(n_36),
.B2(n_40),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_6),
.A2(n_40),
.B1(n_53),
.B2(n_54),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_6),
.A2(n_40),
.B1(n_60),
.B2(n_62),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_8),
.A2(n_53),
.B1(n_54),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_8),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_8),
.A2(n_60),
.B1(n_62),
.B2(n_67),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_67),
.Y(n_108)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_10),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g145 ( 
.A1(n_10),
.A2(n_29),
.B1(n_53),
.B2(n_54),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_10),
.A2(n_29),
.B1(n_60),
.B2(n_62),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_11),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_11),
.A2(n_53),
.B1(n_54),
.B2(n_63),
.Y(n_65)
);

OAI32xp33_ASAP7_75t_L g226 ( 
.A1(n_11),
.A2(n_53),
.A3(n_62),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_12),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_132),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_12),
.A2(n_60),
.B1(n_62),
.B2(n_132),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_12),
.A2(n_53),
.B1(n_54),
.B2(n_132),
.Y(n_270)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_14),
.B(n_35),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_14),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_14),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_15),
.A2(n_35),
.B1(n_36),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_15),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_15),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_15),
.A2(n_56),
.B1(n_60),
.B2(n_62),
.Y(n_127)
);

INVx11_ASAP7_75t_SL g61 ( 
.A(n_16),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_17),
.A2(n_27),
.B1(n_28),
.B2(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_17),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_L g187 ( 
.A1(n_17),
.A2(n_35),
.B1(n_36),
.B2(n_149),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_17),
.A2(n_53),
.B1(n_54),
.B2(n_149),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_17),
.A2(n_60),
.B1(n_62),
.B2(n_149),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_113),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_112),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_100),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_22),
.B(n_100),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_71),
.C(n_77),
.Y(n_22)
);

FAx1_ASAP7_75t_SL g133 ( 
.A(n_23),
.B(n_71),
.CI(n_77),
.CON(n_133),
.SN(n_133)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_42),
.B2(n_70),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_24),
.A2(n_25),
.B1(n_102),
.B2(n_110),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_25),
.B(n_43),
.C(n_69),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_39),
.B2(n_41),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_26),
.A2(n_30),
.B1(n_41),
.B2(n_97),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_31)
);

NAND2xp33_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_32),
.Y(n_33)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_28),
.A2(n_38),
.B(n_160),
.C(n_161),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_30),
.A2(n_41),
.B1(n_154),
.B2(n_157),
.Y(n_153)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_31),
.A2(n_34),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_31),
.A2(n_34),
.B1(n_98),
.B2(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_31),
.A2(n_34),
.B1(n_131),
.B2(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_31),
.A2(n_34),
.B1(n_155),
.B2(n_193),
.Y(n_192)
);

AO22x1_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_34)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_49),
.B(n_51),
.C(n_52),
.Y(n_48)
);

OAI32xp33_ASAP7_75t_L g274 ( 
.A1(n_35),
.A2(n_54),
.A3(n_267),
.B1(n_275),
.B2(n_277),
.Y(n_274)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_36),
.B(n_160),
.Y(n_267)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_39),
.Y(n_104)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_58),
.B1(n_68),
.B2(n_69),
.Y(n_42)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B1(n_55),
.B2(n_57),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_48),
.B1(n_52),
.B2(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_47),
.A2(n_55),
.B1(n_57),
.B2(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_47),
.A2(n_57),
.B1(n_74),
.B2(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_47),
.A2(n_57),
.B1(n_124),
.B2(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_47),
.A2(n_57),
.B1(n_187),
.B2(n_198),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_48),
.A2(n_52),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_48),
.A2(n_52),
.B1(n_166),
.B2(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_48),
.A2(n_52),
.B1(n_199),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_53),
.B(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_58),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_58),
.A2(n_69),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_64),
.B(n_66),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_59),
.B(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_59),
.A2(n_64),
.B1(n_66),
.B2(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_59),
.A2(n_64),
.B1(n_83),
.B2(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_59),
.A2(n_64),
.B1(n_129),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_59),
.A2(n_64),
.B1(n_222),
.B2(n_224),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_59),
.A2(n_64),
.B1(n_224),
.B2(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_59),
.B(n_160),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_59),
.A2(n_64),
.B1(n_191),
.B2(n_294),
.Y(n_293)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_60),
.B(n_63),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_60),
.B(n_256),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_71),
.A2(n_72),
.B(n_75),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_76),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_95),
.B(n_96),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_78),
.A2(n_79),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_87),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_80),
.A2(n_81),
.B1(n_87),
.B2(n_95),
.Y(n_171)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_84),
.A2(n_86),
.B1(n_145),
.B2(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_84),
.A2(n_86),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_87),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_95),
.B1(n_96),
.B2(n_118),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_91),
.B(n_94),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_88),
.A2(n_93),
.B1(n_94),
.B2(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_88),
.A2(n_91),
.B1(n_127),
.B2(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_88),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_88),
.A2(n_93),
.B1(n_244),
.B2(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_88),
.A2(n_238),
.B1(n_239),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_89),
.A2(n_142),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_89),
.A2(n_92),
.B1(n_163),
.B2(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_89),
.A2(n_92),
.B1(n_243),
.B2(n_245),
.Y(n_242)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_91),
.Y(n_164)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx5_ASAP7_75t_SL g239 ( 
.A(n_92),
.Y(n_239)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_111),
.Y(n_100)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_106),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_107),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_134),
.B(n_310),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_133),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_115),
.B(n_133),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.C(n_121),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_116),
.B(n_120),
.Y(n_178)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_121),
.A2(n_122),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_125),
.C(n_130),
.Y(n_122)
);

FAx1_ASAP7_75t_SL g172 ( 
.A(n_123),
.B(n_125),
.CI(n_130),
.CON(n_172),
.SN(n_172)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_128),
.Y(n_168)
);

BUFx24_ASAP7_75t_SL g311 ( 
.A(n_133),
.Y(n_311)
);

AOI321xp33_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_174),
.A3(n_179),
.B1(n_304),
.B2(n_309),
.C(n_314),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_136),
.A2(n_305),
.B(n_308),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_169),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_137),
.B(n_169),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_152),
.C(n_168),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_138),
.B(n_168),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_146),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_147),
.C(n_150),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_140),
.B(n_143),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_148),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_151),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_152),
.B(n_213),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_158),
.C(n_165),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_153),
.B(n_165),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_158),
.B(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_162),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_160),
.B(n_254),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_172),
.C(n_173),
.Y(n_175)
);

BUFx24_ASAP7_75t_SL g313 ( 
.A(n_172),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_175),
.B(n_176),
.Y(n_309)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NOR3xp33_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_209),
.C(n_214),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_203),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_181),
.B(n_203),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_194),
.C(n_195),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_182),
.B(n_301),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_192),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_188),
.B2(n_189),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_189),
.C(n_192),
.Y(n_206)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_302),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_194),
.Y(n_302)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.C(n_202),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_197),
.B(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_200),
.B(n_202),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_201),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_206),
.C(n_207),
.Y(n_211)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AOI21xp33_ASAP7_75t_L g305 ( 
.A1(n_210),
.A2(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_211),
.B(n_212),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_298),
.B(n_303),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_284),
.B(n_297),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_260),
.B(n_283),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_240),
.B(n_259),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_229),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_219),
.B(n_229),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_225),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_220),
.A2(n_221),
.B1(n_225),
.B2(n_226),
.Y(n_246)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_223),
.Y(n_227)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_236),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_234),
.C(n_236),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_235),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_237),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_247),
.B(n_258),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_242),
.B(n_246),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_252),
.B(n_257),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_249),
.B(n_251),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_261),
.B(n_262),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_273),
.B1(n_281),
.B2(n_282),
.Y(n_262)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_268),
.B1(n_271),
.B2(n_272),
.Y(n_263)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_264),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_268),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_272),
.C(n_282),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_270),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_273),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_279),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_279),
.Y(n_292)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_275),
.Y(n_278)
);

INVx8_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_285),
.B(n_286),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_290),
.B2(n_291),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_293),
.C(n_295),
.Y(n_299)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_295),
.B2(n_296),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_292),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_293),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_299),
.B(n_300),
.Y(n_303)
);


endmodule