module real_jpeg_15276_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_0),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_0),
.B(n_51),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_0),
.B(n_98),
.Y(n_97)
);

INVxp33_ASAP7_75t_L g169 ( 
.A(n_0),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_0),
.B(n_228),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_0),
.B(n_245),
.Y(n_244)
);

AND2x2_ASAP7_75t_SL g280 ( 
.A(n_0),
.B(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_1),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_1),
.B(n_40),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_1),
.B(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_2),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_2),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_2),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_3),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_3),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_3),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_3),
.B(n_247),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_3),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_3),
.B(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_3),
.B(n_381),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_3),
.B(n_421),
.Y(n_420)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_4),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_4),
.Y(n_148)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_4),
.Y(n_242)
);

BUFx5_ASAP7_75t_L g245 ( 
.A(n_4),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_4),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_5),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_5),
.B(n_51),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_5),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_5),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_5),
.B(n_187),
.Y(n_186)
);

AOI22x1_ASAP7_75t_L g213 ( 
.A1(n_5),
.A2(n_8),
.B1(n_214),
.B2(n_218),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_5),
.Y(n_325)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g217 ( 
.A(n_6),
.Y(n_217)
);

BUFx5_ASAP7_75t_L g384 ( 
.A(n_6),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_7),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_7),
.Y(n_130)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_7),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_7),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_8),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_8),
.B(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_8),
.B(n_284),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_8),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_8),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_8),
.B(n_405),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_8),
.B(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_8),
.B(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_9),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_9),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_9),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_9),
.B(n_40),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_9),
.B(n_192),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_10),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_10),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_11),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_11),
.B(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_11),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_11),
.B(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_11),
.B(n_437),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_11),
.B(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_11),
.B(n_461),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_12),
.B(n_28),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_12),
.B(n_133),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g150 ( 
.A(n_12),
.B(n_32),
.Y(n_150)
);

AND2x4_ASAP7_75t_L g234 ( 
.A(n_12),
.B(n_235),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_12),
.B(n_245),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_12),
.B(n_142),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_12),
.B(n_384),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_13),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_14),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_14),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_14),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_14),
.B(n_183),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_14),
.B(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_14),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_14),
.B(n_217),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g84 ( 
.A(n_15),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_15),
.Y(n_144)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_15),
.Y(n_230)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_16),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_202),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_200),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_155),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_21),
.B(n_155),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_89),
.C(n_116),
.Y(n_21)
);

XNOR2x1_ASAP7_75t_L g297 ( 
.A(n_22),
.B(n_89),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_66),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_48),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_24),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_34),
.B1(n_46),
.B2(n_47),
.Y(n_24)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_26),
.Y(n_180)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_27),
.B(n_140),
.C(n_141),
.Y(n_139)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_30),
.Y(n_184)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_31),
.A2(n_62),
.B1(n_65),
.B2(n_154),
.Y(n_153)
);

MAJx2_ASAP7_75t_L g179 ( 
.A(n_31),
.B(n_47),
.C(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_32),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_34),
.Y(n_47)
);

MAJx2_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_39),
.C(n_42),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_35),
.B(n_39),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_35),
.A2(n_92),
.B1(n_93),
.B2(n_96),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_35),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_36),
.B(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_38),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_39),
.B(n_78),
.C(n_81),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_39),
.B(n_81),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_40),
.Y(n_281)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_41),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_42),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_42),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_42),
.A2(n_86),
.B1(n_227),
.B2(n_273),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_48),
.B(n_157),
.C(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_62),
.C(n_65),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_49),
.B(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_55),
.C(n_58),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_50),
.B(n_58),
.Y(n_137)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_55),
.B(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_62),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_64),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_66),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_77),
.C(n_85),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_67),
.B(n_77),
.Y(n_256)
);

XNOR2x1_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_71),
.C(n_72),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2x1_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_120),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_83),
.Y(n_419)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_84),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_85),
.B(n_256),
.Y(n_255)
);

MAJx2_ASAP7_75t_L g222 ( 
.A(n_86),
.B(n_223),
.C(n_227),
.Y(n_222)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_104),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_90),
.B(n_105),
.C(n_106),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_97),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_92),
.A2(n_93),
.B1(n_163),
.B2(n_167),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_93),
.B(n_96),
.C(n_97),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_103),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g221 ( 
.A(n_103),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_103),
.Y(n_323)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_103),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_107),
.B(n_111),
.C(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_109),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_115),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_116),
.B(n_297),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_138),
.C(n_151),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_118),
.B(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_121),
.C(n_136),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_119),
.B(n_121),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_127),
.C(n_131),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_122),
.A2(n_131),
.B1(n_132),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_122),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_127),
.B(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g438 ( 
.A(n_130),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_131),
.B(n_351),
.C(n_355),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_131),
.A2(n_132),
.B1(n_355),
.B2(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_136),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_138),
.B(n_152),
.Y(n_254)
);

MAJx2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_145),
.C(n_149),
.Y(n_138)
);

XNOR2x1_ASAP7_75t_SL g249 ( 
.A(n_139),
.B(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_140),
.B(n_141),
.Y(n_211)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_145),
.A2(n_149),
.B1(n_150),
.B2(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_145),
.Y(n_251)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_149),
.A2(n_150),
.B1(n_334),
.B2(n_335),
.Y(n_387)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_150),
.B(n_331),
.C(n_334),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_177),
.B1(n_198),
.B2(n_199),
.Y(n_159)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

XNOR2x1_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_173),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_168),
.Y(n_161)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_166),
.Y(n_237)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_166),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_197),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_211),
.Y(n_210)
);

XNOR2x1_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.Y(n_181)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_190),
.B1(n_191),
.B2(n_196),
.Y(n_185)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_186),
.Y(n_196)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_195),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AO21x2_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_301),
.B(n_471),
.Y(n_203)
);

NOR2xp67_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_295),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_259),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_206),
.B(n_259),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_252),
.Y(n_206)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_207),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_231),
.C(n_248),
.Y(n_207)
);

INVxp33_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XNOR2x1_ASAP7_75t_SL g261 ( 
.A(n_209),
.B(n_262),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.C(n_222),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_210),
.B(n_338),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_212),
.A2(n_213),
.B1(n_222),
.B2(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_213),
.A2(n_316),
.B(n_324),
.Y(n_315)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_222),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_223),
.B(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_226),
.Y(n_285)
);

INVx11_ASAP7_75t_SL g273 ( 
.A(n_227),
.Y(n_273)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_232),
.A2(n_248),
.B1(n_249),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_243),
.C(n_246),
.Y(n_232)
);

XOR2x2_ASAP7_75t_L g289 ( 
.A(n_233),
.B(n_290),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_238),
.C(n_240),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_234),
.A2(n_240),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_234),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_234),
.B(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_238),
.B(n_312),
.Y(n_311)
);

INVx13_ASAP7_75t_SL g314 ( 
.A(n_240),
.Y(n_314)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_242),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_243),
.A2(n_244),
.B1(n_246),
.B2(n_291),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_245),
.Y(n_377)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_246),
.Y(n_291)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_255),
.B1(n_257),
.B2(n_258),
.Y(n_252)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_253),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_255),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_255),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_257),
.B(n_299),
.C(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_264),
.C(n_267),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_261),
.B(n_264),
.Y(n_305)
);

XOR2x2_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_268),
.B(n_305),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_289),
.C(n_292),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_269),
.B(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_274),
.C(n_282),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_271),
.B(n_362),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_274),
.B(n_282),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_280),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_275),
.B(n_280),
.Y(n_360)
);

NOR2x1_ASAP7_75t_R g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_279),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_286),
.C(n_287),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_283),
.A2(n_286),
.B1(n_347),
.B2(n_348),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_283),
.Y(n_347)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_286),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_286),
.B(n_433),
.C(n_435),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_286),
.A2(n_348),
.B1(n_435),
.B2(n_436),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_287),
.B(n_346),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_292),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_295),
.A2(n_472),
.B(n_473),
.Y(n_471)
);

AND2x2_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_298),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_296),
.B(n_298),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_365),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_306),
.C(n_340),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_304),
.B(n_307),
.Y(n_470)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_310),
.C(n_337),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_308),
.B(n_364),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_310),
.B(n_337),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_315),
.C(n_330),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_311),
.B(n_315),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_313),
.B(n_400),
.C(n_404),
.Y(n_399)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_330),
.B(n_343),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g386 ( 
.A(n_331),
.B(n_387),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_332),
.B(n_333),
.Y(n_374)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_332),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_332),
.A2(n_442),
.B1(n_443),
.B2(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

NOR2xp67_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_363),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_341),
.B(n_363),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_344),
.C(n_361),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_342),
.B(n_389),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_344),
.B(n_361),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_349),
.C(n_359),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_345),
.B(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_360),
.Y(n_372)
);

XOR2x2_ASAP7_75t_L g408 ( 
.A(n_351),
.B(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_355),
.Y(n_410)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

NAND3xp33_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.C(n_470),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_368),
.A2(n_390),
.B(n_469),
.Y(n_367)
);

NOR2xp67_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_388),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_369),
.B(n_388),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_373),
.C(n_385),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_370),
.A2(n_371),
.B1(n_393),
.B2(n_394),
.Y(n_392)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_373),
.A2(n_385),
.B1(n_386),
.B2(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_373),
.Y(n_395)
);

MAJx2_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.C(n_378),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_375),
.Y(n_398)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_378),
.B(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_383),
.Y(n_378)
);

AO22x1_ASAP7_75t_SL g423 ( 
.A1(n_379),
.A2(n_380),
.B1(n_383),
.B2(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_383),
.Y(n_424)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_384),
.Y(n_422)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_384),
.Y(n_445)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_391),
.A2(n_411),
.B(n_468),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_392),
.B(n_396),
.Y(n_391)
);

NOR2xp67_ASAP7_75t_SL g468 ( 
.A(n_392),
.B(n_396),
.Y(n_468)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_399),
.C(n_407),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_397),
.B(n_426),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_399),
.B(n_408),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_400),
.B(n_404),
.Y(n_415)
);

INVx8_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx6_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx8_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

OAI21x1_ASAP7_75t_SL g411 ( 
.A1(n_412),
.A2(n_427),
.B(n_467),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_425),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_413),
.B(n_425),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_416),
.C(n_423),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_414),
.B(n_430),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_416),
.A2(n_417),
.B1(n_423),
.B2(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_420),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_418),
.B(n_420),
.Y(n_434)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_423),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_424),
.B(n_460),
.Y(n_459)
);

AOI21x1_ASAP7_75t_SL g427 ( 
.A1(n_428),
.A2(n_439),
.B(n_466),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_429),
.B(n_432),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_429),
.B(n_432),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_433),
.A2(n_434),
.B1(n_447),
.B2(n_448),
.Y(n_446)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_440),
.A2(n_449),
.B(n_465),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_446),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_441),
.B(n_446),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_442),
.B(n_443),
.Y(n_441)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_443),
.Y(n_458)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_450),
.A2(n_459),
.B(n_464),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_457),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_451),
.B(n_457),
.Y(n_464)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx8_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);


endmodule