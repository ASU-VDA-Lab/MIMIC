module fake_jpeg_28356_n_67 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_67);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_67;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;
wire n_66;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

AND2x2_ASAP7_75t_L g8 ( 
.A(n_4),
.B(n_5),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_5),
.B(n_0),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_16),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_17),
.B(n_18),
.Y(n_22)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_17),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_19),
.A2(n_20),
.B1(n_11),
.B2(n_10),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_15),
.A2(n_11),
.B1(n_12),
.B2(n_7),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_23),
.B(n_9),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_25),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_23),
.B(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_22),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_27),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_23),
.B(n_22),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_20),
.Y(n_34)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_8),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_20),
.C(n_13),
.Y(n_33)
);

MAJx2_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_28),
.C(n_20),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_35),
.B(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_39),
.Y(n_43)
);

A2O1A1O1Ixp25_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_8),
.B(n_16),
.C(n_21),
.D(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_21),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_41),
.B(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_37),
.C(n_7),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_8),
.B(n_1),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_46),
.B1(n_47),
.B2(n_21),
.Y(n_50)
);

OAI22x1_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_21),
.B1(n_7),
.B2(n_2),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_50),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_52),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_1),
.B(n_2),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_56),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_1),
.C(n_3),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_49),
.C(n_3),
.Y(n_59)
);

OAI21xp33_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_5),
.B(n_6),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_49),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_59),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_55),
.B(n_4),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_SL g63 ( 
.A(n_60),
.B(n_62),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_SL g64 ( 
.A(n_61),
.B(n_6),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_63),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_0),
.Y(n_67)
);


endmodule